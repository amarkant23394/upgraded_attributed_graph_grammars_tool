module Benchmark_testing45000(I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1295,I1303,I1311,I1319,I1327,I1335,I1343,I1351,I1359,I1367,I1375,I1383,I1391,I1399,I1407,I1415,I1423,I1431,I1439,I1447,I1455,I1463,I1471,I1479,I1487,I1495,I1503,I1511,I1519,I1527,I1535,I1543,I1551,I1559,I1567,I1575,I1583,I1591,I1599,I1607,I1615,I1623,I1631,I1639,I1647,I1655,I1663,I1671,I1679,I1687,I1695,I1703,I1711,I1719,I1727,I1735,I1743,I1751,I1759,I1767,I1775,I1783,I1791,I1799,I1807,I1815,I1823,I1831,I1839,I1847,I1855,I1863,I1871,I1879,I1887,I1895,I1903,I1911,I1919,I1927,I1935,I1943,I1951,I1959,I1967,I1975,I1983,I1991,I1999,I2007,I2015,I2023,I2031,I2039,I2047,I2055,I2063,I2071,I2079,I2087,I2095,I2103,I2111,I2119,I2127,I2135,I2143,I2151,I2159,I2167,I2175,I2183,I2191,I2199,I2207,I2215,I2223,I2231,I2239,I2247,I2255,I2263,I2271,I2279,I2287,I2295,I2303,I2311,I2319,I2327,I2335,I2343,I2351,I2359,I2367,I2375,I2383,I2391,I2399,I2407,I2415,I2423,I2431,I2439,I2447,I2455,I2463,I2471,I2479,I2487,I2495,I2503,I2511,I2519,I2527,I2535,I2543,I2551,I2559,I2567,I2575,I2583,I2591,I2599,I2607,I2615,I2623,I2631,I2639,I2647,I2655,I2663,I2671,I2679,I2687,I2695,I2702,I2709,I45930,I45918,I45927,I45936,I45915,I45933,I45924,I45939,I45912,I45921,I45909,I71081,I71096,I71078,I71093,I71075,I71072,I71087,I71084,I71090,I71099,I71069,I100797,I100812,I100794,I100809,I100791,I100788,I100803,I100800,I100806,I100815,I100785,I239169,I239148,I239175,I239178,I239163,I239166,I239160,I239154,I239172,I239157,I239151,I245119,I245098,I245125,I245128,I245113,I245116,I245110,I245104,I245122,I245107,I245101,I281454,I281439,I281436,I281433,I281451,I281448,I281427,I281430,I281457,I281442,I281445,I390644,I390641,I390635,I390665,I390638,I390662,I390659,I390656,I390650,I390653,I390647,I435011,I435014,I435008,I435017,I435023,I435026,I435005,I435035,I435032,I435020,I435029,I440791,I440794,I440788,I440797,I440803,I440806,I440785,I440815,I440812,I440800,I440809,I573865,I573868,I573850,I573871,I573862,I573853,I573844,I573874,I573859,I573856,I573847,I581588,I581585,I581579,I581606,I581597,I581591,I581594,I581609,I581603,I581600,I581582,I629427,I629400,I629421,I629406,I629403,I629409,I629415,I629430,I629418,I629424,I629412,I640749,I640722,I640743,I640728,I640725,I640731,I640737,I640752,I640740,I640746,I640734,I680376,I680349,I680370,I680355,I680352,I680358,I680364,I680379,I680367,I680373,I680361,I691545,I691533,I691536,I691521,I691527,I691539,I691548,I691518,I691542,I691530,I691524,I692123,I692111,I692114,I692099,I692105,I692117,I692126,I692096,I692120,I692108,I692102,I714665,I714653,I714656,I714641,I714647,I714659,I714668,I714638,I714662,I714650,I714644);
input I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1295,I1303,I1311,I1319,I1327,I1335,I1343,I1351,I1359,I1367,I1375,I1383,I1391,I1399,I1407,I1415,I1423,I1431,I1439,I1447,I1455,I1463,I1471,I1479,I1487,I1495,I1503,I1511,I1519,I1527,I1535,I1543,I1551,I1559,I1567,I1575,I1583,I1591,I1599,I1607,I1615,I1623,I1631,I1639,I1647,I1655,I1663,I1671,I1679,I1687,I1695,I1703,I1711,I1719,I1727,I1735,I1743,I1751,I1759,I1767,I1775,I1783,I1791,I1799,I1807,I1815,I1823,I1831,I1839,I1847,I1855,I1863,I1871,I1879,I1887,I1895,I1903,I1911,I1919,I1927,I1935,I1943,I1951,I1959,I1967,I1975,I1983,I1991,I1999,I2007,I2015,I2023,I2031,I2039,I2047,I2055,I2063,I2071,I2079,I2087,I2095,I2103,I2111,I2119,I2127,I2135,I2143,I2151,I2159,I2167,I2175,I2183,I2191,I2199,I2207,I2215,I2223,I2231,I2239,I2247,I2255,I2263,I2271,I2279,I2287,I2295,I2303,I2311,I2319,I2327,I2335,I2343,I2351,I2359,I2367,I2375,I2383,I2391,I2399,I2407,I2415,I2423,I2431,I2439,I2447,I2455,I2463,I2471,I2479,I2487,I2495,I2503,I2511,I2519,I2527,I2535,I2543,I2551,I2559,I2567,I2575,I2583,I2591,I2599,I2607,I2615,I2623,I2631,I2639,I2647,I2655,I2663,I2671,I2679,I2687,I2695,I2702,I2709;
output I45930,I45918,I45927,I45936,I45915,I45933,I45924,I45939,I45912,I45921,I45909,I71081,I71096,I71078,I71093,I71075,I71072,I71087,I71084,I71090,I71099,I71069,I100797,I100812,I100794,I100809,I100791,I100788,I100803,I100800,I100806,I100815,I100785,I239169,I239148,I239175,I239178,I239163,I239166,I239160,I239154,I239172,I239157,I239151,I245119,I245098,I245125,I245128,I245113,I245116,I245110,I245104,I245122,I245107,I245101,I281454,I281439,I281436,I281433,I281451,I281448,I281427,I281430,I281457,I281442,I281445,I390644,I390641,I390635,I390665,I390638,I390662,I390659,I390656,I390650,I390653,I390647,I435011,I435014,I435008,I435017,I435023,I435026,I435005,I435035,I435032,I435020,I435029,I440791,I440794,I440788,I440797,I440803,I440806,I440785,I440815,I440812,I440800,I440809,I573865,I573868,I573850,I573871,I573862,I573853,I573844,I573874,I573859,I573856,I573847,I581588,I581585,I581579,I581606,I581597,I581591,I581594,I581609,I581603,I581600,I581582,I629427,I629400,I629421,I629406,I629403,I629409,I629415,I629430,I629418,I629424,I629412,I640749,I640722,I640743,I640728,I640725,I640731,I640737,I640752,I640740,I640746,I640734,I680376,I680349,I680370,I680355,I680352,I680358,I680364,I680379,I680367,I680373,I680361,I691545,I691533,I691536,I691521,I691527,I691539,I691548,I691518,I691542,I691530,I691524,I692123,I692111,I692114,I692099,I692105,I692117,I692126,I692096,I692120,I692108,I692102,I714665,I714653,I714656,I714641,I714647,I714659,I714668,I714638,I714662,I714650,I714644;
wire I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1295,I1303,I1311,I1319,I1327,I1335,I1343,I1351,I1359,I1367,I1375,I1383,I1391,I1399,I1407,I1415,I1423,I1431,I1439,I1447,I1455,I1463,I1471,I1479,I1487,I1495,I1503,I1511,I1519,I1527,I1535,I1543,I1551,I1559,I1567,I1575,I1583,I1591,I1599,I1607,I1615,I1623,I1631,I1639,I1647,I1655,I1663,I1671,I1679,I1687,I1695,I1703,I1711,I1719,I1727,I1735,I1743,I1751,I1759,I1767,I1775,I1783,I1791,I1799,I1807,I1815,I1823,I1831,I1839,I1847,I1855,I1863,I1871,I1879,I1887,I1895,I1903,I1911,I1919,I1927,I1935,I1943,I1951,I1959,I1967,I1975,I1983,I1991,I1999,I2007,I2015,I2023,I2031,I2039,I2047,I2055,I2063,I2071,I2079,I2087,I2095,I2103,I2111,I2119,I2127,I2135,I2143,I2151,I2159,I2167,I2175,I2183,I2191,I2199,I2207,I2215,I2223,I2231,I2239,I2247,I2255,I2263,I2271,I2279,I2287,I2295,I2303,I2311,I2319,I2327,I2335,I2343,I2351,I2359,I2367,I2375,I2383,I2391,I2399,I2407,I2415,I2423,I2431,I2439,I2447,I2455,I2463,I2471,I2479,I2487,I2495,I2503,I2511,I2519,I2527,I2535,I2543,I2551,I2559,I2567,I2575,I2583,I2591,I2599,I2607,I2615,I2623,I2631,I2639,I2647,I2655,I2663,I2671,I2679,I2687,I2695,I2702,I2709,I2750,I2767,I109204,I109207,I2784,I109189,I2801,I2818,I2835,I109186,I2733,I2721,I2880,I109210,I2897,I2914,I109195,I109201,I2931,I109213,I2948,I2730,I2979,I2996,I3013,I109192,I3030,I109183,I2739,I2718,I3075,I109198,I3092,I2736,I3123,I2727,I2742,I3168,I3185,I3202,I3219,I2715,I2724,I2712,I3311,I3328,I554212,I554215,I3345,I554227,I3362,I3379,I3396,I554221,I3294,I3282,I3441,I554224,I3458,I3475,I554218,I554236,I3492,I554239,I3509,I3291,I3540,I3557,I3574,I554209,I3591,I554230,I3300,I3279,I3636,I554233,I3653,I3297,I3684,I3288,I3303,I3729,I3746,I3763,I3780,I3276,I3285,I3273,I3872,I3889,I484147,I484144,I3906,I484138,I3923,I3940,I3957,I484150,I3855,I3843,I4002,I484162,I4019,I4036,I484153,I484135,I4053,I484165,I4070,I3852,I4101,I4118,I4135,I484141,I4152,I484159,I3861,I3840,I4197,I484156,I4214,I3858,I4245,I3849,I3864,I4290,I4307,I4324,I4341,I3837,I3846,I3834,I4433,I4450,I199224,I199221,I4467,I199218,I4484,I4501,I4518,I199242,I4416,I4404,I4563,I199236,I4580,I4597,I199215,I199227,I4614,I199230,I4631,I4413,I4662,I4679,I4696,I199239,I4713,I199245,I4422,I4401,I4758,I199233,I4775,I4419,I4806,I4410,I4425,I4851,I4868,I4885,I4902,I4398,I4407,I4395,I4994,I5011,I386143,I386134,I5028,I386137,I5045,I5062,I5079,I386113,I4977,I4965,I5124,I386128,I5141,I5158,I386116,I386131,I5175,I386125,I5192,I4974,I5223,I5240,I5257,I386140,I5274,I386119,I4983,I4962,I5319,I386122,I5336,I4980,I5367,I4971,I4986,I5412,I5429,I5446,I5463,I4959,I4968,I4956,I5555,I5572,I282114,I282105,I5589,I282120,I5606,I5623,I5640,I282090,I5538,I5526,I5685,I282093,I5702,I5719,I282111,I282108,I5736,I282096,I5753,I5535,I5784,I5801,I5818,I282117,I5835,I282102,I5544,I5523,I5880,I282099,I5897,I5541,I5928,I5532,I5547,I5973,I5990,I6007,I6024,I5520,I5529,I5517,I6116,I6133,I74966,I74969,I6150,I74951,I6167,I6184,I6201,I74948,I6099,I6087,I6246,I74972,I6263,I6280,I74957,I74963,I6297,I74975,I6314,I6096,I6345,I6362,I6379,I74954,I6396,I74945,I6105,I6084,I6441,I74960,I6458,I6102,I6489,I6093,I6108,I6534,I6551,I6568,I6585,I6081,I6090,I6078,I6677,I6694,I621852,I621855,I6711,I621861,I6728,I6745,I6762,I621873,I6660,I6648,I6807,I621882,I6824,I6841,I621870,I621867,I6858,I621879,I6875,I6657,I6906,I6923,I6940,I621876,I6957,I621864,I6666,I6645,I7002,I621858,I7019,I6663,I7050,I6654,I6669,I7095,I7112,I7129,I7146,I6642,I6651,I6639,I7238,I7255,I432705,I432702,I7272,I432696,I7289,I7306,I7323,I432708,I7221,I7209,I7368,I432720,I7385,I7402,I432711,I432693,I7419,I432723,I7436,I7218,I7467,I7484,I7501,I432699,I7518,I432717,I7227,I7206,I7563,I432714,I7580,I7224,I7611,I7215,I7230,I7656,I7673,I7690,I7707,I7203,I7212,I7200,I7799,I7816,I586955,I586943,I7833,I586940,I7850,I7867,I7884,I586961,I7782,I7770,I7929,I586964,I7946,I7963,I586934,I586952,I7980,I586949,I7997,I7779,I8028,I8045,I8062,I586958,I8079,I586946,I7788,I7767,I8124,I586937,I8141,I7785,I8172,I7776,I7791,I8217,I8234,I8251,I8268,I7764,I7773,I7761,I8360,I8377,I624997,I625000,I8394,I625006,I8411,I8428,I8445,I625018,I8343,I8331,I8490,I625027,I8507,I8524,I625015,I625012,I8541,I625024,I8558,I8340,I8589,I8606,I8623,I625021,I8640,I625009,I8349,I8328,I8685,I625003,I8702,I8346,I8733,I8337,I8352,I8778,I8795,I8812,I8829,I8325,I8334,I8322,I8921,I8938,I142206,I142203,I8955,I142200,I8972,I8989,I9006,I142224,I8904,I8892,I9051,I142218,I9068,I9085,I142197,I142209,I9102,I142212,I9119,I8901,I9150,I9167,I9184,I142221,I9201,I142227,I8910,I8889,I9246,I142215,I9263,I8907,I9294,I8898,I8913,I9339,I9356,I9373,I9390,I8886,I8895,I8883,I9482,I9499,I54294,I54297,I9516,I54279,I9533,I9550,I9567,I54276,I9465,I9453,I9612,I54300,I9629,I9646,I54285,I54291,I9663,I54303,I9680,I9462,I9711,I9728,I9745,I54282,I9762,I54273,I9471,I9450,I9807,I54288,I9824,I9468,I9855,I9459,I9474,I9900,I9917,I9934,I9951,I9447,I9456,I9444,I10043,I10060,I721005,I721026,I10077,I721014,I10094,I10111,I10128,I721020,I10026,I10014,I10173,I721008,I10190,I10207,I720999,I721017,I10224,I721011,I10241,I10023,I10272,I10289,I10306,I721023,I10323,I720996,I10032,I10011,I10368,I721002,I10385,I10029,I10416,I10020,I10035,I10461,I10478,I10495,I10512,I10008,I10017,I10005,I10604,I10621,I497935,I497929,I10638,I497920,I10655,I10672,I10689,I497911,I10587,I10575,I10734,I497926,I10751,I10768,I497917,I497932,I10785,I497914,I10802,I10584,I10833,I10850,I10867,I497923,I10884,I497905,I10593,I10572,I10929,I497908,I10946,I10590,I10977,I10581,I10596,I11022,I11039,I11056,I11073,I10569,I10578,I10566,I11165,I11182,I321894,I321885,I11199,I321900,I11216,I11233,I11250,I321870,I11148,I11136,I11295,I321873,I11312,I11329,I321891,I321888,I11346,I321876,I11363,I11145,I11394,I11411,I11428,I321897,I11445,I321882,I11154,I11133,I11490,I321879,I11507,I11151,I11538,I11142,I11157,I11583,I11600,I11617,I11634,I11130,I11139,I11127,I11726,I11743,I689793,I689814,I11760,I689802,I11777,I11794,I11811,I689808,I11709,I11697,I11856,I689796,I11873,I11890,I689787,I689805,I11907,I689799,I11924,I11706,I11955,I11972,I11989,I689811,I12006,I689784,I11715,I11694,I12051,I689790,I12068,I11712,I12099,I11703,I11718,I12144,I12161,I12178,I12195,I11691,I11700,I11688,I12287,I12304,I227855,I227849,I12321,I227843,I12338,I12355,I12372,I227870,I12270,I12258,I12417,I227867,I12434,I12451,I227873,I227861,I12468,I227858,I12485,I12267,I12516,I12533,I12550,I227846,I12567,I227864,I12276,I12255,I12612,I227852,I12629,I12273,I12660,I12264,I12279,I12705,I12722,I12739,I12756,I12252,I12261,I12249,I12848,I12865,I374515,I374506,I12882,I374509,I12899,I12916,I12933,I374485,I12831,I12819,I12978,I374500,I12995,I13012,I374488,I374503,I13029,I374497,I13046,I12828,I13077,I13094,I13111,I374512,I13128,I374491,I12837,I12816,I13173,I374494,I13190,I12834,I13221,I12825,I12840,I13266,I13283,I13300,I13317,I12813,I12822,I12810,I13409,I13426,I523867,I523870,I13443,I523882,I13460,I13477,I13494,I523876,I13392,I13380,I13539,I523879,I13556,I13573,I523873,I523891,I13590,I523894,I13607,I13389,I13638,I13655,I13672,I523864,I13689,I523885,I13398,I13377,I13734,I523888,I13751,I13395,I13782,I13386,I13401,I13827,I13844,I13861,I13878,I13374,I13383,I13371,I13970,I13987,I408753,I408744,I14004,I408747,I14021,I14038,I14055,I408723,I13953,I13941,I14100,I408738,I14117,I14134,I408726,I408741,I14151,I408735,I14168,I13950,I14199,I14216,I14233,I408750,I14250,I408729,I13959,I13938,I14295,I408732,I14312,I13956,I14343,I13947,I13962,I14388,I14405,I14422,I14439,I13935,I13944,I13932,I14531,I14548,I538147,I538150,I14565,I538162,I14582,I14599,I14616,I538156,I14514,I14502,I14661,I538159,I14678,I14695,I538153,I538171,I14712,I538174,I14729,I14511,I14760,I14777,I14794,I538144,I14811,I538165,I14520,I14499,I14856,I538168,I14873,I14517,I14904,I14508,I14523,I14949,I14966,I14983,I15000,I14496,I14505,I14493,I15092,I15109,I404877,I404868,I15126,I404871,I15143,I15160,I15177,I404847,I15075,I15063,I15222,I404862,I15239,I15256,I404850,I404865,I15273,I404859,I15290,I15072,I15321,I15338,I15355,I404874,I15372,I404853,I15081,I15060,I15417,I404856,I15434,I15078,I15465,I15069,I15084,I15510,I15527,I15544,I15561,I15057,I15066,I15054,I15653,I15670,I15687,I15704,I15721,I15738,I15636,I15624,I15783,I15800,I15817,I15834,I15851,I15633,I15882,I15899,I15916,I15933,I15642,I15621,I15978,I15995,I15639,I16026,I15630,I15645,I16071,I16088,I16105,I16122,I15618,I15627,I15615,I16214,I16231,I264213,I264204,I16248,I264219,I16265,I16282,I16299,I264189,I16197,I16185,I16344,I264192,I16361,I16378,I264210,I264207,I16395,I264195,I16412,I16194,I16443,I16460,I16477,I264216,I16494,I264201,I16203,I16182,I16539,I264198,I16556,I16200,I16587,I16191,I16206,I16632,I16649,I16666,I16683,I16179,I16188,I16176,I16775,I16792,I382267,I382258,I16809,I382261,I16826,I16843,I16860,I382237,I16758,I16746,I16905,I382252,I16922,I16939,I382240,I382255,I16956,I382249,I16973,I16755,I17004,I17021,I17038,I382264,I17055,I382243,I16764,I16743,I17100,I382246,I17117,I16761,I17148,I16752,I16767,I17193,I17210,I17227,I17244,I16740,I16749,I16737,I17336,I17353,I156792,I156789,I17370,I156786,I17387,I17404,I17421,I156810,I17319,I17307,I17466,I156804,I17483,I17500,I156783,I156795,I17517,I156798,I17534,I17316,I17565,I17582,I17599,I156807,I17616,I156813,I17325,I17304,I17661,I156801,I17678,I17322,I17709,I17313,I17328,I17754,I17771,I17788,I17805,I17301,I17310,I17298,I17897,I17914,I454091,I454088,I17931,I454082,I17948,I17965,I17982,I454094,I17880,I17868,I18027,I454106,I18044,I18061,I454097,I454079,I18078,I454109,I18095,I17877,I18126,I18143,I18160,I454085,I18177,I454103,I17886,I17865,I18222,I454100,I18239,I17883,I18270,I17874,I17889,I18315,I18332,I18349,I18366,I17862,I17871,I17859,I18458,I18475,I212397,I212400,I18492,I212394,I18509,I18526,I18543,I212385,I18441,I18429,I18588,I212373,I18605,I18622,I212382,I212376,I18639,I212388,I18656,I18438,I18687,I18704,I18721,I212403,I18738,I212391,I18447,I18426,I18783,I212379,I18800,I18444,I18831,I18435,I18450,I18876,I18893,I18910,I18927,I18423,I18432,I18420,I19019,I19036,I470275,I470272,I19053,I470266,I19070,I19087,I19104,I470278,I19002,I18990,I19149,I470290,I19166,I19183,I470281,I470263,I19200,I470293,I19217,I18999,I19248,I19265,I19282,I470269,I19299,I470287,I19008,I18987,I19344,I470284,I19361,I19005,I19392,I18996,I19011,I19437,I19454,I19471,I19488,I18984,I18993,I18981,I19580,I19597,I692683,I692704,I19614,I692692,I19631,I19648,I19665,I692698,I19563,I19551,I19710,I692686,I19727,I19744,I692677,I692695,I19761,I692689,I19778,I19560,I19809,I19826,I19843,I692701,I19860,I692674,I19569,I19548,I19905,I692680,I19922,I19566,I19953,I19557,I19572,I19998,I20015,I20032,I20049,I19545,I19554,I19542,I20141,I20158,I227272,I227275,I20175,I227269,I20192,I20209,I20226,I227260,I20124,I20112,I20271,I227248,I20288,I20305,I227257,I227251,I20322,I227263,I20339,I20121,I20370,I20387,I20404,I227278,I20421,I227266,I20130,I20109,I20466,I227254,I20483,I20127,I20514,I20118,I20133,I20559,I20576,I20593,I20610,I20106,I20115,I20103,I20702,I20719,I719271,I719292,I20736,I719280,I20753,I20770,I20787,I719286,I20685,I20673,I20832,I719274,I20849,I20866,I719265,I719283,I20883,I719277,I20900,I20682,I20931,I20948,I20965,I719289,I20982,I719262,I20691,I20670,I21027,I719268,I21044,I20688,I21075,I20679,I20694,I21120,I21137,I21154,I21171,I20667,I20676,I20664,I21263,I21280,I288744,I288735,I21297,I288750,I21314,I21331,I21348,I288720,I21246,I21234,I21393,I288723,I21410,I21427,I288741,I288738,I21444,I288726,I21461,I21243,I21492,I21509,I21526,I288747,I21543,I288732,I21252,I21231,I21588,I288729,I21605,I21249,I21636,I21240,I21255,I21681,I21698,I21715,I21732,I21228,I21237,I21225,I21824,I21841,I591715,I591703,I21858,I591700,I21875,I21892,I21909,I591721,I21807,I21795,I21954,I591724,I21971,I21988,I591694,I591712,I22005,I591709,I22022,I21804,I22053,I22070,I22087,I591718,I22104,I591706,I21813,I21792,I22149,I591697,I22166,I21810,I22197,I21801,I21816,I22242,I22259,I22276,I22293,I21789,I21798,I21786,I22385,I22402,I525057,I525060,I22419,I525072,I22436,I22453,I22470,I525066,I22368,I22356,I22515,I525069,I22532,I22549,I525063,I525081,I22566,I525084,I22583,I22365,I22614,I22631,I22648,I525054,I22665,I525075,I22374,I22353,I22710,I525078,I22727,I22371,I22758,I22362,I22377,I22803,I22820,I22837,I22854,I22350,I22359,I22347,I22946,I22963,I303330,I303321,I22980,I303336,I22997,I23014,I23031,I303306,I22929,I22917,I23076,I303309,I23093,I23110,I303327,I303324,I23127,I303312,I23144,I22926,I23175,I23192,I23209,I303333,I23226,I303318,I22935,I22914,I23271,I303315,I23288,I22932,I23319,I22923,I22938,I23364,I23381,I23398,I23415,I22911,I22920,I22908,I23507,I23524,I517322,I517325,I23541,I517337,I23558,I23575,I23592,I517331,I23490,I23478,I23637,I517334,I23654,I23671,I517328,I517346,I23688,I517349,I23705,I23487,I23736,I23753,I23770,I517319,I23787,I517340,I23496,I23475,I23832,I517343,I23849,I23493,I23880,I23484,I23499,I23925,I23942,I23959,I23976,I23472,I23481,I23469,I24068,I24085,I377745,I377736,I24102,I377739,I24119,I24136,I24153,I377715,I24051,I24039,I24198,I377730,I24215,I24232,I377718,I377733,I24249,I377727,I24266,I24048,I24297,I24314,I24331,I377742,I24348,I377721,I24057,I24036,I24393,I377724,I24410,I24054,I24441,I24045,I24060,I24486,I24503,I24520,I24537,I24033,I24042,I24030,I24629,I24646,I131168,I131171,I24663,I131153,I24680,I24697,I24714,I131150,I24612,I24600,I24759,I131174,I24776,I24793,I131159,I131165,I24810,I131177,I24827,I24609,I24858,I24875,I24892,I131156,I24909,I131147,I24618,I24597,I24954,I131162,I24971,I24615,I25002,I24606,I24621,I25047,I25064,I25081,I25098,I24594,I24603,I24591,I25190,I25207,I146847,I146844,I25224,I146841,I25241,I25258,I25275,I146865,I25173,I25161,I25320,I146859,I25337,I25354,I146838,I146850,I25371,I146853,I25388,I25170,I25419,I25436,I25453,I146862,I25470,I146868,I25179,I25158,I25515,I146856,I25532,I25176,I25563,I25167,I25182,I25608,I25625,I25642,I25659,I25155,I25164,I25152,I25751,I25768,I694417,I694438,I25785,I694426,I25802,I25819,I25836,I694432,I25734,I25722,I25881,I694420,I25898,I25915,I694411,I694429,I25932,I694423,I25949,I25731,I25980,I25997,I26014,I694435,I26031,I694408,I25740,I25719,I26076,I694414,I26093,I25737,I26124,I25728,I25743,I26169,I26186,I26203,I26220,I25716,I25725,I25713,I26312,I26329,I205257,I205260,I26346,I205254,I26363,I26380,I26397,I205245,I26295,I26283,I26442,I205233,I26459,I26476,I205242,I205236,I26493,I205248,I26510,I26292,I26541,I26558,I26575,I205263,I26592,I205251,I26301,I26280,I26637,I205239,I26654,I26298,I26685,I26289,I26304,I26730,I26747,I26764,I26781,I26277,I26286,I26274,I26873,I26890,I350613,I350604,I26907,I350607,I26924,I26941,I26958,I350583,I26856,I26844,I27003,I350598,I27020,I27037,I350586,I350601,I27054,I350595,I27071,I26853,I27102,I27119,I27136,I350610,I27153,I350589,I26862,I26841,I27198,I350592,I27215,I26859,I27246,I26850,I26865,I27291,I27308,I27325,I27342,I26838,I26847,I26835,I27434,I27451,I635690,I635693,I27468,I635699,I27485,I27502,I27519,I635711,I27417,I27405,I27564,I635720,I27581,I27598,I635708,I635705,I27615,I635717,I27632,I27414,I27663,I27680,I27697,I635714,I27714,I635702,I27423,I27402,I27759,I635696,I27776,I27420,I27807,I27411,I27426,I27852,I27869,I27886,I27903,I27399,I27408,I27396,I27995,I28012,I422990,I422984,I28029,I422996,I28046,I28063,I28080,I422993,I27978,I27966,I28125,I422972,I28142,I28159,I422978,I422987,I28176,I422975,I28193,I27975,I28224,I28241,I28258,I422999,I28275,I422969,I27984,I27963,I28320,I422981,I28337,I27981,I28368,I27972,I27987,I28413,I28430,I28447,I28464,I27960,I27969,I27957,I28556,I28573,I316590,I316581,I28590,I316596,I28607,I28624,I28641,I316566,I28539,I28527,I28686,I316569,I28703,I28720,I316587,I316584,I28737,I316572,I28754,I28536,I28785,I28802,I28819,I316593,I28836,I316578,I28545,I28524,I28881,I316575,I28898,I28542,I28929,I28533,I28548,I28974,I28991,I29008,I29025,I28521,I28530,I28518,I29117,I29134,I700197,I700218,I29151,I700206,I29168,I29185,I29202,I700212,I29100,I29088,I29247,I700200,I29264,I29281,I700191,I700209,I29298,I700203,I29315,I29097,I29346,I29363,I29380,I700215,I29397,I700188,I29106,I29085,I29442,I700194,I29459,I29103,I29490,I29094,I29109,I29535,I29552,I29569,I29586,I29082,I29091,I29079,I29678,I29695,I230235,I230229,I29712,I230223,I29729,I29746,I29763,I230250,I29661,I29649,I29808,I230247,I29825,I29842,I230253,I230241,I29859,I230238,I29876,I29658,I29907,I29924,I29941,I230226,I29958,I230244,I29667,I29646,I30003,I230232,I30020,I29664,I30051,I29655,I29670,I30096,I30113,I30130,I30147,I29643,I29652,I29640,I30239,I30256,I448311,I448308,I30273,I448302,I30290,I30307,I30324,I448314,I30222,I30210,I30369,I448326,I30386,I30403,I448317,I448299,I30420,I448329,I30437,I30219,I30468,I30485,I30502,I448305,I30519,I448323,I30228,I30207,I30564,I448320,I30581,I30225,I30612,I30216,I30231,I30657,I30674,I30691,I30708,I30204,I30213,I30201,I30800,I30817,I94992,I94995,I30834,I94977,I30851,I30868,I30885,I94974,I30783,I30771,I30930,I94998,I30947,I30964,I94983,I94989,I30981,I95001,I30998,I30780,I31029,I31046,I31063,I94980,I31080,I94971,I30789,I30768,I31125,I94986,I31142,I30786,I31173,I30777,I30792,I31218,I31235,I31252,I31269,I30765,I30774,I30762,I31361,I31378,I598855,I598843,I31395,I598840,I31412,I31429,I31446,I598861,I31344,I31332,I31491,I598864,I31508,I31525,I598834,I598852,I31542,I598849,I31559,I31341,I31590,I31607,I31624,I598858,I31641,I598846,I31350,I31329,I31686,I598837,I31703,I31347,I31734,I31338,I31353,I31779,I31796,I31813,I31830,I31326,I31335,I31323,I31922,I31939,I108558,I108561,I31956,I108543,I31973,I31990,I32007,I108540,I31905,I31893,I32052,I108564,I32069,I32086,I108549,I108555,I32103,I108567,I32120,I31902,I32151,I32168,I32185,I108546,I32202,I108537,I31911,I31890,I32247,I108552,I32264,I31908,I32295,I31899,I31914,I32340,I32357,I32374,I32391,I31887,I31896,I31884,I32483,I32500,I612540,I612528,I32517,I612525,I32534,I32551,I32568,I612546,I32466,I32454,I32613,I612549,I32630,I32647,I612519,I612537,I32664,I612534,I32681,I32463,I32712,I32729,I32746,I612543,I32763,I612531,I32472,I32451,I32808,I612522,I32825,I32469,I32856,I32460,I32475,I32901,I32918,I32935,I32952,I32448,I32457,I32445,I33044,I33061,I314601,I314592,I33078,I314607,I33095,I33112,I33129,I314577,I33027,I33015,I33174,I314580,I33191,I33208,I314598,I314595,I33225,I314583,I33242,I33024,I33273,I33290,I33307,I314604,I33324,I314589,I33033,I33012,I33369,I314586,I33386,I33030,I33417,I33021,I33036,I33462,I33479,I33496,I33513,I33009,I33018,I33006,I33605,I33622,I718693,I718714,I33639,I718702,I33656,I33673,I33690,I718708,I33588,I33576,I33735,I718696,I33752,I33769,I718687,I718705,I33786,I718699,I33803,I33585,I33834,I33851,I33868,I718711,I33885,I718684,I33594,I33573,I33930,I718690,I33947,I33591,I33978,I33582,I33597,I34023,I34040,I34057,I34074,I33570,I33579,I33567,I34166,I34183,I679091,I679094,I34200,I679100,I34217,I34234,I34251,I679112,I34149,I34137,I34296,I679121,I34313,I34330,I679109,I679106,I34347,I679118,I34364,I34146,I34395,I34412,I34429,I679115,I34446,I679103,I34155,I34134,I34491,I679097,I34508,I34152,I34539,I34143,I34158,I34584,I34601,I34618,I34635,I34131,I34140,I34128,I34727,I34744,I583385,I583373,I34761,I583370,I34778,I34795,I34812,I583391,I34710,I34698,I34857,I583394,I34874,I34891,I583364,I583382,I34908,I583379,I34925,I34707,I34956,I34973,I34990,I583388,I35007,I583376,I34716,I34695,I35052,I583367,I35069,I34713,I35100,I34704,I34719,I35145,I35162,I35179,I35196,I34692,I34701,I34689,I35288,I35305,I596475,I596463,I35322,I596460,I35339,I35356,I35373,I596481,I35271,I35259,I35418,I596484,I35435,I35452,I596454,I596472,I35469,I596469,I35486,I35268,I35517,I35534,I35551,I596478,I35568,I596466,I35277,I35256,I35613,I596457,I35630,I35274,I35661,I35265,I35280,I35706,I35723,I35740,I35757,I35253,I35262,I35250,I35849,I35866,I491951,I491933,I35883,I491942,I35900,I35917,I35934,I491927,I35832,I35820,I35979,I491936,I35996,I36013,I491924,I491930,I36030,I491939,I36047,I35829,I36078,I36095,I36112,I491948,I36129,I491921,I35838,I35817,I36174,I491945,I36191,I35835,I36222,I35826,I35841,I36267,I36284,I36301,I36318,I35814,I35823,I35811,I36410,I36427,I197235,I197232,I36444,I197229,I36461,I36478,I36495,I197253,I36393,I36381,I36540,I197247,I36557,I36574,I197226,I197238,I36591,I197241,I36608,I36390,I36639,I36656,I36673,I197250,I36690,I197256,I36399,I36378,I36735,I197244,I36752,I36396,I36783,I36387,I36402,I36828,I36845,I36862,I36879,I36375,I36384,I36372,I36971,I36988,I467385,I467382,I37005,I467376,I37022,I37039,I37056,I467388,I36954,I36942,I37101,I467400,I37118,I37135,I467391,I467373,I37152,I467403,I37169,I36951,I37200,I37217,I37234,I467379,I37251,I467397,I36960,I36939,I37296,I467394,I37313,I36957,I37344,I36948,I36963,I37389,I37406,I37423,I37440,I36936,I36945,I36933,I37532,I37549,I457559,I457556,I37566,I457550,I37583,I37600,I37617,I457562,I37515,I37503,I37662,I457574,I37679,I37696,I457565,I457547,I37713,I457577,I37730,I37512,I37761,I37778,I37795,I457553,I37812,I457571,I37521,I37500,I37857,I457568,I37874,I37518,I37905,I37509,I37524,I37950,I37967,I37984,I38001,I37497,I37506,I37494,I38093,I38110,I415646,I415640,I38127,I415652,I38144,I38161,I38178,I415649,I38076,I38064,I38223,I415628,I38240,I38257,I415634,I415643,I38274,I415631,I38291,I38073,I38322,I38339,I38356,I415655,I38373,I415625,I38082,I38061,I38418,I415637,I38435,I38079,I38466,I38070,I38085,I38511,I38528,I38545,I38562,I38058,I38067,I38055,I38654,I38671,I167400,I167397,I38688,I167394,I38705,I38722,I38739,I167418,I38637,I38625,I38784,I167412,I38801,I38818,I167391,I167403,I38835,I167406,I38852,I38634,I38883,I38900,I38917,I167415,I38934,I167421,I38643,I38622,I38979,I167409,I38996,I38640,I39027,I38631,I38646,I39072,I39089,I39106,I39123,I38619,I38628,I38616,I39215,I39232,I203472,I203475,I39249,I203469,I39266,I39283,I39300,I203460,I39198,I39186,I39345,I203448,I39362,I39379,I203457,I203451,I39396,I203463,I39413,I39195,I39444,I39461,I39478,I203478,I39495,I203466,I39204,I39183,I39540,I203454,I39557,I39201,I39588,I39192,I39207,I39633,I39650,I39667,I39684,I39180,I39189,I39177,I39776,I39793,I518512,I518515,I39810,I518527,I39827,I39844,I39861,I518521,I39759,I39747,I39906,I518524,I39923,I39940,I518518,I518536,I39957,I518539,I39974,I39756,I40005,I40022,I40039,I518509,I40056,I518530,I39765,I39744,I40101,I518533,I40118,I39762,I40149,I39753,I39768,I40194,I40211,I40228,I40245,I39741,I39750,I39738,I40337,I40354,I324546,I324537,I40371,I324552,I40388,I40405,I40422,I324522,I40320,I40308,I40467,I324525,I40484,I40501,I324543,I324540,I40518,I324528,I40535,I40317,I40566,I40583,I40600,I324549,I40617,I324534,I40326,I40305,I40662,I324531,I40679,I40323,I40710,I40314,I40329,I40755,I40772,I40789,I40806,I40302,I40311,I40299,I40898,I40915,I243920,I243914,I40932,I243908,I40949,I40966,I40983,I243935,I40881,I40869,I41028,I243932,I41045,I41062,I243938,I243926,I41079,I243923,I41096,I40878,I41127,I41144,I41161,I243911,I41178,I243929,I40887,I40866,I41223,I243917,I41240,I40884,I41271,I40875,I40890,I41316,I41333,I41350,I41367,I40863,I40872,I40860,I41459,I41476,I501981,I501975,I41493,I501966,I41510,I41527,I41544,I501957,I41442,I41430,I41589,I501972,I41606,I41623,I501963,I501978,I41640,I501960,I41657,I41439,I41688,I41705,I41722,I501969,I41739,I501951,I41448,I41427,I41784,I501954,I41801,I41445,I41832,I41436,I41451,I41877,I41894,I41911,I41928,I41424,I41433,I41421,I42020,I42037,I589930,I589918,I42054,I589915,I42071,I42088,I42105,I589936,I42003,I41991,I42150,I589939,I42167,I42184,I589909,I589927,I42201,I589924,I42218,I42000,I42249,I42266,I42283,I589933,I42300,I589921,I42009,I41988,I42345,I589912,I42362,I42006,I42393,I41997,I42012,I42438,I42455,I42472,I42489,I41985,I41994,I41982,I42581,I42598,I698463,I698484,I42615,I698472,I42632,I42649,I42666,I698478,I42564,I42552,I42711,I698466,I42728,I42745,I698457,I698475,I42762,I698469,I42779,I42561,I42810,I42827,I42844,I698481,I42861,I698454,I42570,I42549,I42906,I698460,I42923,I42567,I42954,I42558,I42573,I42999,I43016,I43033,I43050,I42546,I42555,I42543,I43142,I43159,I666511,I666514,I43176,I666520,I43193,I43210,I43227,I666532,I43125,I43113,I43272,I666541,I43289,I43306,I666529,I666526,I43323,I666538,I43340,I43122,I43371,I43388,I43405,I666535,I43422,I666523,I43131,I43110,I43467,I666517,I43484,I43128,I43515,I43119,I43134,I43560,I43577,I43594,I43611,I43107,I43116,I43104,I43703,I43720,I159444,I159441,I43737,I159438,I43754,I43771,I43788,I159462,I43686,I43674,I43833,I159456,I43850,I43867,I159435,I159447,I43884,I159450,I43901,I43683,I43932,I43949,I43966,I159459,I43983,I159465,I43692,I43671,I44028,I159453,I44045,I43689,I44076,I43680,I43695,I44121,I44138,I44155,I44172,I43668,I43677,I43665,I44264,I44281,I424826,I424820,I44298,I424832,I44315,I44332,I44349,I424829,I44247,I44235,I44394,I424808,I44411,I44428,I424814,I424823,I44445,I424811,I44462,I44244,I44493,I44510,I44527,I424835,I44544,I424805,I44253,I44232,I44589,I424817,I44606,I44250,I44637,I44241,I44256,I44682,I44699,I44716,I44733,I44229,I44238,I44226,I44825,I44842,I331839,I331830,I44859,I331845,I44876,I44893,I44910,I331815,I44808,I44796,I44955,I331818,I44972,I44989,I331836,I331833,I45006,I331821,I45023,I44805,I45054,I45071,I45088,I331842,I45105,I331827,I44814,I44793,I45150,I331824,I45167,I44811,I45198,I44802,I44817,I45243,I45260,I45277,I45294,I44790,I44799,I44787,I45386,I45403,I587550,I587538,I45420,I587535,I45437,I45454,I45471,I587556,I45369,I45357,I45516,I587559,I45533,I45550,I587529,I587547,I45567,I587544,I45584,I45366,I45615,I45632,I45649,I587553,I45666,I587541,I45375,I45354,I45711,I587532,I45728,I45372,I45759,I45363,I45378,I45804,I45821,I45838,I45855,I45351,I45360,I45348,I45947,I45964,I499669,I499663,I45981,I499654,I45998,I46015,I46032,I499645,I46077,I499660,I46094,I46111,I499651,I499666,I46128,I499648,I46145,I46176,I46193,I46210,I499657,I46227,I499639,I46272,I499642,I46289,I46320,I46365,I46382,I46399,I46416,I46508,I46525,I515537,I515540,I46542,I515552,I46559,I46576,I46593,I515546,I46491,I46479,I46638,I515549,I46655,I46672,I515543,I515561,I46689,I515564,I46706,I46488,I46737,I46754,I46771,I515534,I46788,I515555,I46497,I46476,I46833,I515558,I46850,I46494,I46881,I46485,I46500,I46926,I46943,I46960,I46977,I46473,I46482,I46470,I47069,I47086,I201092,I201095,I47103,I201089,I47120,I47137,I47154,I201080,I47052,I47040,I47199,I201068,I47216,I47233,I201077,I201071,I47250,I201083,I47267,I47049,I47298,I47315,I47332,I201098,I47349,I201086,I47058,I47037,I47394,I201074,I47411,I47055,I47442,I47046,I47061,I47487,I47504,I47521,I47538,I47034,I47043,I47031,I47630,I47647,I614304,I614307,I47664,I614313,I47681,I47698,I47715,I614325,I47613,I47601,I47760,I614334,I47777,I47794,I614322,I614319,I47811,I614331,I47828,I47610,I47859,I47876,I47893,I614328,I47910,I614316,I47619,I47598,I47955,I614310,I47972,I47616,I48003,I47607,I47622,I48048,I48065,I48082,I48099,I47595,I47604,I47592,I48191,I48208,I426662,I426656,I48225,I426668,I48242,I48259,I48276,I426665,I48174,I48162,I48321,I426644,I48338,I48355,I426650,I426659,I48372,I426647,I48389,I48171,I48420,I48437,I48454,I426671,I48471,I426641,I48180,I48159,I48516,I426653,I48533,I48177,I48564,I48168,I48183,I48609,I48626,I48643,I48660,I48156,I48165,I48153,I48752,I48769,I434439,I434436,I48786,I434430,I48803,I48820,I48837,I434442,I48735,I48723,I48882,I434454,I48899,I48916,I434445,I434427,I48933,I434457,I48950,I48732,I48981,I48998,I49015,I434433,I49032,I434451,I48741,I48720,I49077,I434448,I49094,I48738,I49125,I48729,I48744,I49170,I49187,I49204,I49221,I48717,I48726,I48714,I49313,I49330,I190605,I190602,I49347,I190599,I49364,I49381,I49398,I190623,I49296,I49284,I49443,I190617,I49460,I49477,I190596,I190608,I49494,I190611,I49511,I49293,I49542,I49559,I49576,I190620,I49593,I190626,I49302,I49281,I49638,I190614,I49655,I49299,I49686,I49290,I49305,I49731,I49748,I49765,I49782,I49278,I49287,I49275,I49874,I49891,I711757,I711778,I49908,I711766,I49925,I49942,I49959,I711772,I49857,I49845,I50004,I711760,I50021,I50038,I711751,I711769,I50055,I711763,I50072,I49854,I50103,I50120,I50137,I711775,I50154,I711748,I49863,I49842,I50199,I711754,I50216,I49860,I50247,I49851,I49866,I50292,I50309,I50326,I50343,I49839,I49848,I49836,I50435,I50452,I707133,I50469,I707130,I707127,I50486,I707148,I50409,I50517,I50534,I707151,I50424,I50406,I50579,I50596,I50613,I707124,I50630,I707136,I50647,I707145,I50664,I707139,I50681,I50698,I50715,I50421,I50746,I50763,I50780,I50403,I50811,I50400,I50842,I707154,I50859,I50876,I50893,I50415,I50924,I50412,I50955,I707142,I50972,I50989,I50418,I50427,I50397,I51081,I51098,I418091,I51115,I418073,I418088,I51132,I418097,I51055,I51163,I51180,I418100,I51070,I51052,I51225,I51242,I51259,I418103,I51276,I418079,I51293,I418082,I51310,I418076,I51327,I51344,I51361,I51067,I51392,I51409,I51426,I51049,I51457,I51046,I51488,I418085,I51505,I51522,I51539,I51061,I51570,I51058,I51601,I418094,I51618,I51635,I51064,I51073,I51043,I51727,I51744,I379025,I51761,I379037,I379019,I51778,I379034,I51701,I51809,I51826,I379022,I51716,I51698,I51871,I51888,I51905,I379031,I51922,I379010,I51939,I379013,I51956,I379016,I51973,I51990,I52007,I51713,I52038,I52055,I52072,I51695,I52103,I51692,I52134,I379007,I52151,I52168,I52185,I51707,I52216,I51704,I52247,I379028,I52264,I52281,I51710,I51719,I51689,I52373,I52390,I52407,I52424,I52347,I52455,I52472,I52362,I52344,I52517,I52534,I52551,I52568,I52585,I52602,I52619,I52636,I52653,I52359,I52684,I52701,I52718,I52341,I52749,I52338,I52780,I52797,I52814,I52831,I52353,I52862,I52350,I52893,I52910,I52927,I52356,I52365,I52335,I53019,I53036,I361583,I53053,I361595,I361577,I53070,I361592,I52993,I53101,I53118,I361580,I53008,I52990,I53163,I53180,I53197,I361589,I53214,I361568,I53231,I361571,I53248,I361574,I53265,I53282,I53299,I53005,I53330,I53347,I53364,I52987,I53395,I52984,I53426,I361565,I53443,I53460,I53477,I52999,I53508,I52996,I53539,I361586,I53556,I53573,I53002,I53011,I52981,I53665,I53682,I455828,I53699,I455816,I455822,I53716,I455813,I53639,I53747,I53764,I455819,I53654,I53636,I53809,I53826,I53843,I455831,I53860,I455843,I53877,I455825,I53894,I455840,I53911,I53928,I53945,I53651,I53976,I53993,I54010,I53633,I54041,I53630,I54072,I455834,I54089,I54106,I54123,I53645,I54154,I53642,I54185,I455837,I54202,I54219,I53648,I53657,I53627,I54311,I54328,I646383,I54345,I646398,I646413,I54362,I646401,I54393,I54410,I646404,I54455,I54472,I54489,I646410,I54506,I646407,I54523,I646386,I54540,I646395,I54557,I54574,I54591,I54622,I54639,I54656,I54687,I54718,I646392,I54735,I54752,I54769,I54800,I54831,I646389,I54848,I54865,I54957,I54974,I238559,I54991,I238580,I238553,I55008,I238568,I54931,I55039,I55056,I238583,I54946,I54928,I55101,I55118,I55135,I238556,I55152,I238574,I55169,I238562,I55186,I238565,I55203,I55220,I55237,I54943,I55268,I55285,I55302,I54925,I55333,I54922,I55364,I238577,I55381,I55398,I55415,I54937,I55446,I54934,I55477,I238571,I55494,I55511,I54940,I54949,I54919,I55603,I55620,I675317,I55637,I675332,I675347,I55654,I675335,I55577,I55685,I55702,I675338,I55592,I55574,I55747,I55764,I55781,I675344,I55798,I675341,I55815,I675320,I55832,I675329,I55849,I55866,I55883,I55589,I55914,I55931,I55948,I55571,I55979,I55568,I56010,I675326,I56027,I56044,I56061,I55583,I56092,I55580,I56123,I675323,I56140,I56157,I55586,I55595,I55565,I56249,I56266,I556021,I56283,I555997,I556003,I56300,I556006,I56223,I56331,I56348,I556015,I56238,I56220,I56393,I56410,I56427,I555994,I56444,I556009,I56461,I556000,I56478,I556012,I56495,I56512,I56529,I56235,I56560,I56577,I56594,I56217,I56625,I56214,I56656,I556024,I56673,I56690,I56707,I56229,I56738,I56226,I56769,I556018,I56786,I56803,I56232,I56241,I56211,I56895,I56912,I570896,I56929,I570872,I570878,I56946,I570881,I56869,I56977,I56994,I570890,I56884,I56866,I57039,I57056,I57073,I570869,I57090,I570884,I57107,I570875,I57124,I570887,I57141,I57158,I57175,I56881,I57206,I57223,I57240,I56863,I57271,I56860,I57302,I570899,I57319,I57336,I57353,I56875,I57384,I56872,I57415,I570893,I57432,I57449,I56878,I56887,I56857,I57541,I57558,I505446,I57575,I505422,I505428,I57592,I505431,I57515,I57623,I57640,I505440,I57530,I57512,I57685,I57702,I57719,I505419,I57736,I505434,I57753,I505425,I57770,I505437,I57787,I57804,I57821,I57527,I57852,I57869,I57886,I57509,I57917,I57506,I57948,I505449,I57965,I57982,I57999,I57521,I58030,I57518,I58061,I505443,I58078,I58095,I57524,I57533,I57503,I58187,I58204,I424211,I58221,I424193,I424208,I58238,I424217,I58161,I58269,I58286,I424220,I58176,I58158,I58331,I58348,I58365,I424223,I58382,I424199,I58399,I424202,I58416,I424196,I58433,I58450,I58467,I58173,I58498,I58515,I58532,I58155,I58563,I58152,I58594,I424205,I58611,I58628,I58645,I58167,I58676,I58164,I58707,I424214,I58724,I58741,I58170,I58179,I58149,I58833,I58850,I504859,I58867,I504871,I504853,I58884,I504862,I58807,I58915,I58932,I504868,I58822,I58804,I58977,I58994,I59011,I504841,I59028,I504844,I59045,I504850,I59062,I504865,I59079,I59096,I59113,I58819,I59144,I59161,I59178,I58801,I59209,I58798,I59240,I504847,I59257,I59274,I59291,I58813,I59322,I58810,I59353,I504856,I59370,I59387,I58816,I58825,I58795,I59479,I59496,I244509,I59513,I244530,I244503,I59530,I244518,I59453,I59561,I59578,I244533,I59468,I59450,I59623,I59640,I59657,I244506,I59674,I244524,I59691,I244512,I59708,I244515,I59725,I59742,I59759,I59465,I59790,I59807,I59824,I59447,I59855,I59444,I59886,I244527,I59903,I59920,I59937,I59459,I59968,I59456,I59999,I244521,I60016,I60033,I59462,I59471,I59441,I60125,I60142,I60159,I60176,I60099,I60207,I60224,I60114,I60096,I60269,I60286,I60303,I60320,I60337,I60354,I60371,I60388,I60405,I60111,I60436,I60453,I60470,I60093,I60501,I60090,I60532,I60549,I60566,I60583,I60105,I60614,I60102,I60645,I60662,I60679,I60108,I60117,I60087,I60771,I60788,I340265,I60805,I340277,I340259,I60822,I340274,I60745,I60853,I60870,I340262,I60760,I60742,I60915,I60932,I60949,I340271,I60966,I340250,I60983,I340253,I61000,I340256,I61017,I61034,I61051,I60757,I61082,I61099,I61116,I60739,I61147,I60736,I61178,I340247,I61195,I61212,I61229,I60751,I61260,I60748,I61291,I340268,I61308,I61325,I60754,I60763,I60733,I61417,I61434,I204638,I61451,I204668,I204647,I61468,I204659,I61391,I61499,I61516,I204641,I61406,I61388,I61561,I61578,I61595,I204644,I61612,I204662,I61629,I204653,I61646,I204650,I61663,I61680,I61697,I61403,I61728,I61745,I61762,I61385,I61793,I61382,I61824,I204656,I61841,I61858,I61875,I61397,I61906,I61394,I61937,I204665,I61954,I61971,I61400,I61409,I61379,I62063,I62080,I709445,I62097,I709442,I709439,I62114,I709460,I62037,I62145,I62162,I709463,I62052,I62034,I62207,I62224,I62241,I709436,I62258,I709448,I62275,I709457,I62292,I709451,I62309,I62326,I62343,I62049,I62374,I62391,I62408,I62031,I62439,I62028,I62470,I709466,I62487,I62504,I62521,I62043,I62552,I62040,I62583,I709454,I62600,I62617,I62046,I62055,I62025,I62709,I62726,I444268,I62743,I444256,I444262,I62760,I444253,I62683,I62791,I62808,I444259,I62698,I62680,I62853,I62870,I62887,I444271,I62904,I444283,I62921,I444265,I62938,I444280,I62955,I62972,I62989,I62695,I63020,I63037,I63054,I62677,I63085,I62674,I63116,I444274,I63133,I63150,I63167,I62689,I63198,I62686,I63229,I444277,I63246,I63263,I62692,I62701,I62671,I63355,I63372,I668398,I63389,I668413,I668428,I63406,I668416,I63329,I63437,I63454,I668419,I63344,I63326,I63499,I63516,I63533,I668425,I63550,I668422,I63567,I668401,I63584,I668410,I63601,I63618,I63635,I63341,I63666,I63683,I63700,I63323,I63731,I63320,I63762,I668407,I63779,I63796,I63813,I63335,I63844,I63332,I63875,I668404,I63892,I63909,I63338,I63347,I63317,I64001,I64018,I357707,I64035,I357719,I357701,I64052,I357716,I63975,I64083,I64100,I357704,I63990,I63972,I64145,I64162,I64179,I357713,I64196,I357692,I64213,I357695,I64230,I357698,I64247,I64264,I64281,I63987,I64312,I64329,I64346,I63969,I64377,I63966,I64408,I357689,I64425,I64442,I64459,I63981,I64490,I63978,I64521,I357710,I64538,I64555,I63984,I63993,I63963,I64647,I64664,I266196,I64681,I266193,I266181,I64698,I266184,I64621,I64729,I64746,I266190,I64636,I64618,I64791,I64808,I64825,I266202,I64842,I266178,I64859,I266199,I64876,I266187,I64893,I64910,I64927,I64633,I64958,I64975,I64992,I64615,I65023,I64612,I65054,I266208,I65071,I65088,I65105,I64627,I65136,I64624,I65167,I266205,I65184,I65201,I64630,I64639,I64609,I65293,I65310,I409387,I65327,I409399,I409381,I65344,I409396,I65267,I65375,I65392,I409384,I65282,I65264,I65437,I65454,I65471,I409393,I65488,I409372,I65505,I409375,I65522,I409378,I65539,I65556,I65573,I65279,I65604,I65621,I65638,I65261,I65669,I65258,I65700,I409369,I65717,I65734,I65751,I65273,I65782,I65270,I65813,I409390,I65830,I65847,I65276,I65285,I65255,I65939,I65956,I708867,I65973,I708864,I708861,I65990,I708882,I65913,I66021,I66038,I708885,I65928,I65910,I66083,I66100,I66117,I708858,I66134,I708870,I66151,I708879,I66168,I708873,I66185,I66202,I66219,I65925,I66250,I66267,I66284,I65907,I66315,I65904,I66346,I708888,I66363,I66380,I66397,I65919,I66428,I65916,I66459,I708876,I66476,I66493,I65922,I65931,I65901,I66585,I66602,I613129,I66619,I613114,I613141,I66636,I613117,I66559,I66667,I66684,I613132,I66574,I66556,I66729,I66746,I66763,I613144,I66780,I613126,I66797,I613135,I66814,I613120,I66831,I66848,I66865,I66571,I66896,I66913,I66930,I66553,I66961,I66550,I66992,I613123,I67009,I67026,I67043,I66565,I67074,I66562,I67105,I613138,I67122,I67139,I66568,I66577,I66547,I67231,I67248,I289401,I67265,I289398,I289386,I67282,I289389,I67205,I67313,I67330,I289395,I67220,I67202,I67375,I67392,I67409,I289407,I67426,I289383,I67443,I289404,I67460,I289392,I67477,I67494,I67511,I67217,I67542,I67559,I67576,I67199,I67607,I67196,I67638,I289413,I67655,I67672,I67689,I67211,I67720,I67208,I67751,I289410,I67768,I67785,I67214,I67223,I67193,I67877,I67894,I503703,I67911,I503715,I503697,I67928,I503706,I67851,I67959,I67976,I503712,I67866,I67848,I68021,I68038,I68055,I503685,I68072,I503688,I68089,I503694,I68106,I503709,I68123,I68140,I68157,I67863,I68188,I68205,I68222,I67845,I68253,I67842,I68284,I503691,I68301,I68318,I68335,I67857,I68366,I67854,I68397,I503700,I68414,I68431,I67860,I67869,I67839,I68523,I68540,I397759,I68557,I397771,I397753,I68574,I397768,I68497,I68605,I68622,I397756,I68512,I68494,I68667,I68684,I68701,I397765,I68718,I397744,I68735,I397747,I68752,I397750,I68769,I68786,I68803,I68509,I68834,I68851,I68868,I68491,I68899,I68488,I68930,I397741,I68947,I68964,I68981,I68503,I69012,I68500,I69043,I397762,I69060,I69077,I68506,I68515,I68485,I69169,I69186,I693261,I69203,I693258,I693255,I69220,I693276,I69143,I69251,I69268,I693279,I69158,I69140,I69313,I69330,I69347,I693252,I69364,I693264,I69381,I693273,I69398,I693267,I69415,I69432,I69449,I69155,I69480,I69497,I69514,I69137,I69545,I69134,I69576,I693282,I69593,I69610,I69627,I69149,I69658,I69146,I69689,I693270,I69706,I69723,I69152,I69161,I69131,I69815,I69832,I69849,I69866,I69789,I69897,I69914,I69804,I69786,I69959,I69976,I69993,I70010,I70027,I70044,I70061,I70078,I70095,I69801,I70126,I70143,I70160,I69783,I70191,I69780,I70222,I70239,I70256,I70273,I69795,I70304,I69792,I70335,I70352,I70369,I69798,I69807,I69777,I70461,I70478,I465654,I70495,I465642,I465648,I70512,I465639,I70435,I70543,I70560,I465645,I70450,I70432,I70605,I70622,I70639,I465657,I70656,I465669,I70673,I465651,I70690,I465666,I70707,I70724,I70741,I70447,I70772,I70789,I70806,I70429,I70837,I70426,I70868,I465660,I70885,I70902,I70919,I70441,I70950,I70438,I70981,I465663,I70998,I71015,I70444,I70453,I70423,I71107,I71124,I365459,I71141,I365471,I365453,I71158,I365468,I71189,I71206,I365456,I71251,I71268,I71285,I365465,I71302,I365444,I71319,I365447,I71336,I365450,I71353,I71370,I71387,I71418,I71435,I71452,I71483,I71514,I365441,I71531,I71548,I71565,I71596,I71627,I365462,I71644,I71661,I71753,I71770,I466232,I71787,I466220,I466226,I71804,I466217,I71727,I71835,I71852,I466223,I71742,I71724,I71897,I71914,I71931,I466235,I71948,I466247,I71965,I466229,I71982,I466244,I71999,I72016,I72033,I71739,I72064,I72081,I72098,I71721,I72129,I71718,I72160,I466238,I72177,I72194,I72211,I71733,I72242,I71730,I72273,I466241,I72290,I72307,I71736,I71745,I71715,I72399,I72416,I610154,I72433,I610139,I610166,I72450,I610142,I72373,I72481,I72498,I610157,I72388,I72370,I72543,I72560,I72577,I610169,I72594,I610151,I72611,I610160,I72628,I610145,I72645,I72662,I72679,I72385,I72710,I72727,I72744,I72367,I72775,I72364,I72806,I610148,I72823,I72840,I72857,I72379,I72888,I72376,I72919,I610163,I72936,I72953,I72382,I72391,I72361,I73045,I73062,I73079,I73096,I73019,I73127,I73144,I73034,I73016,I73189,I73206,I73223,I73240,I73257,I73274,I73291,I73308,I73325,I73031,I73356,I73373,I73390,I73013,I73421,I73010,I73452,I73469,I73486,I73503,I73025,I73534,I73022,I73565,I73582,I73599,I73028,I73037,I73007,I73691,I73708,I497345,I73725,I497357,I497339,I73742,I497348,I73665,I73773,I73790,I497354,I73680,I73662,I73835,I73852,I73869,I497327,I73886,I497330,I73903,I497336,I73920,I497351,I73937,I73954,I73971,I73677,I74002,I74019,I74036,I73659,I74067,I73656,I74098,I497333,I74115,I74132,I74149,I73671,I74180,I73668,I74211,I497342,I74228,I74245,I73674,I73683,I73653,I74337,I74354,I309291,I74371,I309288,I309276,I74388,I309279,I74311,I74419,I74436,I309285,I74326,I74308,I74481,I74498,I74515,I309297,I74532,I309273,I74549,I309294,I74566,I309282,I74583,I74600,I74617,I74323,I74648,I74665,I74682,I74305,I74713,I74302,I74744,I309303,I74761,I74778,I74795,I74317,I74826,I74314,I74857,I309300,I74874,I74891,I74320,I74329,I74299,I74983,I75000,I75017,I75034,I75065,I75082,I75127,I75144,I75161,I75178,I75195,I75212,I75229,I75246,I75263,I75294,I75311,I75328,I75359,I75390,I75407,I75424,I75441,I75472,I75503,I75520,I75537,I75629,I75646,I213563,I75663,I213593,I213572,I75680,I213584,I75603,I75711,I75728,I213566,I75618,I75600,I75773,I75790,I75807,I213569,I75824,I213587,I75841,I213578,I75858,I213575,I75875,I75892,I75909,I75615,I75940,I75957,I75974,I75597,I76005,I75594,I76036,I213581,I76053,I76070,I76087,I75609,I76118,I75606,I76149,I213590,I76166,I76183,I75612,I75621,I75591,I76275,I76292,I362875,I76309,I362887,I362869,I76326,I362884,I76249,I76357,I76374,I362872,I76264,I76246,I76419,I76436,I76453,I362881,I76470,I362860,I76487,I362863,I76504,I362866,I76521,I76538,I76555,I76261,I76586,I76603,I76620,I76243,I76651,I76240,I76682,I362857,I76699,I76716,I76733,I76255,I76764,I76252,I76795,I362878,I76812,I76829,I76258,I76267,I76237,I76921,I76938,I270837,I76955,I270834,I270822,I76972,I270825,I76895,I77003,I77020,I270831,I76910,I76892,I77065,I77082,I77099,I270843,I77116,I270819,I77133,I270840,I77150,I270828,I77167,I77184,I77201,I76907,I77232,I77249,I77266,I76889,I77297,I76886,I77328,I270849,I77345,I77362,I77379,I76901,I77410,I76898,I77441,I270846,I77458,I77475,I76904,I76913,I76883,I77567,I77584,I622481,I77601,I622496,I622511,I77618,I622499,I77541,I77649,I77666,I622502,I77556,I77538,I77711,I77728,I77745,I622508,I77762,I622505,I77779,I622484,I77796,I622493,I77813,I77830,I77847,I77553,I77878,I77895,I77912,I77535,I77943,I77532,I77974,I622490,I77991,I78008,I78025,I77547,I78056,I77544,I78087,I622487,I78104,I78121,I77550,I77559,I77529,I78213,I78230,I473746,I78247,I473734,I473740,I78264,I473731,I78187,I78295,I78312,I473737,I78202,I78184,I78357,I78374,I78391,I473749,I78408,I473761,I78425,I473743,I78442,I473758,I78459,I78476,I78493,I78199,I78524,I78541,I78558,I78181,I78589,I78178,I78620,I473752,I78637,I78654,I78671,I78193,I78702,I78190,I78733,I473755,I78750,I78767,I78196,I78205,I78175,I78859,I78876,I504281,I78893,I504293,I504275,I78910,I504284,I78833,I78941,I78958,I504290,I78848,I78830,I79003,I79020,I79037,I504263,I79054,I504266,I79071,I504272,I79088,I504287,I79105,I79122,I79139,I78845,I79170,I79187,I79204,I78827,I79235,I78824,I79266,I504269,I79283,I79300,I79317,I78839,I79348,I78836,I79379,I504278,I79396,I79413,I78842,I78851,I78821,I79505,I79522,I262881,I79539,I262878,I262866,I79556,I262869,I79479,I79587,I79604,I262875,I79494,I79476,I79649,I79666,I79683,I262887,I79700,I262863,I79717,I262884,I79734,I262872,I79751,I79768,I79785,I79491,I79816,I79833,I79850,I79473,I79881,I79470,I79912,I262893,I79929,I79946,I79963,I79485,I79994,I79482,I80025,I262890,I80042,I80059,I79488,I79497,I79467,I80151,I80168,I547096,I80185,I547072,I547078,I80202,I547081,I80125,I80233,I80250,I547090,I80140,I80122,I80295,I80312,I80329,I547069,I80346,I547084,I80363,I547075,I80380,I547087,I80397,I80414,I80431,I80137,I80462,I80479,I80496,I80119,I80527,I80116,I80558,I547099,I80575,I80592,I80609,I80131,I80640,I80128,I80671,I547093,I80688,I80705,I80134,I80143,I80113,I80797,I80814,I151497,I80831,I151485,I151491,I80848,I151500,I80771,I80879,I80896,I151488,I80786,I80768,I80941,I80958,I80975,I151509,I80992,I151482,I81009,I151503,I81026,I151494,I81043,I81060,I81077,I80783,I81108,I81125,I81142,I80765,I81173,I80762,I81204,I151479,I81221,I81238,I81255,I80777,I81286,I80774,I81317,I151506,I81334,I81351,I80780,I80789,I80759,I81443,I81460,I433286,I81477,I433274,I433280,I81494,I433271,I81417,I81525,I81542,I433277,I81432,I81414,I81587,I81604,I81621,I433289,I81638,I433301,I81655,I433283,I81672,I433298,I81689,I81706,I81723,I81429,I81754,I81771,I81788,I81411,I81819,I81408,I81850,I433292,I81867,I81884,I81901,I81423,I81932,I81420,I81963,I433295,I81980,I81997,I81426,I81435,I81405,I82089,I82106,I280782,I82123,I280779,I280767,I82140,I280770,I82063,I82171,I82188,I280776,I82078,I82060,I82233,I82250,I82267,I280788,I82284,I280764,I82301,I280785,I82318,I280773,I82335,I82352,I82369,I82075,I82400,I82417,I82434,I82057,I82465,I82054,I82496,I280794,I82513,I82530,I82547,I82069,I82578,I82066,I82609,I280791,I82626,I82643,I82072,I82081,I82051,I82735,I82752,I352539,I82769,I352551,I352533,I82786,I352548,I82709,I82817,I82834,I352536,I82724,I82706,I82879,I82896,I82913,I352545,I82930,I352524,I82947,I352527,I82964,I352530,I82981,I82998,I83015,I82721,I83046,I83063,I83080,I82703,I83111,I82700,I83142,I352521,I83159,I83176,I83193,I82715,I83224,I82712,I83255,I352542,I83272,I83289,I82718,I82727,I82697,I83381,I83398,I148845,I83415,I148833,I148839,I83432,I148848,I83355,I83463,I83480,I148836,I83370,I83352,I83525,I83542,I83559,I148857,I83576,I148830,I83593,I148851,I83610,I148842,I83627,I83644,I83661,I83367,I83692,I83709,I83726,I83349,I83757,I83346,I83788,I148827,I83805,I83822,I83839,I83361,I83870,I83358,I83901,I148854,I83918,I83935,I83364,I83373,I83343,I84027,I84044,I84061,I84078,I84001,I84109,I84126,I84016,I83998,I84171,I84188,I84205,I84222,I84239,I84256,I84273,I84290,I84307,I84013,I84338,I84355,I84372,I83995,I84403,I83992,I84434,I84451,I84468,I84485,I84007,I84516,I84004,I84547,I84564,I84581,I84010,I84019,I83989,I84673,I84690,I608964,I84707,I608949,I608976,I84724,I608952,I84647,I84755,I84772,I608967,I84662,I84644,I84817,I84834,I84851,I608979,I84868,I608961,I84885,I608970,I84902,I608955,I84919,I84936,I84953,I84659,I84984,I85001,I85018,I84641,I85049,I84638,I85080,I608958,I85097,I85114,I85131,I84653,I85162,I84650,I85193,I608973,I85210,I85227,I84656,I84665,I84635,I85319,I85336,I689155,I85353,I689170,I689185,I85370,I689173,I85293,I85401,I85418,I689176,I85308,I85290,I85463,I85480,I85497,I689182,I85514,I689179,I85531,I689158,I85548,I689167,I85565,I85582,I85599,I85305,I85630,I85647,I85664,I85287,I85695,I85284,I85726,I689164,I85743,I85760,I85777,I85299,I85808,I85296,I85839,I689161,I85856,I85873,I85302,I85311,I85281,I85965,I85982,I664624,I85999,I664639,I664654,I86016,I664642,I85939,I86047,I86064,I664645,I85954,I85936,I86109,I86126,I86143,I664651,I86160,I664648,I86177,I664627,I86194,I664636,I86211,I86228,I86245,I85951,I86276,I86293,I86310,I85933,I86341,I85930,I86372,I664633,I86389,I86406,I86423,I85945,I86454,I85942,I86485,I664630,I86502,I86519,I85948,I85957,I85927,I86611,I86628,I602419,I86645,I602404,I602431,I86662,I602407,I86585,I86693,I86710,I602422,I86600,I86582,I86755,I86772,I86789,I602434,I86806,I602416,I86823,I602425,I86840,I602410,I86857,I86874,I86891,I86597,I86922,I86939,I86956,I86579,I86987,I86576,I87018,I602413,I87035,I87052,I87069,I86591,I87100,I86588,I87131,I602428,I87148,I87165,I86594,I86603,I86573,I87257,I87274,I388069,I87291,I388081,I388063,I87308,I388078,I87231,I87339,I87356,I388066,I87246,I87228,I87401,I87418,I87435,I388075,I87452,I388054,I87469,I388057,I87486,I388060,I87503,I87520,I87537,I87243,I87568,I87585,I87602,I87225,I87633,I87222,I87664,I388051,I87681,I87698,I87715,I87237,I87746,I87234,I87777,I388072,I87794,I87811,I87240,I87249,I87219,I87903,I87920,I247632,I87937,I247629,I247617,I87954,I247620,I87877,I87985,I88002,I247626,I87892,I87874,I88047,I88064,I88081,I247638,I88098,I247614,I88115,I247635,I88132,I247623,I88149,I88166,I88183,I87889,I88214,I88231,I88248,I87871,I88279,I87868,I88310,I247644,I88327,I88344,I88361,I87883,I88392,I87880,I88423,I247641,I88440,I88457,I87886,I87895,I87865,I88549,I88566,I410033,I88583,I410045,I410027,I88600,I410042,I88523,I88631,I88648,I410030,I88538,I88520,I88693,I88710,I88727,I410039,I88744,I410018,I88761,I410021,I88778,I410024,I88795,I88812,I88829,I88535,I88860,I88877,I88894,I88517,I88925,I88514,I88956,I410015,I88973,I88990,I89007,I88529,I89038,I88526,I89069,I410036,I89086,I89103,I88532,I88541,I88511,I89195,I89212,I478370,I89229,I478358,I478364,I89246,I478355,I89169,I89277,I89294,I478361,I89184,I89166,I89339,I89356,I89373,I478373,I89390,I478385,I89407,I478367,I89424,I478382,I89441,I89458,I89475,I89181,I89506,I89523,I89540,I89163,I89571,I89160,I89602,I478376,I89619,I89636,I89653,I89175,I89684,I89172,I89715,I478379,I89732,I89749,I89178,I89187,I89157,I89841,I89858,I139563,I89875,I139551,I139557,I89892,I139566,I89815,I89923,I89940,I139554,I89830,I89812,I89985,I90002,I90019,I139575,I90036,I139548,I90053,I139569,I90070,I139560,I90087,I90104,I90121,I89827,I90152,I90169,I90186,I89809,I90217,I89806,I90248,I139545,I90265,I90282,I90299,I89821,I90330,I89818,I90361,I139572,I90378,I90395,I89824,I89833,I89803,I90487,I90504,I570301,I90521,I570277,I570283,I90538,I570286,I90461,I90569,I90586,I570295,I90476,I90458,I90631,I90648,I90665,I570274,I90682,I570289,I90699,I570280,I90716,I570292,I90733,I90750,I90767,I90473,I90798,I90815,I90832,I90455,I90863,I90452,I90894,I570304,I90911,I90928,I90945,I90467,I90976,I90464,I91007,I570298,I91024,I91041,I90470,I90479,I90449,I91133,I91150,I703665,I91167,I703662,I703659,I91184,I703680,I91107,I91215,I91232,I703683,I91122,I91104,I91277,I91294,I91311,I703656,I91328,I703668,I91345,I703677,I91362,I703671,I91379,I91396,I91413,I91119,I91444,I91461,I91478,I91101,I91509,I91098,I91540,I703686,I91557,I91574,I91591,I91113,I91622,I91110,I91653,I703674,I91670,I91687,I91116,I91125,I91095,I91779,I91796,I144867,I91813,I144855,I144861,I91830,I144870,I91753,I91861,I91878,I144858,I91768,I91750,I91923,I91940,I91957,I144879,I91974,I144852,I91991,I144873,I92008,I144864,I92025,I92042,I92059,I91765,I92090,I92107,I92124,I91747,I92155,I91744,I92186,I144849,I92203,I92220,I92237,I91759,I92268,I91756,I92299,I144876,I92316,I92333,I91762,I91771,I91741,I92425,I92442,I717537,I92459,I717534,I717531,I92476,I717552,I92399,I92507,I92524,I717555,I92414,I92396,I92569,I92586,I92603,I717528,I92620,I717540,I92637,I717549,I92654,I717543,I92671,I92688,I92705,I92411,I92736,I92753,I92770,I92393,I92801,I92390,I92832,I717558,I92849,I92866,I92883,I92405,I92914,I92402,I92945,I717546,I92962,I92979,I92408,I92417,I92387,I93071,I93088,I296694,I93105,I296691,I296679,I93122,I296682,I93045,I93153,I93170,I296688,I93060,I93042,I93215,I93232,I93249,I296700,I93266,I296676,I93283,I296697,I93300,I296685,I93317,I93334,I93351,I93057,I93382,I93399,I93416,I93039,I93447,I93036,I93478,I296706,I93495,I93512,I93529,I93051,I93560,I93048,I93591,I296703,I93608,I93625,I93054,I93063,I93033,I93717,I93734,I346725,I93751,I346737,I346719,I93768,I346734,I93691,I93799,I93816,I346722,I93706,I93688,I93861,I93878,I93895,I346731,I93912,I346710,I93929,I346713,I93946,I346716,I93963,I93980,I93997,I93703,I94028,I94045,I94062,I93685,I94093,I93682,I94124,I346707,I94141,I94158,I94175,I93697,I94206,I93694,I94237,I346728,I94254,I94271,I93700,I93709,I93679,I94363,I94380,I443112,I94397,I443100,I443106,I94414,I443097,I94337,I94445,I94462,I443103,I94352,I94334,I94507,I94524,I94541,I443115,I94558,I443127,I94575,I443109,I94592,I443124,I94609,I94626,I94643,I94349,I94674,I94691,I94708,I94331,I94739,I94328,I94770,I443118,I94787,I94804,I94821,I94343,I94852,I94340,I94883,I443121,I94900,I94917,I94346,I94355,I94325,I95009,I95026,I255588,I95043,I255585,I255573,I95060,I255576,I95091,I95108,I255582,I95153,I95170,I95187,I255594,I95204,I255570,I95221,I255591,I95238,I255579,I95255,I95272,I95289,I95320,I95337,I95354,I95385,I95416,I255600,I95433,I95450,I95467,I95498,I95529,I255597,I95546,I95563,I95655,I95672,I95689,I95706,I95629,I95737,I95754,I95644,I95626,I95799,I95816,I95833,I95850,I95867,I95884,I95901,I95918,I95935,I95641,I95966,I95983,I96000,I95623,I96031,I95620,I96062,I96079,I96096,I96113,I95635,I96144,I95632,I96175,I96192,I96209,I95638,I95647,I95617,I96301,I96318,I173376,I96335,I173364,I173370,I96352,I173379,I96275,I96383,I96400,I173367,I96290,I96272,I96445,I96462,I96479,I173388,I96496,I173361,I96513,I173382,I96530,I173373,I96547,I96564,I96581,I96287,I96612,I96629,I96646,I96269,I96677,I96266,I96708,I173358,I96725,I96742,I96759,I96281,I96790,I96278,I96821,I173385,I96838,I96855,I96284,I96293,I96263,I96947,I96964,I353185,I96981,I353197,I353179,I96998,I353194,I96921,I97029,I97046,I353182,I96936,I96918,I97091,I97108,I97125,I353191,I97142,I353170,I97159,I353173,I97176,I353176,I97193,I97210,I97227,I96933,I97258,I97275,I97292,I96915,I97323,I96912,I97354,I353167,I97371,I97388,I97405,I96927,I97436,I96924,I97467,I353188,I97484,I97501,I96930,I96939,I96909,I97593,I97610,I342203,I97627,I342215,I342197,I97644,I342212,I97567,I97675,I97692,I342200,I97582,I97564,I97737,I97754,I97771,I342209,I97788,I342188,I97805,I342191,I97822,I342194,I97839,I97856,I97873,I97579,I97904,I97921,I97938,I97561,I97969,I97558,I98000,I342185,I98017,I98034,I98051,I97573,I98082,I97570,I98113,I342206,I98130,I98147,I97576,I97585,I97555,I98239,I98256,I315921,I98273,I315918,I315906,I98290,I315909,I98213,I98321,I98338,I315915,I98228,I98210,I98383,I98400,I98417,I315927,I98434,I315903,I98451,I315924,I98468,I315912,I98485,I98502,I98519,I98225,I98550,I98567,I98584,I98207,I98615,I98204,I98646,I315933,I98663,I98680,I98697,I98219,I98728,I98216,I98759,I315930,I98776,I98793,I98222,I98231,I98201,I98885,I98902,I576251,I98919,I576227,I576233,I98936,I576236,I98859,I98967,I98984,I576245,I98874,I98856,I99029,I99046,I99063,I576224,I99080,I576239,I99097,I576230,I99114,I576242,I99131,I99148,I99165,I98871,I99196,I99213,I99230,I98853,I99261,I98850,I99292,I576254,I99309,I99326,I99343,I98865,I99374,I98862,I99405,I576248,I99422,I99439,I98868,I98877,I98847,I99531,I99548,I461030,I99565,I461018,I461024,I99582,I461015,I99505,I99613,I99630,I461021,I99520,I99502,I99675,I99692,I99709,I461033,I99726,I461045,I99743,I461027,I99760,I461042,I99777,I99794,I99811,I99517,I99842,I99859,I99876,I99499,I99907,I99496,I99938,I461036,I99955,I99972,I99989,I99511,I100020,I99508,I100051,I461039,I100068,I100085,I99514,I99523,I99493,I100177,I100194,I399697,I100211,I399709,I399691,I100228,I399706,I100151,I100259,I100276,I399694,I100166,I100148,I100321,I100338,I100355,I399703,I100372,I399682,I100389,I399685,I100406,I399688,I100423,I100440,I100457,I100163,I100488,I100505,I100522,I100145,I100553,I100142,I100584,I399679,I100601,I100618,I100635,I100157,I100666,I100154,I100697,I399700,I100714,I100731,I100160,I100169,I100139,I100823,I100840,I419315,I100857,I419297,I419312,I100874,I419321,I100905,I100922,I419324,I100967,I100984,I101001,I419327,I101018,I419303,I101035,I419306,I101052,I419300,I101069,I101086,I101103,I101134,I101151,I101168,I101199,I101230,I419309,I101247,I101264,I101281,I101312,I101343,I419318,I101360,I101377,I101469,I101486,I218918,I101503,I218948,I218927,I101520,I218939,I101443,I101551,I101568,I218921,I101458,I101440,I101613,I101630,I101647,I218924,I101664,I218942,I101681,I218933,I101698,I218930,I101715,I101732,I101749,I101455,I101780,I101797,I101814,I101437,I101845,I101434,I101876,I218936,I101893,I101910,I101927,I101449,I101958,I101446,I101989,I218945,I102006,I102023,I101452,I101461,I101431,I102115,I102132,I158127,I102149,I158115,I158121,I102166,I158130,I102089,I102197,I102214,I158118,I102104,I102086,I102259,I102276,I102293,I158139,I102310,I158112,I102327,I158133,I102344,I158124,I102361,I102378,I102395,I102101,I102426,I102443,I102460,I102083,I102491,I102080,I102522,I158109,I102539,I102556,I102573,I102095,I102604,I102092,I102635,I158136,I102652,I102669,I102098,I102107,I102077,I102761,I102778,I368043,I102795,I368055,I368037,I102812,I368052,I102735,I102843,I102860,I368040,I102750,I102732,I102905,I102922,I102939,I368049,I102956,I368028,I102973,I368031,I102990,I368034,I103007,I103024,I103041,I102747,I103072,I103089,I103106,I102729,I103137,I102726,I103168,I368025,I103185,I103202,I103219,I102741,I103250,I102738,I103281,I368046,I103298,I103315,I102744,I102753,I102723,I103407,I103424,I103441,I103458,I103381,I103489,I103506,I103396,I103378,I103551,I103568,I103585,I103602,I103619,I103636,I103653,I103670,I103687,I103393,I103718,I103735,I103752,I103375,I103783,I103372,I103814,I103831,I103848,I103865,I103387,I103896,I103384,I103927,I103944,I103961,I103390,I103399,I103369,I104053,I104070,I436176,I104087,I436164,I436170,I104104,I436161,I104027,I104135,I104152,I436167,I104042,I104024,I104197,I104214,I104231,I436179,I104248,I436191,I104265,I436173,I104282,I436188,I104299,I104316,I104333,I104039,I104364,I104381,I104398,I104021,I104429,I104018,I104460,I436182,I104477,I104494,I104511,I104033,I104542,I104030,I104573,I436185,I104590,I104607,I104036,I104045,I104015,I104699,I104716,I284760,I104733,I284757,I284745,I104750,I284748,I104673,I104781,I104798,I284754,I104688,I104670,I104843,I104860,I104877,I284766,I104894,I284742,I104911,I284763,I104928,I284751,I104945,I104962,I104979,I104685,I105010,I105027,I105044,I104667,I105075,I104664,I105106,I284772,I105123,I105140,I105157,I104679,I105188,I104676,I105219,I284769,I105236,I105253,I104682,I104691,I104661,I105345,I105362,I510801,I105379,I510777,I510783,I105396,I510786,I105319,I105427,I105444,I510795,I105334,I105316,I105489,I105506,I105523,I510774,I105540,I510789,I105557,I510780,I105574,I510792,I105591,I105608,I105625,I105331,I105656,I105673,I105690,I105313,I105721,I105310,I105752,I510804,I105769,I105786,I105803,I105325,I105834,I105322,I105865,I510798,I105882,I105899,I105328,I105337,I105307,I105991,I106008,I575061,I106025,I575037,I575043,I106042,I575046,I105965,I106073,I106090,I575055,I105980,I105962,I106135,I106152,I106169,I575034,I106186,I575049,I106203,I575040,I106220,I575052,I106237,I106254,I106271,I105977,I106302,I106319,I106336,I105959,I106367,I105956,I106398,I575064,I106415,I106432,I106449,I105971,I106480,I105968,I106511,I575058,I106528,I106545,I105974,I105983,I105953,I106637,I106654,I248295,I106671,I248292,I248280,I106688,I248283,I106611,I106719,I106736,I248289,I106626,I106608,I106781,I106798,I106815,I248301,I106832,I248277,I106849,I248298,I106866,I248286,I106883,I106900,I106917,I106623,I106948,I106965,I106982,I106605,I107013,I106602,I107044,I248307,I107061,I107078,I107095,I106617,I107126,I106614,I107157,I248304,I107174,I107191,I106620,I106629,I106599,I107283,I107300,I649528,I107317,I649543,I649558,I107334,I649546,I107257,I107365,I107382,I649549,I107272,I107254,I107427,I107444,I107461,I649555,I107478,I649552,I107495,I649531,I107512,I649540,I107529,I107546,I107563,I107269,I107594,I107611,I107628,I107251,I107659,I107248,I107690,I649537,I107707,I107724,I107741,I107263,I107772,I107260,I107803,I649534,I107820,I107837,I107266,I107275,I107245,I107929,I107946,I329181,I107963,I329178,I329166,I107980,I329169,I107903,I108011,I108028,I329175,I107918,I107900,I108073,I108090,I108107,I329187,I108124,I329163,I108141,I329184,I108158,I329172,I108175,I108192,I108209,I107915,I108240,I108257,I108274,I107897,I108305,I107894,I108336,I329193,I108353,I108370,I108387,I107909,I108418,I107906,I108449,I329190,I108466,I108483,I107912,I107921,I107891,I108575,I108592,I181332,I108609,I181320,I181326,I108626,I181335,I108657,I108674,I181323,I108719,I108736,I108753,I181344,I108770,I181317,I108787,I181338,I108804,I181329,I108821,I108838,I108855,I108886,I108903,I108920,I108951,I108982,I181314,I108999,I109016,I109033,I109064,I109095,I181341,I109112,I109129,I109221,I109238,I500235,I109255,I500247,I500229,I109272,I500238,I109303,I109320,I500244,I109365,I109382,I109399,I500217,I109416,I500220,I109433,I500226,I109450,I500241,I109467,I109484,I109501,I109532,I109549,I109566,I109597,I109628,I500223,I109645,I109662,I109679,I109710,I109741,I500232,I109758,I109775,I109867,I109884,I216538,I109901,I216568,I216547,I109918,I216559,I109841,I109949,I109966,I216541,I109856,I109838,I110011,I110028,I110045,I216544,I110062,I216562,I110079,I216553,I110096,I216550,I110113,I110130,I110147,I109853,I110178,I110195,I110212,I109835,I110243,I109832,I110274,I216556,I110291,I110308,I110325,I109847,I110356,I109844,I110387,I216565,I110404,I110421,I109850,I109859,I109829,I110513,I110530,I592304,I110547,I592289,I592316,I110564,I592292,I110487,I110595,I110612,I592307,I110502,I110484,I110657,I110674,I110691,I592319,I110708,I592301,I110725,I592310,I110742,I592295,I110759,I110776,I110793,I110499,I110824,I110841,I110858,I110481,I110889,I110478,I110920,I592298,I110937,I110954,I110971,I110493,I111002,I110490,I111033,I592313,I111050,I111067,I110496,I110505,I110475,I111159,I111176,I619965,I111193,I619980,I619995,I111210,I619983,I111133,I111241,I111258,I619986,I111148,I111130,I111303,I111320,I111337,I619992,I111354,I619989,I111371,I619968,I111388,I619977,I111405,I111422,I111439,I111145,I111470,I111487,I111504,I111127,I111535,I111124,I111566,I619974,I111583,I111600,I111617,I111139,I111648,I111136,I111679,I619971,I111696,I111713,I111142,I111151,I111121,I111805,I111822,I111839,I111856,I111779,I111887,I111904,I111794,I111776,I111949,I111966,I111983,I112000,I112017,I112034,I112051,I112068,I112085,I111791,I112116,I112133,I112150,I111773,I112181,I111770,I112212,I112229,I112246,I112263,I111785,I112294,I111782,I112325,I112342,I112359,I111788,I111797,I111767,I112451,I112468,I261555,I112485,I261552,I261540,I112502,I261543,I112425,I112533,I112550,I261549,I112440,I112422,I112595,I112612,I112629,I261561,I112646,I261537,I112663,I261558,I112680,I261546,I112697,I112714,I112731,I112437,I112762,I112779,I112796,I112419,I112827,I112416,I112858,I261567,I112875,I112892,I112909,I112431,I112940,I112428,I112971,I261564,I112988,I113005,I112434,I112443,I112413,I113097,I113114,I183984,I113131,I183972,I183978,I113148,I183987,I113071,I113179,I113196,I183975,I113086,I113068,I113241,I113258,I113275,I183996,I113292,I183969,I113309,I183990,I113326,I183981,I113343,I113360,I113377,I113083,I113408,I113425,I113442,I113065,I113473,I113062,I113504,I183966,I113521,I113538,I113555,I113077,I113586,I113074,I113617,I183993,I113634,I113651,I113080,I113089,I113059,I113743,I113760,I400343,I113777,I400355,I400337,I113794,I400352,I113717,I113825,I113842,I400340,I113732,I113714,I113887,I113904,I113921,I400349,I113938,I400328,I113955,I400331,I113972,I400334,I113989,I114006,I114023,I113729,I114054,I114071,I114088,I113711,I114119,I113708,I114150,I400325,I114167,I114184,I114201,I113723,I114232,I113720,I114263,I400346,I114280,I114297,I113726,I113735,I113705,I114389,I114406,I242724,I114423,I242745,I242718,I114440,I242733,I114363,I114471,I114488,I242748,I114378,I114360,I114533,I114550,I114567,I242721,I114584,I242739,I114601,I242727,I114618,I242730,I114635,I114652,I114669,I114375,I114700,I114717,I114734,I114357,I114765,I114354,I114796,I242742,I114813,I114830,I114847,I114369,I114878,I114366,I114909,I242736,I114926,I114943,I114372,I114381,I114351,I115035,I115052,I565541,I115069,I565517,I565523,I115086,I565526,I115009,I115117,I115134,I565535,I115024,I115006,I115179,I115196,I115213,I565514,I115230,I565529,I115247,I565520,I115264,I565532,I115281,I115298,I115315,I115021,I115346,I115363,I115380,I115003,I115411,I115000,I115442,I565544,I115459,I115476,I115493,I115015,I115524,I115012,I115555,I565538,I115572,I115589,I115018,I115027,I114997,I115681,I115698,I438488,I115715,I438476,I438482,I115732,I438473,I115655,I115763,I115780,I438479,I115670,I115652,I115825,I115842,I115859,I438491,I115876,I438503,I115893,I438485,I115910,I438500,I115927,I115944,I115961,I115667,I115992,I116009,I116026,I115649,I116057,I115646,I116088,I438494,I116105,I116122,I116139,I115661,I116170,I115658,I116201,I438497,I116218,I116235,I115664,I115673,I115643,I116327,I116344,I360291,I116361,I360303,I360285,I116378,I360300,I116301,I116409,I116426,I360288,I116316,I116298,I116471,I116488,I116505,I360297,I116522,I360276,I116539,I360279,I116556,I360282,I116573,I116590,I116607,I116313,I116638,I116655,I116672,I116295,I116703,I116292,I116734,I360273,I116751,I116768,I116785,I116307,I116816,I116304,I116847,I360294,I116864,I116881,I116310,I116319,I116289,I116973,I116990,I375149,I117007,I375161,I375143,I117024,I375158,I116947,I117055,I117072,I375146,I116962,I116944,I117117,I117134,I117151,I375155,I117168,I375134,I117185,I375137,I117202,I375140,I117219,I117236,I117253,I116959,I117284,I117301,I117318,I116941,I117349,I116938,I117380,I375131,I117397,I117414,I117431,I116953,I117462,I116950,I117493,I375152,I117510,I117527,I116956,I116965,I116935,I117619,I117636,I512586,I117653,I512562,I512568,I117670,I512571,I117593,I117701,I117718,I512580,I117608,I117590,I117763,I117780,I117797,I512559,I117814,I512574,I117831,I512565,I117848,I512577,I117865,I117882,I117899,I117605,I117930,I117947,I117964,I117587,I117995,I117584,I118026,I512589,I118043,I118060,I118077,I117599,I118108,I117596,I118139,I512583,I118156,I118173,I117602,I117611,I117581,I118265,I118282,I118299,I118316,I118239,I118347,I118364,I118254,I118236,I118409,I118426,I118443,I118460,I118477,I118494,I118511,I118528,I118545,I118251,I118576,I118593,I118610,I118233,I118641,I118230,I118672,I118689,I118706,I118723,I118245,I118754,I118242,I118785,I118802,I118819,I118248,I118257,I118227,I118911,I118928,I665882,I118945,I665897,I665912,I118962,I665900,I118885,I118993,I119010,I665903,I118900,I118882,I119055,I119072,I119089,I665909,I119106,I665906,I119123,I665885,I119140,I665894,I119157,I119174,I119191,I118897,I119222,I119239,I119256,I118879,I119287,I118876,I119318,I665891,I119335,I119352,I119369,I118891,I119400,I118888,I119431,I665888,I119448,I119465,I118894,I118903,I118873,I119557,I119574,I152160,I119591,I152148,I152154,I119608,I152163,I119531,I119639,I119656,I152151,I119546,I119528,I119701,I119718,I119735,I152172,I119752,I152145,I119769,I152166,I119786,I152157,I119803,I119820,I119837,I119543,I119868,I119885,I119902,I119525,I119933,I119522,I119964,I152142,I119981,I119998,I120015,I119537,I120046,I119534,I120077,I152169,I120094,I120111,I119540,I119549,I119519,I120203,I120220,I358353,I120237,I358365,I358347,I120254,I358362,I120177,I120285,I120302,I358350,I120192,I120174,I120347,I120364,I120381,I358359,I120398,I358338,I120415,I358341,I120432,I358344,I120449,I120466,I120483,I120189,I120514,I120531,I120548,I120171,I120579,I120168,I120610,I358335,I120627,I120644,I120661,I120183,I120692,I120180,I120723,I358356,I120740,I120757,I120186,I120195,I120165,I120849,I120866,I607774,I120883,I607759,I607786,I120900,I607762,I120823,I120931,I120948,I607777,I120838,I120820,I120993,I121010,I121027,I607789,I121044,I607771,I121061,I607780,I121078,I607765,I121095,I121112,I121129,I120835,I121160,I121177,I121194,I120817,I121225,I120814,I121256,I607768,I121273,I121290,I121307,I120829,I121338,I120826,I121369,I607783,I121386,I121403,I120832,I120841,I120811,I121495,I121512,I339619,I121529,I339631,I339613,I121546,I339628,I121469,I121577,I121594,I339616,I121484,I121466,I121639,I121656,I121673,I339625,I121690,I339604,I121707,I339607,I121724,I339610,I121741,I121758,I121775,I121481,I121806,I121823,I121840,I121463,I121871,I121460,I121902,I339601,I121919,I121936,I121953,I121475,I121984,I121472,I122015,I339622,I122032,I122049,I121478,I121487,I121457,I122141,I122158,I122175,I122192,I122115,I122223,I122240,I122130,I122112,I122285,I122302,I122319,I122336,I122353,I122370,I122387,I122404,I122421,I122127,I122452,I122469,I122486,I122109,I122517,I122106,I122548,I122565,I122582,I122599,I122121,I122630,I122118,I122661,I122678,I122695,I122124,I122133,I122103,I122787,I122804,I432130,I122821,I432118,I432124,I122838,I432115,I122761,I122869,I122886,I432121,I122776,I122758,I122931,I122948,I122965,I432133,I122982,I432145,I122999,I432127,I123016,I432142,I123033,I123050,I123067,I122773,I123098,I123115,I123132,I122755,I123163,I122752,I123194,I432136,I123211,I123228,I123245,I122767,I123276,I122764,I123307,I432139,I123324,I123341,I122770,I122779,I122749,I123433,I123450,I290064,I123467,I290061,I290049,I123484,I290052,I123407,I123515,I123532,I290058,I123422,I123404,I123577,I123594,I123611,I290070,I123628,I290046,I123645,I290067,I123662,I290055,I123679,I123696,I123713,I123419,I123744,I123761,I123778,I123401,I123809,I123398,I123840,I290076,I123857,I123874,I123891,I123413,I123922,I123410,I123953,I290073,I123970,I123987,I123416,I123425,I123395,I124079,I124096,I162105,I124113,I162093,I162099,I124130,I162108,I124053,I124161,I124178,I162096,I124068,I124050,I124223,I124240,I124257,I162117,I124274,I162090,I124291,I162111,I124308,I162102,I124325,I124342,I124359,I124065,I124390,I124407,I124424,I124047,I124455,I124044,I124486,I162087,I124503,I124520,I124537,I124059,I124568,I124056,I124599,I162114,I124616,I124633,I124062,I124071,I124041,I124725,I124742,I313932,I124759,I313929,I313917,I124776,I313920,I124699,I124807,I124824,I313926,I124714,I124696,I124869,I124886,I124903,I313938,I124920,I313914,I124937,I313935,I124954,I313923,I124971,I124988,I125005,I124711,I125036,I125053,I125070,I124693,I125101,I124690,I125132,I313944,I125149,I125166,I125183,I124705,I125214,I124702,I125245,I313941,I125262,I125279,I124708,I124717,I124687,I125371,I125388,I493169,I125405,I493151,I493160,I125422,I493172,I125345,I125453,I125470,I493157,I125360,I125342,I125515,I125532,I125549,I493148,I125566,I493166,I125583,I493154,I125600,I493175,I125617,I125634,I125651,I125357,I125682,I125699,I125716,I125339,I125747,I125336,I125778,I493163,I125795,I125812,I125829,I125351,I125860,I125348,I125891,I493145,I125908,I125925,I125354,I125363,I125333,I126017,I126034,I417479,I126051,I417461,I417476,I126068,I417485,I125991,I126099,I126116,I417488,I126006,I125988,I126161,I126178,I126195,I417491,I126212,I417467,I126229,I417470,I126246,I417464,I126263,I126280,I126297,I126003,I126328,I126345,I126362,I125985,I126393,I125982,I126424,I417473,I126441,I126458,I126475,I125997,I126506,I125994,I126537,I417482,I126554,I126571,I126000,I126009,I125979,I126663,I126680,I334451,I126697,I334463,I334445,I126714,I334460,I126637,I126745,I126762,I334448,I126652,I126634,I126807,I126824,I126841,I334457,I126858,I334436,I126875,I334439,I126892,I334442,I126909,I126926,I126943,I126649,I126974,I126991,I127008,I126631,I127039,I126628,I127070,I334433,I127087,I127104,I127121,I126643,I127152,I126640,I127183,I334454,I127200,I127217,I126646,I126655,I126625,I127309,I127326,I127343,I127360,I127283,I127391,I127408,I127298,I127280,I127453,I127470,I127487,I127504,I127521,I127538,I127555,I127572,I127589,I127295,I127620,I127637,I127654,I127277,I127685,I127274,I127716,I127733,I127750,I127767,I127289,I127798,I127286,I127829,I127846,I127863,I127292,I127301,I127271,I127955,I127972,I662108,I127989,I662123,I662138,I128006,I662126,I127929,I128037,I128054,I662129,I127944,I127926,I128099,I128116,I128133,I662135,I128150,I662132,I128167,I662111,I128184,I662120,I128201,I128218,I128235,I127941,I128266,I128283,I128300,I127923,I128331,I127920,I128362,I662117,I128379,I128396,I128413,I127935,I128444,I127932,I128475,I662114,I128492,I128509,I127938,I127947,I127917,I128601,I128618,I191277,I128635,I191265,I191271,I128652,I191280,I128575,I128683,I128700,I191268,I128590,I128572,I128745,I128762,I128779,I191289,I128796,I191262,I128813,I191283,I128830,I191274,I128847,I128864,I128881,I128587,I128912,I128929,I128946,I128569,I128977,I128566,I129008,I191259,I129025,I129042,I129059,I128581,I129090,I128578,I129121,I191286,I129138,I129155,I128584,I128593,I128563,I129247,I129264,I641980,I129281,I641995,I642010,I129298,I641998,I129221,I129329,I129346,I642001,I129236,I129218,I129391,I129408,I129425,I642007,I129442,I642004,I129459,I641983,I129476,I641992,I129493,I129510,I129527,I129233,I129558,I129575,I129592,I129215,I129623,I129212,I129654,I641989,I129671,I129688,I129705,I129227,I129736,I129224,I129767,I641986,I129784,I129801,I129230,I129239,I129209,I129893,I129910,I170724,I129927,I170712,I170718,I129944,I170727,I129867,I129975,I129992,I170715,I129882,I129864,I130037,I130054,I130071,I170736,I130088,I170709,I130105,I170730,I130122,I170721,I130139,I130156,I130173,I129879,I130204,I130221,I130238,I129861,I130269,I129858,I130300,I170706,I130317,I130334,I130351,I129873,I130382,I129870,I130413,I170733,I130430,I130447,I129876,I129885,I129855,I130539,I130556,I427883,I130573,I427865,I427880,I130590,I427889,I130513,I130621,I130638,I427892,I130528,I130510,I130683,I130700,I130717,I427895,I130734,I427871,I130751,I427874,I130768,I427868,I130785,I130802,I130819,I130525,I130850,I130867,I130884,I130507,I130915,I130504,I130946,I427877,I130963,I130980,I130997,I130519,I131028,I130516,I131059,I427886,I131076,I131093,I130522,I130531,I130501,I131185,I131202,I633174,I131219,I633189,I633204,I131236,I633192,I131267,I131284,I633195,I131329,I131346,I131363,I633201,I131380,I633198,I131397,I633177,I131414,I633186,I131431,I131448,I131465,I131496,I131513,I131530,I131561,I131592,I633183,I131609,I131626,I131643,I131674,I131705,I633180,I131722,I131739,I131831,I131848,I616191,I131865,I616206,I616221,I131882,I616209,I131805,I131913,I131930,I616212,I131820,I131802,I131975,I131992,I132009,I616218,I132026,I616215,I132043,I616194,I132060,I616203,I132077,I132094,I132111,I131817,I132142,I132159,I132176,I131799,I132207,I131796,I132238,I616200,I132255,I132272,I132289,I131811,I132320,I131808,I132351,I616197,I132368,I132385,I131814,I131823,I131793,I132477,I132494,I651415,I132511,I651430,I651445,I132528,I651433,I132451,I132559,I132576,I651436,I132466,I132448,I132621,I132638,I132655,I651442,I132672,I651439,I132689,I651418,I132706,I651427,I132723,I132740,I132757,I132463,I132788,I132805,I132822,I132445,I132853,I132442,I132884,I651424,I132901,I132918,I132935,I132457,I132966,I132454,I132997,I651421,I133014,I133031,I132460,I132469,I132439,I133123,I133140,I364167,I133157,I364179,I364161,I133174,I364176,I133097,I133205,I133222,I364164,I133112,I133094,I133267,I133284,I133301,I364173,I133318,I364152,I133335,I364155,I133352,I364158,I133369,I133386,I133403,I133109,I133434,I133451,I133468,I133091,I133499,I133088,I133530,I364149,I133547,I133564,I133581,I133103,I133612,I133100,I133643,I364170,I133660,I133677,I133106,I133115,I133085,I133769,I133786,I133803,I133820,I133743,I133851,I133868,I133758,I133740,I133913,I133930,I133947,I133964,I133981,I133998,I134015,I134032,I134049,I133755,I134080,I134097,I134114,I133737,I134145,I133734,I134176,I134193,I134210,I134227,I133749,I134258,I133746,I134289,I134306,I134323,I133752,I133761,I133731,I134415,I134432,I469700,I134449,I469688,I469694,I134466,I469685,I134389,I134497,I134514,I469691,I134404,I134386,I134559,I134576,I134593,I469703,I134610,I469715,I134627,I469697,I134644,I469712,I134661,I134678,I134695,I134401,I134726,I134743,I134760,I134383,I134791,I134380,I134822,I469706,I134839,I134856,I134873,I134395,I134904,I134392,I134935,I469709,I134952,I134969,I134398,I134407,I134377,I135061,I135078,I347371,I135095,I347383,I347365,I135112,I347380,I135035,I135143,I135160,I347368,I135050,I135032,I135205,I135222,I135239,I347377,I135256,I347356,I135273,I347359,I135290,I347362,I135307,I135324,I135341,I135047,I135372,I135389,I135406,I135029,I135437,I135026,I135468,I347353,I135485,I135502,I135519,I135041,I135550,I135038,I135581,I347374,I135598,I135615,I135044,I135053,I135023,I135707,I135724,I199878,I135741,I199908,I199887,I135758,I199899,I135681,I135789,I135806,I199881,I135696,I135678,I135851,I135868,I135885,I199884,I135902,I199902,I135919,I199893,I135936,I199890,I135953,I135970,I135987,I135693,I136018,I136035,I136052,I135675,I136083,I135672,I136114,I199896,I136131,I136148,I136165,I135687,I136196,I135684,I136227,I199905,I136244,I136261,I135690,I135699,I135669,I136353,I136370,I566136,I136387,I566112,I566118,I136404,I566121,I136327,I136435,I136452,I566130,I136342,I136324,I136497,I136514,I136531,I566109,I136548,I566124,I136565,I566115,I136582,I566127,I136599,I136616,I136633,I136339,I136664,I136681,I136698,I136321,I136729,I136318,I136760,I566139,I136777,I136794,I136811,I136333,I136842,I136330,I136873,I566133,I136890,I136907,I136336,I136345,I136315,I136999,I137016,I516751,I137033,I516727,I516733,I137050,I516736,I136973,I137081,I137098,I516745,I136988,I136970,I137143,I137160,I137177,I516724,I137194,I516739,I137211,I516730,I137228,I516742,I137245,I137262,I137279,I136985,I137310,I137327,I137344,I136967,I137375,I136964,I137406,I516754,I137423,I137440,I137457,I136979,I137488,I136976,I137519,I516748,I137536,I137553,I136982,I136991,I136961,I137645,I137662,I671543,I137679,I671558,I671573,I137696,I671561,I137619,I137727,I137744,I671564,I137634,I137616,I137789,I137806,I137823,I671570,I137840,I671567,I137857,I671546,I137874,I671555,I137891,I137908,I137925,I137631,I137956,I137973,I137990,I137613,I138021,I137610,I138052,I671552,I138069,I138086,I138103,I137625,I138134,I137622,I138165,I671549,I138182,I138199,I137628,I137637,I137607,I138291,I138308,I300672,I138325,I300669,I300657,I138342,I300660,I138265,I138373,I138390,I300666,I138280,I138262,I138435,I138452,I138469,I300678,I138486,I300654,I138503,I300675,I138520,I300663,I138537,I138554,I138571,I138277,I138602,I138619,I138636,I138259,I138667,I138256,I138698,I300684,I138715,I138732,I138749,I138271,I138780,I138268,I138811,I300681,I138828,I138845,I138274,I138283,I138253,I138937,I138954,I138971,I138988,I138911,I139019,I139036,I138926,I138908,I139081,I139098,I139115,I139132,I139149,I139166,I139183,I139200,I139217,I138923,I139248,I139265,I139282,I138905,I139313,I138902,I139344,I139361,I139378,I139395,I138917,I139426,I138914,I139457,I139474,I139491,I138920,I138929,I138899,I139583,I139600,I528044,I139617,I528056,I528059,I139634,I528047,I139665,I139682,I528032,I139699,I139716,I139733,I528035,I139750,I528038,I139767,I528041,I139784,I528050,I139801,I139818,I139863,I139894,I139925,I139942,I139959,I139976,I528053,I139993,I140010,I140041,I140086,I528029,I140103,I140134,I140151,I140168,I140246,I140263,I415025,I140280,I415043,I415031,I140297,I415037,I140217,I140328,I140345,I415040,I140362,I140379,I140396,I415019,I140413,I415013,I140430,I415022,I140447,I415034,I140464,I140481,I140232,I140229,I140526,I140214,I140557,I140211,I140588,I140605,I140622,I140639,I415028,I140656,I140673,I140238,I140704,I140226,I140220,I140749,I415016,I140766,I140235,I140797,I140814,I140831,I140223,I140208,I140909,I140926,I494987,I140943,I494993,I494984,I140960,I495002,I140880,I140991,I141008,I494981,I141025,I141042,I141059,I495011,I141076,I494990,I141093,I494999,I141110,I495005,I141127,I141144,I140895,I140892,I141189,I140877,I141220,I140874,I141251,I141268,I141285,I141302,I494996,I141319,I141336,I140901,I141367,I140889,I140883,I141412,I495008,I141429,I140898,I141460,I141477,I141494,I140886,I140871,I141572,I141589,I604790,I141606,I604805,I604787,I141623,I604799,I141543,I141654,I141671,I604796,I141688,I141705,I141722,I604814,I141739,I604784,I141756,I604793,I141773,I604811,I141790,I141807,I141558,I141555,I141852,I141540,I141883,I141537,I141914,I141931,I141948,I141965,I604802,I141982,I141999,I141564,I142030,I141552,I141546,I142075,I604808,I142092,I141561,I142123,I142140,I142157,I141549,I141534,I142235,I142252,I503107,I142269,I503119,I503122,I142286,I503128,I142317,I142334,I503131,I142351,I142368,I142385,I503110,I142402,I503125,I142419,I503134,I142436,I503137,I142453,I142470,I142515,I142546,I142577,I142594,I142611,I142628,I503113,I142645,I142662,I142693,I142738,I503116,I142755,I142786,I142803,I142820,I142898,I142915,I506624,I142932,I506636,I506639,I142949,I506627,I142869,I142980,I142997,I506612,I143014,I143031,I143048,I506615,I143065,I506618,I143082,I506621,I143099,I506630,I143116,I143133,I142884,I142881,I143178,I142866,I143209,I142863,I143240,I143257,I143274,I143291,I506633,I143308,I143325,I142890,I143356,I142878,I142872,I143401,I506609,I143418,I142887,I143449,I143466,I143483,I142875,I142860,I143561,I143578,I143595,I143612,I143532,I143643,I143660,I143677,I143694,I143711,I143728,I143745,I143762,I143779,I143796,I143547,I143544,I143841,I143529,I143872,I143526,I143903,I143920,I143937,I143954,I143971,I143988,I143553,I144019,I143541,I143535,I144064,I144081,I143550,I144112,I144129,I144146,I143538,I143523,I144224,I144241,I221917,I144258,I221899,I221893,I144275,I221896,I144195,I144306,I144323,I221905,I144340,I144357,I144374,I221914,I144391,I221902,I144408,I221908,I144425,I221923,I144442,I144459,I144210,I144207,I144504,I144192,I144535,I144189,I144566,I144583,I144600,I144617,I221911,I144634,I144651,I144216,I144682,I144204,I144198,I144727,I221920,I144744,I144213,I144775,I144792,I144809,I144201,I144186,I144887,I144904,I338973,I144921,I338982,I338955,I144938,I338967,I144969,I144986,I338979,I145003,I145020,I145037,I338958,I145054,I338964,I145071,I338976,I145088,I338961,I145105,I145122,I145167,I145198,I145229,I145246,I145263,I145280,I338985,I145297,I145314,I145345,I145390,I338970,I145407,I145438,I145455,I145472,I145550,I145567,I145584,I145601,I145521,I145632,I145649,I145666,I145683,I145700,I145717,I145734,I145751,I145768,I145785,I145536,I145533,I145830,I145518,I145861,I145515,I145892,I145909,I145926,I145943,I145960,I145977,I145542,I146008,I145530,I145524,I146053,I146070,I145539,I146101,I146118,I146135,I145527,I145512,I146213,I146230,I146247,I146264,I146184,I146295,I146312,I146329,I146346,I146363,I146380,I146397,I146414,I146431,I146448,I146199,I146196,I146493,I146181,I146524,I146178,I146555,I146572,I146589,I146606,I146623,I146640,I146205,I146671,I146193,I146187,I146716,I146733,I146202,I146764,I146781,I146798,I146190,I146175,I146876,I146893,I366105,I146910,I366114,I366087,I146927,I366099,I146958,I146975,I366111,I146992,I147009,I147026,I366090,I147043,I366096,I147060,I366108,I147077,I366093,I147094,I147111,I147156,I147187,I147218,I147235,I147252,I147269,I366117,I147286,I147303,I147334,I147379,I366102,I147396,I147427,I147444,I147461,I147539,I147556,I520904,I147573,I520916,I520919,I147590,I520907,I147510,I147621,I147638,I520892,I147655,I147672,I147689,I520895,I147706,I520898,I147723,I520901,I147740,I520910,I147757,I147774,I147525,I147522,I147819,I147507,I147850,I147504,I147881,I147898,I147915,I147932,I520913,I147949,I147966,I147531,I147997,I147519,I147513,I148042,I520889,I148059,I147528,I148090,I148107,I148124,I147516,I147501,I148202,I148219,I513764,I148236,I513776,I513779,I148253,I513767,I148173,I148284,I148301,I513752,I148318,I148335,I148352,I513755,I148369,I513758,I148386,I513761,I148403,I513770,I148420,I148437,I148188,I148185,I148482,I148170,I148513,I148167,I148544,I148561,I148578,I148595,I513773,I148612,I148629,I148194,I148660,I148182,I148176,I148705,I513749,I148722,I148191,I148753,I148770,I148787,I148179,I148164,I148865,I148882,I386777,I148899,I386786,I386759,I148916,I386771,I148947,I148964,I386783,I148981,I148998,I149015,I386762,I149032,I386768,I149049,I386780,I149066,I386765,I149083,I149100,I149145,I149176,I149207,I149224,I149241,I149258,I386789,I149275,I149292,I149323,I149368,I386774,I149385,I149416,I149433,I149450,I149528,I149545,I327174,I149562,I327183,I327195,I149579,I327186,I149499,I149610,I149627,I327198,I149644,I149661,I149678,I327204,I149695,I327180,I149712,I327189,I149729,I327177,I149746,I149763,I149514,I149511,I149808,I149496,I149839,I149493,I149870,I149887,I149904,I149921,I327201,I149938,I149955,I149520,I149986,I149508,I149502,I150031,I327192,I150048,I149517,I150079,I150096,I150113,I149505,I149490,I150191,I150208,I475465,I150225,I475471,I475468,I150242,I475486,I150162,I150273,I150290,I475495,I150307,I150324,I150341,I475489,I150358,I475480,I150375,I475483,I150392,I475474,I150409,I150426,I150177,I150174,I150471,I150159,I150502,I150156,I150533,I150550,I150567,I150584,I475492,I150601,I150618,I150183,I150649,I150171,I150165,I150694,I475477,I150711,I150180,I150742,I150759,I150776,I150168,I150153,I150854,I150871,I716974,I150888,I716953,I716965,I150905,I716959,I150825,I150936,I150953,I716980,I150970,I150987,I151004,I716956,I151021,I716968,I151038,I716971,I151055,I716977,I151072,I151089,I150840,I150837,I151134,I150822,I151165,I150819,I151196,I151213,I151230,I151247,I716950,I151264,I151281,I150846,I151312,I150834,I150828,I151357,I716962,I151374,I150843,I151405,I151422,I151439,I150831,I150816,I151517,I151534,I529234,I151551,I529246,I529249,I151568,I529237,I151599,I151616,I529222,I151633,I151650,I151667,I529225,I151684,I529228,I151701,I529231,I151718,I529240,I151735,I151752,I151797,I151828,I151859,I151876,I151893,I151910,I529243,I151927,I151944,I151975,I152020,I529219,I152037,I152068,I152085,I152102,I152180,I152197,I252918,I152214,I252927,I252939,I152231,I252930,I152262,I152279,I252942,I152296,I152313,I152330,I252948,I152347,I252924,I152364,I252933,I152381,I252921,I152398,I152415,I152460,I152491,I152522,I152539,I152556,I152573,I252945,I152590,I152607,I152638,I152683,I252936,I152700,I152731,I152748,I152765,I152843,I152860,I251592,I152877,I251601,I251613,I152894,I251604,I152814,I152925,I152942,I251616,I152959,I152976,I152993,I251622,I153010,I251598,I153027,I251607,I153044,I251595,I153061,I153078,I152829,I152826,I153123,I152811,I153154,I152808,I153185,I153202,I153219,I153236,I251619,I153253,I153270,I152835,I153301,I152823,I152817,I153346,I251610,I153363,I152832,I153394,I153411,I153428,I152820,I152805,I153506,I153523,I680990,I153540,I680996,I681008,I153557,I680999,I153477,I153588,I153605,I680978,I153622,I153639,I153656,I680993,I153673,I680981,I153690,I681002,I153707,I680984,I153724,I153741,I153492,I153489,I153786,I153474,I153817,I153471,I153848,I153865,I153882,I153899,I681005,I153916,I153933,I153498,I153964,I153486,I153480,I154009,I680987,I154026,I153495,I154057,I154074,I154091,I153483,I153468,I154169,I154186,I713506,I154203,I713485,I713497,I154220,I713491,I154140,I154251,I154268,I713512,I154285,I154302,I154319,I713488,I154336,I713500,I154353,I713503,I154370,I713509,I154387,I154404,I154155,I154152,I154449,I154137,I154480,I154134,I154511,I154528,I154545,I154562,I713482,I154579,I154596,I154161,I154627,I154149,I154143,I154672,I713494,I154689,I154158,I154720,I154737,I154754,I154146,I154131,I154832,I154849,I588725,I154866,I588740,I588722,I154883,I588734,I154803,I154914,I154931,I588731,I154948,I154965,I154982,I588749,I154999,I588719,I155016,I588728,I155033,I588746,I155050,I155067,I154818,I154815,I155112,I154800,I155143,I154797,I155174,I155191,I155208,I155225,I588737,I155242,I155259,I154824,I155290,I154812,I154806,I155335,I588743,I155352,I154821,I155383,I155400,I155417,I154809,I154794,I155495,I155512,I155529,I155546,I155466,I155577,I155594,I155611,I155628,I155645,I155662,I155679,I155696,I155713,I155730,I155481,I155478,I155775,I155463,I155806,I155460,I155837,I155854,I155871,I155888,I155905,I155922,I155487,I155953,I155475,I155469,I155998,I156015,I155484,I156046,I156063,I156080,I155472,I155457,I156158,I156175,I236780,I156192,I236774,I236792,I156209,I236768,I156129,I156240,I156257,I236783,I156274,I156291,I156308,I236798,I156325,I236789,I156342,I236777,I156359,I236795,I156376,I156393,I156144,I156141,I156438,I156126,I156469,I156123,I156500,I156517,I156534,I156551,I236786,I156568,I156585,I156150,I156616,I156138,I156132,I156661,I236771,I156678,I156147,I156709,I156726,I156743,I156135,I156120,I156821,I156838,I683506,I156855,I683512,I683524,I156872,I683515,I156903,I156920,I683494,I156937,I156954,I156971,I683509,I156988,I683497,I157005,I683518,I157022,I683500,I157039,I157056,I157101,I157132,I157163,I157180,I157197,I157214,I683521,I157231,I157248,I157279,I157324,I683503,I157341,I157372,I157389,I157406,I157484,I157501,I657088,I157518,I657094,I657106,I157535,I657097,I157455,I157566,I157583,I657076,I157600,I157617,I157634,I657091,I157651,I657079,I157668,I657100,I157685,I657082,I157702,I157719,I157470,I157467,I157764,I157452,I157795,I157449,I157826,I157843,I157860,I157877,I657103,I157894,I157911,I157476,I157942,I157464,I157458,I157987,I657085,I158004,I157473,I158035,I158052,I158069,I157461,I157446,I158147,I158164,I211802,I158181,I211784,I211778,I158198,I211781,I158229,I158246,I211790,I158263,I158280,I158297,I211799,I158314,I211787,I158331,I211793,I158348,I211808,I158365,I158382,I158427,I158458,I158489,I158506,I158523,I158540,I211796,I158557,I158574,I158605,I158650,I211805,I158667,I158698,I158715,I158732,I158810,I158827,I459859,I158844,I459865,I459862,I158861,I459880,I158781,I158892,I158909,I459889,I158926,I158943,I158960,I459883,I158977,I459874,I158994,I459877,I159011,I459868,I159028,I159045,I158796,I158793,I159090,I158778,I159121,I158775,I159152,I159169,I159186,I159203,I459886,I159220,I159237,I158802,I159268,I158790,I158784,I159313,I459871,I159330,I158799,I159361,I159378,I159395,I158787,I158772,I159473,I159490,I516144,I159507,I516156,I516159,I159524,I516147,I159555,I159572,I516132,I159589,I159606,I159623,I516135,I159640,I516138,I159657,I516141,I159674,I516150,I159691,I159708,I159753,I159784,I159815,I159832,I159849,I159866,I516153,I159883,I159900,I159931,I159976,I516129,I159993,I160024,I160041,I160058,I160136,I160153,I660862,I160170,I660868,I660880,I160187,I660871,I160107,I160218,I160235,I660850,I160252,I160269,I160286,I660865,I160303,I660853,I160320,I660874,I160337,I660856,I160354,I160371,I160122,I160119,I160416,I160104,I160447,I160101,I160478,I160495,I160512,I160529,I660877,I160546,I160563,I160128,I160594,I160116,I160110,I160639,I660859,I160656,I160125,I160687,I160704,I160721,I160113,I160098,I160799,I160816,I160833,I160850,I160770,I160881,I160898,I160915,I160932,I160949,I160966,I160983,I161000,I161017,I161034,I160785,I160782,I161079,I160767,I161110,I160764,I161141,I161158,I161175,I161192,I161209,I161226,I160791,I161257,I160779,I160773,I161302,I161319,I160788,I161350,I161367,I161384,I160776,I160761,I161462,I161479,I566719,I161496,I566731,I566734,I161513,I566722,I161433,I161544,I161561,I566707,I161578,I161595,I161612,I566710,I161629,I566713,I161646,I566716,I161663,I566725,I161680,I161697,I161448,I161445,I161742,I161430,I161773,I161427,I161804,I161821,I161838,I161855,I566728,I161872,I161889,I161454,I161920,I161442,I161436,I161965,I566704,I161982,I161451,I162013,I162030,I162047,I161439,I161424,I162125,I162142,I162159,I162176,I162207,I162224,I162241,I162258,I162275,I162292,I162309,I162326,I162343,I162360,I162405,I162436,I162467,I162484,I162501,I162518,I162535,I162552,I162583,I162628,I162645,I162676,I162693,I162710,I162788,I162805,I640105,I162822,I640111,I640123,I162839,I640114,I162759,I162870,I162887,I640093,I162904,I162921,I162938,I640108,I162955,I640096,I162972,I640117,I162989,I640099,I163006,I163023,I162774,I162771,I163068,I162756,I163099,I162753,I163130,I163147,I163164,I163181,I640120,I163198,I163215,I162780,I163246,I162768,I162762,I163291,I640102,I163308,I162777,I163339,I163356,I163373,I162765,I162750,I163451,I163468,I367397,I163485,I367406,I367379,I163502,I367391,I163422,I163533,I163550,I367403,I163567,I163584,I163601,I367382,I163618,I367388,I163635,I367400,I163652,I367385,I163669,I163686,I163437,I163434,I163731,I163419,I163762,I163416,I163793,I163810,I163827,I163844,I367409,I163861,I163878,I163443,I163909,I163431,I163425,I163954,I367394,I163971,I163440,I164002,I164019,I164036,I163428,I163413,I164114,I164131,I276123,I164148,I276132,I276144,I164165,I276135,I164085,I164196,I164213,I276147,I164230,I164247,I164264,I276153,I164281,I276129,I164298,I276138,I164315,I276126,I164332,I164349,I164100,I164097,I164394,I164082,I164425,I164079,I164456,I164473,I164490,I164507,I276150,I164524,I164541,I164106,I164572,I164094,I164088,I164617,I276141,I164634,I164103,I164665,I164682,I164699,I164091,I164076,I164777,I164794,I164811,I164828,I164748,I164859,I164876,I164893,I164910,I164927,I164944,I164961,I164978,I164995,I165012,I164763,I164760,I165057,I164745,I165088,I164742,I165119,I165136,I165153,I165170,I165187,I165204,I164769,I165235,I164757,I164751,I165280,I165297,I164766,I165328,I165345,I165362,I164754,I164739,I165440,I165457,I657717,I165474,I657723,I657735,I165491,I657726,I165411,I165522,I165539,I657705,I165556,I165573,I165590,I657720,I165607,I657708,I165624,I657729,I165641,I657711,I165658,I165675,I165426,I165423,I165720,I165408,I165751,I165405,I165782,I165799,I165816,I165833,I657732,I165850,I165867,I165432,I165898,I165420,I165414,I165943,I657714,I165960,I165429,I165991,I166008,I166025,I165417,I165402,I166103,I166120,I384839,I166137,I384848,I384821,I166154,I384833,I166074,I166185,I166202,I384845,I166219,I166236,I166253,I384824,I166270,I384830,I166287,I384842,I166304,I384827,I166321,I166338,I166089,I166086,I166383,I166071,I166414,I166068,I166445,I166462,I166479,I166496,I384851,I166513,I166530,I166095,I166561,I166083,I166077,I166606,I384836,I166623,I166092,I166654,I166671,I166688,I166080,I166065,I166766,I166783,I647653,I166800,I647659,I647671,I166817,I647662,I166737,I166848,I166865,I647641,I166882,I166899,I166916,I647656,I166933,I647644,I166950,I647665,I166967,I647647,I166984,I167001,I166752,I166749,I167046,I166734,I167077,I166731,I167108,I167125,I167142,I167159,I647668,I167176,I167193,I166758,I167224,I166746,I166740,I167269,I647650,I167286,I166755,I167317,I167334,I167351,I166743,I166728,I167429,I167446,I585750,I167463,I585765,I585747,I167480,I585759,I167511,I167528,I585756,I167545,I167562,I167579,I585774,I167596,I585744,I167613,I585753,I167630,I585771,I167647,I167664,I167709,I167740,I167771,I167788,I167805,I167822,I585762,I167839,I167856,I167887,I167932,I585768,I167949,I167980,I167997,I168014,I168092,I168109,I168126,I168143,I168063,I168174,I168191,I168208,I168225,I168242,I168259,I168276,I168293,I168310,I168327,I168078,I168075,I168372,I168060,I168403,I168057,I168434,I168451,I168468,I168485,I168502,I168519,I168084,I168550,I168072,I168066,I168595,I168612,I168081,I168643,I168660,I168677,I168069,I168054,I168755,I168772,I353831,I168789,I353840,I353813,I168806,I353825,I168726,I168837,I168854,I353837,I168871,I168888,I168905,I353816,I168922,I353822,I168939,I353834,I168956,I353819,I168973,I168990,I168741,I168738,I169035,I168723,I169066,I168720,I169097,I169114,I169131,I169148,I353843,I169165,I169182,I168747,I169213,I168735,I168729,I169258,I353828,I169275,I168744,I169306,I169323,I169340,I168732,I168717,I169418,I169435,I169452,I169469,I169389,I169500,I169517,I169534,I169551,I169568,I169585,I169602,I169619,I169636,I169653,I169404,I169401,I169698,I169386,I169729,I169383,I169760,I169777,I169794,I169811,I169828,I169845,I169410,I169876,I169398,I169392,I169921,I169938,I169407,I169969,I169986,I170003,I169395,I169380,I170081,I170098,I659604,I170115,I659610,I659622,I170132,I659613,I170052,I170163,I170180,I659592,I170197,I170214,I170231,I659607,I170248,I659595,I170265,I659616,I170282,I659598,I170299,I170316,I170067,I170064,I170361,I170049,I170392,I170046,I170423,I170440,I170457,I170474,I659619,I170491,I170508,I170073,I170539,I170061,I170055,I170584,I659601,I170601,I170070,I170632,I170649,I170666,I170058,I170043,I170744,I170761,I223702,I170778,I223684,I223678,I170795,I223681,I170826,I170843,I223690,I170860,I170877,I170894,I223699,I170911,I223687,I170928,I223693,I170945,I223708,I170962,I170979,I171024,I171055,I171086,I171103,I171120,I171137,I223696,I171154,I171171,I171202,I171247,I223705,I171264,I171295,I171312,I171329,I171407,I171424,I171441,I171458,I171378,I171489,I171506,I171523,I171540,I171557,I171574,I171591,I171608,I171625,I171642,I171393,I171390,I171687,I171375,I171718,I171372,I171749,I171766,I171783,I171800,I171817,I171834,I171399,I171865,I171387,I171381,I171910,I171927,I171396,I171958,I171975,I171992,I171384,I171369,I172070,I172087,I519119,I172104,I519131,I519134,I172121,I519122,I172041,I172152,I172169,I519107,I172186,I172203,I172220,I519110,I172237,I519113,I172254,I519116,I172271,I519125,I172288,I172305,I172056,I172053,I172350,I172038,I172381,I172035,I172412,I172429,I172446,I172463,I519128,I172480,I172497,I172062,I172528,I172050,I172044,I172573,I519104,I172590,I172059,I172621,I172638,I172655,I172047,I172032,I172733,I172750,I297339,I172767,I297348,I297360,I172784,I297351,I172704,I172815,I172832,I297363,I172849,I172866,I172883,I297369,I172900,I297345,I172917,I297354,I172934,I297342,I172951,I172968,I172719,I172716,I173013,I172701,I173044,I172698,I173075,I173092,I173109,I173126,I297366,I173143,I173160,I172725,I173191,I172713,I172707,I173236,I297357,I173253,I172722,I173284,I173301,I173318,I172710,I172695,I173396,I173413,I560174,I173430,I560186,I560189,I173447,I560177,I173478,I173495,I560162,I173512,I173529,I173546,I560165,I173563,I560168,I173580,I560171,I173597,I560180,I173614,I173631,I173676,I173707,I173738,I173755,I173772,I173789,I560183,I173806,I173823,I173854,I173899,I560159,I173916,I173947,I173964,I173981,I174059,I174076,I537564,I174093,I537576,I537579,I174110,I537567,I174030,I174141,I174158,I537552,I174175,I174192,I174209,I537555,I174226,I537558,I174243,I537561,I174260,I537570,I174277,I174294,I174045,I174042,I174339,I174027,I174370,I174024,I174401,I174418,I174435,I174452,I537573,I174469,I174486,I174051,I174517,I174039,I174033,I174562,I537549,I174579,I174048,I174610,I174627,I174644,I174036,I174021,I174722,I174739,I482401,I174756,I482407,I482404,I174773,I482422,I174693,I174804,I174821,I482431,I174838,I174855,I174872,I482425,I174889,I482416,I174906,I482419,I174923,I482410,I174940,I174957,I174708,I174705,I175002,I174690,I175033,I174687,I175064,I175081,I175098,I175115,I482428,I175132,I175149,I174714,I175180,I174702,I174696,I175225,I482413,I175242,I174711,I175273,I175290,I175307,I174699,I174684,I175385,I175402,I419921,I175419,I419939,I419927,I175436,I419933,I175356,I175467,I175484,I419936,I175501,I175518,I175535,I419915,I175552,I419909,I175569,I419918,I175586,I419930,I175603,I175620,I175371,I175368,I175665,I175353,I175696,I175350,I175727,I175744,I175761,I175778,I419924,I175795,I175812,I175377,I175843,I175365,I175359,I175888,I419912,I175905,I175374,I175936,I175953,I175970,I175362,I175347,I176048,I176065,I623751,I176082,I623757,I623769,I176099,I623760,I176019,I176130,I176147,I623739,I176164,I176181,I176198,I623754,I176215,I623742,I176232,I623763,I176249,I623745,I176266,I176283,I176034,I176031,I176328,I176016,I176359,I176013,I176390,I176407,I176424,I176441,I623766,I176458,I176475,I176040,I176506,I176028,I176022,I176551,I623748,I176568,I176037,I176599,I176616,I176633,I176025,I176010,I176711,I176728,I621235,I176745,I621241,I621253,I176762,I621244,I176682,I176793,I176810,I621223,I176827,I176844,I176861,I621238,I176878,I621226,I176895,I621247,I176912,I621229,I176929,I176946,I176697,I176694,I176991,I176679,I177022,I176676,I177053,I177070,I177087,I177104,I621250,I177121,I177138,I176703,I177169,I176691,I176685,I177214,I621232,I177231,I176700,I177262,I177279,I177296,I176688,I176673,I177374,I177391,I635073,I177408,I635079,I635091,I177425,I635082,I177345,I177456,I177473,I635061,I177490,I177507,I177524,I635076,I177541,I635064,I177558,I635085,I177575,I635067,I177592,I177609,I177360,I177357,I177654,I177342,I177685,I177339,I177716,I177733,I177750,I177767,I635088,I177784,I177801,I177366,I177832,I177354,I177348,I177877,I635070,I177894,I177363,I177925,I177942,I177959,I177351,I177336,I178037,I178054,I460437,I178071,I460443,I460440,I178088,I460458,I178008,I178119,I178136,I460467,I178153,I178170,I178187,I460461,I178204,I460452,I178221,I460455,I178238,I460446,I178255,I178272,I178023,I178020,I178317,I178005,I178348,I178002,I178379,I178396,I178413,I178430,I460464,I178447,I178464,I178029,I178495,I178017,I178011,I178540,I460449,I178557,I178026,I178588,I178605,I178622,I178014,I177999,I178700,I178717,I290709,I178734,I290718,I290730,I178751,I290721,I178671,I178782,I178799,I290733,I178816,I178833,I178850,I290739,I178867,I290715,I178884,I290724,I178901,I290712,I178918,I178935,I178686,I178683,I178980,I178668,I179011,I178665,I179042,I179059,I179076,I179093,I290736,I179110,I179127,I178692,I179158,I178680,I178674,I179203,I290727,I179220,I178689,I179251,I179268,I179285,I178677,I178662,I179363,I179380,I257559,I179397,I257568,I257580,I179414,I257571,I179334,I179445,I179462,I257583,I179479,I179496,I179513,I257589,I179530,I257565,I179547,I257574,I179564,I257562,I179581,I179598,I179349,I179346,I179643,I179331,I179674,I179328,I179705,I179722,I179739,I179756,I257586,I179773,I179790,I179355,I179821,I179343,I179337,I179866,I257577,I179883,I179352,I179914,I179931,I179948,I179340,I179325,I180026,I180043,I557199,I180060,I557211,I557214,I180077,I557202,I179997,I180108,I180125,I557187,I180142,I180159,I180176,I557190,I180193,I557193,I180210,I557196,I180227,I557205,I180244,I180261,I180012,I180009,I180306,I179994,I180337,I179991,I180368,I180385,I180402,I180419,I557208,I180436,I180453,I180018,I180484,I180006,I180000,I180529,I557184,I180546,I180015,I180577,I180594,I180611,I180003,I179988,I180689,I180706,I337035,I180723,I337044,I337017,I180740,I337029,I180660,I180771,I180788,I337041,I180805,I180822,I180839,I337020,I180856,I337026,I180873,I337038,I180890,I337023,I180907,I180924,I180675,I180672,I180969,I180657,I181000,I180654,I181031,I181048,I181065,I181082,I337047,I181099,I181116,I180681,I181147,I180669,I180663,I181192,I337032,I181209,I180678,I181240,I181257,I181274,I180666,I180651,I181352,I181369,I181386,I181403,I181434,I181451,I181468,I181485,I181502,I181519,I181536,I181553,I181570,I181587,I181632,I181663,I181694,I181711,I181728,I181745,I181762,I181779,I181810,I181855,I181872,I181903,I181920,I181937,I182015,I182032,I246951,I182049,I246960,I246972,I182066,I246963,I181986,I182097,I182114,I246975,I182131,I182148,I182165,I246981,I182182,I246957,I182199,I246966,I182216,I246954,I182233,I182250,I182001,I181998,I182295,I181983,I182326,I181980,I182357,I182374,I182391,I182408,I246978,I182425,I182442,I182007,I182473,I181995,I181989,I182518,I246969,I182535,I182004,I182566,I182583,I182600,I181992,I181977,I182678,I182695,I182712,I182729,I182649,I182760,I182777,I182794,I182811,I182828,I182845,I182862,I182879,I182896,I182913,I182664,I182661,I182958,I182646,I182989,I182643,I183020,I183037,I183054,I183071,I183088,I183105,I182670,I183136,I182658,I182652,I183181,I183198,I182667,I183229,I183246,I183263,I182655,I182640,I183341,I183358,I183375,I183392,I183312,I183423,I183440,I183457,I183474,I183491,I183508,I183525,I183542,I183559,I183576,I183327,I183324,I183621,I183309,I183652,I183306,I183683,I183700,I183717,I183734,I183751,I183768,I183333,I183799,I183321,I183315,I183844,I183861,I183330,I183892,I183909,I183926,I183318,I183303,I184004,I184021,I605385,I184038,I605400,I605382,I184055,I605394,I184086,I184103,I605391,I184120,I184137,I184154,I605409,I184171,I605379,I184188,I605388,I184205,I605406,I184222,I184239,I184284,I184315,I184346,I184363,I184380,I184397,I605397,I184414,I184431,I184462,I184507,I605403,I184524,I184555,I184572,I184589,I184667,I184684,I217752,I184701,I217734,I217728,I184718,I217731,I184638,I184749,I184766,I217740,I184783,I184800,I184817,I217749,I184834,I217737,I184851,I217743,I184868,I217758,I184885,I184902,I184653,I184650,I184947,I184635,I184978,I184632,I185009,I185026,I185043,I185060,I217746,I185077,I185094,I184659,I185125,I184647,I184641,I185170,I217755,I185187,I184656,I185218,I185235,I185252,I184644,I184629,I185330,I185347,I539349,I185364,I539361,I539364,I185381,I539352,I185301,I185412,I185429,I539337,I185446,I185463,I185480,I539340,I185497,I539343,I185514,I539346,I185531,I539355,I185548,I185565,I185316,I185313,I185610,I185298,I185641,I185295,I185672,I185689,I185706,I185723,I539358,I185740,I185757,I185322,I185788,I185310,I185304,I185833,I539334,I185850,I185319,I185881,I185898,I185915,I185307,I185292,I185993,I186010,I662749,I186027,I662755,I662767,I186044,I662758,I185964,I186075,I186092,I662737,I186109,I186126,I186143,I662752,I186160,I662740,I186177,I662761,I186194,I662743,I186211,I186228,I185979,I185976,I186273,I185961,I186304,I185958,I186335,I186352,I186369,I186386,I662764,I186403,I186420,I185985,I186451,I185973,I185967,I186496,I662746,I186513,I185982,I186544,I186561,I186578,I185970,I185955,I186656,I186673,I186690,I186707,I186627,I186738,I186755,I186772,I186789,I186806,I186823,I186840,I186857,I186874,I186891,I186642,I186639,I186936,I186624,I186967,I186621,I186998,I187015,I187032,I187049,I187066,I187083,I186648,I187114,I186636,I186630,I187159,I187176,I186645,I187207,I187224,I187241,I186633,I186618,I187319,I187336,I487643,I187353,I487649,I487640,I187370,I487658,I187290,I187401,I187418,I487637,I187435,I187452,I187469,I487667,I187486,I487646,I187503,I487655,I187520,I487661,I187537,I187554,I187305,I187302,I187599,I187287,I187630,I187284,I187661,I187678,I187695,I187712,I487652,I187729,I187746,I187311,I187777,I187299,I187293,I187822,I487664,I187839,I187308,I187870,I187887,I187904,I187296,I187281,I187982,I187999,I452923,I188016,I452929,I452926,I188033,I452944,I187953,I188064,I188081,I452953,I188098,I188115,I188132,I452947,I188149,I452938,I188166,I452941,I188183,I452932,I188200,I188217,I187968,I187965,I188262,I187950,I188293,I187947,I188324,I188341,I188358,I188375,I452950,I188392,I188409,I187974,I188440,I187962,I187956,I188485,I452935,I188502,I187971,I188533,I188550,I188567,I187959,I187944,I188645,I188662,I322533,I188679,I322542,I322554,I188696,I322545,I188616,I188727,I188744,I322557,I188761,I188778,I188795,I322563,I188812,I322539,I188829,I322548,I188846,I322536,I188863,I188880,I188631,I188628,I188925,I188613,I188956,I188610,I188987,I189004,I189021,I189038,I322560,I189055,I189072,I188637,I189103,I188625,I188619,I189148,I322551,I189165,I188634,I189196,I189213,I189230,I188622,I188607,I189308,I189325,I362229,I189342,I362238,I362211,I189359,I362223,I189279,I189390,I189407,I362235,I189424,I189441,I189458,I362214,I189475,I362220,I189492,I362232,I189509,I362217,I189526,I189543,I189294,I189291,I189588,I189276,I189619,I189273,I189650,I189667,I189684,I189701,I362241,I189718,I189735,I189300,I189766,I189288,I189282,I189811,I362226,I189828,I189297,I189859,I189876,I189893,I189285,I189270,I189971,I189988,I476621,I190005,I476627,I476624,I190022,I476642,I189942,I190053,I190070,I476651,I190087,I190104,I190121,I476645,I190138,I476636,I190155,I476639,I190172,I476630,I190189,I190206,I189957,I189954,I190251,I189939,I190282,I189936,I190313,I190330,I190347,I190364,I476648,I190381,I190398,I189963,I190429,I189951,I189945,I190474,I476633,I190491,I189960,I190522,I190539,I190556,I189948,I189933,I190634,I190651,I304632,I190668,I304641,I304653,I190685,I304644,I190716,I190733,I304656,I190750,I190767,I190784,I304662,I190801,I304638,I190818,I304647,I190835,I304635,I190852,I190869,I190914,I190945,I190976,I190993,I191010,I191027,I304659,I191044,I191061,I191092,I191137,I304650,I191154,I191185,I191202,I191219,I191297,I191314,I462171,I191331,I462177,I462174,I191348,I462192,I191379,I191396,I462201,I191413,I191430,I191447,I462195,I191464,I462186,I191481,I462189,I191498,I462180,I191515,I191532,I191577,I191608,I191639,I191656,I191673,I191690,I462198,I191707,I191724,I191755,I191800,I462183,I191817,I191848,I191865,I191882,I191960,I191977,I377087,I191994,I377096,I377069,I192011,I377081,I191931,I192042,I192059,I377093,I192076,I192093,I192110,I377072,I192127,I377078,I192144,I377090,I192161,I377075,I192178,I192195,I191946,I191943,I192240,I191928,I192271,I191925,I192302,I192319,I192336,I192353,I377099,I192370,I192387,I191952,I192418,I191940,I191934,I192463,I377084,I192480,I191949,I192511,I192528,I192545,I191937,I191922,I192623,I192640,I256896,I192657,I256905,I256917,I192674,I256908,I192594,I192705,I192722,I256920,I192739,I192756,I192773,I256926,I192790,I256902,I192807,I256911,I192824,I256899,I192841,I192858,I192609,I192606,I192903,I192591,I192934,I192588,I192965,I192982,I192999,I193016,I256923,I193033,I193050,I192615,I193081,I192603,I192597,I193126,I256914,I193143,I192612,I193174,I193191,I193208,I192600,I192585,I193286,I193303,I572074,I193320,I572086,I572089,I193337,I572077,I193257,I193368,I193385,I572062,I193402,I193419,I193436,I572065,I193453,I572068,I193470,I572071,I193487,I572080,I193504,I193521,I193272,I193269,I193566,I193254,I193597,I193251,I193628,I193645,I193662,I193679,I572083,I193696,I193713,I193278,I193744,I193266,I193260,I193789,I572059,I193806,I193275,I193837,I193854,I193871,I193263,I193248,I193949,I193966,I385485,I193983,I385494,I385467,I194000,I385479,I193920,I194031,I194048,I385491,I194065,I194082,I194099,I385470,I194116,I385476,I194133,I385488,I194150,I385473,I194167,I194184,I193935,I193932,I194229,I193917,I194260,I193914,I194291,I194308,I194325,I194342,I385497,I194359,I194376,I193941,I194407,I193929,I193923,I194452,I385482,I194469,I193938,I194500,I194517,I194534,I193926,I193911,I194612,I194629,I248940,I194646,I248949,I248961,I194663,I248952,I194583,I194694,I194711,I248964,I194728,I194745,I194762,I248970,I194779,I248946,I194796,I248955,I194813,I248943,I194830,I194847,I194598,I194595,I194892,I194580,I194923,I194577,I194954,I194971,I194988,I195005,I248967,I195022,I195039,I194604,I195070,I194592,I194586,I195115,I248958,I195132,I194601,I195163,I195180,I195197,I194589,I194574,I195275,I195292,I448877,I195309,I448883,I448880,I195326,I448898,I195246,I195357,I195374,I448907,I195391,I195408,I195425,I448901,I195442,I448892,I195459,I448895,I195476,I448886,I195493,I195510,I195261,I195258,I195555,I195243,I195586,I195240,I195617,I195634,I195651,I195668,I448904,I195685,I195702,I195267,I195733,I195255,I195249,I195778,I448889,I195795,I195264,I195826,I195843,I195860,I195252,I195237,I195938,I195955,I532804,I195972,I532816,I532819,I195989,I532807,I195909,I196020,I196037,I532792,I196054,I196071,I196088,I532795,I196105,I532798,I196122,I532801,I196139,I532810,I196156,I196173,I195924,I195921,I196218,I195906,I196249,I195903,I196280,I196297,I196314,I196331,I532813,I196348,I196365,I195930,I196396,I195918,I195912,I196441,I532789,I196458,I195927,I196489,I196506,I196523,I195915,I195900,I196601,I196618,I320544,I196635,I320553,I320565,I196652,I320556,I196572,I196683,I196700,I320568,I196717,I196734,I196751,I320574,I196768,I320550,I196785,I320559,I196802,I320547,I196819,I196836,I196587,I196584,I196881,I196569,I196912,I196566,I196943,I196960,I196977,I196994,I320571,I197011,I197028,I196593,I197059,I196581,I196575,I197104,I320562,I197121,I196590,I197152,I197169,I197186,I196578,I196563,I197264,I197281,I576825,I197298,I576840,I576822,I197315,I576834,I197346,I197363,I576831,I197380,I197397,I197414,I576849,I197431,I576819,I197448,I576828,I197465,I576846,I197482,I197499,I197544,I197575,I197606,I197623,I197640,I197657,I576837,I197674,I197691,I197722,I197767,I576843,I197784,I197815,I197832,I197849,I197927,I197944,I197961,I197978,I197898,I198009,I198026,I198043,I198060,I198077,I198094,I198111,I198128,I198145,I198162,I197913,I197910,I198207,I197895,I198238,I197892,I198269,I198286,I198303,I198320,I198337,I198354,I197919,I198385,I197907,I197901,I198430,I198447,I197916,I198478,I198495,I198512,I197904,I197889,I198590,I198607,I716396,I198624,I716375,I716387,I198641,I716381,I198561,I198672,I198689,I716402,I198706,I198723,I198740,I716378,I198757,I716390,I198774,I716393,I198791,I716399,I198808,I198825,I198576,I198573,I198870,I198558,I198901,I198555,I198932,I198949,I198966,I198983,I716372,I199000,I199017,I198582,I199048,I198570,I198564,I199093,I716384,I199110,I198579,I199141,I199158,I199175,I198567,I198552,I199253,I199270,I439051,I199287,I439057,I439054,I199304,I439072,I199335,I199352,I439081,I199369,I199386,I199403,I439075,I199420,I439066,I199437,I439069,I199454,I439060,I199471,I199488,I199533,I199564,I199595,I199612,I199629,I199646,I439078,I199663,I199680,I199711,I199756,I439063,I199773,I199804,I199821,I199838,I199916,I199933,I199950,I199981,I199998,I200015,I200032,I200049,I200066,I200083,I200100,I200117,I200148,I200165,I200196,I200213,I200230,I200275,I200292,I200309,I200326,I200343,I200374,I200405,I200511,I200528,I478963,I478948,I200545,I478960,I200485,I200576,I478942,I478933,I200593,I200610,I200627,I478957,I200644,I200661,I478936,I478954,I200678,I200695,I200712,I200479,I200743,I200760,I200476,I200791,I478945,I200808,I478939,I200825,I200488,I200473,I200870,I478951,I200887,I200904,I200921,I200938,I200494,I200969,I200503,I201000,I200497,I200500,I200491,I200482,I201106,I201123,I344787,I344784,I201140,I344769,I201171,I344778,I344781,I201188,I201205,I201222,I344793,I201239,I201256,I344799,I344775,I201273,I201290,I201307,I201338,I201355,I201386,I344790,I201403,I344796,I201420,I201465,I344772,I201482,I201499,I201516,I201533,I201564,I201595,I201701,I201718,I594086,I594080,I201735,I594074,I201675,I201766,I594077,I594083,I201783,I201800,I201817,I594101,I201834,I201851,I594104,I594095,I201868,I201885,I201902,I201669,I201933,I201950,I201666,I201981,I594092,I201998,I594089,I202015,I201678,I201663,I202060,I594098,I202077,I202094,I202111,I202128,I201684,I202159,I201693,I202190,I201687,I201690,I201681,I201672,I202296,I202313,I427268,I427253,I202330,I427262,I202270,I202361,I427274,I427283,I202378,I202395,I202412,I427271,I202429,I202446,I427280,I427256,I202463,I202480,I202497,I202264,I202528,I202545,I202261,I202576,I427265,I202593,I427259,I202610,I202273,I202258,I202655,I427277,I202672,I202689,I202706,I202723,I202279,I202754,I202288,I202785,I202282,I202285,I202276,I202267,I202891,I202908,I202925,I202865,I202956,I202973,I202990,I203007,I203024,I203041,I203058,I203075,I203092,I202859,I203123,I203140,I202856,I203171,I203188,I203205,I202868,I202853,I203250,I203267,I203284,I203301,I203318,I202874,I203349,I202883,I203380,I202877,I202880,I202871,I202862,I203486,I203503,I203520,I203551,I203568,I203585,I203602,I203619,I203636,I203653,I203670,I203687,I203718,I203735,I203766,I203783,I203800,I203845,I203862,I203879,I203896,I203913,I203944,I203975,I204081,I204098,I204115,I204055,I204146,I204163,I204180,I204197,I204214,I204231,I204248,I204265,I204282,I204049,I204313,I204330,I204046,I204361,I204378,I204395,I204058,I204043,I204440,I204457,I204474,I204491,I204508,I204064,I204539,I204073,I204570,I204067,I204070,I204061,I204052,I204676,I204693,I204710,I204741,I204758,I204775,I204792,I204809,I204826,I204843,I204860,I204877,I204908,I204925,I204956,I204973,I204990,I205035,I205052,I205069,I205086,I205103,I205134,I205165,I205271,I205288,I266841,I266856,I205305,I266844,I205336,I266847,I266862,I205353,I205370,I205387,I266850,I205404,I205421,I266853,I266871,I205438,I205455,I205472,I205503,I205520,I205551,I266868,I205568,I266859,I205585,I205630,I266865,I205647,I205664,I205681,I205698,I205729,I205760,I205866,I205883,I325185,I325200,I205900,I325188,I205840,I205931,I325191,I325206,I205948,I205965,I205982,I325194,I205999,I206016,I325197,I325215,I206033,I206050,I206067,I205834,I206098,I206115,I205831,I206146,I325212,I206163,I325203,I206180,I205843,I205828,I206225,I325209,I206242,I206259,I206276,I206293,I205849,I206324,I205858,I206355,I205852,I205855,I205846,I205837,I206461,I206478,I230833,I230824,I206495,I230845,I206435,I206526,I230848,I230827,I206543,I206560,I206577,I230836,I206594,I206611,I230821,I230839,I206628,I206645,I206662,I206429,I206693,I206710,I206426,I206741,I230842,I206758,I230818,I206775,I206438,I206423,I206820,I230830,I206837,I206854,I206871,I206888,I206444,I206919,I206453,I206950,I206447,I206450,I206441,I206432,I207056,I207073,I345433,I345430,I207090,I345415,I207030,I207121,I345424,I345427,I207138,I207155,I207172,I345439,I207189,I207206,I345445,I345421,I207223,I207240,I207257,I207024,I207288,I207305,I207021,I207336,I345436,I207353,I345442,I207370,I207033,I207018,I207415,I345418,I207432,I207449,I207466,I207483,I207039,I207514,I207048,I207545,I207042,I207045,I207036,I207027,I207651,I207668,I546489,I546474,I207685,I546495,I207625,I207716,I546501,I546483,I207733,I207750,I207767,I546480,I207784,I207801,I546477,I546486,I207818,I207835,I207852,I207619,I207883,I207900,I207616,I207931,I546504,I207948,I546492,I207965,I207628,I207613,I208010,I546498,I208027,I208044,I208061,I208078,I207634,I208109,I207643,I208140,I207637,I207640,I207631,I207622,I208246,I208263,I594681,I594675,I208280,I594669,I208220,I208311,I594672,I594678,I208328,I208345,I208362,I594696,I208379,I208396,I594699,I594690,I208413,I208430,I208447,I208214,I208478,I208495,I208211,I208526,I594687,I208543,I594684,I208560,I208223,I208208,I208605,I594693,I208622,I208639,I208656,I208673,I208229,I208704,I208238,I208735,I208232,I208235,I208226,I208217,I208841,I208858,I208875,I208815,I208906,I208923,I208940,I208957,I208974,I208991,I209008,I209025,I209042,I208809,I209073,I209090,I208806,I209121,I209138,I209155,I208818,I208803,I209200,I209217,I209234,I209251,I209268,I208824,I209299,I208833,I209330,I208827,I208830,I208821,I208812,I209436,I209453,I209470,I209410,I209501,I209518,I209535,I209552,I209569,I209586,I209603,I209620,I209637,I209404,I209668,I209685,I209401,I209716,I209733,I209750,I209413,I209398,I209795,I209812,I209829,I209846,I209863,I209419,I209894,I209428,I209925,I209422,I209425,I209416,I209407,I210031,I210048,I210065,I210005,I210096,I210113,I210130,I210147,I210164,I210181,I210198,I210215,I210232,I209999,I210263,I210280,I209996,I210311,I210328,I210345,I210008,I209993,I210390,I210407,I210424,I210441,I210458,I210014,I210489,I210023,I210520,I210017,I210020,I210011,I210002,I210626,I210643,I601821,I601815,I210660,I601809,I210600,I210691,I601812,I601818,I210708,I210725,I210742,I601836,I210759,I210776,I601839,I601830,I210793,I210810,I210827,I210594,I210858,I210875,I210591,I210906,I601827,I210923,I601824,I210940,I210603,I210588,I210985,I601833,I211002,I211019,I211036,I211053,I210609,I211084,I210618,I211115,I210612,I210615,I210606,I210597,I211221,I211238,I555414,I555399,I211255,I555420,I211195,I211286,I555426,I555408,I211303,I211320,I211337,I555405,I211354,I211371,I555402,I555411,I211388,I211405,I211422,I211189,I211453,I211470,I211186,I211501,I555429,I211518,I555417,I211535,I211198,I211183,I211580,I555423,I211597,I211614,I211631,I211648,I211204,I211679,I211213,I211710,I211207,I211210,I211201,I211192,I211816,I211833,I425432,I425417,I211850,I425426,I211881,I425438,I425447,I211898,I211915,I211932,I425435,I211949,I211966,I425444,I425420,I211983,I212000,I212017,I212048,I212065,I212096,I425429,I212113,I425423,I212130,I212175,I425441,I212192,I212209,I212226,I212243,I212274,I212305,I212411,I212428,I403573,I403570,I212445,I403555,I212476,I403564,I403567,I212493,I212510,I212527,I403579,I212544,I212561,I403585,I403561,I212578,I212595,I212612,I212643,I212660,I212691,I403576,I212708,I403582,I212725,I212770,I403558,I212787,I212804,I212821,I212838,I212869,I212900,I213006,I213023,I391299,I391296,I213040,I391281,I212980,I213071,I391290,I391293,I213088,I213105,I213122,I391305,I213139,I213156,I391311,I391287,I213173,I213190,I213207,I212974,I213238,I213255,I212971,I213286,I391302,I213303,I391308,I213320,I212983,I212968,I213365,I391284,I213382,I213399,I213416,I213433,I212989,I213464,I212998,I213495,I212992,I212995,I212986,I212977,I213601,I213618,I496749,I496770,I213635,I496761,I213666,I496779,I496773,I213683,I213700,I213717,I496758,I213734,I213751,I496767,I496752,I213768,I213785,I213802,I213833,I213850,I213881,I496764,I213898,I496755,I213915,I213960,I496776,I213977,I213994,I214011,I214028,I214059,I214090,I214196,I214213,I638838,I638835,I214230,I638865,I214170,I214261,I638844,I638850,I214278,I214295,I214312,I638841,I214329,I214346,I638853,I638862,I214363,I214380,I214397,I214164,I214428,I214445,I214161,I214476,I638856,I214493,I638847,I214510,I214173,I214158,I214555,I638859,I214572,I214589,I214606,I214623,I214179,I214654,I214188,I214685,I214182,I214185,I214176,I214167,I214791,I214808,I214825,I214765,I214856,I214873,I214890,I214907,I214924,I214941,I214958,I214975,I214992,I214759,I215023,I215040,I214756,I215071,I215088,I215105,I214768,I214753,I215150,I215167,I215184,I215201,I215218,I214774,I215249,I214783,I215280,I214777,I214780,I214771,I214762,I215386,I215403,I648273,I648270,I215420,I648300,I215360,I215451,I648279,I648285,I215468,I215485,I215502,I648276,I215519,I215536,I648288,I648297,I215553,I215570,I215587,I215354,I215618,I215635,I215351,I215666,I648291,I215683,I648282,I215700,I215363,I215348,I215745,I648294,I215762,I215779,I215796,I215813,I215369,I215844,I215378,I215875,I215372,I215375,I215366,I215357,I215981,I215998,I378379,I378376,I216015,I378361,I215955,I216046,I378370,I378373,I216063,I216080,I216097,I378385,I216114,I216131,I378391,I378367,I216148,I216165,I216182,I215949,I216213,I216230,I215946,I216261,I378382,I216278,I378388,I216295,I215958,I215943,I216340,I378364,I216357,I216374,I216391,I216408,I215964,I216439,I215973,I216470,I215967,I215970,I215961,I215952,I216576,I216593,I216610,I216641,I216658,I216675,I216692,I216709,I216726,I216743,I216760,I216777,I216808,I216825,I216856,I216873,I216890,I216935,I216952,I216969,I216986,I217003,I217034,I217065,I217171,I217188,I459311,I459296,I217205,I459308,I217145,I217236,I459290,I459281,I217253,I217270,I217287,I459305,I217304,I217321,I459284,I459302,I217338,I217355,I217372,I217139,I217403,I217420,I217136,I217451,I459293,I217468,I459287,I217485,I217148,I217133,I217530,I459299,I217547,I217564,I217581,I217598,I217154,I217629,I217163,I217660,I217157,I217160,I217151,I217142,I217766,I217783,I695564,I695582,I217800,I695567,I217831,I695576,I695579,I217848,I217865,I217882,I695585,I217899,I217916,I695591,I695570,I217933,I217950,I217967,I217998,I218015,I218046,I695594,I218063,I695588,I218080,I218125,I695573,I218142,I218159,I218176,I218193,I218224,I218255,I218361,I218378,I218395,I218335,I218426,I218443,I218460,I218477,I218494,I218511,I218528,I218545,I218562,I218329,I218593,I218610,I218326,I218641,I218658,I218675,I218338,I218323,I218720,I218737,I218754,I218771,I218788,I218344,I218819,I218353,I218850,I218347,I218350,I218341,I218332,I218956,I218973,I464513,I464498,I218990,I464510,I219021,I464492,I464483,I219038,I219055,I219072,I464507,I219089,I219106,I464486,I464504,I219123,I219140,I219157,I219188,I219205,I219236,I464495,I219253,I464489,I219270,I219315,I464501,I219332,I219349,I219366,I219383,I219414,I219445,I219551,I219568,I632548,I632545,I219585,I632575,I219525,I219616,I632554,I632560,I219633,I219650,I219667,I632551,I219684,I219701,I632563,I632572,I219718,I219735,I219752,I219519,I219783,I219800,I219516,I219831,I632566,I219848,I632557,I219865,I219528,I219513,I219910,I632569,I219927,I219944,I219961,I219978,I219534,I220009,I219543,I220040,I219537,I219540,I219531,I219522,I220146,I220163,I220180,I220120,I220211,I220228,I220245,I220262,I220279,I220296,I220313,I220330,I220347,I220114,I220378,I220395,I220111,I220426,I220443,I220460,I220123,I220108,I220505,I220522,I220539,I220556,I220573,I220129,I220604,I220138,I220635,I220132,I220135,I220126,I220117,I220741,I220758,I232023,I232014,I220775,I232035,I220715,I220806,I232038,I232017,I220823,I220840,I220857,I232026,I220874,I220891,I232011,I232029,I220908,I220925,I220942,I220709,I220973,I220990,I220706,I221021,I232032,I221038,I232008,I221055,I220718,I220703,I221100,I232020,I221117,I221134,I221151,I221168,I220724,I221199,I220733,I221230,I220727,I220730,I220721,I220712,I221336,I221353,I562554,I562539,I221370,I562560,I221310,I221401,I562566,I562548,I221418,I221435,I221452,I562545,I221469,I221486,I562542,I562551,I221503,I221520,I221537,I221304,I221568,I221585,I221301,I221616,I562569,I221633,I562557,I221650,I221313,I221298,I221695,I562563,I221712,I221729,I221746,I221763,I221319,I221794,I221328,I221825,I221322,I221325,I221316,I221307,I221931,I221948,I221965,I221996,I222013,I222030,I222047,I222064,I222081,I222098,I222115,I222132,I222163,I222180,I222211,I222228,I222245,I222290,I222307,I222324,I222341,I222358,I222389,I222420,I222526,I222543,I294687,I294702,I222560,I294690,I222500,I222591,I294693,I294708,I222608,I222625,I222642,I294696,I222659,I222676,I294699,I294717,I222693,I222710,I222727,I222494,I222758,I222775,I222491,I222806,I294714,I222823,I294705,I222840,I222503,I222488,I222885,I294711,I222902,I222919,I222936,I222953,I222509,I222984,I222518,I223015,I222512,I222515,I222506,I222497,I223121,I223138,I590516,I590510,I223155,I590504,I223095,I223186,I590507,I590513,I223203,I223220,I223237,I590531,I223254,I223271,I590534,I590525,I223288,I223305,I223322,I223089,I223353,I223370,I223086,I223401,I590522,I223418,I590519,I223435,I223098,I223083,I223480,I590528,I223497,I223514,I223531,I223548,I223104,I223579,I223113,I223610,I223107,I223110,I223101,I223092,I223716,I223733,I388715,I388712,I223750,I388697,I223781,I388706,I388709,I223798,I223815,I223832,I388721,I223849,I223866,I388727,I388703,I223883,I223900,I223917,I223948,I223965,I223996,I388718,I224013,I388724,I224030,I224075,I388700,I224092,I224109,I224126,I224143,I224174,I224205,I224311,I224328,I400989,I400986,I224345,I400971,I224285,I224376,I400980,I400983,I224393,I224410,I224427,I400995,I224444,I224461,I401001,I400977,I224478,I224495,I224512,I224279,I224543,I224560,I224276,I224591,I400992,I224608,I400998,I224625,I224288,I224273,I224670,I400974,I224687,I224704,I224721,I224738,I224294,I224769,I224303,I224800,I224297,I224300,I224291,I224282,I224906,I224923,I265515,I265530,I224940,I265518,I224880,I224971,I265521,I265536,I224988,I225005,I225022,I265524,I225039,I225056,I265527,I265545,I225073,I225090,I225107,I224874,I225138,I225155,I224871,I225186,I265542,I225203,I265533,I225220,I224883,I224868,I225265,I265539,I225282,I225299,I225316,I225333,I224889,I225364,I224898,I225395,I224892,I224895,I224886,I224877,I225501,I225518,I288057,I288072,I225535,I288060,I225475,I225566,I288063,I288078,I225583,I225600,I225617,I288066,I225634,I225651,I288069,I288087,I225668,I225685,I225702,I225469,I225733,I225750,I225466,I225781,I288084,I225798,I288075,I225815,I225478,I225463,I225860,I288081,I225877,I225894,I225911,I225928,I225484,I225959,I225493,I225990,I225487,I225490,I225481,I225472,I226096,I226113,I241543,I241534,I226130,I241555,I226070,I226161,I241558,I241537,I226178,I226195,I226212,I241546,I226229,I226246,I241531,I241549,I226263,I226280,I226297,I226064,I226328,I226345,I226061,I226376,I241552,I226393,I241528,I226410,I226073,I226058,I226455,I241540,I226472,I226489,I226506,I226523,I226079,I226554,I226088,I226585,I226082,I226085,I226076,I226067,I226691,I226708,I226725,I226665,I226756,I226773,I226790,I226807,I226824,I226841,I226858,I226875,I226892,I226659,I226923,I226940,I226656,I226971,I226988,I227005,I226668,I226653,I227050,I227067,I227084,I227101,I227118,I226674,I227149,I226683,I227180,I226677,I226680,I226671,I226662,I227286,I227303,I326511,I326526,I227320,I326514,I227351,I326517,I326532,I227368,I227385,I227402,I326520,I227419,I227436,I326523,I326541,I227453,I227470,I227487,I227518,I227535,I227566,I326538,I227583,I326529,I227600,I227645,I326535,I227662,I227679,I227696,I227713,I227744,I227775,I227881,I227898,I227943,I227960,I227977,I227994,I228011,I228028,I228045,I228062,I228079,I228110,I228127,I228144,I228161,I228192,I228209,I228226,I228243,I228260,I228291,I228308,I228367,I228398,I228476,I228493,I228459,I228438,I228538,I228555,I228572,I228589,I228606,I228623,I228640,I228657,I228674,I228465,I228705,I228722,I228739,I228756,I228468,I228787,I228804,I228821,I228838,I228855,I228453,I228886,I228903,I228456,I228450,I228444,I228962,I228462,I228993,I228447,I228441,I229071,I229088,I229054,I229033,I229133,I229150,I229167,I229184,I229201,I229218,I229235,I229252,I229269,I229060,I229300,I229317,I229334,I229351,I229063,I229382,I229399,I229416,I229433,I229450,I229048,I229481,I229498,I229051,I229045,I229039,I229557,I229057,I229588,I229042,I229036,I229666,I229683,I229649,I229628,I229728,I229745,I229762,I229779,I229796,I229813,I229830,I229847,I229864,I229655,I229895,I229912,I229929,I229946,I229658,I229977,I229994,I230011,I230028,I230045,I229643,I230076,I230093,I229646,I229640,I229634,I230152,I229652,I230183,I229637,I229631,I230261,I230278,I645131,I645140,I230323,I645149,I230340,I645143,I645137,I230357,I230374,I230391,I645146,I230408,I230425,I230442,I645134,I645152,I230459,I230490,I230507,I230524,I230541,I230572,I645155,I230589,I645128,I230606,I230623,I230640,I230671,I230688,I230747,I645125,I230778,I230856,I230873,I380948,I380945,I230918,I380954,I230935,I380969,I380960,I230952,I230969,I230986,I380963,I231003,I231020,I231037,I380975,I380972,I231054,I231085,I231102,I231119,I231136,I231167,I380951,I231184,I380966,I231201,I231218,I231235,I231266,I231283,I231342,I380957,I231373,I231451,I231468,I684129,I684138,I231434,I231413,I231513,I684147,I231530,I684141,I684135,I231547,I231564,I231581,I684144,I231598,I231615,I231632,I684132,I684150,I231649,I231440,I231680,I231697,I231714,I231731,I231443,I231762,I684153,I231779,I684126,I231796,I231813,I231830,I231428,I231861,I231878,I231431,I231425,I231419,I231937,I684123,I231437,I231968,I231422,I231416,I232046,I232063,I548265,I548277,I232108,I548289,I232125,I548283,I548268,I232142,I232159,I232176,I548280,I232193,I232210,I232227,I548274,I548271,I232244,I232275,I232292,I232309,I232326,I232357,I548286,I232374,I548259,I232391,I232408,I232425,I232456,I232473,I232532,I548262,I232563,I232641,I232658,I468529,I468559,I232624,I232603,I232703,I468538,I232720,I468544,I468541,I232737,I232754,I232771,I468550,I232788,I232805,I232822,I468535,I468553,I232839,I232630,I232870,I232887,I232904,I232921,I232633,I232952,I468556,I232969,I468547,I232986,I233003,I233020,I232618,I233051,I233068,I232621,I232615,I232609,I233127,I468532,I232627,I233158,I232612,I232606,I233236,I233253,I233219,I233198,I233298,I233315,I233332,I233349,I233366,I233383,I233400,I233417,I233434,I233225,I233465,I233482,I233499,I233516,I233228,I233547,I233564,I233581,I233598,I233615,I233213,I233646,I233663,I233216,I233210,I233204,I233722,I233222,I233753,I233207,I233201,I233831,I233848,I233814,I233793,I233893,I233910,I233927,I233944,I233961,I233978,I233995,I234012,I234029,I233820,I234060,I234077,I234094,I234111,I233823,I234142,I234159,I234176,I234193,I234210,I233808,I234241,I234258,I233811,I233805,I233799,I234317,I233817,I234348,I233802,I233796,I234426,I234443,I643873,I643882,I234409,I234388,I234488,I643891,I234505,I643885,I643879,I234522,I234539,I234556,I643888,I234573,I234590,I234607,I643876,I643894,I234624,I234415,I234655,I234672,I234689,I234706,I234418,I234737,I643897,I234754,I643870,I234771,I234788,I234805,I234403,I234836,I234853,I234406,I234400,I234394,I234912,I643867,I234412,I234943,I234397,I234391,I235021,I235038,I384178,I384175,I235004,I234983,I235083,I384184,I235100,I384199,I384190,I235117,I235134,I235151,I384193,I235168,I235185,I235202,I384205,I384202,I235219,I235010,I235250,I235267,I235284,I235301,I235013,I235332,I384181,I235349,I384196,I235366,I235383,I235400,I234998,I235431,I235448,I235001,I234995,I234989,I235507,I384187,I235007,I235538,I234992,I234986,I235616,I235633,I598245,I598239,I235599,I235578,I235678,I598266,I235695,I598269,I598254,I235712,I235729,I235746,I598263,I235763,I235780,I235797,I598248,I598251,I235814,I235605,I235845,I235862,I235879,I235896,I235608,I235927,I598260,I235944,I598242,I235961,I235978,I235995,I235593,I236026,I236043,I235596,I235590,I235584,I236102,I598257,I235602,I236133,I235587,I235581,I236211,I236228,I572660,I572672,I236194,I236173,I236273,I572684,I236290,I572678,I572663,I236307,I236324,I236341,I572675,I236358,I236375,I236392,I572669,I572666,I236409,I236200,I236440,I236457,I236474,I236491,I236203,I236522,I572681,I236539,I572654,I236556,I236573,I236590,I236188,I236621,I236638,I236191,I236185,I236179,I236697,I572657,I236197,I236728,I236182,I236176,I236806,I236823,I259563,I259551,I236868,I259548,I236885,I259578,I259569,I236902,I236919,I236936,I259557,I236953,I236970,I236987,I259560,I259554,I237004,I237035,I237052,I237069,I237086,I237117,I259575,I237134,I259572,I237151,I237168,I237185,I237216,I237233,I237292,I259566,I237323,I237401,I237418,I522085,I522097,I237384,I237363,I237463,I522109,I237480,I522103,I522088,I237497,I237514,I237531,I522100,I237548,I237565,I237582,I522094,I522091,I237599,I237390,I237630,I237647,I237664,I237681,I237393,I237712,I522106,I237729,I522079,I237746,I237763,I237780,I237378,I237811,I237828,I237381,I237375,I237369,I237887,I522082,I237387,I237918,I237372,I237366,I237996,I238013,I509590,I509602,I237979,I237958,I238058,I509614,I238075,I509608,I509593,I238092,I238109,I238126,I509605,I238143,I238160,I238177,I509599,I509596,I238194,I237985,I238225,I238242,I238259,I238276,I237988,I238307,I509611,I238324,I509584,I238341,I238358,I238375,I237973,I238406,I238423,I237976,I237970,I237964,I238482,I509587,I237982,I238513,I237967,I237961,I238591,I238608,I580395,I580389,I238653,I580416,I238670,I580419,I580404,I238687,I238704,I238721,I580413,I238738,I238755,I238772,I580398,I580401,I238789,I238820,I238837,I238854,I238871,I238902,I580410,I238919,I580392,I238936,I238953,I238970,I239001,I239018,I239077,I580407,I239108,I239186,I239203,I239248,I239265,I239282,I239299,I239316,I239333,I239350,I239367,I239384,I239415,I239432,I239449,I239466,I239497,I239514,I239531,I239548,I239565,I239596,I239613,I239672,I239703,I239781,I239798,I239764,I239743,I239843,I239860,I239877,I239894,I239911,I239928,I239945,I239962,I239979,I239770,I240010,I240027,I240044,I240061,I239773,I240092,I240109,I240126,I240143,I240160,I239758,I240191,I240208,I239761,I239755,I239749,I240267,I239767,I240298,I239752,I239746,I240376,I240393,I703099,I703081,I240359,I240338,I240438,I703108,I240455,I703090,I703105,I240472,I240489,I240506,I703087,I240523,I240540,I240557,I703102,I703078,I240574,I240365,I240605,I240622,I240639,I240656,I240368,I240687,I703096,I240704,I703084,I240721,I240738,I240755,I240353,I240786,I240803,I240356,I240350,I240344,I240862,I703093,I240362,I240893,I240347,I240341,I240971,I240988,I240954,I240933,I241033,I241050,I241067,I241084,I241101,I241118,I241135,I241152,I241169,I240960,I241200,I241217,I241234,I241251,I240963,I241282,I241299,I241316,I241333,I241350,I240948,I241381,I241398,I240951,I240945,I240939,I241457,I240957,I241488,I240942,I240936,I241566,I241583,I348002,I347999,I241628,I348008,I241645,I348023,I348014,I241662,I241679,I241696,I348017,I241713,I241730,I241747,I348029,I348026,I241764,I241795,I241812,I241829,I241846,I241877,I348005,I241894,I348020,I241911,I241928,I241945,I241976,I241993,I242052,I348011,I242083,I242161,I242178,I631922,I631931,I242144,I242123,I242223,I631940,I242240,I631934,I631928,I242257,I242274,I242291,I631937,I242308,I242325,I242342,I631925,I631943,I242359,I242150,I242390,I242407,I242424,I242441,I242153,I242472,I631946,I242489,I631919,I242506,I242523,I242540,I242138,I242571,I242588,I242141,I242135,I242129,I242647,I631916,I242147,I242678,I242132,I242126,I242756,I242773,I402266,I402263,I242818,I402272,I242835,I402287,I402278,I242852,I242869,I242886,I402281,I242903,I242920,I242937,I402293,I402290,I242954,I242985,I243002,I243019,I243036,I243067,I402269,I243084,I402284,I243101,I243118,I243135,I243166,I243183,I243242,I402275,I243273,I243351,I243368,I394514,I394511,I243334,I243313,I243413,I394520,I243430,I394535,I394526,I243447,I243464,I243481,I394529,I243498,I243515,I243532,I394541,I394538,I243549,I243340,I243580,I243597,I243614,I243631,I243343,I243662,I394517,I243679,I394532,I243696,I243713,I243730,I243328,I243761,I243778,I243331,I243325,I243319,I243837,I394523,I243337,I243868,I243322,I243316,I243946,I243963,I244008,I244025,I244042,I244059,I244076,I244093,I244110,I244127,I244144,I244175,I244192,I244209,I244226,I244257,I244274,I244291,I244308,I244325,I244356,I244373,I244432,I244463,I244541,I244558,I244603,I244620,I244637,I244654,I244671,I244688,I244705,I244722,I244739,I244770,I244787,I244804,I244821,I244852,I244869,I244886,I244903,I244920,I244951,I244968,I245027,I245058,I245136,I245153,I543505,I543517,I245198,I543529,I245215,I543523,I543508,I245232,I245249,I245266,I543520,I245283,I245300,I245317,I543514,I543511,I245334,I245365,I245382,I245399,I245416,I245447,I543526,I245464,I543499,I245481,I245498,I245515,I245546,I245563,I245622,I543502,I245653,I245731,I245748,I245714,I245693,I245793,I245810,I245827,I245844,I245861,I245878,I245895,I245912,I245929,I245720,I245960,I245977,I245994,I246011,I245723,I246042,I246059,I246076,I246093,I246110,I245708,I246141,I246158,I245711,I245705,I245699,I246217,I245717,I246248,I245702,I245696,I246326,I246343,I520312,I246360,I520321,I520303,I246377,I520324,I246394,I246411,I520315,I246428,I246445,I246315,I246476,I246300,I246507,I520309,I246524,I520300,I246541,I520297,I246558,I520294,I246575,I246592,I246609,I246297,I246640,I246657,I246294,I246688,I520318,I246705,I246312,I246736,I246309,I246767,I246784,I246288,I246291,I246829,I520306,I246846,I246863,I246880,I246318,I246911,I246303,I246306,I246989,I247006,I247023,I247040,I247057,I247074,I247091,I247108,I247139,I247170,I247187,I247204,I247221,I247238,I247255,I247272,I247303,I247320,I247351,I247368,I247399,I247430,I247447,I247492,I247509,I247526,I247543,I247574,I247652,I247669,I412571,I247686,I412574,I412580,I247703,I412586,I247720,I247737,I412565,I247754,I247771,I247802,I247833,I412577,I247850,I412592,I247867,I412595,I247884,I412568,I247901,I247918,I247935,I247966,I247983,I248014,I412589,I248031,I248062,I248093,I248110,I248155,I412583,I248172,I248189,I248206,I248237,I248315,I248332,I248349,I248366,I248383,I248400,I248417,I248434,I248465,I248496,I248513,I248530,I248547,I248564,I248581,I248598,I248629,I248646,I248677,I248694,I248725,I248756,I248773,I248818,I248835,I248852,I248869,I248900,I248978,I248995,I435598,I249012,I435610,I435592,I249029,I435613,I249046,I249063,I435604,I249080,I249097,I249128,I249159,I435595,I249176,I435589,I249193,I435601,I249210,I435586,I249227,I249244,I249261,I249292,I249309,I249340,I435583,I249357,I249388,I249419,I249436,I249481,I435607,I249498,I249515,I249532,I249563,I249641,I249658,I507817,I249675,I507826,I507808,I249692,I507829,I249709,I249726,I507820,I249743,I249760,I249630,I249791,I249615,I249822,I507814,I249839,I507805,I249856,I507802,I249873,I507799,I249890,I249907,I249924,I249612,I249955,I249972,I249609,I250003,I507823,I250020,I249627,I250051,I249624,I250082,I250099,I249603,I249606,I250144,I507811,I250161,I250178,I250195,I249633,I250226,I249618,I249621,I250304,I250321,I592902,I250338,I592899,I592890,I250355,I592893,I250372,I250389,I592887,I250406,I250423,I250293,I250454,I250278,I250485,I592908,I250502,I592911,I250519,I592896,I250536,I592884,I250553,I250570,I250587,I250275,I250618,I250635,I250272,I250666,I592905,I250683,I250290,I250714,I250287,I250745,I250762,I250266,I250269,I250807,I592914,I250824,I250841,I250858,I250296,I250889,I250281,I250284,I250967,I250984,I251001,I251018,I251035,I251052,I251069,I251086,I250956,I251117,I250941,I251148,I251165,I251182,I251199,I251216,I251233,I251250,I250938,I251281,I251298,I250935,I251329,I251346,I250953,I251377,I250950,I251408,I251425,I250929,I250932,I251470,I251487,I251504,I251521,I250959,I251552,I250944,I250947,I251630,I251647,I251664,I251681,I251698,I251715,I251732,I251749,I251780,I251811,I251828,I251845,I251862,I251879,I251896,I251913,I251944,I251961,I251992,I252009,I252040,I252071,I252088,I252133,I252150,I252167,I252184,I252215,I252293,I252310,I707714,I252327,I707705,I707711,I252344,I707723,I252361,I252378,I707708,I252395,I252412,I252282,I252443,I252267,I252474,I707732,I252491,I707726,I252508,I707717,I252525,I707702,I252542,I252559,I252576,I252264,I252607,I252624,I252261,I252655,I707720,I252672,I252279,I252703,I252276,I252734,I252751,I252255,I252258,I252796,I707729,I252813,I252830,I252847,I252285,I252878,I252270,I252273,I252956,I252973,I477214,I252990,I477226,I477208,I253007,I477229,I253024,I253041,I477220,I253058,I253075,I253106,I253137,I477211,I253154,I477205,I253171,I477217,I253188,I477202,I253205,I253222,I253239,I253270,I253287,I253318,I477199,I253335,I253366,I253397,I253414,I253459,I477223,I253476,I253493,I253510,I253541,I253619,I253636,I688532,I253653,I688550,I688541,I253670,I688547,I253687,I253704,I688553,I253721,I253738,I253608,I253769,I253593,I253800,I688529,I253817,I688544,I253834,I688526,I253851,I688535,I253868,I253885,I253902,I253590,I253933,I253950,I253587,I253981,I688538,I253998,I253605,I254029,I253602,I254060,I254077,I253581,I253584,I254122,I688556,I254139,I254156,I254173,I253611,I254204,I253596,I253599,I254282,I254299,I544112,I254316,I544121,I544103,I254333,I544124,I254350,I254367,I544115,I254384,I254401,I254271,I254432,I254256,I254463,I544109,I254480,I544100,I254497,I544097,I254514,I544094,I254531,I254548,I254565,I254253,I254596,I254613,I254250,I254644,I544118,I254661,I254268,I254692,I254265,I254723,I254740,I254244,I254247,I254785,I544106,I254802,I254819,I254836,I254274,I254867,I254259,I254262,I254945,I254962,I371267,I254979,I371264,I371282,I254996,I371285,I255013,I255030,I371270,I255047,I255064,I254934,I255095,I254919,I255126,I371279,I255143,I371261,I255160,I371255,I255177,I371273,I255194,I255211,I255228,I254916,I255259,I255276,I254913,I255307,I371258,I255324,I254931,I255355,I254928,I255386,I255403,I254907,I254910,I255448,I371276,I255465,I255482,I255499,I254937,I255530,I254922,I254925,I255608,I255625,I553632,I255642,I553641,I553623,I255659,I553644,I255676,I255693,I553635,I255710,I255727,I255758,I255789,I553629,I255806,I553620,I255823,I553617,I255840,I553614,I255857,I255874,I255891,I255922,I255939,I255970,I553638,I255987,I256018,I256049,I256066,I256111,I553626,I256128,I256145,I256162,I256193,I256271,I256288,I348657,I256305,I348654,I348672,I256322,I348675,I256339,I256356,I348660,I256373,I256390,I256260,I256421,I256245,I256452,I348669,I256469,I348651,I256486,I348645,I256503,I348663,I256520,I256537,I256554,I256242,I256585,I256602,I256239,I256633,I348648,I256650,I256257,I256681,I256254,I256712,I256729,I256233,I256236,I256774,I348666,I256791,I256808,I256825,I256263,I256856,I256248,I256251,I256934,I256951,I256968,I256985,I257002,I257019,I257036,I257053,I257084,I257115,I257132,I257149,I257166,I257183,I257200,I257217,I257248,I257265,I257296,I257313,I257344,I257375,I257392,I257437,I257454,I257471,I257488,I257519,I257597,I257614,I257631,I257648,I257665,I257682,I257699,I257716,I257747,I257778,I257795,I257812,I257829,I257846,I257863,I257880,I257911,I257928,I257959,I257976,I258007,I258038,I258055,I258100,I258117,I258134,I258151,I258182,I258260,I258277,I636954,I258294,I636972,I636963,I258311,I636969,I258328,I258345,I636975,I258362,I258379,I258249,I258410,I258234,I258441,I636951,I258458,I636966,I258475,I636948,I258492,I636957,I258509,I258526,I258543,I258231,I258574,I258591,I258228,I258622,I636960,I258639,I258246,I258670,I258243,I258701,I258718,I258222,I258225,I258763,I636978,I258780,I258797,I258814,I258252,I258845,I258237,I258240,I258923,I258940,I258957,I258974,I258991,I259008,I259025,I259042,I258912,I259073,I258897,I259104,I259121,I259138,I259155,I259172,I259189,I259206,I258894,I259237,I259254,I258891,I259285,I259302,I258909,I259333,I258906,I259364,I259381,I258885,I258888,I259426,I259443,I259460,I259477,I258915,I259508,I258900,I258903,I259586,I259603,I510197,I259620,I510206,I510188,I259637,I510209,I259654,I259671,I510200,I259688,I259705,I259736,I259767,I510194,I259784,I510185,I259801,I510182,I259818,I510179,I259835,I259852,I259869,I259900,I259917,I259948,I510203,I259965,I259996,I260027,I260044,I260089,I510191,I260106,I260123,I260140,I260171,I260249,I260266,I260283,I260300,I260317,I260334,I260351,I260368,I260238,I260399,I260223,I260430,I260447,I260464,I260481,I260498,I260515,I260532,I260220,I260563,I260580,I260217,I260611,I260628,I260235,I260659,I260232,I260690,I260707,I260211,I260214,I260752,I260769,I260786,I260803,I260241,I260834,I260226,I260229,I260912,I260929,I260946,I260963,I260980,I260997,I261014,I261031,I260901,I261062,I260886,I261093,I261110,I261127,I261144,I261161,I261178,I261195,I260883,I261226,I261243,I260880,I261274,I261291,I260898,I261322,I260895,I261353,I261370,I260874,I260877,I261415,I261432,I261449,I261466,I260904,I261497,I260889,I260892,I261575,I261592,I261609,I261626,I261643,I261660,I261677,I261694,I261725,I261756,I261773,I261790,I261807,I261824,I261841,I261858,I261889,I261906,I261937,I261954,I261985,I262016,I262033,I262078,I262095,I262112,I262129,I262160,I262238,I262255,I507222,I262272,I507231,I507213,I262289,I507234,I262306,I262323,I507225,I262340,I262357,I262227,I262388,I262212,I262419,I507219,I262436,I507210,I262453,I507207,I262470,I507204,I262487,I262504,I262521,I262209,I262552,I262569,I262206,I262600,I507228,I262617,I262224,I262648,I262221,I262679,I262696,I262200,I262203,I262741,I507216,I262758,I262775,I262792,I262230,I262823,I262215,I262218,I262901,I262918,I262935,I262952,I262969,I262986,I263003,I263020,I263051,I263082,I263099,I263116,I263133,I263150,I263167,I263184,I263215,I263232,I263263,I263280,I263311,I263342,I263359,I263404,I263421,I263438,I263455,I263486,I263564,I263581,I528642,I263598,I528651,I528633,I263615,I528654,I263632,I263649,I528645,I263666,I263683,I263553,I263714,I263538,I263745,I528639,I263762,I528630,I263779,I528627,I263796,I528624,I263813,I263830,I263847,I263535,I263878,I263895,I263532,I263926,I528648,I263943,I263550,I263974,I263547,I264005,I264022,I263526,I263529,I264067,I528636,I264084,I264101,I264118,I263556,I264149,I263541,I263544,I264227,I264244,I559582,I264261,I559591,I559573,I264278,I559594,I264295,I264312,I559585,I264329,I264346,I264377,I264408,I559579,I264425,I559570,I264442,I559567,I264459,I559564,I264476,I264493,I264510,I264541,I264558,I264589,I559588,I264606,I264637,I264668,I264685,I264730,I559576,I264747,I264764,I264781,I264812,I264890,I264907,I429095,I264924,I429098,I429104,I264941,I429110,I264958,I264975,I429089,I264992,I265009,I264879,I265040,I264864,I265071,I429101,I265088,I429116,I265105,I429119,I265122,I429092,I265139,I265156,I265173,I264861,I265204,I265221,I264858,I265252,I429113,I265269,I264876,I265300,I264873,I265331,I265348,I264852,I264855,I265393,I429107,I265410,I265427,I265444,I264882,I265475,I264867,I264870,I265553,I265570,I670920,I265587,I670938,I670929,I265604,I670935,I265621,I265638,I670941,I265655,I265672,I265703,I265734,I670917,I265751,I670932,I265768,I670914,I265785,I670923,I265802,I265819,I265836,I265867,I265884,I265915,I670926,I265932,I265963,I265994,I266011,I266056,I670944,I266073,I266090,I266107,I266138,I266216,I266233,I266250,I266267,I266284,I266301,I266318,I266335,I266366,I266397,I266414,I266431,I266448,I266465,I266482,I266499,I266530,I266547,I266578,I266595,I266626,I266657,I266674,I266719,I266736,I266753,I266770,I266801,I266879,I266896,I664001,I266913,I664019,I664010,I266930,I664016,I266947,I266964,I664022,I266981,I266998,I267029,I267060,I663998,I267077,I664013,I267094,I663995,I267111,I664004,I267128,I267145,I267162,I267193,I267210,I267241,I664007,I267258,I267289,I267320,I267337,I267382,I664025,I267399,I267416,I267433,I267464,I267542,I267559,I463342,I267576,I463354,I463336,I267593,I463357,I267610,I267627,I463348,I267644,I267661,I267531,I267692,I267516,I267723,I463339,I267740,I463333,I267757,I463345,I267774,I463330,I267791,I267808,I267825,I267513,I267856,I267873,I267510,I267904,I463327,I267921,I267528,I267952,I267525,I267983,I268000,I267504,I267507,I268045,I463351,I268062,I268079,I268096,I267534,I268127,I267519,I267522,I268205,I268222,I550657,I268239,I550666,I550648,I268256,I550669,I268273,I268290,I550660,I268307,I268324,I268194,I268355,I268179,I268386,I550654,I268403,I550645,I268420,I550642,I268437,I550639,I268454,I268471,I268488,I268176,I268519,I268536,I268173,I268567,I550663,I268584,I268191,I268615,I268188,I268646,I268663,I268167,I268170,I268708,I550651,I268725,I268742,I268759,I268197,I268790,I268182,I268185,I268868,I268885,I722742,I268902,I722733,I722739,I268919,I722751,I268936,I268953,I722736,I268970,I268987,I268857,I269018,I268842,I269049,I722760,I269066,I722754,I269083,I722745,I269100,I722730,I269117,I269134,I269151,I268839,I269182,I269199,I268836,I269230,I722748,I269247,I268854,I269278,I268851,I269309,I269326,I268830,I268833,I269371,I722757,I269388,I269405,I269422,I268860,I269453,I268845,I268848,I269531,I269548,I579217,I269565,I579214,I579205,I269582,I579208,I269599,I269616,I579202,I269633,I269650,I269520,I269681,I269505,I269712,I579223,I269729,I579226,I269746,I579211,I269763,I579199,I269780,I269797,I269814,I269502,I269845,I269862,I269499,I269893,I579220,I269910,I269517,I269941,I269514,I269972,I269989,I269493,I269496,I270034,I579229,I270051,I270068,I270085,I269523,I270116,I269508,I269511,I270194,I270211,I270228,I270245,I270262,I270279,I270296,I270313,I270183,I270344,I270168,I270375,I270392,I270409,I270426,I270443,I270460,I270477,I270165,I270508,I270525,I270162,I270556,I270573,I270180,I270604,I270177,I270635,I270652,I270156,I270159,I270697,I270714,I270731,I270748,I270186,I270779,I270171,I270174,I270857,I270874,I270891,I270908,I270925,I270942,I270959,I270976,I271007,I271038,I271055,I271072,I271089,I271106,I271123,I271140,I271171,I271188,I271219,I271236,I271267,I271298,I271315,I271360,I271377,I271394,I271411,I271442,I271520,I271537,I271554,I271571,I271588,I271605,I271622,I271639,I271509,I271670,I271494,I271701,I271718,I271735,I271752,I271769,I271786,I271803,I271491,I271834,I271851,I271488,I271882,I271899,I271506,I271930,I271503,I271961,I271978,I271482,I271485,I272023,I272040,I272057,I272074,I271512,I272105,I271497,I271500,I272183,I272200,I272217,I272234,I272251,I272268,I272285,I272302,I272172,I272333,I272157,I272364,I272381,I272398,I272415,I272432,I272449,I272466,I272154,I272497,I272514,I272151,I272545,I272562,I272169,I272593,I272166,I272624,I272641,I272145,I272148,I272686,I272703,I272720,I272737,I272175,I272768,I272160,I272163,I272846,I272863,I527452,I272880,I527461,I527443,I272897,I527464,I272914,I272931,I527455,I272948,I272965,I272835,I272996,I272820,I273027,I527449,I273044,I527440,I273061,I527437,I273078,I527434,I273095,I273112,I273129,I272817,I273160,I273177,I272814,I273208,I527458,I273225,I272832,I273256,I272829,I273287,I273304,I272808,I272811,I273349,I527446,I273366,I273383,I273400,I272838,I273431,I272823,I272826,I273509,I273526,I273543,I273560,I273577,I273594,I273611,I273628,I273498,I273659,I273483,I273690,I273707,I273724,I273741,I273758,I273775,I273792,I273480,I273823,I273840,I273477,I273871,I273888,I273495,I273919,I273492,I273950,I273967,I273471,I273474,I274012,I274029,I274046,I274063,I273501,I274094,I273486,I273489,I274172,I274189,I454672,I274206,I454684,I454666,I274223,I454687,I274240,I274257,I454678,I274274,I274291,I274161,I274322,I274146,I274353,I454669,I274370,I454663,I274387,I454675,I274404,I454660,I274421,I274438,I274455,I274143,I274486,I274503,I274140,I274534,I454657,I274551,I274158,I274582,I274155,I274613,I274630,I274134,I274137,I274675,I454681,I274692,I274709,I274726,I274164,I274757,I274149,I274152,I274835,I274852,I467966,I274869,I467978,I467960,I274886,I467981,I274903,I274920,I467972,I274937,I274954,I274824,I274985,I274809,I275016,I467963,I275033,I467957,I275050,I467969,I275067,I467954,I275084,I275101,I275118,I274806,I275149,I275166,I274803,I275197,I467951,I275214,I274821,I275245,I274818,I275276,I275293,I274797,I274800,I275338,I467975,I275355,I275372,I275389,I274827,I275420,I274812,I274815,I275498,I275515,I275532,I275549,I275566,I275583,I275600,I275617,I275487,I275648,I275472,I275679,I275696,I275713,I275730,I275747,I275764,I275781,I275469,I275812,I275829,I275466,I275860,I275877,I275484,I275908,I275481,I275939,I275956,I275460,I275463,I276001,I276018,I276035,I276052,I275490,I276083,I275475,I275478,I276161,I276178,I484728,I276195,I484740,I484722,I276212,I484743,I276229,I276246,I484734,I276263,I276280,I276311,I276342,I484725,I276359,I484719,I276376,I484731,I276393,I484716,I276410,I276427,I276444,I276475,I276492,I276523,I484713,I276540,I276571,I276602,I276619,I276664,I484737,I276681,I276698,I276715,I276746,I276824,I276841,I276858,I276875,I276892,I276909,I276926,I276943,I276813,I276974,I276798,I277005,I277022,I277039,I277056,I277073,I277090,I277107,I276795,I277138,I277155,I276792,I277186,I277203,I276810,I277234,I276807,I277265,I277282,I276786,I276789,I277327,I277344,I277361,I277378,I276816,I277409,I276801,I276804,I277487,I277504,I682242,I277521,I682260,I682251,I277538,I682257,I277555,I277572,I682263,I277589,I277606,I277476,I277637,I277461,I277668,I682239,I277685,I682254,I277702,I682236,I277719,I682245,I277736,I277753,I277770,I277458,I277801,I277818,I277455,I277849,I682248,I277866,I277473,I277897,I277470,I277928,I277945,I277449,I277452,I277990,I682266,I278007,I278024,I278041,I277479,I278072,I277464,I277467,I278150,I278167,I335091,I278184,I335088,I335106,I278201,I335109,I278218,I278235,I335094,I278252,I278269,I278139,I278300,I278124,I278331,I335103,I278348,I335085,I278365,I335079,I278382,I335097,I278399,I278416,I278433,I278121,I278464,I278481,I278118,I278512,I335082,I278529,I278136,I278560,I278133,I278591,I278608,I278112,I278115,I278653,I335100,I278670,I278687,I278704,I278142,I278735,I278127,I278130,I278813,I278830,I439644,I278847,I439656,I439638,I278864,I439659,I278881,I278898,I439650,I278915,I278932,I278802,I278963,I278787,I278994,I439641,I279011,I439635,I279028,I439647,I279045,I439632,I279062,I279079,I279096,I278784,I279127,I279144,I278781,I279175,I439629,I279192,I278799,I279223,I278796,I279254,I279271,I278775,I278778,I279316,I439653,I279333,I279350,I279367,I278805,I279398,I278790,I278793,I279476,I279493,I508412,I279510,I508421,I508403,I279527,I508424,I279544,I279561,I508415,I279578,I279595,I279465,I279626,I279450,I279657,I508409,I279674,I508400,I279691,I508397,I279708,I508394,I279725,I279742,I279759,I279447,I279790,I279807,I279444,I279838,I508418,I279855,I279462,I279886,I279459,I279917,I279934,I279438,I279441,I279979,I508406,I279996,I280013,I280030,I279468,I280061,I279453,I279456,I280139,I280156,I552442,I280173,I552451,I552433,I280190,I552454,I280207,I280224,I552445,I280241,I280258,I280128,I280289,I280113,I280320,I552439,I280337,I552430,I280354,I552427,I280371,I552424,I280388,I280405,I280422,I280110,I280453,I280470,I280107,I280501,I552448,I280518,I280125,I280549,I280122,I280580,I280597,I280101,I280104,I280642,I552436,I280659,I280676,I280693,I280131,I280724,I280116,I280119,I280802,I280819,I280836,I280853,I280870,I280887,I280904,I280921,I280952,I280983,I281000,I281017,I281034,I281051,I281068,I281085,I281116,I281133,I281164,I281181,I281212,I281243,I281260,I281305,I281322,I281339,I281356,I281387,I281465,I281482,I281499,I281516,I281533,I281550,I281567,I281584,I281615,I281646,I281663,I281680,I281697,I281714,I281731,I281748,I281779,I281796,I281827,I281844,I281875,I281906,I281923,I281968,I281985,I282002,I282019,I282050,I282128,I282145,I282162,I282179,I282196,I282213,I282230,I282247,I282278,I282309,I282326,I282343,I282360,I282377,I282394,I282411,I282442,I282459,I282490,I282507,I282538,I282569,I282586,I282631,I282648,I282665,I282682,I282713,I282791,I282808,I485884,I282825,I485896,I485878,I282842,I485899,I282859,I282876,I485890,I282893,I282910,I282780,I282941,I282765,I282972,I485881,I282989,I485875,I283006,I485887,I283023,I485872,I283040,I283057,I283074,I282762,I283105,I283122,I282759,I283153,I485869,I283170,I282777,I283201,I282774,I283232,I283249,I282753,I282756,I283294,I485893,I283311,I283328,I283345,I282783,I283376,I282768,I282771,I283454,I283471,I283488,I283505,I283522,I283539,I283556,I283573,I283443,I283604,I283428,I283635,I283652,I283669,I283686,I283703,I283720,I283737,I283425,I283768,I283785,I283422,I283816,I283833,I283440,I283864,I283437,I283895,I283912,I283416,I283419,I283957,I283974,I283991,I284008,I283446,I284039,I283431,I283434,I284117,I284134,I373851,I284151,I373848,I373866,I284168,I373869,I284185,I284202,I373854,I284219,I284236,I284106,I284267,I284091,I284298,I373863,I284315,I373845,I284332,I373839,I284349,I373857,I284366,I284383,I284400,I284088,I284431,I284448,I284085,I284479,I373842,I284496,I284103,I284527,I284100,I284558,I284575,I284079,I284082,I284620,I373860,I284637,I284654,I284671,I284109,I284702,I284094,I284097,I284780,I284797,I550062,I284814,I550071,I550053,I284831,I550074,I284848,I284865,I550065,I284882,I284899,I284930,I284961,I550059,I284978,I550050,I284995,I550047,I285012,I550044,I285029,I285046,I285063,I285094,I285111,I285142,I550068,I285159,I285190,I285221,I285238,I285283,I550056,I285300,I285317,I285334,I285365,I285443,I285460,I584572,I285477,I584569,I584560,I285494,I584563,I285511,I285528,I584557,I285545,I285562,I285432,I285593,I285417,I285624,I584578,I285641,I584581,I285658,I584566,I285675,I584554,I285692,I285709,I285726,I285414,I285757,I285774,I285411,I285805,I584575,I285822,I285429,I285853,I285426,I285884,I285901,I285405,I285408,I285946,I584584,I285963,I285980,I285997,I285435,I286028,I285420,I285423,I286106,I286123,I456984,I286140,I456996,I456978,I286157,I456999,I286174,I286191,I456990,I286208,I286225,I286095,I286256,I286080,I286287,I456981,I286304,I456975,I286321,I456987,I286338,I456972,I286355,I286372,I286389,I286077,I286420,I286437,I286074,I286468,I456969,I286485,I286092,I286516,I286089,I286547,I286564,I286068,I286071,I286609,I456993,I286626,I286643,I286660,I286098,I286691,I286083,I286086,I286769,I286786,I451782,I286803,I451794,I451776,I286820,I451797,I286837,I286854,I451788,I286871,I286888,I286758,I286919,I286743,I286950,I451779,I286967,I451773,I286984,I451785,I287001,I451770,I287018,I287035,I287052,I286740,I287083,I287100,I286737,I287131,I451767,I287148,I286755,I287179,I286752,I287210,I287227,I286731,I286734,I287272,I451791,I287289,I287306,I287323,I286761,I287354,I286746,I286749,I287432,I287449,I351241,I287466,I351238,I351256,I287483,I351259,I287500,I287517,I351244,I287534,I287551,I287421,I287582,I287406,I287613,I351253,I287630,I351235,I287647,I351229,I287664,I351247,I287681,I287698,I287715,I287403,I287746,I287763,I287400,I287794,I351232,I287811,I287418,I287842,I287415,I287873,I287890,I287394,I287397,I287935,I351250,I287952,I287969,I287986,I287424,I288017,I287409,I287412,I288095,I288112,I338321,I288129,I338318,I338336,I288146,I338339,I288163,I288180,I338324,I288197,I288214,I288245,I288276,I338333,I288293,I338315,I288310,I338309,I288327,I338327,I288344,I288361,I288378,I288409,I288426,I288457,I338312,I288474,I288505,I288536,I288553,I288598,I338330,I288615,I288632,I288649,I288680,I288758,I288775,I288792,I288809,I288826,I288843,I288860,I288877,I288908,I288939,I288956,I288973,I288990,I289007,I289024,I289041,I289072,I289089,I289120,I289137,I289168,I289199,I289216,I289261,I289278,I289295,I289312,I289343,I289421,I289438,I487043,I289455,I487040,I487037,I289472,I487025,I289489,I289506,I487046,I289523,I289540,I289571,I289602,I487028,I289619,I487034,I289636,I487031,I289653,I487055,I289670,I289687,I289704,I289735,I289752,I289783,I487052,I289800,I289831,I289862,I289879,I289924,I487049,I289941,I289958,I289975,I290006,I290084,I290101,I290118,I290135,I290152,I290169,I290186,I290203,I290234,I290265,I290282,I290299,I290316,I290333,I290350,I290367,I290398,I290415,I290446,I290463,I290494,I290525,I290542,I290587,I290604,I290621,I290638,I290669,I290747,I290764,I663372,I290781,I663390,I663381,I290798,I663387,I290815,I290832,I663393,I290849,I290866,I290897,I290928,I663369,I290945,I663384,I290962,I663366,I290979,I663375,I290996,I291013,I291030,I291061,I291078,I291109,I663378,I291126,I291157,I291188,I291205,I291250,I663396,I291267,I291284,I291301,I291332,I291410,I291427,I644502,I291444,I644520,I644511,I291461,I644517,I291478,I291495,I644523,I291512,I291529,I291399,I291560,I291384,I291591,I644499,I291608,I644514,I291625,I644496,I291642,I644505,I291659,I291676,I291693,I291381,I291724,I291741,I291378,I291772,I644508,I291789,I291396,I291820,I291393,I291851,I291868,I291372,I291375,I291913,I644526,I291930,I291947,I291964,I291402,I291995,I291387,I291390,I292073,I292090,I292107,I292124,I292141,I292158,I292175,I292192,I292062,I292223,I292047,I292254,I292271,I292288,I292305,I292322,I292339,I292356,I292044,I292387,I292404,I292041,I292435,I292452,I292059,I292483,I292056,I292514,I292531,I292035,I292038,I292576,I292593,I292610,I292627,I292065,I292658,I292050,I292053,I292736,I292753,I292770,I292787,I292804,I292821,I292838,I292855,I292725,I292886,I292710,I292917,I292934,I292951,I292968,I292985,I293002,I293019,I292707,I293050,I293067,I292704,I293098,I293115,I292722,I293146,I292719,I293177,I293194,I292698,I292701,I293239,I293256,I293273,I293290,I292728,I293321,I292713,I292716,I293399,I293416,I399045,I293433,I399042,I399060,I293450,I399063,I293467,I293484,I399048,I293501,I293518,I293388,I293549,I293373,I293580,I399057,I293597,I399039,I293614,I399033,I293631,I399051,I293648,I293665,I293682,I293370,I293713,I293730,I293367,I293761,I399036,I293778,I293385,I293809,I293382,I293840,I293857,I293361,I293364,I293902,I399054,I293919,I293936,I293953,I293391,I293984,I293376,I293379,I294062,I294079,I645760,I294096,I645778,I645769,I294113,I645775,I294130,I294147,I645781,I294164,I294181,I294051,I294212,I294036,I294243,I645757,I294260,I645772,I294277,I645754,I294294,I645763,I294311,I294328,I294345,I294033,I294376,I294393,I294030,I294424,I645766,I294441,I294048,I294472,I294045,I294503,I294520,I294024,I294027,I294565,I645784,I294582,I294599,I294616,I294054,I294647,I294039,I294042,I294725,I294742,I642615,I294759,I642633,I642624,I294776,I642630,I294793,I294810,I642636,I294827,I294844,I294875,I294906,I642612,I294923,I642627,I294940,I642609,I294957,I642618,I294974,I294991,I295008,I295039,I295056,I295087,I642621,I295104,I295135,I295166,I295183,I295228,I642639,I295245,I295262,I295279,I295310,I295388,I295405,I295422,I295439,I295456,I295473,I295490,I295507,I295377,I295538,I295362,I295569,I295586,I295603,I295620,I295637,I295654,I295671,I295359,I295702,I295719,I295356,I295750,I295767,I295374,I295798,I295371,I295829,I295846,I295350,I295353,I295891,I295908,I295925,I295942,I295380,I295973,I295365,I295368,I296051,I296068,I357055,I296085,I357052,I357070,I296102,I357073,I296119,I296136,I357058,I296153,I296170,I296040,I296201,I296025,I296232,I357067,I296249,I357049,I296266,I357043,I296283,I357061,I296300,I296317,I296334,I296022,I296365,I296382,I296019,I296413,I357046,I296430,I296037,I296461,I296034,I296492,I296509,I296013,I296016,I296554,I357064,I296571,I296588,I296605,I296043,I296636,I296028,I296031,I296714,I296731,I591117,I296748,I591114,I591105,I296765,I591108,I296782,I296799,I591102,I296816,I296833,I296864,I296895,I591123,I296912,I591126,I296929,I591111,I296946,I591099,I296963,I296980,I296997,I297028,I297045,I297076,I591120,I297093,I297124,I297155,I297172,I297217,I591129,I297234,I297251,I297268,I297299,I297377,I297394,I297411,I297428,I297445,I297462,I297479,I297496,I297527,I297558,I297575,I297592,I297609,I297626,I297643,I297660,I297691,I297708,I297739,I297756,I297787,I297818,I297835,I297880,I297897,I297914,I297931,I297962,I298040,I298057,I647018,I298074,I647036,I647027,I298091,I647033,I298108,I298125,I647039,I298142,I298159,I298029,I298190,I298014,I298221,I647015,I298238,I647030,I298255,I647012,I298272,I647021,I298289,I298306,I298323,I298011,I298354,I298371,I298008,I298402,I647024,I298419,I298026,I298450,I298023,I298481,I298498,I298002,I298005,I298543,I647042,I298560,I298577,I298594,I298032,I298625,I298017,I298020,I298703,I298720,I491327,I298737,I491324,I491321,I298754,I491309,I298771,I298788,I491330,I298805,I298822,I298692,I298853,I298677,I298884,I491312,I298901,I491318,I298918,I491315,I298935,I491339,I298952,I298969,I298986,I298674,I299017,I299034,I298671,I299065,I491336,I299082,I298689,I299113,I298686,I299144,I299161,I298665,I298668,I299206,I491333,I299223,I299240,I299257,I298695,I299288,I298680,I298683,I299366,I299383,I299400,I299417,I299434,I299451,I299468,I299485,I299355,I299516,I299340,I299547,I299564,I299581,I299598,I299615,I299632,I299649,I299337,I299680,I299697,I299334,I299728,I299745,I299352,I299776,I299349,I299807,I299824,I299328,I299331,I299869,I299886,I299903,I299920,I299358,I299951,I299343,I299346,I300029,I300046,I406797,I300063,I406794,I406812,I300080,I406815,I300097,I300114,I406800,I300131,I300148,I300018,I300179,I300003,I300210,I406809,I300227,I406791,I300244,I406785,I300261,I406803,I300278,I300295,I300312,I300000,I300343,I300360,I299997,I300391,I406788,I300408,I300015,I300439,I300012,I300470,I300487,I299991,I299994,I300532,I406806,I300549,I300566,I300583,I300021,I300614,I300006,I300009,I300692,I300709,I524477,I300726,I524486,I524468,I300743,I524489,I300760,I300777,I524480,I300794,I300811,I300842,I300873,I524474,I300890,I524465,I300907,I524462,I300924,I524459,I300941,I300958,I300975,I301006,I301023,I301054,I524483,I301071,I301102,I301133,I301150,I301195,I524471,I301212,I301229,I301246,I301277,I301355,I301372,I354471,I301389,I354468,I354486,I301406,I354489,I301423,I301440,I354474,I301457,I301474,I301344,I301505,I301329,I301536,I354483,I301553,I354465,I301570,I354459,I301587,I354477,I301604,I301621,I301638,I301326,I301669,I301686,I301323,I301717,I354462,I301734,I301341,I301765,I301338,I301796,I301813,I301317,I301320,I301858,I354480,I301875,I301892,I301909,I301347,I301940,I301332,I301335,I302018,I302035,I690374,I302052,I690365,I690371,I302069,I690383,I302086,I302103,I690368,I302120,I302137,I302007,I302168,I301992,I302199,I690392,I302216,I690386,I302233,I690377,I302250,I690362,I302267,I302284,I302301,I301989,I302332,I302349,I301986,I302380,I690380,I302397,I302004,I302428,I302001,I302459,I302476,I301980,I301983,I302521,I690389,I302538,I302555,I302572,I302010,I302603,I301995,I301998,I302681,I302698,I700778,I302715,I700769,I700775,I302732,I700787,I302749,I302766,I700772,I302783,I302800,I302670,I302831,I302655,I302862,I700796,I302879,I700790,I302896,I700781,I302913,I700766,I302930,I302947,I302964,I302652,I302995,I303012,I302649,I303043,I700784,I303060,I302667,I303091,I302664,I303122,I303139,I302643,I302646,I303184,I700793,I303201,I303218,I303235,I302673,I303266,I302658,I302661,I303344,I303361,I303378,I303395,I303412,I303429,I303446,I303463,I303494,I303525,I303542,I303559,I303576,I303593,I303610,I303627,I303658,I303675,I303706,I303723,I303754,I303785,I303802,I303847,I303864,I303881,I303898,I303929,I304007,I304024,I577432,I304041,I577429,I577420,I304058,I577423,I304075,I304092,I577417,I304109,I304126,I303996,I304157,I303981,I304188,I577438,I304205,I577441,I304222,I577426,I304239,I577414,I304256,I304273,I304290,I303978,I304321,I304338,I303975,I304369,I577435,I304386,I303993,I304417,I303990,I304448,I304465,I303969,I303972,I304510,I577444,I304527,I304544,I304561,I303999,I304592,I303984,I303987,I304670,I304687,I514957,I304704,I514966,I514948,I304721,I514969,I304738,I304755,I514960,I304772,I304789,I304820,I304851,I514954,I304868,I514945,I304885,I514942,I304902,I514939,I304919,I304936,I304953,I304984,I305001,I305032,I514963,I305049,I305080,I305111,I305128,I305173,I514951,I305190,I305207,I305224,I305255,I305333,I305350,I710604,I305367,I710595,I710601,I305384,I710613,I305401,I305418,I710598,I305435,I305452,I305322,I305483,I305307,I305514,I710622,I305531,I710616,I305548,I710607,I305565,I710592,I305582,I305599,I305616,I305304,I305647,I305664,I305301,I305695,I710610,I305712,I305319,I305743,I305316,I305774,I305791,I305295,I305298,I305836,I710619,I305853,I305870,I305887,I305325,I305918,I305310,I305313,I305996,I306013,I306030,I306047,I306064,I306081,I306098,I306115,I305985,I306146,I305970,I306177,I306194,I306211,I306228,I306245,I306262,I306279,I305967,I306310,I306327,I305964,I306358,I306375,I305982,I306406,I305979,I306437,I306454,I305958,I305961,I306499,I306516,I306533,I306550,I305988,I306581,I305973,I305976,I306659,I306676,I420527,I306693,I420530,I420536,I306710,I420542,I306727,I306744,I420521,I306761,I306778,I306648,I306809,I306633,I306840,I420533,I306857,I420548,I306874,I420551,I306891,I420524,I306908,I306925,I306942,I306630,I306973,I306990,I306627,I307021,I420545,I307038,I306645,I307069,I306642,I307100,I307117,I306621,I306624,I307162,I420539,I307179,I307196,I307213,I306651,I307244,I306636,I306639,I307322,I307339,I567317,I307356,I567326,I567308,I307373,I567329,I307390,I307407,I567320,I307424,I307441,I307311,I307472,I307296,I307503,I567314,I307520,I567305,I307537,I567302,I307554,I567299,I307571,I307588,I307605,I307293,I307636,I307653,I307290,I307684,I567323,I307701,I307308,I307732,I307305,I307763,I307780,I307284,I307287,I307825,I567311,I307842,I307859,I307876,I307314,I307907,I307299,I307302,I307985,I308002,I308019,I308036,I308053,I308070,I308087,I308104,I307974,I308135,I307959,I308166,I308183,I308200,I308217,I308234,I308251,I308268,I307956,I308299,I308316,I307953,I308347,I308364,I307971,I308395,I307968,I308426,I308443,I307947,I307950,I308488,I308505,I308522,I308539,I307977,I308570,I307962,I307965,I308648,I308665,I373205,I308682,I373202,I373220,I308699,I373223,I308716,I308733,I373208,I308750,I308767,I308637,I308798,I308622,I308829,I373217,I308846,I373199,I308863,I373193,I308880,I373211,I308897,I308914,I308931,I308619,I308962,I308979,I308616,I309010,I373196,I309027,I308634,I309058,I308631,I309089,I309106,I308610,I308613,I309151,I373214,I309168,I309185,I309202,I308640,I309233,I308625,I308628,I309311,I309328,I569697,I309345,I569706,I569688,I309362,I569709,I309379,I309396,I569700,I309413,I309430,I309461,I309492,I569694,I309509,I569685,I309526,I569682,I309543,I569679,I309560,I309577,I309594,I309625,I309642,I309673,I569703,I309690,I309721,I309752,I309769,I309814,I569691,I309831,I309848,I309865,I309896,I309974,I309991,I310008,I310025,I310042,I310059,I310076,I310093,I309963,I310124,I309948,I310155,I310172,I310189,I310206,I310223,I310240,I310257,I309945,I310288,I310305,I309942,I310336,I310353,I309960,I310384,I309957,I310415,I310432,I309936,I309939,I310477,I310494,I310511,I310528,I309966,I310559,I309951,I309954,I310637,I310654,I447158,I310671,I447170,I447152,I310688,I447173,I310705,I310722,I447164,I310739,I310756,I310626,I310787,I310611,I310818,I447155,I310835,I447149,I310852,I447161,I310869,I447146,I310886,I310903,I310920,I310608,I310951,I310968,I310605,I310999,I447143,I311016,I310623,I311047,I310620,I311078,I311095,I310599,I310602,I311140,I447167,I311157,I311174,I311191,I310629,I311222,I310614,I310617,I311300,I311317,I675952,I311334,I675970,I675961,I311351,I675967,I311368,I311385,I675973,I311402,I311419,I311289,I311450,I311274,I311481,I675949,I311498,I675964,I311515,I675946,I311532,I675955,I311549,I311566,I311583,I311271,I311614,I311631,I311268,I311662,I675958,I311679,I311286,I311710,I311283,I311741,I311758,I311262,I311265,I311803,I675976,I311820,I311837,I311854,I311292,I311885,I311277,I311280,I311963,I311980,I311997,I312014,I312031,I312048,I312065,I312082,I311952,I312113,I311937,I312144,I312161,I312178,I312195,I312212,I312229,I312246,I311934,I312277,I312294,I311931,I312325,I312342,I311949,I312373,I311946,I312404,I312421,I311925,I311928,I312466,I312483,I312500,I312517,I311955,I312548,I311940,I311943,I312626,I312643,I670291,I312660,I670309,I670300,I312677,I670306,I312694,I312711,I670312,I312728,I312745,I312615,I312776,I312600,I312807,I670288,I312824,I670303,I312841,I670285,I312858,I670294,I312875,I312892,I312909,I312597,I312940,I312957,I312594,I312988,I670297,I313005,I312612,I313036,I312609,I313067,I313084,I312588,I312591,I313129,I670315,I313146,I313163,I313180,I312618,I313211,I312603,I312606,I313289,I313306,I519717,I313323,I519726,I519708,I313340,I519729,I313357,I313374,I519720,I313391,I313408,I313278,I313439,I313263,I313470,I519714,I313487,I519705,I313504,I519702,I313521,I519699,I313538,I313555,I313572,I313260,I313603,I313620,I313257,I313651,I519723,I313668,I313275,I313699,I313272,I313730,I313747,I313251,I313254,I313792,I519711,I313809,I313826,I313843,I313281,I313874,I313266,I313269,I313952,I313969,I699044,I313986,I699035,I699041,I314003,I699053,I314020,I314037,I699038,I314054,I314071,I314102,I314133,I699062,I314150,I699056,I314167,I699047,I314184,I699032,I314201,I314218,I314235,I314266,I314283,I314314,I699050,I314331,I314362,I314393,I314410,I314455,I699059,I314472,I314489,I314506,I314537,I314615,I314632,I314649,I314666,I314683,I314700,I314717,I314734,I314765,I314796,I314813,I314830,I314847,I314864,I314881,I314898,I314929,I314946,I314977,I314994,I315025,I315056,I315073,I315118,I315135,I315152,I315169,I315200,I315278,I315295,I315312,I315329,I315346,I315363,I315380,I315397,I315267,I315428,I315252,I315459,I315476,I315493,I315510,I315527,I315544,I315561,I315249,I315592,I315609,I315246,I315640,I315657,I315264,I315688,I315261,I315719,I315736,I315240,I315243,I315781,I315798,I315815,I315832,I315270,I315863,I315255,I315258,I315941,I315958,I355763,I315975,I355760,I355778,I315992,I355781,I316009,I316026,I355766,I316043,I316060,I316091,I316122,I355775,I316139,I355757,I316156,I355751,I316173,I355769,I316190,I316207,I316224,I316255,I316272,I316303,I355754,I316320,I316351,I316382,I316399,I316444,I355772,I316461,I316478,I316495,I316526,I316604,I316621,I316638,I316655,I316672,I316689,I316706,I316723,I316754,I316785,I316802,I316819,I316836,I316853,I316870,I316887,I316918,I316935,I316966,I316983,I317014,I317045,I317062,I317107,I317124,I317141,I317158,I317189,I317267,I317284,I727366,I317301,I727357,I727363,I317318,I727375,I317335,I317352,I727360,I317369,I317386,I317256,I317417,I317241,I317448,I727384,I317465,I727378,I317482,I727369,I317499,I727354,I317516,I317533,I317550,I317238,I317581,I317598,I317235,I317629,I727372,I317646,I317253,I317677,I317250,I317708,I317725,I317229,I317232,I317770,I727381,I317787,I317804,I317821,I317259,I317852,I317244,I317247,I317930,I317947,I317964,I317981,I317998,I318015,I318032,I318049,I317919,I318080,I317904,I318111,I318128,I318145,I318162,I318179,I318196,I318213,I317901,I318244,I318261,I317898,I318292,I318309,I317916,I318340,I317913,I318371,I318388,I317892,I317895,I318433,I318450,I318467,I318484,I317922,I318515,I317907,I317910,I318593,I318610,I624374,I318627,I624392,I624383,I318644,I624389,I318661,I318678,I624395,I318695,I318712,I318582,I318743,I318567,I318774,I624371,I318791,I624386,I318808,I624368,I318825,I624377,I318842,I318859,I318876,I318564,I318907,I318924,I318561,I318955,I624380,I318972,I318579,I319003,I318576,I319034,I319051,I318555,I318558,I319096,I624398,I319113,I319130,I319147,I318585,I319178,I318570,I318573,I319256,I319273,I319290,I319307,I319324,I319341,I319358,I319375,I319245,I319406,I319230,I319437,I319454,I319471,I319488,I319505,I319522,I319539,I319227,I319570,I319587,I319224,I319618,I319635,I319242,I319666,I319239,I319697,I319714,I319218,I319221,I319759,I319776,I319793,I319810,I319248,I319841,I319233,I319236,I319919,I319936,I319953,I319970,I319987,I320004,I320021,I320038,I319908,I320069,I319893,I320100,I320117,I320134,I320151,I320168,I320185,I320202,I319890,I320233,I320250,I319887,I320281,I320298,I319905,I320329,I319902,I320360,I320377,I319881,I319884,I320422,I320439,I320456,I320473,I319911,I320504,I319896,I319899,I320582,I320599,I320616,I320633,I320650,I320667,I320684,I320701,I320732,I320763,I320780,I320797,I320814,I320831,I320848,I320865,I320896,I320913,I320944,I320961,I320992,I321023,I321040,I321085,I321102,I321119,I321136,I321167,I321245,I321262,I321279,I321296,I321313,I321330,I321347,I321364,I321234,I321395,I321219,I321426,I321443,I321460,I321477,I321494,I321511,I321528,I321216,I321559,I321576,I321213,I321607,I321624,I321231,I321655,I321228,I321686,I321703,I321207,I321210,I321748,I321765,I321782,I321799,I321237,I321830,I321222,I321225,I321908,I321925,I398399,I321942,I398396,I398414,I321959,I398417,I321976,I321993,I398402,I322010,I322027,I322058,I322089,I398411,I322106,I398393,I322123,I398387,I322140,I398405,I322157,I322174,I322191,I322222,I322239,I322270,I398390,I322287,I322318,I322349,I322366,I322411,I398408,I322428,I322445,I322462,I322493,I322571,I322588,I322605,I322622,I322639,I322656,I322673,I322690,I322721,I322752,I322769,I322786,I322803,I322820,I322837,I322854,I322885,I322902,I322933,I322950,I322981,I323012,I323029,I323074,I323091,I323108,I323125,I323156,I323234,I323251,I582787,I323268,I582784,I582775,I323285,I582778,I323302,I323319,I582772,I323336,I323353,I323223,I323384,I323208,I323415,I582793,I323432,I582796,I323449,I582781,I323466,I582769,I323483,I323500,I323517,I323205,I323548,I323565,I323202,I323596,I582790,I323613,I323220,I323644,I323217,I323675,I323692,I323196,I323199,I323737,I582799,I323754,I323771,I323788,I323226,I323819,I323211,I323214,I323897,I323914,I323931,I323948,I323965,I323982,I323999,I324016,I323886,I324047,I323871,I324078,I324095,I324112,I324129,I324146,I324163,I324180,I323868,I324211,I324228,I323865,I324259,I324276,I323883,I324307,I323880,I324338,I324355,I323859,I323862,I324400,I324417,I324434,I324451,I323889,I324482,I323874,I323877,I324560,I324577,I324594,I324611,I324628,I324645,I324662,I324679,I324710,I324741,I324758,I324775,I324792,I324809,I324826,I324843,I324874,I324891,I324922,I324939,I324970,I325001,I325018,I325063,I325080,I325097,I325114,I325145,I325223,I325240,I325257,I325274,I325291,I325308,I325325,I325342,I325373,I325404,I325421,I325438,I325455,I325472,I325489,I325506,I325537,I325554,I325585,I325602,I325633,I325664,I325681,I325726,I325743,I325760,I325777,I325808,I325886,I325903,I325920,I325937,I325954,I325971,I325988,I326005,I325875,I326036,I325860,I326067,I326084,I326101,I326118,I326135,I326152,I326169,I325857,I326200,I326217,I325854,I326248,I326265,I325872,I326296,I325869,I326327,I326344,I325848,I325851,I326389,I326406,I326423,I326440,I325878,I326471,I325863,I325866,I326549,I326566,I326583,I326600,I326617,I326634,I326651,I326668,I326699,I326730,I326747,I326764,I326781,I326798,I326815,I326832,I326863,I326880,I326911,I326928,I326959,I326990,I327007,I327052,I327069,I327086,I327103,I327134,I327212,I327229,I633809,I327246,I633827,I633818,I327263,I633824,I327280,I327297,I633830,I327314,I327331,I327362,I327393,I633806,I327410,I633821,I327427,I633803,I327444,I633812,I327461,I327478,I327495,I327526,I327543,I327574,I633815,I327591,I327622,I327653,I327670,I327715,I633833,I327732,I327749,I327766,I327797,I327875,I327892,I626261,I327909,I626279,I626270,I327926,I626276,I327943,I327960,I626282,I327977,I327994,I327864,I328025,I327849,I328056,I626258,I328073,I626273,I328090,I626255,I328107,I626264,I328124,I328141,I328158,I327846,I328189,I328206,I327843,I328237,I626267,I328254,I327861,I328285,I327858,I328316,I328333,I327837,I327840,I328378,I626285,I328395,I328412,I328429,I327867,I328460,I327852,I327855,I328538,I328555,I482994,I328572,I483006,I482988,I328589,I483009,I328606,I328623,I483000,I328640,I328657,I328527,I328688,I328512,I328719,I482991,I328736,I482985,I328753,I482997,I328770,I482982,I328787,I328804,I328821,I328509,I328852,I328869,I328506,I328900,I482979,I328917,I328524,I328948,I328521,I328979,I328996,I328500,I328503,I329041,I483003,I329058,I329075,I329092,I328530,I329123,I328515,I328518,I329201,I329218,I479526,I329235,I479538,I479520,I329252,I479541,I329269,I329286,I479532,I329303,I329320,I329351,I329382,I479523,I329399,I479517,I329416,I479529,I329433,I479514,I329450,I329467,I329484,I329515,I329532,I329563,I479511,I329580,I329611,I329642,I329659,I329704,I479535,I329721,I329738,I329755,I329786,I329864,I329881,I375789,I329898,I375786,I375804,I329915,I375807,I329932,I329949,I375792,I329966,I329983,I329853,I330014,I329838,I330045,I375801,I330062,I375783,I330079,I375777,I330096,I375795,I330113,I330130,I330147,I329835,I330178,I330195,I329832,I330226,I375780,I330243,I329850,I330274,I329847,I330305,I330322,I329826,I329829,I330367,I375798,I330384,I330401,I330418,I329856,I330449,I329841,I329844,I330527,I330544,I330561,I330578,I330595,I330612,I330629,I330646,I330516,I330677,I330501,I330708,I330725,I330742,I330759,I330776,I330793,I330810,I330498,I330841,I330858,I330495,I330889,I330906,I330513,I330937,I330510,I330968,I330985,I330489,I330492,I331030,I331047,I331064,I331081,I330519,I331112,I330504,I330507,I331190,I331207,I477792,I331224,I477804,I477786,I331241,I477807,I331258,I331275,I477798,I331292,I331309,I331179,I331340,I331164,I331371,I477789,I331388,I477783,I331405,I477795,I331422,I477780,I331439,I331456,I331473,I331161,I331504,I331521,I331158,I331552,I477777,I331569,I331176,I331600,I331173,I331631,I331648,I331152,I331155,I331693,I477801,I331710,I331727,I331744,I331182,I331775,I331167,I331170,I331853,I331870,I488267,I331887,I488264,I488261,I331904,I488249,I331921,I331938,I488270,I331955,I331972,I332003,I332034,I488252,I332051,I488258,I332068,I488255,I332085,I488279,I332102,I332119,I332136,I332167,I332184,I332215,I488276,I332232,I332263,I332294,I332311,I332356,I488273,I332373,I332390,I332407,I332438,I332516,I332533,I332550,I332567,I332584,I332601,I332618,I332635,I332505,I332666,I332490,I332697,I332714,I332731,I332748,I332765,I332782,I332799,I332487,I332830,I332847,I332484,I332878,I332895,I332502,I332926,I332499,I332957,I332974,I332478,I332481,I333019,I333036,I333053,I333070,I332508,I333101,I332493,I332496,I333179,I333196,I333213,I333230,I333247,I333264,I333281,I333150,I333312,I333329,I333346,I333363,I333380,I333397,I333414,I333147,I333445,I333141,I333476,I333493,I333510,I333171,I333144,I333555,I333168,I333586,I333165,I333162,I333631,I333648,I333665,I333682,I333699,I333156,I333730,I333747,I333159,I333153,I333825,I333842,I333859,I333876,I333893,I333910,I333927,I333796,I333958,I333975,I333992,I334009,I334026,I334043,I334060,I333793,I334091,I333787,I334122,I334139,I334156,I333817,I333790,I334201,I333814,I334232,I333811,I333808,I334277,I334294,I334311,I334328,I334345,I333802,I334376,I334393,I333805,I333799,I334471,I334488,I334505,I334522,I334539,I334556,I334573,I334604,I334621,I334638,I334655,I334672,I334689,I334706,I334737,I334768,I334785,I334802,I334847,I334878,I334923,I334940,I334957,I334974,I334991,I335022,I335039,I335117,I335134,I335151,I335168,I335185,I335202,I335219,I335250,I335267,I335284,I335301,I335318,I335335,I335352,I335383,I335414,I335431,I335448,I335493,I335524,I335569,I335586,I335603,I335620,I335637,I335668,I335685,I335763,I335780,I636340,I335797,I636337,I636322,I335814,I636331,I335831,I335848,I636346,I335865,I335734,I335896,I335913,I335930,I636319,I335947,I636325,I335964,I636349,I335981,I636343,I335998,I335731,I336029,I335725,I336060,I336077,I336094,I335755,I335728,I336139,I636328,I335752,I336170,I335749,I335746,I336215,I636334,I336232,I336249,I336266,I336283,I335740,I336314,I336331,I335743,I335737,I336409,I336426,I336443,I336460,I336477,I336494,I336511,I336380,I336542,I336559,I336576,I336593,I336610,I336627,I336644,I336377,I336675,I336371,I336706,I336723,I336740,I336401,I336374,I336785,I336398,I336816,I336395,I336392,I336861,I336878,I336895,I336912,I336929,I336386,I336960,I336977,I336389,I336383,I337055,I337072,I337089,I337106,I337123,I337140,I337157,I337188,I337205,I337222,I337239,I337256,I337273,I337290,I337321,I337352,I337369,I337386,I337431,I337462,I337507,I337524,I337541,I337558,I337575,I337606,I337623,I337701,I337718,I337735,I337752,I337769,I337786,I337803,I337672,I337834,I337851,I337868,I337885,I337902,I337919,I337936,I337669,I337967,I337663,I337998,I338015,I338032,I337693,I337666,I338077,I337690,I338108,I337687,I337684,I338153,I338170,I338187,I338204,I338221,I337678,I338252,I338269,I337681,I337675,I338347,I338364,I561358,I338381,I561370,I561364,I338398,I561349,I338415,I338432,I561376,I338449,I338480,I338497,I338514,I561373,I338531,I561355,I338548,I561352,I338565,I561379,I338582,I338613,I338644,I338661,I338678,I338723,I561367,I338754,I338799,I561361,I338816,I338833,I338850,I338867,I338898,I338915,I338993,I339010,I339027,I339044,I339061,I339078,I339095,I339126,I339143,I339160,I339177,I339194,I339211,I339228,I339259,I339290,I339307,I339324,I339369,I339400,I339445,I339462,I339479,I339496,I339513,I339544,I339561,I339639,I339656,I558383,I339673,I558395,I558389,I339690,I558374,I339707,I339724,I558401,I339741,I339772,I339789,I339806,I558398,I339823,I558380,I339840,I558377,I339857,I558404,I339874,I339905,I339936,I339953,I339970,I340015,I558392,I340046,I340091,I558386,I340108,I340125,I340142,I340159,I340190,I340207,I340285,I340302,I340319,I340336,I340353,I340370,I340387,I340418,I340435,I340452,I340469,I340486,I340503,I340520,I340551,I340582,I340599,I340616,I340661,I340692,I340737,I340754,I340771,I340788,I340805,I340836,I340853,I340931,I340948,I340965,I340982,I340999,I341016,I341033,I340902,I341064,I341081,I341098,I341115,I341132,I341149,I341166,I340899,I341197,I340893,I341228,I341245,I341262,I340923,I340896,I341307,I340920,I341338,I340917,I340914,I341383,I341400,I341417,I341434,I341451,I340908,I341482,I341499,I340911,I340905,I341577,I341594,I341611,I341628,I341645,I341662,I341679,I341548,I341710,I341727,I341744,I341761,I341778,I341795,I341812,I341545,I341843,I341539,I341874,I341891,I341908,I341569,I341542,I341953,I341566,I341984,I341563,I341560,I342029,I342046,I342063,I342080,I342097,I341554,I342128,I342145,I341557,I341551,I342223,I342240,I620615,I342257,I620612,I620597,I342274,I620606,I342291,I342308,I620621,I342325,I342356,I342373,I342390,I620594,I342407,I620600,I342424,I620624,I342441,I620618,I342458,I342489,I342520,I342537,I342554,I342599,I620603,I342630,I342675,I620609,I342692,I342709,I342726,I342743,I342774,I342791,I342869,I342886,I342903,I342920,I342937,I342954,I342971,I342840,I343002,I343019,I343036,I343053,I343070,I343087,I343104,I342837,I343135,I342831,I343166,I343183,I343200,I342861,I342834,I343245,I342858,I343276,I342855,I342852,I343321,I343338,I343355,I343372,I343389,I342846,I343420,I343437,I342849,I342843,I343515,I343532,I582192,I343549,I582180,I582189,I343566,I582204,I343583,I343600,I582186,I343617,I343486,I343648,I343665,I343682,I582174,I343699,I582195,I343716,I582177,I343733,I582183,I343750,I343483,I343781,I343477,I343812,I343829,I343846,I343507,I343480,I343891,I582201,I343504,I343922,I343501,I343498,I343967,I582198,I343984,I344001,I344018,I344035,I343492,I344066,I344083,I343495,I343489,I344161,I344178,I344195,I344212,I344229,I344246,I344263,I344132,I344294,I344311,I344328,I344345,I344362,I344379,I344396,I344129,I344427,I344123,I344458,I344475,I344492,I344153,I344126,I344537,I344150,I344568,I344147,I344144,I344613,I344630,I344647,I344664,I344681,I344138,I344712,I344729,I344141,I344135,I344807,I344824,I531608,I344841,I531620,I531614,I344858,I531599,I344875,I344892,I531626,I344909,I344940,I344957,I344974,I531623,I344991,I531605,I345008,I531602,I345025,I531629,I345042,I345073,I345104,I345121,I345138,I345183,I531617,I345214,I345259,I531611,I345276,I345293,I345310,I345327,I345358,I345375,I345453,I345470,I345487,I345504,I345521,I345538,I345555,I345586,I345603,I345620,I345637,I345654,I345671,I345688,I345719,I345750,I345767,I345784,I345829,I345860,I345905,I345922,I345939,I345956,I345973,I346004,I346021,I346099,I346116,I346133,I346150,I346167,I346184,I346201,I346070,I346232,I346249,I346266,I346283,I346300,I346317,I346334,I346067,I346365,I346061,I346396,I346413,I346430,I346091,I346064,I346475,I346088,I346506,I346085,I346082,I346551,I346568,I346585,I346602,I346619,I346076,I346650,I346667,I346079,I346073,I346745,I346762,I556598,I346779,I556610,I556604,I346796,I556589,I346813,I346830,I556616,I346847,I346878,I346895,I346912,I556613,I346929,I556595,I346946,I556592,I346963,I556619,I346980,I347011,I347042,I347059,I347076,I347121,I556607,I347152,I347197,I556601,I347214,I347231,I347248,I347265,I347296,I347313,I347391,I347408,I347425,I347442,I347459,I347476,I347493,I347524,I347541,I347558,I347575,I347592,I347609,I347626,I347657,I347688,I347705,I347722,I347767,I347798,I347843,I347860,I347877,I347894,I347911,I347942,I347959,I348037,I348054,I348071,I348088,I348105,I348122,I348139,I348170,I348187,I348204,I348221,I348238,I348255,I348272,I348303,I348334,I348351,I348368,I348413,I348444,I348489,I348506,I348523,I348540,I348557,I348588,I348605,I348683,I348700,I348717,I348734,I348751,I348768,I348785,I348816,I348833,I348850,I348867,I348884,I348901,I348918,I348949,I348980,I348997,I349014,I349059,I349090,I349135,I349152,I349169,I349186,I349203,I349234,I349251,I349329,I349346,I349363,I349380,I349397,I349414,I349431,I349300,I349462,I349479,I349496,I349513,I349530,I349547,I349564,I349297,I349595,I349291,I349626,I349643,I349660,I349321,I349294,I349705,I349318,I349736,I349315,I349312,I349781,I349798,I349815,I349832,I349849,I349306,I349880,I349897,I349309,I349303,I349975,I349992,I423599,I350009,I423608,I423593,I350026,I423581,I350043,I350060,I423584,I350077,I349946,I350108,I350125,I350142,I423596,I350159,I423590,I350176,I423587,I350193,I423602,I350210,I349943,I350241,I349937,I350272,I350289,I350306,I349967,I349940,I350351,I423611,I349964,I350382,I349961,I349958,I350427,I423605,I350444,I350461,I350478,I350495,I349952,I350526,I350543,I349955,I349949,I350621,I350638,I719858,I350655,I719843,I719849,I350672,I719846,I350689,I350706,I719855,I350723,I350754,I350771,I350788,I719870,I350805,I719864,I350822,I719861,I350839,I719840,I350856,I350887,I350918,I350935,I350952,I350997,I719867,I351028,I351073,I719852,I351090,I351107,I351124,I351141,I351172,I351189,I351267,I351284,I351301,I351318,I351335,I351352,I351369,I351400,I351417,I351434,I351451,I351468,I351485,I351502,I351533,I351564,I351581,I351598,I351643,I351674,I351719,I351736,I351753,I351770,I351787,I351818,I351835,I351913,I351930,I704830,I351947,I704815,I704821,I351964,I704818,I351981,I351998,I704827,I352015,I351884,I352046,I352063,I352080,I704842,I352097,I704836,I352114,I704833,I352131,I704812,I352148,I351881,I352179,I351875,I352210,I352227,I352244,I351905,I351878,I352289,I704839,I351902,I352320,I351899,I351896,I352365,I704824,I352382,I352399,I352416,I352433,I351890,I352464,I352481,I351893,I351887,I352559,I352576,I471434,I352593,I471437,I471419,I352610,I471446,I352627,I352644,I471425,I352661,I352692,I352709,I352726,I471431,I352743,I471443,I352760,I471449,I352777,I471428,I352794,I352825,I352856,I352873,I352890,I352935,I471440,I352966,I353011,I471422,I353028,I353045,I353062,I353079,I353110,I353127,I353205,I353222,I353239,I353256,I353273,I353290,I353307,I353338,I353355,I353372,I353389,I353406,I353423,I353440,I353471,I353502,I353519,I353536,I353581,I353612,I353657,I353674,I353691,I353708,I353725,I353756,I353773,I353851,I353868,I353885,I353902,I353919,I353936,I353953,I353984,I354001,I354018,I354035,I354052,I354069,I354086,I354117,I354148,I354165,I354182,I354227,I354258,I354303,I354320,I354337,I354354,I354371,I354402,I354419,I354497,I354514,I354531,I354548,I354565,I354582,I354599,I354630,I354647,I354664,I354681,I354698,I354715,I354732,I354763,I354794,I354811,I354828,I354873,I354904,I354949,I354966,I354983,I355000,I355017,I355048,I355065,I355143,I355160,I355177,I355194,I355211,I355228,I355245,I355114,I355276,I355293,I355310,I355327,I355344,I355361,I355378,I355111,I355409,I355105,I355440,I355457,I355474,I355135,I355108,I355519,I355132,I355550,I355129,I355126,I355595,I355612,I355629,I355646,I355663,I355120,I355694,I355711,I355123,I355117,I355789,I355806,I355823,I355840,I355857,I355874,I355891,I355922,I355939,I355956,I355973,I355990,I356007,I356024,I356055,I356086,I356103,I356120,I356165,I356196,I356241,I356258,I356275,I356292,I356309,I356340,I356357,I356435,I356452,I356469,I356486,I356503,I356520,I356537,I356406,I356568,I356585,I356602,I356619,I356636,I356653,I356670,I356403,I356701,I356397,I356732,I356749,I356766,I356427,I356400,I356811,I356424,I356842,I356421,I356418,I356887,I356904,I356921,I356938,I356955,I356412,I356986,I357003,I356415,I356409,I357081,I357098,I557788,I357115,I557800,I557794,I357132,I557779,I357149,I357166,I557806,I357183,I357214,I357231,I357248,I557803,I357265,I557785,I357282,I557782,I357299,I557809,I357316,I357347,I357378,I357395,I357412,I357457,I557797,I357488,I357533,I557791,I357550,I357567,I357584,I357601,I357632,I357649,I357727,I357744,I357761,I357778,I357795,I357812,I357829,I357860,I357877,I357894,I357911,I357928,I357945,I357962,I357993,I358024,I358041,I358058,I358103,I358134,I358179,I358196,I358213,I358230,I358247,I358278,I358295,I358373,I358390,I358407,I358424,I358441,I358458,I358475,I358506,I358523,I358540,I358557,I358574,I358591,I358608,I358639,I358670,I358687,I358704,I358749,I358780,I358825,I358842,I358859,I358876,I358893,I358924,I358941,I359019,I359036,I674709,I359053,I674706,I674691,I359070,I674700,I359087,I359104,I674715,I359121,I358990,I359152,I359169,I359186,I674688,I359203,I674694,I359220,I674718,I359237,I674712,I359254,I358987,I359285,I358981,I359316,I359333,I359350,I359011,I358984,I359395,I674697,I359008,I359426,I359005,I359002,I359471,I674703,I359488,I359505,I359522,I359539,I358996,I359570,I359587,I358999,I358993,I359665,I359682,I502547,I359699,I502553,I502538,I359716,I502532,I359733,I359750,I502559,I359767,I359636,I359798,I359815,I359832,I502544,I359849,I502550,I359866,I502556,I359883,I502529,I359900,I359633,I359931,I359627,I359962,I359979,I359996,I359657,I359630,I360041,I502535,I359654,I360072,I359651,I359648,I360117,I502541,I360134,I360151,I360168,I360185,I359642,I360216,I360233,I359645,I359639,I360311,I360328,I360345,I360362,I360379,I360396,I360413,I360444,I360461,I360478,I360495,I360512,I360529,I360546,I360577,I360608,I360625,I360642,I360687,I360718,I360763,I360780,I360797,I360814,I360831,I360862,I360879,I360957,I360974,I456406,I360991,I456409,I456391,I361008,I456418,I361025,I361042,I456397,I361059,I360928,I361090,I361107,I361124,I456403,I361141,I456415,I361158,I456421,I361175,I456400,I361192,I360925,I361223,I360919,I361254,I361271,I361288,I360949,I360922,I361333,I456412,I360946,I361364,I360943,I360940,I361409,I456394,I361426,I361443,I361460,I361477,I360934,I361508,I361525,I360937,I360931,I361603,I361620,I508998,I361637,I509010,I509004,I361654,I508989,I361671,I361688,I509016,I361705,I361736,I361753,I361770,I509013,I361787,I508995,I361804,I508992,I361821,I509019,I361838,I361869,I361900,I361917,I361934,I361979,I509007,I362010,I362055,I509001,I362072,I362089,I362106,I362123,I362154,I362171,I362249,I362266,I362283,I362300,I362317,I362334,I362351,I362382,I362399,I362416,I362433,I362450,I362467,I362484,I362515,I362546,I362563,I362580,I362625,I362656,I362701,I362718,I362735,I362752,I362769,I362800,I362817,I362895,I362912,I362929,I362946,I362963,I362980,I362997,I363028,I363045,I363062,I363079,I363096,I363113,I363130,I363161,I363192,I363209,I363226,I363271,I363302,I363347,I363364,I363381,I363398,I363415,I363446,I363463,I363541,I363558,I363575,I363592,I363609,I363626,I363643,I363512,I363674,I363691,I363708,I363725,I363742,I363759,I363776,I363509,I363807,I363503,I363838,I363855,I363872,I363533,I363506,I363917,I363530,I363948,I363527,I363524,I363993,I364010,I364027,I364044,I364061,I363518,I364092,I364109,I363521,I363515,I364187,I364204,I364221,I364238,I364255,I364272,I364289,I364320,I364337,I364354,I364371,I364388,I364405,I364422,I364453,I364484,I364501,I364518,I364563,I364594,I364639,I364656,I364673,I364690,I364707,I364738,I364755,I364833,I364850,I599447,I364867,I599435,I599444,I364884,I599459,I364901,I364918,I599441,I364935,I364804,I364966,I364983,I365000,I599429,I365017,I599450,I365034,I599432,I365051,I599438,I365068,I364801,I365099,I364795,I365130,I365147,I365164,I364825,I364798,I365209,I599456,I364822,I365240,I364819,I364816,I365285,I599453,I365302,I365319,I365336,I365353,I364810,I365384,I365401,I364813,I364807,I365479,I365496,I365513,I365530,I365547,I365564,I365581,I365612,I365629,I365646,I365663,I365680,I365697,I365714,I365745,I365776,I365793,I365810,I365855,I365886,I365931,I365948,I365965,I365982,I365999,I366030,I366047,I366125,I366142,I416867,I366159,I416876,I416861,I366176,I416849,I366193,I366210,I416852,I366227,I366258,I366275,I366292,I416864,I366309,I416858,I366326,I416855,I366343,I416870,I366360,I366391,I366422,I366439,I366456,I366501,I416879,I366532,I366577,I416873,I366594,I366611,I366628,I366645,I366676,I366693,I366771,I366788,I725638,I366805,I725623,I725629,I366822,I725626,I366839,I366856,I725635,I366873,I366742,I366904,I366921,I366938,I725650,I366955,I725644,I366972,I725641,I366989,I725620,I367006,I366739,I367037,I366733,I367068,I367085,I367102,I366763,I366736,I367147,I725647,I366760,I367178,I366757,I366754,I367223,I725632,I367240,I367257,I367274,I367291,I366748,I367322,I367339,I366751,I366745,I367417,I367434,I526253,I367451,I526265,I526259,I367468,I526244,I367485,I367502,I526271,I367519,I367550,I367567,I367584,I526268,I367601,I526250,I367618,I526247,I367635,I526274,I367652,I367683,I367714,I367731,I367748,I367793,I526262,I367824,I367869,I526256,I367886,I367903,I367920,I367937,I367968,I367985,I368063,I368080,I452360,I368097,I452363,I452345,I368114,I452372,I368131,I368148,I452351,I368165,I368196,I368213,I368230,I452357,I368247,I452369,I368264,I452375,I368281,I452354,I368298,I368329,I368360,I368377,I368394,I368439,I452366,I368470,I368515,I452348,I368532,I368549,I368566,I368583,I368614,I368631,I368709,I368726,I676596,I368743,I676593,I676578,I368760,I676587,I368777,I368794,I676602,I368811,I368680,I368842,I368859,I368876,I676575,I368893,I676581,I368910,I676605,I368927,I676599,I368944,I368677,I368975,I368671,I369006,I369023,I369040,I368701,I368674,I369085,I676584,I368698,I369116,I368695,I368692,I369161,I676590,I369178,I369195,I369212,I369229,I368686,I369260,I369277,I368689,I368683,I369355,I369372,I551838,I369389,I551850,I551844,I369406,I551829,I369423,I369440,I551856,I369457,I369326,I369488,I369505,I369522,I551853,I369539,I551835,I369556,I551832,I369573,I551859,I369590,I369323,I369621,I369317,I369652,I369669,I369686,I369347,I369320,I369731,I551847,I369344,I369762,I369341,I369338,I369807,I551841,I369824,I369841,I369858,I369875,I369332,I369906,I369923,I369335,I369329,I370001,I370018,I370035,I370052,I370069,I370086,I370103,I369972,I370134,I370151,I370168,I370185,I370202,I370219,I370236,I369969,I370267,I369963,I370298,I370315,I370332,I369993,I369966,I370377,I369990,I370408,I369987,I369984,I370453,I370470,I370487,I370504,I370521,I369978,I370552,I370569,I369981,I369975,I370647,I370664,I370681,I370698,I370715,I370732,I370749,I370618,I370780,I370797,I370814,I370831,I370848,I370865,I370882,I370615,I370913,I370609,I370944,I370961,I370978,I370639,I370612,I371023,I370636,I371054,I370633,I370630,I371099,I371116,I371133,I371150,I371167,I370624,I371198,I371215,I370627,I370621,I371293,I371310,I669048,I371327,I669045,I669030,I371344,I669039,I371361,I371378,I669054,I371395,I371426,I371443,I371460,I669027,I371477,I669033,I371494,I669057,I371511,I669051,I371528,I371559,I371590,I371607,I371624,I371669,I669036,I371700,I371745,I669042,I371762,I371779,I371796,I371813,I371844,I371861,I371939,I371956,I619357,I371973,I619354,I619339,I371990,I619348,I372007,I372024,I619363,I372041,I371910,I372072,I372089,I372106,I619336,I372123,I619342,I372140,I619366,I372157,I619360,I372174,I371907,I372205,I371901,I372236,I372253,I372270,I371931,I371904,I372315,I619345,I371928,I372346,I371925,I371922,I372391,I619351,I372408,I372425,I372442,I372459,I371916,I372490,I372507,I371919,I371913,I372585,I372602,I372619,I372636,I372653,I372670,I372687,I372556,I372718,I372735,I372752,I372769,I372786,I372803,I372820,I372553,I372851,I372547,I372882,I372899,I372916,I372577,I372550,I372961,I372574,I372992,I372571,I372568,I373037,I373054,I373071,I373088,I373105,I372562,I373136,I373153,I372565,I372559,I373231,I373248,I588142,I373265,I588130,I588139,I373282,I588154,I373299,I373316,I588136,I373333,I373364,I373381,I373398,I588124,I373415,I588145,I373432,I588127,I373449,I588133,I373466,I373497,I373528,I373545,I373562,I373607,I588151,I373638,I373683,I588148,I373700,I373717,I373734,I373751,I373782,I373799,I373877,I373894,I578027,I373911,I578015,I578024,I373928,I578039,I373945,I373962,I578021,I373979,I374010,I374027,I374044,I578009,I374061,I578030,I374078,I578012,I374095,I578018,I374112,I374143,I374174,I374191,I374208,I374253,I578036,I374284,I374329,I578033,I374346,I374363,I374380,I374397,I374428,I374445,I374523,I374540,I374557,I374574,I374591,I374608,I374625,I374656,I374673,I374690,I374707,I374724,I374741,I374758,I374789,I374820,I374837,I374854,I374899,I374930,I374975,I374992,I375009,I375026,I375043,I375074,I375091,I375169,I375186,I375203,I375220,I375237,I375254,I375271,I375302,I375319,I375336,I375353,I375370,I375387,I375404,I375435,I375466,I375483,I375500,I375545,I375576,I375621,I375638,I375655,I375672,I375689,I375720,I375737,I375815,I375832,I375849,I375866,I375883,I375900,I375917,I375948,I375965,I375982,I375999,I376016,I376033,I376050,I376081,I376112,I376129,I376146,I376191,I376222,I376267,I376284,I376301,I376318,I376335,I376366,I376383,I376461,I376478,I376495,I376512,I376529,I376546,I376563,I376432,I376594,I376611,I376628,I376645,I376662,I376679,I376696,I376429,I376727,I376423,I376758,I376775,I376792,I376453,I376426,I376837,I376450,I376868,I376447,I376444,I376913,I376930,I376947,I376964,I376981,I376438,I377012,I377029,I376441,I376435,I377107,I377124,I697894,I377141,I697879,I697885,I377158,I697882,I377175,I377192,I697891,I377209,I377240,I377257,I377274,I697906,I377291,I697900,I377308,I697897,I377325,I697876,I377342,I377373,I377404,I377421,I377438,I377483,I697903,I377514,I377559,I697888,I377576,I377593,I377610,I377627,I377658,I377675,I377753,I377770,I377787,I377804,I377821,I377838,I377855,I377886,I377903,I377920,I377937,I377954,I377971,I377988,I378019,I378050,I378067,I378084,I378129,I378160,I378205,I378222,I378239,I378256,I378273,I378304,I378321,I378399,I378416,I441378,I378433,I441381,I441363,I378450,I441390,I378467,I378484,I441369,I378501,I378532,I378549,I378566,I441375,I378583,I441387,I378600,I441393,I378617,I441372,I378634,I378665,I378696,I378713,I378730,I378775,I441384,I378806,I378851,I441366,I378868,I378885,I378902,I378919,I378950,I378967,I379045,I379062,I379079,I379096,I379113,I379130,I379147,I379178,I379195,I379212,I379229,I379246,I379263,I379280,I379311,I379342,I379359,I379376,I379421,I379452,I379497,I379514,I379531,I379548,I379565,I379596,I379613,I379691,I379708,I653952,I379725,I653949,I653934,I379742,I653943,I379759,I379776,I653958,I379793,I379662,I379824,I379841,I379858,I653931,I379875,I653937,I379892,I653961,I379909,I653955,I379926,I379659,I379957,I379653,I379988,I380005,I380022,I379683,I379656,I380067,I653940,I379680,I380098,I379677,I379674,I380143,I653946,I380160,I380177,I380194,I380211,I379668,I380242,I380259,I379671,I379665,I380337,I380354,I380371,I380388,I380405,I380422,I380439,I380308,I380470,I380487,I380504,I380521,I380538,I380555,I380572,I380305,I380603,I380299,I380634,I380651,I380668,I380329,I380302,I380713,I380326,I380744,I380323,I380320,I380789,I380806,I380823,I380840,I380857,I380314,I380888,I380905,I380317,I380311,I380983,I381000,I381017,I381034,I381051,I381068,I381085,I381116,I381133,I381150,I381167,I381184,I381201,I381218,I381249,I381280,I381297,I381314,I381359,I381390,I381435,I381452,I381469,I381486,I381503,I381534,I381551,I381629,I381646,I414419,I381663,I414428,I414413,I381680,I414401,I381697,I381714,I414404,I381731,I381600,I381762,I381779,I381796,I414416,I381813,I414410,I381830,I414407,I381847,I414422,I381864,I381597,I381895,I381591,I381926,I381943,I381960,I381621,I381594,I382005,I414431,I381618,I382036,I381615,I381612,I382081,I414425,I382098,I382115,I382132,I382149,I381606,I382180,I382197,I381609,I381603,I382275,I382292,I382309,I382326,I382343,I382360,I382377,I382408,I382425,I382442,I382459,I382476,I382493,I382510,I382541,I382572,I382589,I382606,I382651,I382682,I382727,I382744,I382761,I382778,I382795,I382826,I382843,I382921,I382938,I382955,I382972,I382989,I383006,I383023,I382892,I383054,I383071,I383088,I383105,I383122,I383139,I383156,I382889,I383187,I382883,I383218,I383235,I383252,I382913,I382886,I383297,I382910,I383328,I382907,I382904,I383373,I383390,I383407,I383424,I383441,I382898,I383472,I383489,I382901,I382895,I383567,I383584,I623131,I383601,I623128,I623113,I383618,I623122,I383635,I383652,I623137,I383669,I383538,I383700,I383717,I383734,I623110,I383751,I623116,I383768,I623140,I383785,I623134,I383802,I383535,I383833,I383529,I383864,I383881,I383898,I383559,I383532,I383943,I623119,I383556,I383974,I383553,I383550,I384019,I623125,I384036,I384053,I384070,I384087,I383544,I384118,I384135,I383547,I383541,I384213,I384230,I384247,I384264,I384281,I384298,I384315,I384346,I384363,I384380,I384397,I384414,I384431,I384448,I384479,I384510,I384527,I384544,I384589,I384620,I384665,I384682,I384699,I384716,I384733,I384764,I384781,I384859,I384876,I597662,I384893,I597650,I597659,I384910,I597674,I384927,I384944,I597656,I384961,I384992,I385009,I385026,I597644,I385043,I597665,I385060,I597647,I385077,I597653,I385094,I385125,I385156,I385173,I385190,I385235,I597671,I385266,I385311,I597668,I385328,I385345,I385362,I385379,I385410,I385427,I385505,I385522,I385539,I385556,I385573,I385590,I385607,I385638,I385655,I385672,I385689,I385706,I385723,I385740,I385771,I385802,I385819,I385836,I385881,I385912,I385957,I385974,I385991,I386008,I386025,I386056,I386073,I386151,I386168,I690958,I386185,I690943,I690949,I386202,I690946,I386219,I386236,I690955,I386253,I386284,I386301,I386318,I690970,I386335,I690964,I386352,I690961,I386369,I690940,I386386,I386417,I386448,I386465,I386482,I386527,I690967,I386558,I386603,I690952,I386620,I386637,I386654,I386671,I386702,I386719,I386797,I386814,I386831,I386848,I386865,I386882,I386899,I386930,I386947,I386964,I386981,I386998,I387015,I387032,I387063,I387094,I387111,I387128,I387173,I387204,I387249,I387266,I387283,I387300,I387317,I387348,I387365,I387443,I387460,I547673,I387477,I547685,I547679,I387494,I547664,I387511,I387528,I547691,I387545,I387414,I387576,I387593,I387610,I547688,I387627,I547670,I387644,I547667,I387661,I547694,I387678,I387411,I387709,I387405,I387740,I387757,I387774,I387435,I387408,I387819,I547682,I387432,I387850,I387429,I387426,I387895,I547676,I387912,I387929,I387946,I387963,I387420,I387994,I388011,I387423,I387417,I388089,I388106,I701940,I388123,I701925,I701931,I388140,I701928,I388157,I388174,I701937,I388191,I388222,I388239,I388256,I701952,I388273,I701946,I388290,I701943,I388307,I701922,I388324,I388355,I388386,I388403,I388420,I388465,I701949,I388496,I388541,I701934,I388558,I388575,I388592,I388609,I388640,I388657,I388735,I388752,I523278,I388769,I523290,I523284,I388786,I523269,I388803,I388820,I523296,I388837,I388868,I388885,I388902,I523293,I388919,I523275,I388936,I523272,I388953,I523299,I388970,I389001,I389032,I389049,I389066,I389111,I523287,I389142,I389187,I523281,I389204,I389221,I389238,I389255,I389286,I389303,I389381,I389398,I389415,I389432,I389449,I389466,I389483,I389352,I389514,I389531,I389548,I389565,I389582,I389599,I389616,I389349,I389647,I389343,I389678,I389695,I389712,I389373,I389346,I389757,I389370,I389788,I389367,I389364,I389833,I389850,I389867,I389884,I389901,I389358,I389932,I389949,I389361,I389355,I390027,I390044,I390061,I390078,I390095,I390112,I390129,I389998,I390160,I390177,I390194,I390211,I390228,I390245,I390262,I389995,I390293,I389989,I390324,I390341,I390358,I390019,I389992,I390403,I390016,I390434,I390013,I390010,I390479,I390496,I390513,I390530,I390547,I390004,I390578,I390595,I390007,I390001,I390673,I390690,I472590,I390707,I472593,I472575,I390724,I472602,I390741,I390758,I472581,I390775,I390806,I390823,I390840,I472587,I390857,I472599,I390874,I472605,I390891,I472584,I390908,I390939,I390970,I390987,I391004,I391049,I472596,I391080,I391125,I472578,I391142,I391159,I391176,I391193,I391224,I391241,I391319,I391336,I391353,I391370,I391387,I391404,I391421,I391452,I391469,I391486,I391503,I391520,I391537,I391554,I391585,I391616,I391633,I391650,I391695,I391726,I391771,I391788,I391805,I391822,I391839,I391870,I391887,I391965,I391982,I391999,I392016,I392033,I392050,I392067,I391936,I392098,I392115,I392132,I392149,I392166,I392183,I392200,I391933,I392231,I391927,I392262,I392279,I392296,I391957,I391930,I392341,I391954,I392372,I391951,I391948,I392417,I392434,I392451,I392468,I392485,I391942,I392516,I392533,I391945,I391939,I392611,I392628,I463920,I392645,I463923,I463905,I392662,I463932,I392679,I392696,I463911,I392713,I392582,I392744,I392761,I392778,I463917,I392795,I463929,I392812,I463935,I392829,I463914,I392846,I392579,I392877,I392573,I392908,I392925,I392942,I392603,I392576,I392987,I463926,I392600,I393018,I392597,I392594,I393063,I463908,I393080,I393097,I393114,I393131,I392588,I393162,I393179,I392591,I392585,I393257,I393274,I393291,I393308,I393325,I393342,I393359,I393228,I393390,I393407,I393424,I393441,I393458,I393475,I393492,I393225,I393523,I393219,I393554,I393571,I393588,I393249,I393222,I393633,I393246,I393664,I393243,I393240,I393709,I393726,I393743,I393760,I393777,I393234,I393808,I393825,I393237,I393231,I393903,I393920,I393937,I393954,I393971,I393988,I394005,I393874,I394036,I394053,I394070,I394087,I394104,I394121,I394138,I393871,I394169,I393865,I394200,I394217,I394234,I393895,I393868,I394279,I393892,I394310,I393889,I393886,I394355,I394372,I394389,I394406,I394423,I393880,I394454,I394471,I393883,I393877,I394549,I394566,I394583,I394600,I394617,I394634,I394651,I394682,I394699,I394716,I394733,I394750,I394767,I394784,I394815,I394846,I394863,I394880,I394925,I394956,I395001,I395018,I395035,I395052,I395069,I395100,I395117,I395195,I395212,I395229,I395246,I395263,I395280,I395297,I395166,I395328,I395345,I395362,I395379,I395396,I395413,I395430,I395163,I395461,I395157,I395492,I395509,I395526,I395187,I395160,I395571,I395184,I395602,I395181,I395178,I395647,I395664,I395681,I395698,I395715,I395172,I395746,I395763,I395175,I395169,I395841,I395858,I548863,I395875,I548875,I548869,I395892,I548854,I395909,I395926,I548881,I395943,I395812,I395974,I395991,I396008,I548878,I396025,I548860,I396042,I548857,I396059,I548884,I396076,I395809,I396107,I395803,I396138,I396155,I396172,I395833,I395806,I396217,I548872,I395830,I396248,I395827,I395824,I396293,I548866,I396310,I396327,I396344,I396361,I395818,I396392,I396409,I395821,I395815,I396487,I396504,I396521,I396538,I396555,I396572,I396589,I396458,I396620,I396637,I396654,I396671,I396688,I396705,I396722,I396455,I396753,I396449,I396784,I396801,I396818,I396479,I396452,I396863,I396476,I396894,I396473,I396470,I396939,I396956,I396973,I396990,I397007,I396464,I397038,I397055,I396467,I396461,I397133,I397150,I397167,I397184,I397201,I397218,I397235,I397104,I397266,I397283,I397300,I397317,I397334,I397351,I397368,I397101,I397399,I397095,I397430,I397447,I397464,I397125,I397098,I397509,I397122,I397540,I397119,I397116,I397585,I397602,I397619,I397636,I397653,I397110,I397684,I397701,I397113,I397107,I397779,I397796,I616841,I397813,I616838,I616823,I397830,I616832,I397847,I397864,I616847,I397881,I397912,I397929,I397946,I616820,I397963,I616826,I397980,I616850,I397997,I616844,I398014,I398045,I398076,I398093,I398110,I398155,I616829,I398186,I398231,I616835,I398248,I398265,I398282,I398299,I398330,I398347,I398425,I398442,I687918,I398459,I687915,I687900,I398476,I687909,I398493,I398510,I687924,I398527,I398558,I398575,I398592,I687897,I398609,I687903,I398626,I687927,I398643,I687921,I398660,I398691,I398722,I398739,I398756,I398801,I687906,I398832,I398877,I687912,I398894,I398911,I398928,I398945,I398976,I398993,I399071,I399088,I399105,I399122,I399139,I399156,I399173,I399204,I399221,I399238,I399255,I399272,I399289,I399306,I399337,I399368,I399385,I399402,I399447,I399478,I399523,I399540,I399557,I399574,I399591,I399622,I399639,I399717,I399734,I399751,I399768,I399785,I399802,I399819,I399850,I399867,I399884,I399901,I399918,I399935,I399952,I399983,I400014,I400031,I400048,I400093,I400124,I400169,I400186,I400203,I400220,I400237,I400268,I400285,I400363,I400380,I400397,I400414,I400431,I400448,I400465,I400496,I400513,I400530,I400547,I400564,I400581,I400598,I400629,I400660,I400677,I400694,I400739,I400770,I400815,I400832,I400849,I400866,I400883,I400914,I400931,I401009,I401026,I569093,I401043,I569105,I569099,I401060,I569084,I401077,I401094,I569111,I401111,I401142,I401159,I401176,I569108,I401193,I569090,I401210,I569087,I401227,I569114,I401244,I401275,I401306,I401323,I401340,I401385,I569102,I401416,I401461,I569096,I401478,I401495,I401512,I401529,I401560,I401577,I401655,I401672,I401689,I401706,I401723,I401740,I401757,I401626,I401788,I401805,I401822,I401839,I401856,I401873,I401890,I401623,I401921,I401617,I401952,I401969,I401986,I401647,I401620,I402031,I401644,I402062,I401641,I401638,I402107,I402124,I402141,I402158,I402175,I401632,I402206,I402223,I401635,I401629,I402301,I402318,I483572,I402335,I483575,I483557,I402352,I483584,I402369,I402386,I483563,I402403,I402434,I402451,I402468,I483569,I402485,I483581,I402502,I483587,I402519,I483566,I402536,I402567,I402598,I402615,I402632,I402677,I483578,I402708,I402753,I483560,I402770,I402787,I402804,I402821,I402852,I402869,I402947,I402964,I402981,I402998,I403015,I403032,I403049,I402918,I403080,I403097,I403114,I403131,I403148,I403165,I403182,I402915,I403213,I402909,I403244,I403261,I403278,I402939,I402912,I403323,I402936,I403354,I402933,I402930,I403399,I403416,I403433,I403450,I403467,I402924,I403498,I403515,I402927,I402921,I403593,I403610,I403627,I403644,I403661,I403678,I403695,I403726,I403743,I403760,I403777,I403794,I403811,I403828,I403859,I403890,I403907,I403924,I403969,I404000,I404045,I404062,I404079,I404096,I404113,I404144,I404161,I404239,I404256,I627534,I404273,I627531,I627516,I404290,I627525,I404307,I404324,I627540,I404341,I404210,I404372,I404389,I404406,I627513,I404423,I627519,I404440,I627543,I404457,I627537,I404474,I404207,I404505,I404201,I404536,I404553,I404570,I404231,I404204,I404615,I627522,I404228,I404646,I404225,I404222,I404691,I627528,I404708,I404725,I404742,I404759,I404216,I404790,I404807,I404219,I404213,I404885,I404902,I639485,I404919,I639482,I639467,I404936,I639476,I404953,I404970,I639491,I404987,I405018,I405035,I405052,I639464,I405069,I639470,I405086,I639494,I405103,I639488,I405120,I405151,I405182,I405199,I405216,I405261,I639473,I405292,I405337,I639479,I405354,I405371,I405388,I405405,I405436,I405453,I405531,I405548,I611347,I405565,I611335,I611344,I405582,I611359,I405599,I405616,I611341,I405633,I405502,I405664,I405681,I405698,I611329,I405715,I611350,I405732,I611332,I405749,I611338,I405766,I405499,I405797,I405493,I405828,I405845,I405862,I405523,I405496,I405907,I611356,I405520,I405938,I405517,I405514,I405983,I611353,I406000,I406017,I406034,I406051,I405508,I406082,I406099,I405511,I405505,I406177,I406194,I406211,I406228,I406245,I406262,I406279,I406148,I406310,I406327,I406344,I406361,I406378,I406395,I406412,I406145,I406443,I406139,I406474,I406491,I406508,I406169,I406142,I406553,I406166,I406584,I406163,I406160,I406629,I406646,I406663,I406680,I406697,I406154,I406728,I406745,I406157,I406151,I406823,I406840,I715812,I406857,I715797,I715803,I406874,I715800,I406891,I406908,I715809,I406925,I406956,I406973,I406990,I715824,I407007,I715818,I407024,I715815,I407041,I715794,I407058,I407089,I407120,I407137,I407154,I407199,I715821,I407230,I407275,I715806,I407292,I407309,I407326,I407343,I407374,I407391,I407469,I407486,I407503,I407520,I407537,I407554,I407571,I407440,I407602,I407619,I407636,I407653,I407670,I407687,I407704,I407437,I407735,I407431,I407766,I407783,I407800,I407461,I407434,I407845,I407458,I407876,I407455,I407452,I407921,I407938,I407955,I407972,I407989,I407446,I408020,I408037,I407449,I407443,I408115,I408132,I408149,I408166,I408183,I408200,I408217,I408086,I408248,I408265,I408282,I408299,I408316,I408333,I408350,I408083,I408381,I408077,I408412,I408429,I408446,I408107,I408080,I408491,I408104,I408522,I408101,I408098,I408567,I408584,I408601,I408618,I408635,I408092,I408666,I408683,I408095,I408089,I408761,I408778,I408795,I408812,I408829,I408846,I408863,I408894,I408911,I408928,I408945,I408962,I408979,I408996,I409027,I409058,I409075,I409092,I409137,I409168,I409213,I409230,I409247,I409264,I409281,I409312,I409329,I409407,I409424,I605992,I409441,I605980,I605989,I409458,I606004,I409475,I409492,I605986,I409509,I409540,I409557,I409574,I605974,I409591,I605995,I409608,I605977,I409625,I605983,I409642,I409673,I409704,I409721,I409738,I409783,I606001,I409814,I409859,I605998,I409876,I409893,I409910,I409927,I409958,I409975,I410053,I410070,I597067,I410087,I597055,I597064,I410104,I597079,I410121,I410138,I597061,I410155,I410186,I410203,I410220,I597049,I410237,I597070,I410254,I597052,I410271,I597058,I410288,I410319,I410350,I410367,I410384,I410429,I597076,I410460,I410505,I597073,I410522,I410539,I410556,I410573,I410604,I410621,I410699,I410716,I682886,I410733,I682883,I682868,I410750,I682877,I410767,I410784,I682892,I410801,I410670,I410832,I410849,I410866,I682865,I410883,I682871,I410900,I682895,I410917,I682889,I410934,I410667,I410965,I410661,I410996,I411013,I411030,I410691,I410664,I411075,I682874,I410688,I411106,I410685,I410682,I411151,I682880,I411168,I411185,I411202,I411219,I410676,I411250,I411267,I410679,I410673,I411345,I411362,I411379,I411396,I411413,I411430,I411447,I411316,I411478,I411495,I411512,I411529,I411546,I411563,I411580,I411313,I411611,I411307,I411642,I411659,I411676,I411337,I411310,I411721,I411334,I411752,I411331,I411328,I411797,I411814,I411831,I411848,I411865,I411322,I411896,I411913,I411325,I411319,I411991,I412008,I412025,I412042,I412059,I411953,I412090,I412107,I412124,I412141,I412158,I412175,I411962,I412206,I411956,I412237,I412254,I412271,I412288,I411983,I411980,I412333,I412350,I412367,I411977,I412398,I411974,I411965,I412443,I412460,I412477,I411968,I411971,I412522,I412539,I411959,I412603,I412620,I721598,I721583,I412637,I721580,I412654,I721574,I721586,I412671,I412702,I412719,I721601,I412736,I412753,I721589,I721592,I412770,I412787,I412818,I412849,I721577,I412866,I721595,I412883,I412900,I412945,I412962,I412979,I413010,I413055,I721604,I413072,I413089,I413134,I413151,I413215,I413232,I413249,I413266,I413283,I413177,I413314,I413331,I413348,I413365,I413382,I413399,I413186,I413430,I413180,I413461,I413478,I413495,I413512,I413207,I413204,I413557,I413574,I413591,I413201,I413622,I413198,I413189,I413667,I413684,I413701,I413192,I413195,I413746,I413763,I413183,I413827,I413844,I413861,I413878,I413895,I413789,I413926,I413943,I413960,I413977,I413994,I414011,I413798,I414042,I413792,I414073,I414090,I414107,I414124,I413819,I413816,I414169,I414186,I414203,I413813,I414234,I413810,I413801,I414279,I414296,I414313,I413804,I413807,I414358,I414375,I413795,I414439,I414456,I469107,I469122,I414473,I469137,I414490,I469119,I469110,I414507,I414538,I414555,I469128,I414572,I414589,I469134,I469125,I414606,I414623,I414654,I414685,I469113,I414702,I469116,I414719,I414736,I414781,I414798,I414815,I414846,I414891,I469131,I414908,I414925,I414970,I414987,I415051,I415068,I573258,I573270,I415085,I573273,I415102,I573255,I573249,I415119,I415150,I415167,I573261,I415184,I415201,I573264,I573267,I415218,I415235,I415266,I415297,I573279,I415314,I573252,I415331,I415348,I415393,I415410,I415427,I415458,I415503,I573276,I415520,I415537,I415582,I415599,I415663,I415680,I415697,I415714,I415731,I415762,I415779,I415796,I415813,I415830,I415847,I415878,I415909,I415926,I415943,I415960,I416005,I416022,I416039,I416070,I416115,I416132,I416149,I416194,I416211,I416275,I416292,I488888,I488876,I416309,I488891,I416326,I488873,I488867,I416343,I416237,I416374,I416391,I488885,I416408,I416425,I488879,I488861,I416442,I416459,I416246,I416490,I416240,I416521,I488882,I416538,I488870,I416555,I416572,I416267,I416264,I416617,I416634,I416651,I416261,I416682,I416258,I416249,I416727,I488864,I416744,I416761,I416252,I416255,I416806,I416823,I416243,I416887,I416904,I416921,I416938,I416955,I416986,I417003,I417020,I417037,I417054,I417071,I417102,I417133,I417150,I417167,I417184,I417229,I417246,I417263,I417294,I417339,I417356,I417373,I417418,I417435,I417499,I417516,I417533,I417550,I417567,I417598,I417615,I417632,I417649,I417666,I417683,I417714,I417745,I417762,I417779,I417796,I417841,I417858,I417875,I417906,I417951,I417968,I417985,I418030,I418047,I418111,I418128,I418145,I418162,I418179,I418210,I418227,I418244,I418261,I418278,I418295,I418326,I418357,I418374,I418391,I418408,I418453,I418470,I418487,I418518,I418563,I418580,I418597,I418642,I418659,I418723,I418740,I725066,I725051,I418757,I725048,I418774,I725042,I725054,I418791,I418685,I418822,I418839,I725069,I418856,I418873,I725057,I725060,I418890,I418907,I418694,I418938,I418688,I418969,I725045,I418986,I725063,I419003,I419020,I418715,I418712,I419065,I419082,I419099,I418709,I419130,I418706,I418697,I419175,I725072,I419192,I419209,I418700,I418703,I419254,I419271,I418691,I419335,I419352,I447721,I447736,I419369,I447751,I419386,I447733,I447724,I419403,I419434,I419451,I447742,I419468,I419485,I447748,I447739,I419502,I419519,I419550,I419581,I447727,I419598,I447730,I419615,I419632,I419677,I419694,I419711,I419742,I419787,I447745,I419804,I419821,I419866,I419883,I419947,I419964,I419981,I419998,I420015,I420046,I420063,I420080,I420097,I420114,I420131,I420162,I420193,I420210,I420227,I420244,I420289,I420306,I420323,I420354,I420399,I420416,I420433,I420478,I420495,I420559,I420576,I474309,I474324,I420593,I474339,I420610,I474321,I474312,I420627,I420658,I420675,I474330,I420692,I420709,I474336,I474327,I420726,I420743,I420774,I420805,I474315,I420822,I474318,I420839,I420856,I420901,I420918,I420935,I420966,I421011,I474333,I421028,I421045,I421090,I421107,I421171,I421188,I421205,I421222,I421239,I421133,I421270,I421287,I421304,I421321,I421338,I421355,I421142,I421386,I421136,I421417,I421434,I421451,I421468,I421163,I421160,I421513,I421530,I421547,I421157,I421578,I421154,I421145,I421623,I421640,I421657,I421148,I421151,I421702,I421719,I421139,I421783,I421800,I473153,I473168,I421817,I473183,I421834,I473165,I473156,I421851,I421745,I421882,I421899,I473174,I421916,I421933,I473180,I473171,I421950,I421967,I421754,I421998,I421748,I422029,I473159,I422046,I473162,I422063,I422080,I421775,I421772,I422125,I422142,I422159,I421769,I422190,I421766,I421757,I422235,I473177,I422252,I422269,I421760,I421763,I422314,I422331,I421751,I422395,I422412,I422429,I422446,I422463,I422357,I422494,I422511,I422528,I422545,I422562,I422579,I422366,I422610,I422360,I422641,I422658,I422675,I422692,I422387,I422384,I422737,I422754,I422771,I422381,I422802,I422378,I422369,I422847,I422864,I422881,I422372,I422375,I422926,I422943,I422363,I423007,I423024,I705992,I705977,I423041,I705974,I423058,I705968,I705980,I423075,I423106,I423123,I705995,I423140,I423157,I705983,I705986,I423174,I423191,I423222,I423253,I705971,I423270,I705989,I423287,I423304,I423349,I423366,I423383,I423414,I423459,I705998,I423476,I423493,I423538,I423555,I423619,I423636,I490724,I490712,I423653,I490727,I423670,I490709,I490703,I423687,I423718,I423735,I490721,I423752,I423769,I490715,I490697,I423786,I423803,I423834,I423865,I490718,I423882,I490706,I423899,I423916,I423961,I423978,I423995,I424026,I424071,I490700,I424088,I424105,I424150,I424167,I424231,I424248,I424265,I424282,I424299,I424330,I424347,I424364,I424381,I424398,I424415,I424446,I424477,I424494,I424511,I424528,I424573,I424590,I424607,I424638,I424683,I424700,I424717,I424762,I424779,I424843,I424860,I648920,I648923,I424877,I648929,I424894,I648926,I648902,I424911,I424942,I424959,I648905,I424976,I424993,I648914,I648899,I425010,I425027,I425058,I425089,I648917,I425106,I648911,I425123,I425140,I425185,I425202,I425219,I425250,I425295,I648908,I425312,I425329,I425374,I425391,I425455,I425472,I490112,I490100,I425489,I490115,I425506,I490097,I490091,I425523,I425554,I425571,I490109,I425588,I425605,I490103,I490085,I425622,I425639,I425670,I425701,I490106,I425718,I490094,I425735,I425752,I425797,I425814,I425831,I425862,I425907,I490088,I425924,I425941,I425986,I426003,I426067,I426084,I480089,I480104,I426101,I480119,I426118,I480101,I480092,I426135,I426029,I426166,I426183,I480110,I426200,I426217,I480116,I480107,I426234,I426251,I426038,I426282,I426032,I426313,I480095,I426330,I480098,I426347,I426364,I426059,I426056,I426409,I426426,I426443,I426053,I426474,I426050,I426041,I426519,I480113,I426536,I426553,I426044,I426047,I426598,I426615,I426035,I426679,I426696,I426713,I426730,I426747,I426778,I426795,I426812,I426829,I426846,I426863,I426894,I426925,I426942,I426959,I426976,I427021,I427038,I427055,I427086,I427131,I427148,I427165,I427210,I427227,I427291,I427308,I610740,I610761,I427325,I610746,I427342,I610749,I610737,I427359,I427390,I427407,I610755,I427424,I427441,I610743,I610758,I427458,I427475,I427506,I427537,I610734,I427554,I610764,I427571,I427588,I427633,I427650,I427667,I427698,I427743,I610752,I427760,I427777,I427822,I427839,I427903,I427920,I427937,I427954,I427971,I428002,I428019,I428036,I428053,I428070,I428087,I428118,I428149,I428166,I428183,I428200,I428245,I428262,I428279,I428310,I428355,I428372,I428389,I428434,I428451,I428515,I428532,I428549,I428566,I428583,I428477,I428614,I428631,I428648,I428665,I428682,I428699,I428486,I428730,I428480,I428761,I428778,I428795,I428812,I428507,I428504,I428857,I428874,I428891,I428501,I428922,I428498,I428489,I428967,I428984,I429001,I428492,I428495,I429046,I429063,I428483,I429127,I429144,I708304,I708289,I429161,I708286,I429178,I708280,I708292,I429195,I429226,I429243,I708307,I429260,I429277,I708295,I708298,I429294,I429311,I429342,I429373,I708283,I429390,I708301,I429407,I429424,I429469,I429486,I429503,I429534,I429579,I708310,I429596,I429613,I429658,I429675,I429739,I429756,I705414,I705399,I429773,I705396,I429790,I705390,I705402,I429807,I429701,I429838,I429855,I705417,I429872,I429889,I705405,I705408,I429906,I429923,I429710,I429954,I429704,I429985,I705393,I430002,I705411,I430019,I430036,I429731,I429728,I430081,I430098,I430115,I429725,I430146,I429722,I429713,I430191,I705420,I430208,I430225,I429716,I429719,I430270,I430287,I429707,I430351,I430368,I595865,I595886,I430385,I595871,I430402,I595874,I595862,I430419,I430313,I430450,I430467,I595880,I430484,I430501,I595868,I595883,I430518,I430535,I430322,I430566,I430316,I430597,I595859,I430614,I595889,I430631,I430648,I430343,I430340,I430693,I430710,I430727,I430337,I430758,I430334,I430325,I430803,I595877,I430820,I430837,I430328,I430331,I430882,I430899,I430319,I430963,I430980,I430997,I431014,I431031,I430925,I431062,I431079,I431096,I431113,I431130,I431147,I430934,I431178,I430928,I431209,I431226,I431243,I431260,I430955,I430952,I431305,I431322,I431339,I430949,I431370,I430946,I430937,I431415,I431432,I431449,I430940,I430943,I431494,I431511,I430931,I431575,I431592,I726213,I726225,I431609,I726198,I431626,I431643,I431543,I431674,I726216,I431691,I726207,I431708,I431546,I431739,I431540,I431770,I726204,I726210,I431787,I726222,I431804,I431821,I431838,I431549,I431869,I726228,I431886,I726219,I431903,I431920,I431555,I431558,I431537,I431979,I726201,I431996,I432013,I431567,I431564,I432058,I432075,I431552,I431561,I432153,I432170,I432187,I432204,I432221,I432252,I432269,I432286,I432317,I432348,I432365,I432382,I432399,I432416,I432447,I432464,I432481,I432498,I432557,I432574,I432591,I432636,I432653,I432731,I432748,I432765,I432782,I432799,I432830,I432847,I432864,I432895,I432926,I432943,I432960,I432977,I432994,I433025,I433042,I433059,I433076,I433135,I433152,I433169,I433214,I433231,I433309,I433326,I433343,I433360,I433377,I433408,I433425,I433442,I433473,I433504,I433521,I433538,I433555,I433572,I433603,I433620,I433637,I433654,I433713,I433730,I433747,I433792,I433809,I433887,I433904,I433921,I433938,I433955,I433855,I433986,I434003,I434020,I433858,I434051,I433852,I434082,I434099,I434116,I434133,I434150,I433861,I434181,I434198,I434215,I434232,I433867,I433870,I433849,I434291,I434308,I434325,I433879,I433876,I434370,I434387,I433864,I433873,I434465,I434482,I643256,I643259,I434499,I643265,I434516,I434533,I434564,I643262,I434581,I643241,I434598,I434629,I434660,I643238,I643253,I434677,I643250,I434694,I434711,I434728,I434759,I643268,I434776,I643247,I434793,I434810,I434869,I643244,I434886,I434903,I434948,I434965,I435043,I435060,I600628,I600625,I435077,I600619,I435094,I435111,I435142,I600640,I435159,I600643,I435176,I435207,I435238,I600646,I600637,I435255,I600649,I435272,I435289,I435306,I435337,I600622,I435354,I600631,I435371,I435388,I435447,I600634,I435464,I435481,I435526,I435543,I435621,I435638,I542931,I542919,I435655,I542913,I435672,I435689,I435720,I542910,I435737,I542904,I435754,I435785,I435816,I542907,I542922,I435833,I542934,I435850,I435867,I435884,I435915,I542925,I435932,I542916,I435949,I435966,I436025,I542928,I436042,I436059,I436104,I436121,I436199,I436216,I436233,I436250,I436267,I436298,I436315,I436332,I436363,I436394,I436411,I436428,I436445,I436462,I436493,I436510,I436527,I436544,I436603,I436620,I436637,I436682,I436699,I436777,I436794,I436811,I436828,I436845,I436745,I436876,I436893,I436910,I436748,I436941,I436742,I436972,I436989,I437006,I437023,I437040,I436751,I437071,I437088,I437105,I437122,I436757,I436760,I436739,I437181,I437198,I437215,I436769,I436766,I437260,I437277,I436754,I436763,I437355,I437372,I437389,I437406,I437423,I437323,I437454,I437471,I437488,I437326,I437519,I437320,I437550,I437567,I437584,I437601,I437618,I437329,I437649,I437666,I437683,I437700,I437335,I437338,I437317,I437759,I437776,I437793,I437347,I437344,I437838,I437855,I437332,I437341,I437933,I437950,I541146,I541134,I437967,I541128,I437984,I438001,I437901,I438032,I541125,I438049,I541119,I438066,I437904,I438097,I437898,I438128,I541122,I541137,I438145,I541149,I438162,I438179,I438196,I437907,I438227,I541140,I438244,I541131,I438261,I438278,I437913,I437916,I437895,I438337,I541143,I438354,I438371,I437925,I437922,I438416,I438433,I437910,I437919,I438511,I438528,I660239,I660242,I438545,I660248,I438562,I438579,I438610,I660245,I438627,I660224,I438644,I438675,I438706,I660221,I660236,I438723,I660233,I438740,I438757,I438774,I438805,I660251,I438822,I660230,I438839,I438856,I438915,I660227,I438932,I438949,I438994,I439011,I439089,I439106,I439123,I439140,I439157,I439188,I439205,I439222,I439253,I439284,I439301,I439318,I439335,I439352,I439383,I439400,I439417,I439434,I439493,I439510,I439527,I439572,I439589,I439667,I439684,I535791,I535779,I439701,I535773,I439718,I439735,I439766,I535770,I439783,I535764,I439800,I439831,I439862,I535767,I535782,I439879,I535794,I439896,I439913,I439930,I439961,I535785,I439978,I535776,I439995,I440012,I440071,I535788,I440088,I440105,I440150,I440167,I440245,I440262,I595273,I595270,I440279,I595264,I440296,I440313,I440213,I440344,I595285,I440361,I595288,I440378,I440216,I440409,I440210,I440440,I595291,I595282,I440457,I595294,I440474,I440491,I440508,I440219,I440539,I595267,I440556,I595276,I440573,I440590,I440225,I440228,I440207,I440649,I595279,I440666,I440683,I440237,I440234,I440728,I440745,I440222,I440231,I440823,I440840,I681625,I681628,I440857,I681634,I440874,I440891,I440922,I681631,I440939,I681610,I440956,I440987,I441018,I681607,I681622,I441035,I681619,I441052,I441069,I441086,I441117,I681637,I441134,I681616,I441151,I441168,I441227,I681613,I441244,I441261,I441306,I441323,I441401,I441418,I441435,I441452,I441469,I441500,I441517,I441534,I441565,I441596,I441613,I441630,I441647,I441664,I441695,I441712,I441729,I441746,I441805,I441822,I441839,I441884,I441901,I441979,I441996,I442013,I442030,I442047,I441947,I442078,I442095,I442112,I441950,I442143,I441944,I442174,I442191,I442208,I442225,I442242,I441953,I442273,I442290,I442307,I442324,I441959,I441962,I441941,I442383,I442400,I442417,I441971,I441968,I442462,I442479,I441956,I441965,I442557,I442574,I442591,I442608,I442625,I442525,I442656,I442673,I442690,I442528,I442721,I442522,I442752,I442769,I442786,I442803,I442820,I442531,I442851,I442868,I442885,I442902,I442537,I442540,I442519,I442961,I442978,I442995,I442549,I442546,I443040,I443057,I442534,I442543,I443135,I443152,I630676,I630679,I443169,I630685,I443186,I443203,I443234,I630682,I443251,I630661,I443268,I443299,I443330,I630658,I630673,I443347,I630670,I443364,I443381,I443398,I443429,I630688,I443446,I630667,I443463,I443480,I443539,I630664,I443556,I443573,I443618,I443635,I443713,I443730,I443747,I443764,I443781,I443681,I443812,I443829,I443846,I443684,I443877,I443678,I443908,I443925,I443942,I443959,I443976,I443687,I444007,I444024,I444041,I444058,I443693,I443696,I443675,I444117,I444134,I444151,I443705,I443702,I444196,I444213,I443690,I443699,I444291,I444308,I563161,I563149,I444325,I563143,I444342,I444359,I444390,I563140,I444407,I563134,I444424,I444455,I444486,I563137,I563152,I444503,I563164,I444520,I444537,I444554,I444585,I563155,I444602,I563146,I444619,I444636,I444695,I563158,I444712,I444729,I444774,I444791,I444869,I444886,I444903,I444920,I444937,I444837,I444968,I444985,I445002,I444840,I445033,I444834,I445064,I445081,I445098,I445115,I445132,I444843,I445163,I445180,I445197,I445214,I444849,I444852,I444831,I445273,I445290,I445307,I444861,I444858,I445352,I445369,I444846,I444855,I445447,I445464,I445481,I445498,I445515,I445415,I445546,I445563,I445580,I445418,I445611,I445412,I445642,I445659,I445676,I445693,I445710,I445421,I445741,I445758,I445775,I445792,I445427,I445430,I445409,I445851,I445868,I445885,I445439,I445436,I445930,I445947,I445424,I445433,I446025,I446042,I617467,I617470,I446059,I617476,I446076,I446093,I445993,I446124,I617473,I446141,I617452,I446158,I445996,I446189,I445990,I446220,I617449,I617464,I446237,I617461,I446254,I446271,I446288,I445999,I446319,I617479,I446336,I617458,I446353,I446370,I446005,I446008,I445987,I446429,I617455,I446446,I446463,I446017,I446014,I446508,I446525,I446002,I446011,I446603,I446620,I446637,I446654,I446671,I446571,I446702,I446719,I446736,I446574,I446767,I446568,I446798,I446815,I446832,I446849,I446866,I446577,I446897,I446914,I446931,I446948,I446583,I446586,I446565,I447007,I447024,I447041,I446595,I446592,I447086,I447103,I446580,I446589,I447181,I447198,I530436,I530424,I447215,I530418,I447232,I447249,I447280,I530415,I447297,I530409,I447314,I447345,I447376,I530412,I530427,I447393,I530439,I447410,I447427,I447444,I447475,I530430,I447492,I530421,I447509,I447526,I447585,I530433,I447602,I447619,I447664,I447681,I447759,I447776,I585158,I585155,I447793,I585149,I447810,I447827,I447858,I585170,I447875,I585173,I447892,I447923,I447954,I585176,I585167,I447971,I585179,I447988,I448005,I448022,I448053,I585152,I448070,I585161,I448087,I448104,I448163,I585164,I448180,I448197,I448242,I448259,I448337,I448354,I521511,I521499,I448371,I521493,I448388,I448405,I448436,I521490,I448453,I521484,I448470,I448501,I448532,I521487,I521502,I448549,I521514,I448566,I448583,I448600,I448631,I521505,I448648,I521496,I448665,I448682,I448741,I521508,I448758,I448775,I448820,I448837,I448915,I448932,I448949,I448966,I448983,I449014,I449031,I449048,I449079,I449110,I449127,I449144,I449161,I449178,I449209,I449226,I449243,I449260,I449319,I449336,I449353,I449398,I449415,I449493,I449510,I449527,I449544,I449561,I449461,I449592,I449609,I449626,I449464,I449657,I449458,I449688,I449705,I449722,I449739,I449756,I449467,I449787,I449804,I449821,I449838,I449473,I449476,I449455,I449897,I449914,I449931,I449485,I449482,I449976,I449993,I449470,I449479,I450071,I450088,I450105,I450122,I450139,I450039,I450170,I450187,I450204,I450042,I450235,I450036,I450266,I450283,I450300,I450317,I450334,I450045,I450365,I450382,I450399,I450416,I450051,I450054,I450033,I450475,I450492,I450509,I450063,I450060,I450554,I450571,I450048,I450057,I450649,I450666,I496171,I496198,I450683,I496186,I450700,I450717,I450617,I450748,I496177,I450765,I496174,I450782,I450620,I450813,I450614,I450844,I496192,I496195,I450861,I496183,I450878,I450895,I450912,I450623,I450943,I496180,I450960,I496201,I450977,I450994,I450629,I450632,I450611,I451053,I496189,I451070,I451087,I450641,I450638,I451132,I451149,I450626,I450635,I451227,I451244,I661497,I661500,I451261,I661506,I451278,I451295,I451195,I451326,I661503,I451343,I661482,I451360,I451198,I451391,I451192,I451422,I661479,I661494,I451439,I661491,I451456,I451473,I451490,I451201,I451521,I661509,I451538,I661488,I451555,I451572,I451207,I451210,I451189,I451631,I661485,I451648,I451665,I451219,I451216,I451710,I451727,I451204,I451213,I451805,I451822,I451839,I451856,I451873,I451904,I451921,I451938,I451969,I452000,I452017,I452034,I452051,I452068,I452099,I452116,I452133,I452150,I452209,I452226,I452243,I452288,I452305,I452383,I452400,I452417,I452434,I452451,I452482,I452499,I452516,I452547,I452578,I452595,I452612,I452629,I452646,I452677,I452694,I452711,I452728,I452787,I452804,I452821,I452866,I452883,I452961,I452978,I452995,I453012,I453029,I453060,I453077,I453094,I453125,I453156,I453173,I453190,I453207,I453224,I453255,I453272,I453289,I453306,I453365,I453382,I453399,I453444,I453461,I453539,I453556,I453573,I453590,I453607,I453507,I453638,I453655,I453672,I453510,I453703,I453504,I453734,I453751,I453768,I453785,I453802,I453513,I453833,I453850,I453867,I453884,I453519,I453522,I453501,I453943,I453960,I453977,I453531,I453528,I454022,I454039,I453516,I453525,I454117,I454134,I628160,I628163,I454151,I628169,I454168,I454185,I454216,I628166,I454233,I628145,I454250,I454281,I454312,I628142,I628157,I454329,I628154,I454346,I454363,I454380,I454411,I628172,I454428,I628151,I454445,I454462,I454521,I628148,I454538,I454555,I454600,I454617,I454695,I454712,I611933,I611930,I454729,I611924,I454746,I454763,I454794,I611945,I454811,I611948,I454828,I454859,I454890,I611951,I611942,I454907,I611954,I454924,I454941,I454958,I454989,I611927,I455006,I611936,I455023,I455040,I455099,I611939,I455116,I455133,I455178,I455195,I455273,I455290,I580993,I580990,I455307,I580984,I455324,I455341,I455241,I455372,I581005,I455389,I581008,I455406,I455244,I455437,I455238,I455468,I581011,I581002,I455485,I581014,I455502,I455519,I455536,I455247,I455567,I580987,I455584,I580996,I455601,I455618,I455253,I455256,I455235,I455677,I580999,I455694,I455711,I455265,I455262,I455756,I455773,I455250,I455259,I455851,I455868,I712919,I712931,I455885,I712904,I455902,I455919,I455950,I712922,I455967,I712913,I455984,I456015,I456046,I712910,I712916,I456063,I712928,I456080,I456097,I456114,I456145,I712934,I456162,I712925,I456179,I456196,I456255,I712907,I456272,I456289,I456334,I456351,I456429,I456446,I534601,I534589,I456463,I534583,I456480,I456497,I456528,I534580,I456545,I534574,I456562,I456593,I456624,I534577,I534592,I456641,I534604,I456658,I456675,I456692,I456723,I534595,I456740,I534586,I456757,I456774,I456833,I534598,I456850,I456867,I456912,I456929,I457007,I457024,I511396,I511384,I457041,I511378,I457058,I457075,I457106,I511375,I457123,I511369,I457140,I457171,I457202,I511372,I511387,I457219,I511399,I457236,I457253,I457270,I457301,I511390,I457318,I511381,I457335,I457352,I457411,I511393,I457428,I457445,I457490,I457507,I457585,I457602,I684770,I684773,I457619,I684779,I457636,I457653,I457684,I684776,I457701,I684755,I457718,I457749,I457780,I684752,I684767,I457797,I684764,I457814,I457831,I457848,I457879,I684782,I457896,I684761,I457913,I457930,I457989,I684758,I458006,I458023,I458068,I458085,I458163,I458180,I679738,I679741,I458197,I679747,I458214,I458231,I458131,I458262,I679744,I458279,I679723,I458296,I458134,I458327,I458128,I458358,I679720,I679735,I458375,I679732,I458392,I458409,I458426,I458137,I458457,I679750,I458474,I679729,I458491,I458508,I458143,I458146,I458125,I458567,I679726,I458584,I458601,I458155,I458152,I458646,I458663,I458140,I458149,I458741,I458758,I458775,I458792,I458809,I458709,I458840,I458857,I458874,I458712,I458905,I458706,I458936,I458953,I458970,I458987,I459004,I458715,I459035,I459052,I459069,I459086,I458721,I458724,I458703,I459145,I459162,I459179,I458733,I458730,I459224,I459241,I458718,I458727,I459319,I459336,I459353,I459370,I459387,I459418,I459435,I459452,I459483,I459514,I459531,I459548,I459565,I459582,I459613,I459630,I459647,I459664,I459723,I459740,I459757,I459802,I459819,I459897,I459914,I459931,I459948,I459965,I459996,I460013,I460030,I460061,I460092,I460109,I460126,I460143,I460160,I460191,I460208,I460225,I460242,I460301,I460318,I460335,I460380,I460397,I460475,I460492,I460509,I460526,I460543,I460574,I460591,I460608,I460639,I460670,I460687,I460704,I460721,I460738,I460769,I460786,I460803,I460820,I460879,I460896,I460913,I460958,I460975,I461053,I461070,I461087,I461104,I461121,I461152,I461169,I461186,I461217,I461248,I461265,I461282,I461299,I461316,I461347,I461364,I461381,I461398,I461457,I461474,I461491,I461536,I461553,I461631,I461648,I544716,I544704,I461665,I544698,I461682,I461699,I461599,I461730,I544695,I461747,I544689,I461764,I461602,I461795,I461596,I461826,I544692,I544707,I461843,I544719,I461860,I461877,I461894,I461605,I461925,I544710,I461942,I544701,I461959,I461976,I461611,I461614,I461593,I462035,I544713,I462052,I462069,I461623,I461620,I462114,I462131,I461608,I461617,I462209,I462226,I462243,I462260,I462277,I462308,I462325,I462342,I462373,I462404,I462421,I462438,I462455,I462472,I462503,I462520,I462537,I462554,I462613,I462630,I462647,I462692,I462709,I462787,I462804,I462821,I462838,I462855,I462755,I462886,I462903,I462920,I462758,I462951,I462752,I462982,I462999,I463016,I463033,I463050,I462761,I463081,I463098,I463115,I463132,I462767,I462770,I462749,I463191,I463208,I463225,I462779,I462776,I463270,I463287,I462764,I462773,I463365,I463382,I463399,I463416,I463433,I463464,I463481,I463498,I463529,I463560,I463577,I463594,I463611,I463628,I463659,I463676,I463693,I463710,I463769,I463786,I463803,I463848,I463865,I463943,I463960,I463977,I463994,I464011,I464042,I464059,I464076,I464107,I464138,I464155,I464172,I464189,I464206,I464237,I464254,I464271,I464288,I464347,I464364,I464381,I464426,I464443,I464521,I464538,I464555,I464572,I464589,I464620,I464637,I464654,I464685,I464716,I464733,I464750,I464767,I464784,I464815,I464832,I464849,I464866,I464925,I464942,I464959,I465004,I465021,I465099,I465116,I626902,I626905,I465133,I626911,I465150,I465167,I465067,I465198,I626908,I465215,I626887,I465232,I465070,I465263,I465064,I465294,I626884,I626899,I465311,I626896,I465328,I465345,I465362,I465073,I465393,I626914,I465410,I626893,I465427,I465444,I465079,I465082,I465061,I465503,I626890,I465520,I465537,I465091,I465088,I465582,I465599,I465076,I465085,I465677,I465694,I465711,I465728,I465745,I465776,I465793,I465810,I465841,I465872,I465889,I465906,I465923,I465940,I465971,I465988,I466005,I466022,I466081,I466098,I466115,I466160,I466177,I466255,I466272,I466289,I466306,I466323,I466354,I466371,I466388,I466419,I466450,I466467,I466484,I466501,I466518,I466549,I466566,I466583,I466600,I466659,I466676,I466693,I466738,I466755,I466833,I466850,I534006,I533994,I466867,I533988,I466884,I466901,I466801,I466932,I533985,I466949,I533979,I466966,I466804,I466997,I466798,I467028,I533982,I533997,I467045,I534009,I467062,I467079,I467096,I466807,I467127,I534000,I467144,I533991,I467161,I467178,I466813,I466816,I466795,I467237,I534003,I467254,I467271,I466825,I466822,I467316,I467333,I466810,I466819,I467411,I467428,I467445,I467462,I467479,I467510,I467527,I467544,I467575,I467606,I467623,I467640,I467657,I467674,I467705,I467722,I467739,I467756,I467815,I467832,I467849,I467894,I467911,I467989,I468006,I492539,I492563,I468023,I492545,I468040,I468057,I468088,I492533,I468105,I492548,I468122,I468153,I468184,I492554,I492536,I468201,I492557,I468218,I468235,I468252,I468283,I492542,I468300,I492551,I468317,I468334,I468393,I492560,I468410,I468427,I468472,I468489,I468567,I468584,I468601,I468618,I468635,I468666,I468683,I468700,I468731,I468762,I468779,I468796,I468813,I468830,I468861,I468878,I468895,I468912,I468971,I468988,I469005,I469050,I469067,I469145,I469162,I469179,I469196,I469213,I469244,I469261,I469278,I469309,I469340,I469357,I469374,I469391,I469408,I469439,I469456,I469473,I469490,I469549,I469566,I469583,I469628,I469645,I469723,I469740,I469757,I469774,I469791,I469822,I469839,I469856,I469887,I469918,I469935,I469952,I469969,I469986,I470017,I470034,I470051,I470068,I470127,I470144,I470161,I470206,I470223,I470301,I470318,I470335,I470352,I470369,I470400,I470417,I470434,I470465,I470496,I470513,I470530,I470547,I470564,I470595,I470612,I470629,I470646,I470705,I470722,I470739,I470784,I470801,I470879,I470896,I568516,I568504,I470913,I568498,I470930,I470947,I470847,I470978,I568495,I470995,I568489,I471012,I470850,I471043,I470844,I471074,I568492,I568507,I471091,I568519,I471108,I471125,I471142,I470853,I471173,I568510,I471190,I568501,I471207,I471224,I470859,I470862,I470841,I471283,I568513,I471300,I471317,I470871,I470868,I471362,I471379,I470856,I470865,I471457,I471474,I471491,I471508,I471525,I471556,I471573,I471590,I471621,I471652,I471669,I471686,I471703,I471720,I471751,I471768,I471785,I471802,I471861,I471878,I471895,I471940,I471957,I472035,I472052,I472069,I472086,I472103,I472003,I472134,I472151,I472168,I472006,I472199,I472000,I472230,I472247,I472264,I472281,I472298,I472009,I472329,I472346,I472363,I472380,I472015,I472018,I471997,I472439,I472456,I472473,I472027,I472024,I472518,I472535,I472012,I472021,I472613,I472630,I677222,I677225,I472647,I677231,I472664,I472681,I472712,I677228,I472729,I677207,I472746,I472777,I472808,I677204,I677219,I472825,I677216,I472842,I472859,I472876,I472907,I677234,I472924,I677213,I472941,I472958,I473017,I677210,I473034,I473051,I473096,I473113,I473191,I473208,I473225,I473242,I473259,I473290,I473307,I473324,I473355,I473386,I473403,I473420,I473437,I473454,I473485,I473502,I473519,I473536,I473595,I473612,I473629,I473674,I473691,I473769,I473786,I551261,I551249,I473803,I551243,I473820,I473837,I473868,I551240,I473885,I551234,I473902,I473933,I473964,I551237,I551252,I473981,I551264,I473998,I474015,I474032,I474063,I551255,I474080,I551246,I474097,I474114,I474173,I551258,I474190,I474207,I474252,I474269,I474347,I474364,I474381,I474398,I474415,I474446,I474463,I474480,I474511,I474542,I474559,I474576,I474593,I474610,I474641,I474658,I474675,I474692,I474751,I474768,I474785,I474830,I474847,I474925,I474942,I678480,I678483,I474959,I678489,I474976,I474993,I474893,I475024,I678486,I475041,I678465,I475058,I474896,I475089,I474890,I475120,I678462,I678477,I475137,I678474,I475154,I475171,I475188,I474899,I475219,I678492,I475236,I678471,I475253,I475270,I474905,I474908,I474887,I475329,I678468,I475346,I475363,I474917,I474914,I475408,I475425,I474902,I474911,I475503,I475520,I606578,I606575,I475537,I606569,I475554,I475571,I475602,I606590,I475619,I606593,I475636,I475667,I475698,I606596,I606587,I475715,I606599,I475732,I475749,I475766,I475797,I606572,I475814,I606581,I475831,I475848,I475907,I606584,I475924,I475941,I475986,I476003,I476081,I476098,I618725,I618728,I476115,I618734,I476132,I476149,I476049,I476180,I618731,I476197,I618710,I476214,I476052,I476245,I476046,I476276,I618707,I618722,I476293,I618719,I476310,I476327,I476344,I476055,I476375,I618737,I476392,I618716,I476409,I476426,I476061,I476064,I476043,I476485,I618713,I476502,I476519,I476073,I476070,I476564,I476581,I476058,I476067,I476659,I476676,I476693,I476710,I476727,I476758,I476775,I476792,I476823,I476854,I476871,I476888,I476905,I476922,I476953,I476970,I476987,I477004,I477063,I477080,I477097,I477142,I477159,I477237,I477254,I477271,I477288,I477305,I477336,I477353,I477370,I477401,I477432,I477449,I477466,I477483,I477500,I477531,I477548,I477565,I477582,I477641,I477658,I477675,I477720,I477737,I477815,I477832,I538766,I538754,I477849,I538748,I477866,I477883,I477914,I538745,I477931,I538739,I477948,I477979,I478010,I538742,I538757,I478027,I538769,I478044,I478061,I478078,I478109,I538760,I478126,I538751,I478143,I478160,I478219,I538763,I478236,I478253,I478298,I478315,I478393,I478410,I628789,I628792,I478427,I628798,I478444,I478461,I478492,I628795,I478509,I628774,I478526,I478557,I478588,I628771,I628786,I478605,I628783,I478622,I478639,I478656,I478687,I628801,I478704,I628780,I478721,I478738,I478797,I628777,I478814,I478831,I478876,I478893,I478971,I478988,I479005,I479022,I479039,I479070,I479087,I479104,I479135,I479166,I479183,I479200,I479217,I479234,I479265,I479282,I479299,I479316,I479375,I479392,I479409,I479454,I479471,I479549,I479566,I479583,I479600,I479617,I479648,I479665,I479682,I479713,I479744,I479761,I479778,I479795,I479812,I479843,I479860,I479877,I479894,I479953,I479970,I479987,I480032,I480049,I480127,I480144,I480161,I480178,I480195,I480226,I480243,I480260,I480291,I480322,I480339,I480356,I480373,I480390,I480421,I480438,I480455,I480472,I480531,I480548,I480565,I480610,I480627,I480705,I480722,I658352,I658355,I480739,I658361,I480756,I480773,I480673,I480804,I658358,I480821,I658337,I480838,I480676,I480869,I480670,I480900,I658334,I658349,I480917,I658346,I480934,I480951,I480968,I480679,I480999,I658364,I481016,I658343,I481033,I481050,I480685,I480688,I480667,I481109,I658340,I481126,I481143,I480697,I480694,I481188,I481205,I480682,I480691,I481283,I481300,I609553,I609550,I481317,I609544,I481334,I481351,I481251,I481382,I609565,I481399,I609568,I481416,I481254,I481447,I481248,I481478,I609571,I609562,I481495,I609574,I481512,I481529,I481546,I481257,I481577,I609547,I481594,I609556,I481611,I481628,I481263,I481266,I481245,I481687,I609559,I481704,I481721,I481275,I481272,I481766,I481783,I481260,I481269,I481861,I481878,I481895,I481912,I481929,I481829,I481960,I481977,I481994,I481832,I482025,I481826,I482056,I482073,I482090,I482107,I482124,I481835,I482155,I482172,I482189,I482206,I481841,I481844,I481823,I482265,I482282,I482299,I481853,I481850,I482344,I482361,I481838,I481847,I482439,I482456,I652062,I652065,I482473,I652071,I482490,I482507,I482538,I652068,I482555,I652047,I482572,I482603,I482634,I652044,I652059,I482651,I652056,I482668,I482685,I482702,I482733,I652074,I482750,I652053,I482767,I482784,I482843,I652050,I482860,I482877,I482922,I482939,I483017,I483034,I513181,I513169,I483051,I513163,I483068,I483085,I483116,I513160,I483133,I513154,I483150,I483181,I483212,I513157,I513172,I483229,I513184,I483246,I483263,I483280,I483311,I513175,I483328,I513166,I483345,I483362,I483421,I513178,I483438,I483455,I483500,I483517,I483595,I483612,I483629,I483646,I483663,I483694,I483711,I483728,I483759,I483790,I483807,I483824,I483841,I483858,I483889,I483906,I483923,I483940,I483999,I484016,I484033,I484078,I484095,I484173,I484190,I484207,I484224,I484241,I484272,I484289,I484306,I484337,I484368,I484385,I484402,I484419,I484436,I484467,I484484,I484501,I484518,I484577,I484594,I484611,I484656,I484673,I484751,I484768,I484785,I484802,I484819,I484850,I484867,I484884,I484915,I484946,I484963,I484980,I484997,I485014,I485045,I485062,I485079,I485096,I485155,I485172,I485189,I485234,I485251,I485329,I485346,I485363,I485380,I485397,I485297,I485428,I485445,I485462,I485300,I485493,I485294,I485524,I485541,I485558,I485575,I485592,I485303,I485623,I485640,I485657,I485674,I485309,I485312,I485291,I485733,I485750,I485767,I485321,I485318,I485812,I485829,I485306,I485315,I485907,I485924,I702515,I702527,I485941,I702500,I485958,I485975,I486006,I702518,I486023,I702509,I486040,I486071,I486102,I702506,I702512,I486119,I702524,I486136,I486153,I486170,I486201,I702530,I486218,I702521,I486235,I486252,I486311,I702503,I486328,I486345,I486390,I486407,I486485,I486502,I486519,I486536,I486553,I486453,I486584,I486601,I486618,I486456,I486649,I486450,I486680,I486697,I486714,I486731,I486748,I486459,I486779,I486796,I486813,I486830,I486465,I486468,I486447,I486889,I486906,I486923,I486477,I486474,I486968,I486985,I486462,I486471,I487063,I487080,I487097,I487114,I487131,I487162,I487179,I487196,I487213,I487230,I487247,I487264,I487281,I487326,I487343,I487374,I487391,I487422,I487439,I487470,I487501,I487532,I487549,I487580,I487611,I487675,I487692,I625653,I625647,I487709,I625656,I487726,I625650,I625632,I487743,I487774,I487791,I487808,I625629,I487825,I487842,I625644,I625626,I487859,I487876,I487893,I487938,I487955,I487986,I488003,I488034,I625638,I488051,I625641,I488082,I488113,I488144,I625635,I488161,I488192,I488223,I488287,I488304,I488321,I488338,I488355,I488386,I488403,I488420,I488437,I488454,I488471,I488488,I488505,I488550,I488567,I488598,I488615,I488646,I488663,I488694,I488725,I488756,I488773,I488804,I488835,I488899,I488916,I488933,I488950,I488967,I488998,I489015,I489032,I489049,I489066,I489083,I489100,I489117,I489162,I489179,I489210,I489227,I489258,I489275,I489306,I489337,I489368,I489385,I489416,I489447,I489511,I489528,I560778,I560784,I489545,I560781,I489562,I560754,I560772,I489579,I489479,I489610,I489627,I489644,I560766,I489661,I489678,I560769,I560757,I489695,I489712,I489729,I489485,I489476,I489774,I489791,I489500,I489822,I489839,I489488,I489870,I560760,I489887,I560775,I489494,I489918,I489482,I489949,I489473,I489980,I560763,I489997,I489503,I490028,I489497,I490059,I489491,I490123,I490140,I490157,I490174,I490191,I490222,I490239,I490256,I490273,I490290,I490307,I490324,I490341,I490386,I490403,I490434,I490451,I490482,I490499,I490530,I490561,I490592,I490609,I490640,I490671,I490735,I490752,I704234,I704249,I490769,I704243,I490786,I704240,I704237,I490803,I490834,I490851,I490868,I704255,I490885,I490902,I704246,I704252,I490919,I490936,I490953,I490998,I491015,I491046,I491063,I491094,I704264,I491111,I704261,I491142,I491173,I491204,I704258,I491221,I491252,I491283,I491347,I491364,I536383,I536389,I491381,I536386,I491398,I536359,I536377,I491415,I491446,I491463,I491480,I536371,I491497,I491514,I536374,I536362,I491531,I491548,I491565,I491610,I491627,I491658,I491675,I491706,I536365,I491723,I536380,I491754,I491785,I491816,I536368,I491833,I491864,I491895,I491959,I491976,I714060,I714075,I491993,I714069,I492010,I714066,I714063,I492027,I492058,I492075,I492092,I714081,I492109,I492126,I714072,I714078,I492143,I492160,I492177,I492222,I492239,I492270,I492287,I492318,I714090,I492335,I714087,I492366,I492397,I492428,I714084,I492445,I492476,I492507,I492571,I492588,I498510,I498489,I492605,I498492,I492622,I498486,I498498,I492639,I492670,I492687,I492704,I498495,I492721,I492738,I498507,I498513,I492755,I492772,I492789,I492834,I492851,I492882,I492899,I492930,I498483,I492947,I498501,I492978,I493009,I493040,I498504,I493057,I493088,I493119,I493183,I493200,I493217,I493234,I493251,I493282,I493299,I493316,I493333,I493350,I493367,I493384,I493401,I493446,I493463,I493494,I493511,I493542,I493559,I493590,I493621,I493652,I493669,I493700,I493731,I493795,I493812,I493829,I493846,I493863,I493763,I493894,I493911,I493928,I493945,I493962,I493979,I493996,I494013,I493769,I493760,I494058,I494075,I493784,I494106,I494123,I493772,I494154,I494171,I493778,I494202,I493766,I494233,I493757,I494264,I494281,I493787,I494312,I493781,I494343,I493775,I494407,I494424,I494441,I494458,I494475,I494375,I494506,I494523,I494540,I494557,I494574,I494591,I494608,I494625,I494381,I494372,I494670,I494687,I494396,I494718,I494735,I494384,I494766,I494783,I494390,I494814,I494378,I494845,I494369,I494876,I494893,I494399,I494924,I494393,I494955,I494387,I495019,I495036,I495053,I495070,I495087,I495118,I495135,I495152,I495169,I495186,I495203,I495220,I495237,I495282,I495299,I495330,I495347,I495378,I495395,I495426,I495457,I495488,I495505,I495536,I495567,I495631,I495648,I495665,I495682,I495620,I495713,I495730,I495747,I495764,I495781,I495798,I495815,I495605,I495846,I495602,I495877,I495614,I495908,I495925,I495942,I495608,I495623,I495987,I496004,I495593,I496035,I495611,I496066,I496083,I495617,I496114,I496131,I495596,I495599,I496209,I496226,I604210,I604207,I496243,I604195,I496260,I604189,I604216,I496291,I496308,I604201,I496325,I496342,I496359,I604192,I604213,I496376,I496393,I496424,I496455,I496486,I604204,I496503,I604198,I496520,I496565,I496582,I496613,I604219,I496644,I496661,I496692,I496709,I496787,I496804,I669659,I669662,I496821,I669680,I496838,I669674,I669683,I496869,I496886,I669686,I496903,I496920,I496937,I669671,I669656,I496954,I496971,I497002,I497033,I497064,I669668,I497081,I669677,I497098,I497143,I497160,I497191,I669665,I497222,I497239,I497270,I497287,I497365,I497382,I497399,I497416,I497447,I497464,I497481,I497498,I497515,I497532,I497549,I497580,I497611,I497642,I497659,I497676,I497721,I497738,I497769,I497800,I497817,I497848,I497865,I497943,I497960,I497977,I497994,I498025,I498042,I498059,I498076,I498093,I498110,I498127,I498158,I498189,I498220,I498237,I498254,I498299,I498316,I498347,I498378,I498395,I498426,I498443,I498521,I498538,I498555,I498572,I498603,I498620,I498637,I498654,I498671,I498688,I498705,I498736,I498767,I498798,I498815,I498832,I498877,I498894,I498925,I498956,I498973,I499004,I499021,I499099,I499116,I549470,I549464,I499133,I549458,I499150,I549479,I549467,I499088,I499181,I499198,I549452,I499215,I499232,I499249,I549455,I549449,I499266,I499283,I499073,I499314,I499070,I499345,I499082,I499376,I549476,I499393,I549473,I499410,I499076,I499091,I499455,I499472,I499061,I499503,I549461,I499079,I499534,I499551,I499085,I499582,I499599,I499064,I499067,I499677,I499694,I499711,I499728,I499759,I499776,I499793,I499810,I499827,I499844,I499861,I499892,I499923,I499954,I499971,I499988,I500033,I500050,I500081,I500112,I500129,I500160,I500177,I500255,I500272,I650160,I650163,I500289,I650181,I500306,I650175,I650184,I500337,I500354,I650187,I500371,I500388,I500405,I650172,I650157,I500422,I500439,I500470,I500501,I500532,I650169,I500549,I650178,I500566,I500611,I500628,I500659,I650166,I500690,I500707,I500738,I500755,I500833,I500850,I500867,I500884,I500822,I500915,I500932,I500949,I500966,I500983,I501000,I501017,I500807,I501048,I500804,I501079,I500816,I501110,I501127,I501144,I500810,I500825,I501189,I501206,I500795,I501237,I500813,I501268,I501285,I500819,I501316,I501333,I500798,I500801,I501411,I501428,I501445,I501462,I501400,I501493,I501510,I501527,I501544,I501561,I501578,I501595,I501385,I501626,I501382,I501657,I501394,I501688,I501705,I501722,I501388,I501403,I501767,I501784,I501373,I501815,I501391,I501846,I501863,I501397,I501894,I501911,I501376,I501379,I501989,I502006,I638209,I638212,I502023,I638230,I502040,I638224,I638233,I502071,I502088,I638236,I502105,I502122,I502139,I638221,I638206,I502156,I502173,I502204,I502235,I502266,I638218,I502283,I638227,I502300,I502345,I502362,I502393,I638215,I502424,I502441,I502472,I502489,I502567,I502584,I502601,I502618,I502649,I502666,I502683,I502700,I502717,I502734,I502751,I502782,I502813,I502844,I502861,I502878,I502923,I502940,I502971,I503002,I503019,I503050,I503067,I503145,I503162,I503179,I503196,I503227,I503244,I503261,I503278,I503295,I503312,I503329,I503360,I503391,I503422,I503439,I503456,I503501,I503518,I503549,I503580,I503597,I503628,I503645,I503723,I503740,I503757,I503774,I503805,I503822,I503839,I503856,I503873,I503890,I503907,I503938,I503969,I504000,I504017,I504034,I504079,I504096,I504127,I504158,I504175,I504206,I504223,I504301,I504318,I504335,I504352,I504383,I504400,I504417,I504434,I504451,I504468,I504485,I504516,I504547,I504578,I504595,I504612,I504657,I504674,I504705,I504736,I504753,I504784,I504801,I504879,I504896,I504913,I504930,I504961,I504978,I504995,I505012,I505029,I505046,I505063,I505094,I505125,I505156,I505173,I505190,I505235,I505252,I505283,I505314,I505331,I505362,I505379,I505457,I505474,I505491,I505508,I505525,I505542,I505573,I505590,I505607,I505652,I505669,I505686,I505731,I505748,I505765,I505796,I505813,I505844,I505861,I505878,I505909,I505926,I505943,I505960,I506052,I506069,I506086,I506103,I506120,I506137,I506035,I506168,I506185,I506202,I506038,I506020,I506247,I506264,I506281,I506041,I506032,I506326,I506343,I506360,I506023,I506391,I506408,I506014,I506439,I506456,I506473,I506044,I506504,I506521,I506538,I506555,I506029,I506026,I506017,I506647,I506664,I506681,I506698,I506715,I506732,I506763,I506780,I506797,I506842,I506859,I506876,I506921,I506938,I506955,I506986,I507003,I507034,I507051,I507068,I507099,I507116,I507133,I507150,I507242,I507259,I507276,I507293,I507310,I507327,I507358,I507375,I507392,I507437,I507454,I507471,I507516,I507533,I507550,I507581,I507598,I507629,I507646,I507663,I507694,I507711,I507728,I507745,I507837,I507854,I507871,I507888,I507905,I507922,I507953,I507970,I507987,I508032,I508049,I508066,I508111,I508128,I508145,I508176,I508193,I508224,I508241,I508258,I508289,I508306,I508323,I508340,I508432,I508449,I508466,I508483,I508500,I508517,I508548,I508565,I508582,I508627,I508644,I508661,I508706,I508723,I508740,I508771,I508788,I508819,I508836,I508853,I508884,I508901,I508918,I508935,I509027,I509044,I614951,I614942,I509061,I614960,I509078,I509095,I614957,I509112,I509143,I614939,I509160,I509177,I509222,I614948,I614963,I509239,I614954,I509256,I509301,I614936,I509318,I614945,I509335,I509366,I509383,I509414,I614933,I509431,I509448,I509479,I509496,I509513,I509530,I509622,I509639,I509656,I509673,I509690,I509707,I509738,I509755,I509772,I509817,I509834,I509851,I509896,I509913,I509930,I509961,I509978,I510009,I510026,I510043,I510074,I510091,I510108,I510125,I510217,I510234,I510251,I510268,I510285,I510302,I510333,I510350,I510367,I510412,I510429,I510446,I510491,I510508,I510525,I510556,I510573,I510604,I510621,I510638,I510669,I510686,I510703,I510720,I510812,I510829,I510846,I510863,I510880,I510897,I510928,I510945,I510962,I511007,I511024,I511041,I511086,I511103,I511120,I511151,I511168,I511199,I511216,I511233,I511264,I511281,I511298,I511315,I511407,I511424,I511441,I511458,I511475,I511492,I511523,I511540,I511557,I511602,I511619,I511636,I511681,I511698,I511715,I511746,I511763,I511794,I511811,I511828,I511859,I511876,I511893,I511910,I512002,I512019,I512036,I512053,I512070,I512087,I511985,I512118,I512135,I512152,I511988,I511970,I512197,I512214,I512231,I511991,I511982,I512276,I512293,I512310,I511973,I512341,I512358,I511964,I512389,I512406,I512423,I511994,I512454,I512471,I512488,I512505,I511979,I511976,I511967,I512597,I512614,I712338,I712344,I512631,I712335,I512648,I512665,I712347,I512682,I512713,I712326,I512730,I512747,I512792,I712350,I712332,I512809,I712341,I512826,I512871,I712356,I512888,I712329,I512905,I512936,I512953,I512984,I712353,I513001,I513018,I513049,I513066,I513083,I513100,I513192,I513209,I513226,I513243,I513260,I513277,I513308,I513325,I513342,I513387,I513404,I513421,I513466,I513483,I513500,I513531,I513548,I513579,I513596,I513613,I513644,I513661,I513678,I513695,I513787,I513804,I513821,I513838,I513855,I513872,I513903,I513920,I513937,I513982,I513999,I514016,I514061,I514078,I514095,I514126,I514143,I514174,I514191,I514208,I514239,I514256,I514273,I514290,I514382,I514399,I514416,I514433,I514450,I514467,I514365,I514498,I514515,I514532,I514368,I514350,I514577,I514594,I514611,I514371,I514362,I514656,I514673,I514690,I514353,I514721,I514738,I514344,I514769,I514786,I514803,I514374,I514834,I514851,I514868,I514885,I514359,I514356,I514347,I514977,I514994,I515011,I515028,I515045,I515062,I515093,I515110,I515127,I515172,I515189,I515206,I515251,I515268,I515285,I515316,I515333,I515364,I515381,I515398,I515429,I515446,I515463,I515480,I515572,I515589,I515606,I515623,I515640,I515657,I515688,I515705,I515722,I515767,I515784,I515801,I515846,I515863,I515880,I515911,I515928,I515959,I515976,I515993,I516024,I516041,I516058,I516075,I516167,I516184,I516201,I516218,I516235,I516252,I516283,I516300,I516317,I516362,I516379,I516396,I516441,I516458,I516475,I516506,I516523,I516554,I516571,I516588,I516619,I516636,I516653,I516670,I516762,I516779,I516796,I516813,I516830,I516847,I516878,I516895,I516912,I516957,I516974,I516991,I517036,I517053,I517070,I517101,I517118,I517149,I517166,I517183,I517214,I517231,I517248,I517265,I517357,I517374,I517391,I517408,I517425,I517442,I517473,I517490,I517507,I517552,I517569,I517586,I517631,I517648,I517665,I517696,I517713,I517744,I517761,I517778,I517809,I517826,I517843,I517860,I517952,I517969,I517986,I518003,I518020,I518037,I517935,I518068,I518085,I518102,I517938,I517920,I518147,I518164,I518181,I517941,I517932,I518226,I518243,I518260,I517923,I518291,I518308,I517914,I518339,I518356,I518373,I517944,I518404,I518421,I518438,I518455,I517929,I517926,I517917,I518547,I518564,I518581,I518598,I518615,I518632,I518663,I518680,I518697,I518742,I518759,I518776,I518821,I518838,I518855,I518886,I518903,I518934,I518951,I518968,I518999,I519016,I519033,I519050,I519142,I519159,I519176,I519193,I519210,I519227,I519258,I519275,I519292,I519337,I519354,I519371,I519416,I519433,I519450,I519481,I519498,I519529,I519546,I519563,I519594,I519611,I519628,I519645,I519737,I519754,I693842,I693848,I519771,I693839,I519788,I519805,I693851,I519822,I519853,I693830,I519870,I519887,I519932,I693854,I693836,I519949,I693845,I519966,I520011,I693860,I520028,I693833,I520045,I520076,I520093,I520124,I693857,I520141,I520158,I520189,I520206,I520223,I520240,I520332,I520349,I520366,I520383,I520400,I520417,I520448,I520465,I520482,I520527,I520544,I520561,I520606,I520623,I520640,I520671,I520688,I520719,I520736,I520753,I520784,I520801,I520818,I520835,I520927,I520944,I520961,I520978,I520995,I521012,I521043,I521060,I521077,I521122,I521139,I521156,I521201,I521218,I521235,I521266,I521283,I521314,I521331,I521348,I521379,I521396,I521413,I521430,I521522,I521539,I672190,I672181,I521556,I672199,I521573,I521590,I672196,I521607,I521638,I672178,I521655,I521672,I521717,I672187,I672202,I521734,I672193,I521751,I521796,I672175,I521813,I672184,I521830,I521861,I521878,I521909,I672172,I521926,I521943,I521974,I521991,I522008,I522025,I522117,I522134,I723320,I723326,I522151,I723317,I522168,I522185,I723329,I522202,I522233,I723308,I522250,I522267,I522312,I723332,I723314,I522329,I723323,I522346,I522391,I723338,I522408,I723311,I522425,I522456,I522473,I522504,I723335,I522521,I522538,I522569,I522586,I522603,I522620,I522712,I522729,I522746,I522763,I522780,I522797,I522695,I522828,I522845,I522862,I522698,I522680,I522907,I522924,I522941,I522701,I522692,I522986,I523003,I523020,I522683,I523051,I523068,I522674,I523099,I523116,I523133,I522704,I523164,I523181,I523198,I523215,I522689,I522686,I522677,I523307,I523324,I720430,I720436,I523341,I720427,I523358,I523375,I720439,I523392,I523423,I720418,I523440,I523457,I523502,I720442,I720424,I523519,I720433,I523536,I523581,I720448,I523598,I720421,I523615,I523646,I523663,I523694,I720445,I523711,I523728,I523759,I523776,I523793,I523810,I523902,I523919,I523936,I523953,I523970,I523987,I524018,I524035,I524052,I524097,I524114,I524131,I524176,I524193,I524210,I524241,I524258,I524289,I524306,I524323,I524354,I524371,I524388,I524405,I524497,I524514,I524531,I524548,I524565,I524582,I524613,I524630,I524647,I524692,I524709,I524726,I524771,I524788,I524805,I524836,I524853,I524884,I524901,I524918,I524949,I524966,I524983,I525000,I525092,I525109,I618096,I618087,I525126,I618105,I525143,I525160,I618102,I525177,I525208,I618084,I525225,I525242,I525287,I618093,I618108,I525304,I618099,I525321,I525366,I618081,I525383,I618090,I525400,I525431,I525448,I525479,I618078,I525496,I525513,I525544,I525561,I525578,I525595,I525687,I525704,I525721,I525738,I525755,I525772,I525670,I525803,I525820,I525837,I525673,I525655,I525882,I525899,I525916,I525676,I525667,I525961,I525978,I525995,I525658,I526026,I526043,I525649,I526074,I526091,I526108,I525679,I526139,I526156,I526173,I526190,I525664,I525661,I525652,I526282,I526299,I526316,I526333,I526350,I526367,I526398,I526415,I526432,I526477,I526494,I526511,I526556,I526573,I526590,I526621,I526638,I526669,I526686,I526703,I526734,I526751,I526768,I526785,I526877,I526894,I526911,I526928,I526945,I526962,I526860,I526993,I527010,I527027,I526863,I526845,I527072,I527089,I527106,I526866,I526857,I527151,I527168,I527185,I526848,I527216,I527233,I526839,I527264,I527281,I527298,I526869,I527329,I527346,I527363,I527380,I526854,I526851,I526842,I527472,I527489,I593494,I593485,I527506,I593503,I527523,I527540,I593482,I527557,I527588,I593491,I527605,I527622,I527667,I593506,I593488,I527684,I593509,I527701,I527746,I593497,I527763,I593479,I527780,I527811,I527828,I527859,I593500,I527876,I527893,I527924,I527941,I527958,I527975,I528067,I528084,I528101,I528118,I528135,I528152,I528183,I528200,I528217,I528262,I528279,I528296,I528341,I528358,I528375,I528406,I528423,I528454,I528471,I528488,I528519,I528536,I528553,I528570,I528662,I528679,I603609,I603600,I528696,I603618,I528713,I528730,I603597,I528747,I528778,I603606,I528795,I528812,I528857,I603621,I603603,I528874,I603624,I528891,I528936,I603612,I528953,I603594,I528970,I529001,I529018,I529049,I603615,I529066,I529083,I529114,I529131,I529148,I529165,I529257,I529274,I529291,I529308,I529325,I529342,I529373,I529390,I529407,I529452,I529469,I529486,I529531,I529548,I529565,I529596,I529613,I529644,I529661,I529678,I529709,I529726,I529743,I529760,I529852,I529869,I529886,I529903,I529920,I529937,I529835,I529968,I529985,I530002,I529838,I529820,I530047,I530064,I530081,I529841,I529832,I530126,I530143,I530160,I529823,I530191,I530208,I529814,I530239,I530256,I530273,I529844,I530304,I530321,I530338,I530355,I529829,I529826,I529817,I530447,I530464,I530481,I530498,I530515,I530532,I530563,I530580,I530597,I530642,I530659,I530676,I530721,I530738,I530755,I530786,I530803,I530834,I530851,I530868,I530899,I530916,I530933,I530950,I531042,I531059,I531076,I531093,I531110,I531127,I531025,I531158,I531175,I531192,I531028,I531010,I531237,I531254,I531271,I531031,I531022,I531316,I531333,I531350,I531013,I531381,I531398,I531004,I531429,I531446,I531463,I531034,I531494,I531511,I531528,I531545,I531019,I531016,I531007,I531637,I531654,I531671,I531688,I531705,I531722,I531753,I531770,I531787,I531832,I531849,I531866,I531911,I531928,I531945,I531976,I531993,I532024,I532041,I532058,I532089,I532106,I532123,I532140,I532232,I532249,I532266,I532283,I532300,I532317,I532215,I532348,I532365,I532382,I532218,I532200,I532427,I532444,I532461,I532221,I532212,I532506,I532523,I532540,I532203,I532571,I532588,I532194,I532619,I532636,I532653,I532224,I532684,I532701,I532718,I532735,I532209,I532206,I532197,I532827,I532844,I532861,I532878,I532895,I532912,I532943,I532960,I532977,I533022,I533039,I533056,I533101,I533118,I533135,I533166,I533183,I533214,I533231,I533248,I533279,I533296,I533313,I533330,I533422,I533439,I533456,I533473,I533490,I533507,I533405,I533538,I533555,I533572,I533408,I533390,I533617,I533634,I533651,I533411,I533402,I533696,I533713,I533730,I533393,I533761,I533778,I533384,I533809,I533826,I533843,I533414,I533874,I533891,I533908,I533925,I533399,I533396,I533387,I534017,I534034,I534051,I534068,I534085,I534102,I534133,I534150,I534167,I534212,I534229,I534246,I534291,I534308,I534325,I534356,I534373,I534404,I534421,I534438,I534469,I534486,I534503,I534520,I534612,I534629,I534646,I534663,I534680,I534697,I534728,I534745,I534762,I534807,I534824,I534841,I534886,I534903,I534920,I534951,I534968,I534999,I535016,I535033,I535064,I535081,I535098,I535115,I535207,I535224,I535241,I535258,I535275,I535292,I535190,I535323,I535340,I535357,I535193,I535175,I535402,I535419,I535436,I535196,I535187,I535481,I535498,I535515,I535178,I535546,I535563,I535169,I535594,I535611,I535628,I535199,I535659,I535676,I535693,I535710,I535184,I535181,I535172,I535802,I535819,I535836,I535853,I535870,I535887,I535918,I535935,I535952,I535997,I536014,I536031,I536076,I536093,I536110,I536141,I536158,I536189,I536206,I536223,I536254,I536271,I536288,I536305,I536397,I536414,I536431,I536448,I536465,I536482,I536513,I536530,I536547,I536592,I536609,I536626,I536671,I536688,I536705,I536736,I536753,I536784,I536801,I536818,I536849,I536866,I536883,I536900,I536992,I537009,I537026,I537043,I537060,I537077,I536975,I537108,I537125,I537142,I536978,I536960,I537187,I537204,I537221,I536981,I536972,I537266,I537283,I537300,I536963,I537331,I537348,I536954,I537379,I537396,I537413,I536984,I537444,I537461,I537478,I537495,I536969,I536966,I536957,I537587,I537604,I537621,I537638,I537655,I537672,I537703,I537720,I537737,I537782,I537799,I537816,I537861,I537878,I537895,I537926,I537943,I537974,I537991,I538008,I538039,I538056,I538073,I538090,I538182,I538199,I538216,I538233,I538250,I538267,I538298,I538315,I538332,I538377,I538394,I538411,I538456,I538473,I538490,I538521,I538538,I538569,I538586,I538603,I538634,I538651,I538668,I538685,I538777,I538794,I538811,I538828,I538845,I538862,I538893,I538910,I538927,I538972,I538989,I539006,I539051,I539068,I539085,I539116,I539133,I539164,I539181,I539198,I539229,I539246,I539263,I539280,I539372,I539389,I686028,I686019,I539406,I686037,I539423,I539440,I686034,I539457,I539488,I686016,I539505,I539522,I539567,I686025,I686040,I539584,I686031,I539601,I539646,I686013,I539663,I686022,I539680,I539711,I539728,I539759,I686010,I539776,I539793,I539824,I539841,I539858,I539875,I539967,I539984,I540001,I540018,I540035,I540052,I539950,I540083,I540100,I540117,I539953,I539935,I540162,I540179,I540196,I539956,I539947,I540241,I540258,I540275,I539938,I540306,I540323,I539929,I540354,I540371,I540388,I539959,I540419,I540436,I540453,I540470,I539944,I539941,I539932,I540562,I540579,I540596,I540613,I540630,I540647,I540545,I540678,I540695,I540712,I540548,I540530,I540757,I540774,I540791,I540551,I540542,I540836,I540853,I540870,I540533,I540901,I540918,I540524,I540949,I540966,I540983,I540554,I541014,I541031,I541048,I541065,I540539,I540536,I540527,I541157,I541174,I672819,I672810,I541191,I672828,I541208,I541225,I672825,I541242,I541273,I672807,I541290,I541307,I541352,I672816,I672831,I541369,I672822,I541386,I541431,I672804,I541448,I672813,I541465,I541496,I541513,I541544,I672801,I541561,I541578,I541609,I541626,I541643,I541660,I541752,I541769,I541786,I541803,I541820,I541837,I541735,I541868,I541885,I541902,I541738,I541720,I541947,I541964,I541981,I541741,I541732,I542026,I542043,I542060,I541723,I542091,I542108,I541714,I542139,I542156,I542173,I541744,I542204,I542221,I542238,I542255,I541729,I541726,I541717,I542347,I542364,I542381,I542398,I542415,I542432,I542330,I542463,I542480,I542497,I542333,I542315,I542542,I542559,I542576,I542336,I542327,I542621,I542638,I542655,I542318,I542686,I542703,I542309,I542734,I542751,I542768,I542339,I542799,I542816,I542833,I542850,I542324,I542321,I542312,I542942,I542959,I542976,I542993,I543010,I543027,I543058,I543075,I543092,I543137,I543154,I543171,I543216,I543233,I543250,I543281,I543298,I543329,I543346,I543363,I543394,I543411,I543428,I543445,I543537,I543554,I543571,I543588,I543605,I543622,I543653,I543670,I543687,I543732,I543749,I543766,I543811,I543828,I543845,I543876,I543893,I543924,I543941,I543958,I543989,I544006,I544023,I544040,I544132,I544149,I544166,I544183,I544200,I544217,I544248,I544265,I544282,I544327,I544344,I544361,I544406,I544423,I544440,I544471,I544488,I544519,I544536,I544553,I544584,I544601,I544618,I544635,I544727,I544744,I544761,I544778,I544795,I544812,I544843,I544860,I544877,I544922,I544939,I544956,I545001,I545018,I545035,I545066,I545083,I545114,I545131,I545148,I545179,I545196,I545213,I545230,I545322,I545339,I545356,I545373,I545390,I545407,I545305,I545438,I545455,I545472,I545308,I545290,I545517,I545534,I545551,I545311,I545302,I545596,I545613,I545630,I545293,I545661,I545678,I545284,I545709,I545726,I545743,I545314,I545774,I545791,I545808,I545825,I545299,I545296,I545287,I545917,I545934,I545951,I545968,I545985,I546002,I545900,I546033,I546050,I546067,I545903,I545885,I546112,I546129,I546146,I545906,I545897,I546191,I546208,I546225,I545888,I546256,I546273,I545879,I546304,I546321,I546338,I545909,I546369,I546386,I546403,I546420,I545894,I545891,I545882,I546512,I546529,I546546,I546563,I546580,I546597,I546628,I546645,I546662,I546707,I546724,I546741,I546786,I546803,I546820,I546851,I546868,I546899,I546916,I546933,I546964,I546981,I546998,I547015,I547107,I547124,I547141,I547158,I547175,I547192,I547223,I547240,I547257,I547302,I547319,I547336,I547381,I547398,I547415,I547446,I547463,I547494,I547511,I547528,I547559,I547576,I547593,I547610,I547702,I547719,I615580,I615571,I547736,I615589,I547753,I547770,I615586,I547787,I547818,I615568,I547835,I547852,I547897,I615577,I615592,I547914,I615583,I547931,I547976,I615565,I547993,I615574,I548010,I548041,I548058,I548089,I615562,I548106,I548123,I548154,I548171,I548188,I548205,I548297,I548314,I548331,I548348,I548365,I548382,I548413,I548430,I548447,I548492,I548509,I548526,I548571,I548588,I548605,I548636,I548653,I548684,I548701,I548718,I548749,I548766,I548783,I548800,I548892,I548909,I548926,I548943,I548960,I548977,I549008,I549025,I549042,I549087,I549104,I549121,I549166,I549183,I549200,I549231,I549248,I549279,I549296,I549313,I549344,I549361,I549378,I549395,I549487,I549504,I699622,I699628,I549521,I699619,I549538,I549555,I699631,I549572,I549603,I699610,I549620,I549637,I549682,I699634,I699616,I549699,I699625,I549716,I549761,I699640,I549778,I699613,I549795,I549826,I549843,I549874,I699637,I549891,I549908,I549939,I549956,I549973,I549990,I550082,I550099,I583974,I583965,I550116,I583983,I550133,I550150,I583962,I550167,I550198,I583971,I550215,I550232,I550277,I583986,I583968,I550294,I583989,I550311,I550356,I583977,I550373,I583959,I550390,I550421,I550438,I550469,I583980,I550486,I550503,I550534,I550551,I550568,I550585,I550677,I550694,I550711,I550728,I550745,I550762,I550793,I550810,I550827,I550872,I550889,I550906,I550951,I550968,I550985,I551016,I551033,I551064,I551081,I551098,I551129,I551146,I551163,I551180,I551272,I551289,I650804,I650795,I551306,I650813,I551323,I551340,I650810,I551357,I551388,I650792,I551405,I551422,I551467,I650801,I650816,I551484,I650807,I551501,I551546,I650789,I551563,I650798,I551580,I551611,I551628,I551659,I650786,I551676,I551693,I551724,I551741,I551758,I551775,I551867,I551884,I551901,I551918,I551935,I551952,I551983,I552000,I552017,I552062,I552079,I552096,I552141,I552158,I552175,I552206,I552223,I552254,I552271,I552288,I552319,I552336,I552353,I552370,I552462,I552479,I552496,I552513,I552530,I552547,I552578,I552595,I552612,I552657,I552674,I552691,I552736,I552753,I552770,I552801,I552818,I552849,I552866,I552883,I552914,I552931,I552948,I552965,I553057,I553074,I553091,I553108,I553125,I553142,I553040,I553173,I553190,I553207,I553043,I553025,I553252,I553269,I553286,I553046,I553037,I553331,I553348,I553365,I553028,I553396,I553413,I553019,I553444,I553461,I553478,I553049,I553509,I553526,I553543,I553560,I553034,I553031,I553022,I553652,I553669,I553686,I553703,I553720,I553737,I553768,I553785,I553802,I553847,I553864,I553881,I553926,I553943,I553960,I553991,I554008,I554039,I554056,I554073,I554104,I554121,I554138,I554155,I554247,I554264,I554281,I554298,I554315,I554332,I554363,I554380,I554397,I554442,I554459,I554476,I554521,I554538,I554555,I554586,I554603,I554634,I554651,I554668,I554699,I554716,I554733,I554750,I554842,I554859,I554876,I554893,I554910,I554927,I554825,I554958,I554975,I554992,I554828,I554810,I555037,I555054,I555071,I554831,I554822,I555116,I555133,I555150,I554813,I555181,I555198,I554804,I555229,I555246,I555263,I554834,I555294,I555311,I555328,I555345,I554819,I554816,I554807,I555437,I555454,I667158,I667149,I555471,I667167,I555488,I555505,I667164,I555522,I555553,I667146,I555570,I555587,I555632,I667155,I667170,I555649,I667161,I555666,I555711,I667143,I555728,I667152,I555745,I555776,I555793,I555824,I667140,I555841,I555858,I555889,I555906,I555923,I555940,I556032,I556049,I556066,I556083,I556100,I556117,I556148,I556165,I556182,I556227,I556244,I556261,I556306,I556323,I556340,I556371,I556388,I556419,I556436,I556453,I556484,I556501,I556518,I556535,I556627,I556644,I556661,I556678,I556695,I556712,I556743,I556760,I556777,I556822,I556839,I556856,I556901,I556918,I556935,I556966,I556983,I557014,I557031,I557048,I557079,I557096,I557113,I557130,I557222,I557239,I557256,I557273,I557290,I557307,I557338,I557355,I557372,I557417,I557434,I557451,I557496,I557513,I557530,I557561,I557578,I557609,I557626,I557643,I557674,I557691,I557708,I557725,I557817,I557834,I557851,I557868,I557885,I557902,I557933,I557950,I557967,I558012,I558029,I558046,I558091,I558108,I558125,I558156,I558173,I558204,I558221,I558238,I558269,I558286,I558303,I558320,I558412,I558429,I558446,I558463,I558480,I558497,I558528,I558545,I558562,I558607,I558624,I558641,I558686,I558703,I558720,I558751,I558768,I558799,I558816,I558833,I558864,I558881,I558898,I558915,I559007,I559024,I674077,I674068,I559041,I674086,I559058,I559075,I674083,I559092,I558990,I559123,I674065,I559140,I559157,I558993,I558975,I559202,I674074,I674089,I559219,I674080,I559236,I558996,I558987,I559281,I674062,I559298,I674071,I559315,I558978,I559346,I559363,I558969,I559394,I674059,I559411,I559428,I558999,I559459,I559476,I559493,I559510,I558984,I558981,I558972,I559602,I559619,I559636,I559653,I559670,I559687,I559718,I559735,I559752,I559797,I559814,I559831,I559876,I559893,I559910,I559941,I559958,I559989,I560006,I560023,I560054,I560071,I560088,I560105,I560197,I560214,I560231,I560248,I560265,I560282,I560313,I560330,I560347,I560392,I560409,I560426,I560471,I560488,I560505,I560536,I560553,I560584,I560601,I560618,I560649,I560666,I560683,I560700,I560792,I560809,I653320,I653311,I560826,I653329,I560843,I560860,I653326,I560877,I560908,I653308,I560925,I560942,I560987,I653317,I653332,I561004,I653323,I561021,I561066,I653305,I561083,I653314,I561100,I561131,I561148,I561179,I653302,I561196,I561213,I561244,I561261,I561278,I561295,I561387,I561404,I561421,I561438,I561455,I561472,I561503,I561520,I561537,I561582,I561599,I561616,I561661,I561678,I561695,I561726,I561743,I561774,I561791,I561808,I561839,I561856,I561873,I561890,I561982,I561999,I562016,I562033,I562050,I562067,I561965,I562098,I562115,I562132,I561968,I561950,I562177,I562194,I562211,I561971,I561962,I562256,I562273,I562290,I561953,I562321,I562338,I561944,I562369,I562386,I562403,I561974,I562434,I562451,I562468,I562485,I561959,I561956,I561947,I562577,I562594,I562611,I562628,I562645,I562662,I562693,I562710,I562727,I562772,I562789,I562806,I562851,I562868,I562885,I562916,I562933,I562964,I562981,I562998,I563029,I563046,I563063,I563080,I563172,I563189,I563206,I563223,I563240,I563257,I563288,I563305,I563322,I563367,I563384,I563401,I563446,I563463,I563480,I563511,I563528,I563559,I563576,I563593,I563624,I563641,I563658,I563675,I563767,I563784,I563801,I563818,I563835,I563852,I563750,I563883,I563900,I563917,I563753,I563735,I563962,I563979,I563996,I563756,I563747,I564041,I564058,I564075,I563738,I564106,I564123,I563729,I564154,I564171,I564188,I563759,I564219,I564236,I564253,I564270,I563744,I563741,I563732,I564362,I564379,I564396,I564413,I564430,I564447,I564345,I564478,I564495,I564512,I564348,I564330,I564557,I564574,I564591,I564351,I564342,I564636,I564653,I564670,I564333,I564701,I564718,I564324,I564749,I564766,I564783,I564354,I564814,I564831,I564848,I564865,I564339,I564336,I564327,I564957,I564974,I564991,I565008,I565025,I565042,I564940,I565073,I565090,I565107,I564943,I564925,I565152,I565169,I565186,I564946,I564937,I565231,I565248,I565265,I564928,I565296,I565313,I564919,I565344,I565361,I565378,I564949,I565409,I565426,I565443,I565460,I564934,I564931,I564922,I565552,I565569,I565586,I565603,I565620,I565637,I565668,I565685,I565702,I565747,I565764,I565781,I565826,I565843,I565860,I565891,I565908,I565939,I565956,I565973,I566004,I566021,I566038,I566055,I566147,I566164,I652691,I652682,I566181,I652700,I566198,I566215,I652697,I566232,I566263,I652679,I566280,I566297,I566342,I652688,I652703,I566359,I652694,I566376,I566421,I652676,I566438,I652685,I566455,I566486,I566503,I566534,I652673,I566551,I566568,I566599,I566616,I566633,I566650,I566742,I566759,I601229,I601220,I566776,I601238,I566793,I566810,I601217,I566827,I566858,I601226,I566875,I566892,I566937,I601241,I601223,I566954,I601244,I566971,I567016,I601232,I567033,I601214,I567050,I567081,I567098,I567129,I601235,I567146,I567163,I567194,I567211,I567228,I567245,I567337,I567354,I567371,I567388,I567405,I567422,I567453,I567470,I567487,I567532,I567549,I567566,I567611,I567628,I567645,I567676,I567693,I567724,I567741,I567758,I567789,I567806,I567823,I567840,I567932,I567949,I656465,I656456,I567966,I656474,I567983,I568000,I656471,I568017,I567915,I568048,I656453,I568065,I568082,I567918,I567900,I568127,I656462,I656477,I568144,I656468,I568161,I567921,I567912,I568206,I656450,I568223,I656459,I568240,I567903,I568271,I568288,I567894,I568319,I656447,I568336,I568353,I567924,I568384,I568401,I568418,I568435,I567909,I567906,I567897,I568527,I568544,I607179,I607170,I568561,I607188,I568578,I568595,I607167,I568612,I568643,I607176,I568660,I568677,I568722,I607191,I607173,I568739,I607194,I568756,I568801,I607182,I568818,I607164,I568835,I568866,I568883,I568914,I607185,I568931,I568948,I568979,I568996,I569013,I569030,I569122,I569139,I569156,I569173,I569190,I569207,I569238,I569255,I569272,I569317,I569334,I569351,I569396,I569413,I569430,I569461,I569478,I569509,I569526,I569543,I569574,I569591,I569608,I569625,I569717,I569734,I569751,I569768,I569785,I569802,I569833,I569850,I569867,I569912,I569929,I569946,I569991,I570008,I570025,I570056,I570073,I570104,I570121,I570138,I570169,I570186,I570203,I570220,I570312,I570329,I570346,I570363,I570380,I570397,I570428,I570445,I570462,I570507,I570524,I570541,I570586,I570603,I570620,I570651,I570668,I570699,I570716,I570733,I570764,I570781,I570798,I570815,I570907,I570924,I715228,I715234,I570941,I715225,I570958,I570975,I715237,I570992,I571023,I715216,I571040,I571057,I571102,I715240,I715222,I571119,I715231,I571136,I571181,I715246,I571198,I715219,I571215,I571246,I571263,I571294,I715243,I571311,I571328,I571359,I571376,I571393,I571410,I571502,I571519,I571536,I571553,I571570,I571587,I571485,I571618,I571635,I571652,I571488,I571470,I571697,I571714,I571731,I571491,I571482,I571776,I571793,I571810,I571473,I571841,I571858,I571464,I571889,I571906,I571923,I571494,I571954,I571971,I571988,I572005,I571479,I571476,I571467,I572097,I572114,I697310,I697316,I572131,I697307,I572148,I572165,I697319,I572182,I572213,I697298,I572230,I572247,I572292,I697322,I697304,I572309,I697313,I572326,I572371,I697328,I572388,I697301,I572405,I572436,I572453,I572484,I697325,I572501,I572518,I572549,I572566,I572583,I572600,I572692,I572709,I572726,I572743,I572760,I572777,I572808,I572825,I572842,I572887,I572904,I572921,I572966,I572983,I573000,I573031,I573048,I573079,I573096,I573113,I573144,I573161,I573178,I573195,I573287,I573304,I573321,I573338,I573355,I573372,I573403,I573420,I573437,I573482,I573499,I573516,I573561,I573578,I573595,I573626,I573643,I573674,I573691,I573708,I573739,I573756,I573773,I573790,I573882,I573899,I573916,I573933,I573950,I573967,I573998,I574015,I574032,I574077,I574094,I574111,I574156,I574173,I574190,I574221,I574238,I574269,I574286,I574303,I574334,I574351,I574368,I574385,I574477,I574494,I574511,I574528,I574545,I574562,I574460,I574593,I574610,I574627,I574463,I574445,I574672,I574689,I574706,I574466,I574457,I574751,I574768,I574785,I574448,I574816,I574833,I574439,I574864,I574881,I574898,I574469,I574929,I574946,I574963,I574980,I574454,I574451,I574442,I575072,I575089,I575106,I575123,I575140,I575157,I575188,I575205,I575222,I575267,I575284,I575301,I575346,I575363,I575380,I575411,I575428,I575459,I575476,I575493,I575524,I575541,I575558,I575575,I575667,I575684,I575701,I575718,I575735,I575752,I575650,I575783,I575800,I575817,I575653,I575635,I575862,I575879,I575896,I575656,I575647,I575941,I575958,I575975,I575638,I576006,I576023,I575629,I576054,I576071,I576088,I575659,I576119,I576136,I576153,I576170,I575644,I575641,I575632,I576262,I576279,I576296,I576313,I576330,I576347,I576378,I576395,I576412,I576457,I576474,I576491,I576536,I576553,I576570,I576601,I576618,I576649,I576666,I576683,I576714,I576731,I576748,I576765,I576857,I576874,I576891,I576908,I576925,I576942,I576959,I576990,I577007,I577024,I577041,I577058,I577075,I577092,I577137,I577154,I577171,I577202,I577219,I577264,I577295,I577312,I577343,I577388,I577452,I577469,I577486,I577503,I577520,I577537,I577554,I577585,I577602,I577619,I577636,I577653,I577670,I577687,I577732,I577749,I577766,I577797,I577814,I577859,I577890,I577907,I577938,I577983,I578047,I578064,I578081,I578098,I578115,I578132,I578149,I578180,I578197,I578214,I578231,I578248,I578265,I578282,I578327,I578344,I578361,I578392,I578409,I578454,I578485,I578502,I578533,I578578,I578642,I578659,I578676,I578693,I578710,I578727,I578744,I578613,I578775,I578792,I578809,I578826,I578843,I578860,I578877,I578610,I578604,I578922,I578939,I578956,I578631,I578987,I579004,I578622,I578616,I579049,I578619,I579080,I579097,I578634,I579128,I578628,I578625,I579173,I578607,I579237,I579254,I579271,I579288,I579305,I579322,I579339,I579370,I579387,I579404,I579421,I579438,I579455,I579472,I579517,I579534,I579551,I579582,I579599,I579644,I579675,I579692,I579723,I579768,I579832,I579849,I579866,I579883,I579900,I579917,I579934,I579803,I579965,I579982,I579999,I580016,I580033,I580050,I580067,I579800,I579794,I580112,I580129,I580146,I579821,I580177,I580194,I579812,I579806,I580239,I579809,I580270,I580287,I579824,I580318,I579818,I579815,I580363,I579797,I580427,I580444,I580461,I580478,I580495,I580512,I580529,I580560,I580577,I580594,I580611,I580628,I580645,I580662,I580707,I580724,I580741,I580772,I580789,I580834,I580865,I580882,I580913,I580958,I581022,I581039,I581056,I581073,I581090,I581107,I581124,I581155,I581172,I581189,I581206,I581223,I581240,I581257,I581302,I581319,I581336,I581367,I581384,I581429,I581460,I581477,I581508,I581553,I581617,I581634,I581651,I581668,I581685,I581702,I581719,I581750,I581767,I581784,I581801,I581818,I581835,I581852,I581897,I581914,I581931,I581962,I581979,I582024,I582055,I582072,I582103,I582148,I582212,I582229,I582246,I582263,I582280,I582297,I582314,I582345,I582362,I582379,I582396,I582413,I582430,I582447,I582492,I582509,I582526,I582557,I582574,I582619,I582650,I582667,I582698,I582743,I582807,I582824,I582841,I582858,I582875,I582892,I582909,I582940,I582957,I582974,I582991,I583008,I583025,I583042,I583087,I583104,I583121,I583152,I583169,I583214,I583245,I583262,I583293,I583338,I583402,I583419,I583436,I583453,I583470,I583487,I583504,I583535,I583552,I583569,I583586,I583603,I583620,I583637,I583682,I583699,I583716,I583747,I583764,I583809,I583840,I583857,I583888,I583933,I583997,I584014,I584031,I584048,I584065,I584082,I584099,I584130,I584147,I584164,I584181,I584198,I584215,I584232,I584277,I584294,I584311,I584342,I584359,I584404,I584435,I584452,I584483,I584528,I584592,I584609,I584626,I584643,I584660,I584677,I584694,I584725,I584742,I584759,I584776,I584793,I584810,I584827,I584872,I584889,I584906,I584937,I584954,I584999,I585030,I585047,I585078,I585123,I585187,I585204,I585221,I585238,I585255,I585272,I585289,I585320,I585337,I585354,I585371,I585388,I585405,I585422,I585467,I585484,I585501,I585532,I585549,I585594,I585625,I585642,I585673,I585718,I585782,I585799,I585816,I585833,I585850,I585867,I585884,I585915,I585932,I585949,I585966,I585983,I586000,I586017,I586062,I586079,I586096,I586127,I586144,I586189,I586220,I586237,I586268,I586313,I586377,I586394,I586411,I586428,I586445,I586462,I586479,I586348,I586510,I586527,I586544,I586561,I586578,I586595,I586612,I586345,I586339,I586657,I586674,I586691,I586366,I586722,I586739,I586357,I586351,I586784,I586354,I586815,I586832,I586369,I586863,I586363,I586360,I586908,I586342,I586972,I586989,I587006,I587023,I587040,I587057,I587074,I587105,I587122,I587139,I587156,I587173,I587190,I587207,I587252,I587269,I587286,I587317,I587334,I587379,I587410,I587427,I587458,I587503,I587567,I587584,I587601,I587618,I587635,I587652,I587669,I587700,I587717,I587734,I587751,I587768,I587785,I587802,I587847,I587864,I587881,I587912,I587929,I587974,I588005,I588022,I588053,I588098,I588162,I588179,I588196,I588213,I588230,I588247,I588264,I588295,I588312,I588329,I588346,I588363,I588380,I588397,I588442,I588459,I588476,I588507,I588524,I588569,I588600,I588617,I588648,I588693,I588757,I588774,I701344,I701347,I588791,I701356,I588808,I588825,I701350,I588842,I701371,I588859,I588890,I701368,I701374,I588907,I701359,I588924,I588941,I588958,I588975,I588992,I589037,I701362,I589054,I701365,I589071,I589102,I589119,I589164,I589195,I701353,I589212,I589243,I589288,I589352,I589369,I589386,I589403,I589420,I589437,I589454,I589323,I589485,I589502,I589519,I589536,I589553,I589570,I589587,I589320,I589314,I589632,I589649,I589666,I589341,I589697,I589714,I589332,I589326,I589759,I589329,I589790,I589807,I589344,I589838,I589338,I589335,I589883,I589317,I589947,I589964,I589981,I589998,I590015,I590032,I590049,I590080,I590097,I590114,I590131,I590148,I590165,I590182,I590227,I590244,I590261,I590292,I590309,I590354,I590385,I590402,I590433,I590478,I590542,I590559,I590576,I590593,I590610,I590627,I590644,I590675,I590692,I590709,I590726,I590743,I590760,I590777,I590822,I590839,I590856,I590887,I590904,I590949,I590980,I590997,I591028,I591073,I591137,I591154,I591171,I591188,I591205,I591222,I591239,I591270,I591287,I591304,I591321,I591338,I591355,I591372,I591417,I591434,I591451,I591482,I591499,I591544,I591575,I591592,I591623,I591668,I591732,I591749,I591766,I591783,I591800,I591817,I591834,I591865,I591882,I591899,I591916,I591933,I591950,I591967,I592012,I592029,I592046,I592077,I592094,I592139,I592170,I592187,I592218,I592263,I592327,I592344,I592361,I592378,I592395,I592412,I592429,I592460,I592477,I592494,I592511,I592528,I592545,I592562,I592607,I592624,I592641,I592672,I592689,I592734,I592765,I592782,I592813,I592858,I592922,I592939,I592956,I592973,I592990,I593007,I593024,I593055,I593072,I593089,I593106,I593123,I593140,I593157,I593202,I593219,I593236,I593267,I593284,I593329,I593360,I593377,I593408,I593453,I593517,I593534,I685411,I685399,I593551,I685384,I593568,I593585,I685396,I593602,I685408,I593619,I593650,I685381,I685405,I593667,I685390,I593684,I593701,I593718,I593735,I593752,I593797,I685393,I593814,I685402,I593831,I593862,I593879,I593924,I593955,I685387,I593972,I594003,I594048,I594112,I594129,I594146,I594163,I594180,I594197,I594214,I594245,I594262,I594279,I594296,I594313,I594330,I594347,I594392,I594409,I594426,I594457,I594474,I594519,I594550,I594567,I594598,I594643,I594707,I594724,I726776,I726779,I594741,I726788,I594758,I594775,I726782,I594792,I726803,I594809,I594840,I726800,I726806,I594857,I726791,I594874,I594891,I594908,I594925,I594942,I594987,I726794,I595004,I726797,I595021,I595052,I595069,I595114,I595145,I726785,I595162,I595193,I595238,I595302,I595319,I595336,I595353,I595370,I595387,I595404,I595435,I595452,I595469,I595486,I595503,I595520,I595537,I595582,I595599,I595616,I595647,I595664,I595709,I595740,I595757,I595788,I595833,I595897,I595914,I595931,I595948,I595965,I595982,I595999,I596030,I596047,I596064,I596081,I596098,I596115,I596132,I596177,I596194,I596211,I596242,I596259,I596304,I596335,I596352,I596383,I596428,I596492,I596509,I596526,I596543,I596560,I596577,I596594,I596625,I596642,I596659,I596676,I596693,I596710,I596727,I596772,I596789,I596806,I596837,I596854,I596899,I596930,I596947,I596978,I597023,I597087,I597104,I597121,I597138,I597155,I597172,I597189,I597220,I597237,I597254,I597271,I597288,I597305,I597322,I597367,I597384,I597401,I597432,I597449,I597494,I597525,I597542,I597573,I597618,I597682,I597699,I710014,I710017,I597716,I710026,I597733,I597750,I710020,I597767,I710041,I597784,I597815,I710038,I710044,I597832,I710029,I597849,I597866,I597883,I597900,I597917,I597962,I710032,I597979,I710035,I597996,I598027,I598044,I598089,I598120,I710023,I598137,I598168,I598213,I598277,I598294,I598311,I598328,I598345,I598362,I598379,I598410,I598427,I598444,I598461,I598478,I598495,I598512,I598557,I598574,I598591,I598622,I598639,I598684,I598715,I598732,I598763,I598808,I598872,I598889,I598906,I598923,I598940,I598957,I598974,I599005,I599022,I599039,I599056,I599073,I599090,I599107,I599152,I599169,I599186,I599217,I599234,I599279,I599310,I599327,I599358,I599403,I599467,I599484,I631317,I631305,I599501,I631290,I599518,I599535,I631302,I599552,I631314,I599569,I599600,I631287,I631311,I599617,I631296,I599634,I599651,I599668,I599685,I599702,I599747,I631299,I599764,I631308,I599781,I599812,I599829,I599874,I599905,I631293,I599922,I599953,I599998,I600062,I600079,I724464,I724467,I600096,I724476,I600113,I600130,I724470,I600147,I724491,I600164,I600033,I600195,I724488,I724494,I600212,I724479,I600229,I600246,I600263,I600280,I600297,I600030,I600024,I600342,I724482,I600359,I724485,I600376,I600051,I600407,I600424,I600042,I600036,I600469,I600039,I600500,I724473,I600517,I600054,I600548,I600048,I600045,I600593,I600027,I600657,I600674,I600691,I600708,I600725,I600742,I600759,I600790,I600807,I600824,I600841,I600858,I600875,I600892,I600937,I600954,I600971,I601002,I601019,I601064,I601095,I601112,I601143,I601188,I601252,I601269,I686669,I686657,I601286,I686642,I601303,I601320,I686654,I601337,I686666,I601354,I601385,I686639,I686663,I601402,I686648,I601419,I601436,I601453,I601470,I601487,I601532,I686651,I601549,I686660,I601566,I601597,I601614,I601659,I601690,I686645,I601707,I601738,I601783,I601847,I601864,I601881,I601898,I601915,I601932,I601949,I601980,I601997,I602014,I602031,I602048,I602065,I602082,I602127,I602144,I602161,I602192,I602209,I602254,I602285,I602302,I602333,I602378,I602442,I602459,I602476,I602493,I602510,I602527,I602544,I602575,I602592,I602609,I602626,I602643,I602660,I602677,I602722,I602739,I602756,I602787,I602804,I602849,I602880,I602897,I602928,I602973,I603037,I603054,I603071,I603088,I603105,I603122,I603139,I603008,I603170,I603187,I603204,I603221,I603238,I603255,I603272,I603005,I602999,I603317,I603334,I603351,I603026,I603382,I603399,I603017,I603011,I603444,I603014,I603475,I603492,I603029,I603523,I603023,I603020,I603568,I603002,I603632,I603649,I603666,I603683,I603700,I603717,I603734,I603765,I603782,I603799,I603816,I603833,I603850,I603867,I603912,I603929,I603946,I603977,I603994,I604039,I604070,I604087,I604118,I604163,I604227,I604244,I637607,I637595,I604261,I637580,I604278,I604295,I637592,I604312,I637604,I604329,I604360,I637577,I637601,I604377,I637586,I604394,I604411,I604428,I604445,I604462,I604507,I637589,I604524,I637598,I604541,I604572,I604589,I604634,I604665,I637583,I604682,I604713,I604758,I604822,I604839,I604856,I604873,I604890,I604907,I604924,I604955,I604972,I604989,I605006,I605023,I605040,I605057,I605102,I605119,I605136,I605167,I605184,I605229,I605260,I605277,I605308,I605353,I605417,I605434,I655848,I655836,I605451,I655821,I605468,I605485,I655833,I605502,I655845,I605519,I605550,I655818,I655842,I605567,I655827,I605584,I605601,I605618,I605635,I605652,I605697,I655830,I605714,I655839,I605731,I605762,I605779,I605824,I605855,I655824,I605872,I605903,I605948,I606012,I606029,I606046,I606063,I606080,I606097,I606114,I606145,I606162,I606179,I606196,I606213,I606230,I606247,I606292,I606309,I606326,I606357,I606374,I606419,I606450,I606467,I606498,I606543,I606607,I606624,I606641,I606658,I606675,I606692,I606709,I606740,I606757,I606774,I606791,I606808,I606825,I606842,I606887,I606904,I606921,I606952,I606969,I607014,I607045,I607062,I607093,I607138,I607202,I607219,I607236,I607253,I607270,I607287,I607304,I607335,I607352,I607369,I607386,I607403,I607420,I607437,I607482,I607499,I607516,I607547,I607564,I607609,I607640,I607657,I607688,I607733,I607797,I607814,I607831,I607848,I607865,I607882,I607899,I607930,I607947,I607964,I607981,I607998,I608015,I608032,I608077,I608094,I608111,I608142,I608159,I608204,I608235,I608252,I608283,I608328,I608392,I608409,I608426,I608443,I608460,I608477,I608494,I608363,I608525,I608542,I608559,I608576,I608593,I608610,I608627,I608360,I608354,I608672,I608689,I608706,I608381,I608737,I608754,I608372,I608366,I608799,I608369,I608830,I608847,I608384,I608878,I608378,I608375,I608923,I608357,I608987,I609004,I609021,I609038,I609055,I609072,I609089,I609120,I609137,I609154,I609171,I609188,I609205,I609222,I609267,I609284,I609301,I609332,I609349,I609394,I609425,I609442,I609473,I609518,I609582,I609599,I609616,I609633,I609650,I609667,I609684,I609715,I609732,I609749,I609766,I609783,I609800,I609817,I609862,I609879,I609896,I609927,I609944,I609989,I610020,I610037,I610068,I610113,I610177,I610194,I677863,I677851,I610211,I677836,I610228,I610245,I677848,I610262,I677860,I610279,I610310,I677833,I677857,I610327,I677842,I610344,I610361,I610378,I610395,I610412,I610457,I677845,I610474,I677854,I610491,I610522,I610539,I610584,I610615,I677839,I610632,I610663,I610708,I610772,I610789,I610806,I610823,I610840,I610857,I610874,I610905,I610922,I610939,I610956,I610973,I610990,I611007,I611052,I611069,I611086,I611117,I611134,I611179,I611210,I611227,I611258,I611303,I611367,I611384,I611401,I611418,I611435,I611452,I611469,I611500,I611517,I611534,I611551,I611568,I611585,I611602,I611647,I611664,I611681,I611712,I611729,I611774,I611805,I611822,I611853,I611898,I611962,I611979,I611996,I612013,I612030,I612047,I612064,I612095,I612112,I612129,I612146,I612163,I612180,I612197,I612242,I612259,I612276,I612307,I612324,I612369,I612400,I612417,I612448,I612493,I612557,I612574,I612591,I612608,I612625,I612642,I612659,I612690,I612707,I612724,I612741,I612758,I612775,I612792,I612837,I612854,I612871,I612902,I612919,I612964,I612995,I613012,I613043,I613088,I613152,I613169,I613186,I613203,I613220,I613237,I613254,I613285,I613302,I613319,I613336,I613353,I613370,I613387,I613432,I613449,I613466,I613497,I613514,I613559,I613590,I613607,I613638,I613683,I613747,I613764,I613781,I613798,I613815,I613832,I613849,I613718,I613880,I613897,I613914,I613931,I613948,I613965,I613982,I613715,I613709,I614027,I614044,I614061,I613736,I614092,I614109,I613727,I613721,I614154,I613724,I614185,I614202,I613739,I614233,I613733,I613730,I614278,I613712,I614342,I614359,I614376,I614393,I614410,I614427,I614444,I614461,I614478,I614495,I614512,I614529,I614546,I614563,I614594,I614611,I614628,I614659,I614690,I614707,I614738,I614783,I614800,I614817,I614876,I614893,I614971,I614988,I615005,I615022,I615039,I615056,I615073,I615090,I615107,I615124,I615141,I615158,I615175,I615192,I615223,I615240,I615257,I615288,I615319,I615336,I615367,I615412,I615429,I615446,I615505,I615522,I615600,I615617,I615634,I615651,I615668,I615685,I615702,I615719,I615736,I615753,I615770,I615787,I615804,I615821,I615852,I615869,I615886,I615917,I615948,I615965,I615996,I616041,I616058,I616075,I616134,I616151,I616229,I616246,I616263,I616280,I616297,I616314,I616331,I616348,I616365,I616382,I616399,I616416,I616433,I616450,I616481,I616498,I616515,I616546,I616577,I616594,I616625,I616670,I616687,I616704,I616763,I616780,I616858,I616875,I616892,I616909,I616926,I616943,I616960,I616977,I616994,I617011,I617028,I617045,I617062,I617079,I617110,I617127,I617144,I617175,I617206,I617223,I617254,I617299,I617316,I617333,I617392,I617409,I617487,I617504,I617521,I617538,I617555,I617572,I617589,I617606,I617623,I617640,I617657,I617674,I617691,I617708,I617739,I617756,I617773,I617804,I617835,I617852,I617883,I617928,I617945,I617962,I618021,I618038,I618116,I618133,I618150,I618167,I618184,I618201,I618218,I618235,I618252,I618269,I618286,I618303,I618320,I618337,I618368,I618385,I618402,I618433,I618464,I618481,I618512,I618557,I618574,I618591,I618650,I618667,I618745,I618762,I618779,I618796,I618813,I618830,I618847,I618864,I618881,I618898,I618915,I618932,I618949,I618966,I618997,I619014,I619031,I619062,I619093,I619110,I619141,I619186,I619203,I619220,I619279,I619296,I619374,I619391,I722158,I619408,I722182,I722167,I619425,I722152,I619442,I619459,I722179,I619476,I619493,I619510,I722161,I619527,I722155,I619544,I722176,I619561,I722164,I619578,I619595,I619626,I619643,I619660,I619691,I722173,I619722,I619739,I619770,I619815,I722170,I619832,I619849,I619908,I619925,I620003,I620020,I620037,I620054,I620071,I620088,I620105,I620122,I620139,I620156,I620173,I620190,I620207,I620224,I620255,I620272,I620289,I620320,I620351,I620368,I620399,I620444,I620461,I620478,I620537,I620554,I620632,I620649,I620666,I620683,I620700,I620717,I620734,I620751,I620768,I620785,I620802,I620819,I620836,I620853,I620884,I620901,I620918,I620949,I620980,I620997,I621028,I621073,I621090,I621107,I621166,I621183,I621261,I621278,I621295,I621312,I621329,I621346,I621363,I621380,I621397,I621414,I621431,I621448,I621465,I621482,I621513,I621530,I621547,I621578,I621609,I621626,I621657,I621702,I621719,I621736,I621795,I621812,I621890,I621907,I621924,I621941,I621958,I621975,I621992,I622009,I622026,I622043,I622060,I622077,I622094,I622111,I622142,I622159,I622176,I622207,I622238,I622255,I622286,I622331,I622348,I622365,I622424,I622441,I622519,I622536,I622553,I622570,I622587,I622604,I622621,I622638,I622655,I622672,I622689,I622706,I622723,I622740,I622771,I622788,I622805,I622836,I622867,I622884,I622915,I622960,I622977,I622994,I623053,I623070,I623148,I623165,I623182,I623199,I623216,I623233,I623250,I623267,I623284,I623301,I623318,I623335,I623352,I623369,I623400,I623417,I623434,I623465,I623496,I623513,I623544,I623589,I623606,I623623,I623682,I623699,I623777,I623794,I623811,I623828,I623845,I623862,I623879,I623896,I623913,I623930,I623947,I623964,I623981,I623998,I624029,I624046,I624063,I624094,I624125,I624142,I624173,I624218,I624235,I624252,I624311,I624328,I624406,I624423,I624440,I624457,I624474,I624491,I624508,I624525,I624542,I624559,I624576,I624593,I624610,I624627,I624658,I624675,I624692,I624723,I624754,I624771,I624802,I624847,I624864,I624881,I624940,I624957,I625035,I625052,I625069,I625086,I625103,I625120,I625137,I625154,I625171,I625188,I625205,I625222,I625239,I625256,I625287,I625304,I625321,I625352,I625383,I625400,I625431,I625476,I625493,I625510,I625569,I625586,I625664,I625681,I625698,I625715,I625732,I625749,I625766,I625783,I625800,I625817,I625834,I625851,I625868,I625885,I625916,I625933,I625950,I625981,I626012,I626029,I626060,I626105,I626122,I626139,I626198,I626215,I626293,I626310,I626327,I626344,I626361,I626378,I626395,I626412,I626429,I626446,I626463,I626480,I626497,I626514,I626545,I626562,I626579,I626610,I626641,I626658,I626689,I626734,I626751,I626768,I626827,I626844,I626922,I626939,I711176,I626956,I711200,I711185,I626973,I711170,I626990,I627007,I711197,I627024,I627041,I627058,I711179,I627075,I711173,I627092,I711194,I627109,I711182,I627126,I627143,I627174,I627191,I627208,I627239,I711191,I627270,I627287,I627318,I627363,I711188,I627380,I627397,I627456,I627473,I627551,I627568,I627585,I627602,I627619,I627636,I627653,I627670,I627687,I627704,I627721,I627738,I627755,I627772,I627803,I627820,I627837,I627868,I627899,I627916,I627947,I627992,I628009,I628026,I628085,I628102,I628180,I628197,I628214,I628231,I628248,I628265,I628282,I628299,I628316,I628333,I628350,I628367,I628384,I628401,I628432,I628449,I628466,I628497,I628528,I628545,I628576,I628621,I628638,I628655,I628714,I628731,I628809,I628826,I628843,I628860,I628877,I628894,I628911,I628928,I628945,I628962,I628979,I628996,I629013,I629030,I629061,I629078,I629095,I629126,I629157,I629174,I629205,I629250,I629267,I629284,I629343,I629360,I629438,I629455,I629472,I629489,I629506,I629523,I629540,I629557,I629574,I629591,I629608,I629625,I629642,I629659,I629690,I629707,I629724,I629755,I629786,I629803,I629834,I629879,I629896,I629913,I629972,I629989,I630067,I630084,I630101,I630118,I630135,I630152,I630169,I630186,I630203,I630220,I630237,I630254,I630271,I630288,I630056,I630319,I630336,I630353,I630029,I630384,I630050,I630415,I630432,I630035,I630463,I630032,I630038,I630508,I630525,I630542,I630044,I630059,I630047,I630601,I630618,I630053,I630041,I630696,I630713,I630730,I630747,I630764,I630781,I630798,I630815,I630832,I630849,I630866,I630883,I630900,I630917,I630948,I630965,I630982,I631013,I631044,I631061,I631092,I631137,I631154,I631171,I631230,I631247,I631325,I631342,I631359,I631376,I631393,I631410,I631427,I631444,I631461,I631478,I631495,I631512,I631529,I631546,I631577,I631594,I631611,I631642,I631673,I631690,I631721,I631766,I631783,I631800,I631859,I631876,I631954,I631971,I631988,I632005,I632022,I632039,I632056,I632073,I632090,I632107,I632124,I632141,I632158,I632175,I632206,I632223,I632240,I632271,I632302,I632319,I632350,I632395,I632412,I632429,I632488,I632505,I632583,I632600,I632617,I632634,I632651,I632668,I632685,I632702,I632719,I632736,I632753,I632770,I632787,I632804,I632835,I632852,I632869,I632900,I632931,I632948,I632979,I633024,I633041,I633058,I633117,I633134,I633212,I633229,I633246,I633263,I633280,I633297,I633314,I633331,I633348,I633365,I633382,I633399,I633416,I633433,I633464,I633481,I633498,I633529,I633560,I633577,I633608,I633653,I633670,I633687,I633746,I633763,I633841,I633858,I633875,I633892,I633909,I633926,I633943,I633960,I633977,I633994,I634011,I634028,I634045,I634062,I634093,I634110,I634127,I634158,I634189,I634206,I634237,I634282,I634299,I634316,I634375,I634392,I634470,I634487,I634504,I634521,I634538,I634555,I634572,I634589,I634606,I634623,I634640,I634657,I634674,I634691,I634459,I634722,I634739,I634756,I634432,I634787,I634453,I634818,I634835,I634438,I634866,I634435,I634441,I634911,I634928,I634945,I634447,I634462,I634450,I635004,I635021,I634456,I634444,I635099,I635116,I635133,I635150,I635167,I635184,I635201,I635218,I635235,I635252,I635269,I635286,I635303,I635320,I635351,I635368,I635385,I635416,I635447,I635464,I635495,I635540,I635557,I635574,I635633,I635650,I635728,I635745,I635762,I635779,I635796,I635813,I635830,I635847,I635864,I635881,I635898,I635915,I635932,I635949,I635980,I635997,I636014,I636045,I636076,I636093,I636124,I636169,I636186,I636203,I636262,I636279,I636357,I636374,I636391,I636408,I636425,I636442,I636459,I636476,I636493,I636510,I636527,I636544,I636561,I636578,I636609,I636626,I636643,I636674,I636705,I636722,I636753,I636798,I636815,I636832,I636891,I636908,I636986,I637003,I637020,I637037,I637054,I637071,I637088,I637105,I637122,I637139,I637156,I637173,I637190,I637207,I637238,I637255,I637272,I637303,I637334,I637351,I637382,I637427,I637444,I637461,I637520,I637537,I637615,I637632,I637649,I637666,I637683,I637700,I637717,I637734,I637751,I637768,I637785,I637802,I637819,I637836,I637867,I637884,I637901,I637932,I637963,I637980,I638011,I638056,I638073,I638090,I638149,I638166,I638244,I638261,I638278,I638295,I638312,I638329,I638346,I638363,I638380,I638397,I638414,I638431,I638448,I638465,I638496,I638513,I638530,I638561,I638592,I638609,I638640,I638685,I638702,I638719,I638778,I638795,I638873,I638890,I638907,I638924,I638941,I638958,I638975,I638992,I639009,I639026,I639043,I639060,I639077,I639094,I639125,I639142,I639159,I639190,I639221,I639238,I639269,I639314,I639331,I639348,I639407,I639424,I639502,I639519,I639536,I639553,I639570,I639587,I639604,I639621,I639638,I639655,I639672,I639689,I639706,I639723,I639754,I639771,I639788,I639819,I639850,I639867,I639898,I639943,I639960,I639977,I640036,I640053,I640131,I640148,I640165,I640182,I640199,I640216,I640233,I640250,I640267,I640284,I640301,I640318,I640335,I640352,I640383,I640400,I640417,I640448,I640479,I640496,I640527,I640572,I640589,I640606,I640665,I640682,I640760,I640777,I640794,I640811,I640828,I640845,I640862,I640879,I640896,I640913,I640930,I640947,I640964,I640981,I641012,I641029,I641046,I641077,I641108,I641125,I641156,I641201,I641218,I641235,I641294,I641311,I641389,I641406,I706552,I641423,I706576,I706561,I641440,I706546,I641457,I641474,I706573,I641491,I641508,I641525,I706555,I641542,I706549,I641559,I706570,I641576,I706558,I641593,I641610,I641378,I641641,I641658,I641675,I641351,I641706,I706567,I641372,I641737,I641754,I641357,I641785,I641354,I641360,I641830,I706564,I641847,I641864,I641366,I641381,I641369,I641923,I641940,I641375,I641363,I642018,I642035,I642052,I642069,I642086,I642103,I642120,I642137,I642154,I642171,I642188,I642205,I642222,I642239,I642270,I642287,I642304,I642335,I642366,I642383,I642414,I642459,I642476,I642493,I642552,I642569,I642647,I642664,I696726,I642681,I696750,I696735,I642698,I696720,I642715,I642732,I696747,I642749,I642766,I642783,I696729,I642800,I696723,I642817,I696744,I642834,I696732,I642851,I642868,I642899,I642916,I642933,I642964,I696741,I642995,I643012,I643043,I643088,I696738,I643105,I643122,I643181,I643198,I643276,I643293,I643310,I643327,I643344,I643361,I643378,I643395,I643412,I643429,I643446,I643463,I643480,I643497,I643528,I643545,I643562,I643593,I643624,I643641,I643672,I643717,I643734,I643751,I643810,I643827,I643905,I643922,I643939,I643956,I643973,I643990,I644007,I644024,I644041,I644058,I644075,I644092,I644109,I644126,I644157,I644174,I644191,I644222,I644253,I644270,I644301,I644346,I644363,I644380,I644439,I644456,I644534,I644551,I644568,I644585,I644602,I644619,I644636,I644653,I644670,I644687,I644704,I644721,I644738,I644755,I644786,I644803,I644820,I644851,I644882,I644899,I644930,I644975,I644992,I645009,I645068,I645085,I645163,I645180,I645197,I645214,I645231,I645248,I645265,I645282,I645299,I645316,I645333,I645350,I645367,I645384,I645415,I645432,I645449,I645480,I645511,I645528,I645559,I645604,I645621,I645638,I645697,I645714,I645792,I645809,I645826,I645843,I645860,I645877,I645894,I645911,I645928,I645945,I645962,I645979,I645996,I646013,I646044,I646061,I646078,I646109,I646140,I646157,I646188,I646233,I646250,I646267,I646326,I646343,I646421,I646438,I646455,I646472,I646489,I646506,I646523,I646540,I646557,I646574,I646591,I646608,I646625,I646642,I646673,I646690,I646707,I646738,I646769,I646786,I646817,I646862,I646879,I646896,I646955,I646972,I647050,I647067,I647084,I647101,I647118,I647135,I647152,I647169,I647186,I647203,I647220,I647237,I647254,I647271,I647302,I647319,I647336,I647367,I647398,I647415,I647446,I647491,I647508,I647525,I647584,I647601,I647679,I647696,I647713,I647730,I647747,I647764,I647781,I647798,I647815,I647832,I647849,I647866,I647883,I647900,I647931,I647948,I647965,I647996,I648027,I648044,I648075,I648120,I648137,I648154,I648213,I648230,I648308,I648325,I648342,I648359,I648376,I648393,I648410,I648427,I648444,I648461,I648478,I648495,I648512,I648529,I648560,I648577,I648594,I648625,I648656,I648673,I648704,I648749,I648766,I648783,I648842,I648859,I648937,I648954,I648971,I648988,I649005,I649022,I649039,I649056,I649073,I649090,I649107,I649124,I649141,I649158,I649189,I649206,I649223,I649254,I649285,I649302,I649333,I649378,I649395,I649412,I649471,I649488,I649566,I649583,I649600,I649617,I649634,I649651,I649668,I649685,I649702,I649719,I649736,I649753,I649770,I649787,I649818,I649835,I649852,I649883,I649914,I649931,I649962,I650007,I650024,I650041,I650100,I650117,I650195,I650212,I723892,I650229,I723916,I723901,I650246,I723886,I650263,I650280,I723913,I650297,I650314,I650331,I723895,I650348,I723889,I650365,I723910,I650382,I723898,I650399,I650416,I650447,I650464,I650481,I650512,I723907,I650543,I650560,I650591,I650636,I723904,I650653,I650670,I650729,I650746,I650824,I650841,I650858,I650875,I650892,I650909,I650926,I650943,I650960,I650977,I650994,I651011,I651028,I651045,I651076,I651093,I651110,I651141,I651172,I651189,I651220,I651265,I651282,I651299,I651358,I651375,I651453,I651470,I651487,I651504,I651521,I651538,I651555,I651572,I651589,I651606,I651623,I651640,I651657,I651674,I651705,I651722,I651739,I651770,I651801,I651818,I651849,I651894,I651911,I651928,I651987,I652004,I652082,I652099,I652116,I652133,I652150,I652167,I652184,I652201,I652218,I652235,I652252,I652269,I652286,I652303,I652334,I652351,I652368,I652399,I652430,I652447,I652478,I652523,I652540,I652557,I652616,I652633,I652711,I652728,I652745,I652762,I652779,I652796,I652813,I652830,I652847,I652864,I652881,I652898,I652915,I652932,I652963,I652980,I652997,I653028,I653059,I653076,I653107,I653152,I653169,I653186,I653245,I653262,I653340,I653357,I653374,I653391,I653408,I653425,I653442,I653459,I653476,I653493,I653510,I653527,I653544,I653561,I653592,I653609,I653626,I653657,I653688,I653705,I653736,I653781,I653798,I653815,I653874,I653891,I653969,I653986,I654003,I654020,I654037,I654054,I654071,I654088,I654105,I654122,I654139,I654156,I654173,I654190,I654221,I654238,I654255,I654286,I654317,I654334,I654365,I654410,I654427,I654444,I654503,I654520,I654598,I654615,I654632,I654649,I654666,I654683,I654700,I654717,I654734,I654751,I654768,I654785,I654802,I654819,I654587,I654850,I654867,I654884,I654560,I654915,I654581,I654946,I654963,I654566,I654994,I654563,I654569,I655039,I655056,I655073,I654575,I654590,I654578,I655132,I655149,I654584,I654572,I655227,I655244,I655261,I655278,I655295,I655312,I655329,I655346,I655363,I655380,I655397,I655414,I655431,I655448,I655216,I655479,I655496,I655513,I655189,I655544,I655210,I655575,I655592,I655195,I655623,I655192,I655198,I655668,I655685,I655702,I655204,I655219,I655207,I655761,I655778,I655213,I655201,I655856,I655873,I655890,I655907,I655924,I655941,I655958,I655975,I655992,I656009,I656026,I656043,I656060,I656077,I656108,I656125,I656142,I656173,I656204,I656221,I656252,I656297,I656314,I656331,I656390,I656407,I656485,I656502,I656519,I656536,I656553,I656570,I656587,I656604,I656621,I656638,I656655,I656672,I656689,I656706,I656737,I656754,I656771,I656802,I656833,I656850,I656881,I656926,I656943,I656960,I657019,I657036,I657114,I657131,I657148,I657165,I657182,I657199,I657216,I657233,I657250,I657267,I657284,I657301,I657318,I657335,I657366,I657383,I657400,I657431,I657462,I657479,I657510,I657555,I657572,I657589,I657648,I657665,I657743,I657760,I657777,I657794,I657811,I657828,I657845,I657862,I657879,I657896,I657913,I657930,I657947,I657964,I657995,I658012,I658029,I658060,I658091,I658108,I658139,I658184,I658201,I658218,I658277,I658294,I658372,I658389,I658406,I658423,I658440,I658457,I658474,I658491,I658508,I658525,I658542,I658559,I658576,I658593,I658624,I658641,I658658,I658689,I658720,I658737,I658768,I658813,I658830,I658847,I658906,I658923,I659001,I659018,I659035,I659052,I659069,I659086,I659103,I659120,I659137,I659154,I659171,I659188,I659205,I659222,I658990,I659253,I659270,I659287,I658963,I659318,I658984,I659349,I659366,I658969,I659397,I658966,I658972,I659442,I659459,I659476,I658978,I658993,I658981,I659535,I659552,I658987,I658975,I659630,I659647,I659664,I659681,I659698,I659715,I659732,I659749,I659766,I659783,I659800,I659817,I659834,I659851,I659882,I659899,I659916,I659947,I659978,I659995,I660026,I660071,I660088,I660105,I660164,I660181,I660259,I660276,I660293,I660310,I660327,I660344,I660361,I660378,I660395,I660412,I660429,I660446,I660463,I660480,I660511,I660528,I660545,I660576,I660607,I660624,I660655,I660700,I660717,I660734,I660793,I660810,I660888,I660905,I660922,I660939,I660956,I660973,I660990,I661007,I661024,I661041,I661058,I661075,I661092,I661109,I661140,I661157,I661174,I661205,I661236,I661253,I661284,I661329,I661346,I661363,I661422,I661439,I661517,I661534,I661551,I661568,I661585,I661602,I661619,I661636,I661653,I661670,I661687,I661704,I661721,I661738,I661769,I661786,I661803,I661834,I661865,I661882,I661913,I661958,I661975,I661992,I662051,I662068,I662146,I662163,I662180,I662197,I662214,I662231,I662248,I662265,I662282,I662299,I662316,I662333,I662350,I662367,I662398,I662415,I662432,I662463,I662494,I662511,I662542,I662587,I662604,I662621,I662680,I662697,I662775,I662792,I662809,I662826,I662843,I662860,I662877,I662894,I662911,I662928,I662945,I662962,I662979,I662996,I663027,I663044,I663061,I663092,I663123,I663140,I663171,I663216,I663233,I663250,I663309,I663326,I663404,I663421,I663438,I663455,I663472,I663489,I663506,I663523,I663540,I663557,I663574,I663591,I663608,I663625,I663656,I663673,I663690,I663721,I663752,I663769,I663800,I663845,I663862,I663879,I663938,I663955,I664033,I664050,I664067,I664084,I664101,I664118,I664135,I664152,I664169,I664186,I664203,I664220,I664237,I664254,I664285,I664302,I664319,I664350,I664381,I664398,I664429,I664474,I664491,I664508,I664567,I664584,I664662,I664679,I664696,I664713,I664730,I664747,I664764,I664781,I664798,I664815,I664832,I664849,I664866,I664883,I664914,I664931,I664948,I664979,I665010,I665027,I665058,I665103,I665120,I665137,I665196,I665213,I665291,I665308,I696148,I665325,I696172,I696157,I665342,I696142,I665359,I665376,I696169,I665393,I665410,I665427,I696151,I665444,I696145,I665461,I696166,I665478,I696154,I665495,I665512,I665280,I665543,I665560,I665577,I665253,I665608,I696163,I665274,I665639,I665656,I665259,I665687,I665256,I665262,I665732,I696160,I665749,I665766,I665268,I665283,I665271,I665825,I665842,I665277,I665265,I665920,I665937,I665954,I665971,I665988,I666005,I666022,I666039,I666056,I666073,I666090,I666107,I666124,I666141,I666172,I666189,I666206,I666237,I666268,I666285,I666316,I666361,I666378,I666395,I666454,I666471,I666549,I666566,I666583,I666600,I666617,I666634,I666651,I666668,I666685,I666702,I666719,I666736,I666753,I666770,I666801,I666818,I666835,I666866,I666897,I666914,I666945,I666990,I667007,I667024,I667083,I667100,I667178,I667195,I667212,I667229,I667246,I667263,I667280,I667297,I667314,I667331,I667348,I667365,I667382,I667399,I667430,I667447,I667464,I667495,I667526,I667543,I667574,I667619,I667636,I667653,I667712,I667729,I667807,I667824,I667841,I667858,I667875,I667892,I667909,I667926,I667943,I667960,I667977,I667994,I668011,I668028,I667796,I668059,I668076,I668093,I667769,I668124,I667790,I668155,I668172,I667775,I668203,I667772,I667778,I668248,I668265,I668282,I667784,I667799,I667787,I668341,I668358,I667793,I667781,I668436,I668453,I694992,I668470,I695016,I695001,I668487,I694986,I668504,I668521,I695013,I668538,I668555,I668572,I694995,I668589,I694989,I668606,I695010,I668623,I694998,I668640,I668657,I668688,I668705,I668722,I668753,I695007,I668784,I668801,I668832,I668877,I695004,I668894,I668911,I668970,I668987,I669065,I669082,I669099,I669116,I669133,I669150,I669167,I669184,I669201,I669218,I669235,I669252,I669269,I669286,I669317,I669334,I669351,I669382,I669413,I669430,I669461,I669506,I669523,I669540,I669599,I669616,I669694,I669711,I669728,I669745,I669762,I669779,I669796,I669813,I669830,I669847,I669864,I669881,I669898,I669915,I669946,I669963,I669980,I670011,I670042,I670059,I670090,I670135,I670152,I670169,I670228,I670245,I670323,I670340,I670357,I670374,I670391,I670408,I670425,I670442,I670459,I670476,I670493,I670510,I670527,I670544,I670575,I670592,I670609,I670640,I670671,I670688,I670719,I670764,I670781,I670798,I670857,I670874,I670952,I670969,I670986,I671003,I671020,I671037,I671054,I671071,I671088,I671105,I671122,I671139,I671156,I671173,I671204,I671221,I671238,I671269,I671300,I671317,I671348,I671393,I671410,I671427,I671486,I671503,I671581,I671598,I671615,I671632,I671649,I671666,I671683,I671700,I671717,I671734,I671751,I671768,I671785,I671802,I671833,I671850,I671867,I671898,I671929,I671946,I671977,I672022,I672039,I672056,I672115,I672132,I672210,I672227,I672244,I672261,I672278,I672295,I672312,I672329,I672346,I672363,I672380,I672397,I672414,I672431,I672462,I672479,I672496,I672527,I672558,I672575,I672606,I672651,I672668,I672685,I672744,I672761,I672839,I672856,I672873,I672890,I672907,I672924,I672941,I672958,I672975,I672992,I673009,I673026,I673043,I673060,I673091,I673108,I673125,I673156,I673187,I673204,I673235,I673280,I673297,I673314,I673373,I673390,I673468,I673485,I673502,I673519,I673536,I673553,I673570,I673587,I673604,I673621,I673638,I673655,I673672,I673689,I673457,I673720,I673737,I673754,I673430,I673785,I673451,I673816,I673833,I673436,I673864,I673433,I673439,I673909,I673926,I673943,I673445,I673460,I673448,I674002,I674019,I673454,I673442,I674097,I674114,I674131,I674148,I674165,I674182,I674199,I674216,I674233,I674250,I674267,I674284,I674301,I674318,I674349,I674366,I674383,I674414,I674445,I674462,I674493,I674538,I674555,I674572,I674631,I674648,I674726,I674743,I674760,I674777,I674794,I674811,I674828,I674845,I674862,I674879,I674896,I674913,I674930,I674947,I674978,I674995,I675012,I675043,I675074,I675091,I675122,I675167,I675184,I675201,I675260,I675277,I675355,I675372,I675389,I675406,I675423,I675440,I675457,I675474,I675491,I675508,I675525,I675542,I675559,I675576,I675607,I675624,I675641,I675672,I675703,I675720,I675751,I675796,I675813,I675830,I675889,I675906,I675984,I676001,I676018,I676035,I676052,I676069,I676086,I676103,I676120,I676137,I676154,I676171,I676188,I676205,I676236,I676253,I676270,I676301,I676332,I676349,I676380,I676425,I676442,I676459,I676518,I676535,I676613,I676630,I676647,I676664,I676681,I676698,I676715,I676732,I676749,I676766,I676783,I676800,I676817,I676834,I676865,I676882,I676899,I676930,I676961,I676978,I677009,I677054,I677071,I677088,I677147,I677164,I677242,I677259,I718112,I677276,I718136,I718121,I677293,I718106,I677310,I677327,I718133,I677344,I677361,I677378,I718115,I677395,I718109,I677412,I718130,I677429,I718118,I677446,I677463,I677494,I677511,I677528,I677559,I718127,I677590,I677607,I677638,I677683,I718124,I677700,I677717,I677776,I677793,I677871,I677888,I677905,I677922,I677939,I677956,I677973,I677990,I678007,I678024,I678041,I678058,I678075,I678092,I678123,I678140,I678157,I678188,I678219,I678236,I678267,I678312,I678329,I678346,I678405,I678422,I678500,I678517,I678534,I678551,I678568,I678585,I678602,I678619,I678636,I678653,I678670,I678687,I678704,I678721,I678752,I678769,I678786,I678817,I678848,I678865,I678896,I678941,I678958,I678975,I679034,I679051,I679129,I679146,I679163,I679180,I679197,I679214,I679231,I679248,I679265,I679282,I679299,I679316,I679333,I679350,I679381,I679398,I679415,I679446,I679477,I679494,I679525,I679570,I679587,I679604,I679663,I679680,I679758,I679775,I679792,I679809,I679826,I679843,I679860,I679877,I679894,I679911,I679928,I679945,I679962,I679979,I680010,I680027,I680044,I680075,I680106,I680123,I680154,I680199,I680216,I680233,I680292,I680309,I680387,I680404,I680421,I680438,I680455,I680472,I680489,I680506,I680523,I680540,I680557,I680574,I680591,I680608,I680639,I680656,I680673,I680704,I680735,I680752,I680783,I680828,I680845,I680862,I680921,I680938,I681016,I681033,I681050,I681067,I681084,I681101,I681118,I681135,I681152,I681169,I681186,I681203,I681220,I681237,I681268,I681285,I681302,I681333,I681364,I681381,I681412,I681457,I681474,I681491,I681550,I681567,I681645,I681662,I681679,I681696,I681713,I681730,I681747,I681764,I681781,I681798,I681815,I681832,I681849,I681866,I681897,I681914,I681931,I681962,I681993,I682010,I682041,I682086,I682103,I682120,I682179,I682196,I682274,I682291,I682308,I682325,I682342,I682359,I682376,I682393,I682410,I682427,I682444,I682461,I682478,I682495,I682526,I682543,I682560,I682591,I682622,I682639,I682670,I682715,I682732,I682749,I682808,I682825,I682903,I682920,I682937,I682954,I682971,I682988,I683005,I683022,I683039,I683056,I683073,I683090,I683107,I683124,I683155,I683172,I683189,I683220,I683251,I683268,I683299,I683344,I683361,I683378,I683437,I683454,I683532,I683549,I683566,I683583,I683600,I683617,I683634,I683651,I683668,I683685,I683702,I683719,I683736,I683753,I683784,I683801,I683818,I683849,I683880,I683897,I683928,I683973,I683990,I684007,I684066,I684083,I684161,I684178,I684195,I684212,I684229,I684246,I684263,I684280,I684297,I684314,I684331,I684348,I684365,I684382,I684413,I684430,I684447,I684478,I684509,I684526,I684557,I684602,I684619,I684636,I684695,I684712,I684790,I684807,I684824,I684841,I684858,I684875,I684892,I684909,I684926,I684943,I684960,I684977,I684994,I685011,I685042,I685059,I685076,I685107,I685138,I685155,I685186,I685231,I685248,I685265,I685324,I685341,I685419,I685436,I685453,I685470,I685487,I685504,I685521,I685538,I685555,I685572,I685589,I685606,I685623,I685640,I685671,I685688,I685705,I685736,I685767,I685784,I685815,I685860,I685877,I685894,I685953,I685970,I686048,I686065,I686082,I686099,I686116,I686133,I686150,I686167,I686184,I686201,I686218,I686235,I686252,I686269,I686300,I686317,I686334,I686365,I686396,I686413,I686444,I686489,I686506,I686523,I686582,I686599,I686677,I686694,I686711,I686728,I686745,I686762,I686779,I686796,I686813,I686830,I686847,I686864,I686881,I686898,I686929,I686946,I686963,I686994,I687025,I687042,I687073,I687118,I687135,I687152,I687211,I687228,I687306,I687323,I687340,I687357,I687374,I687391,I687408,I687425,I687442,I687459,I687476,I687493,I687510,I687527,I687295,I687558,I687575,I687592,I687268,I687623,I687289,I687654,I687671,I687274,I687702,I687271,I687277,I687747,I687764,I687781,I687283,I687298,I687286,I687840,I687857,I687292,I687280,I687935,I687952,I687969,I687986,I688003,I688020,I688037,I688054,I688071,I688088,I688105,I688122,I688139,I688156,I688187,I688204,I688221,I688252,I688283,I688300,I688331,I688376,I688393,I688410,I688469,I688486,I688564,I688581,I688598,I688615,I688632,I688649,I688666,I688683,I688700,I688717,I688734,I688751,I688768,I688785,I688816,I688833,I688850,I688881,I688912,I688929,I688960,I689005,I689022,I689039,I689098,I689115,I689193,I689210,I689227,I689244,I689261,I689278,I689295,I689312,I689329,I689346,I689363,I689380,I689397,I689414,I689445,I689462,I689479,I689510,I689541,I689558,I689589,I689634,I689651,I689668,I689727,I689744,I689822,I689839,I689856,I689873,I689904,I689935,I689952,I689969,I689986,I690003,I690034,I690065,I690082,I690099,I690116,I690133,I690150,I690181,I690198,I690215,I690274,I690319,I690336,I690400,I690417,I690434,I690451,I690482,I690513,I690530,I690547,I690564,I690581,I690612,I690643,I690660,I690677,I690694,I690711,I690728,I690759,I690776,I690793,I690852,I690897,I690914,I690978,I690995,I691012,I691029,I691060,I691091,I691108,I691125,I691142,I691159,I691190,I691221,I691238,I691255,I691272,I691289,I691306,I691337,I691354,I691371,I691430,I691475,I691492,I691556,I691573,I691590,I691607,I691638,I691669,I691686,I691703,I691720,I691737,I691768,I691799,I691816,I691833,I691850,I691867,I691884,I691915,I691932,I691949,I692008,I692053,I692070,I692134,I692151,I692168,I692185,I692216,I692247,I692264,I692281,I692298,I692315,I692346,I692377,I692394,I692411,I692428,I692445,I692462,I692493,I692510,I692527,I692586,I692631,I692648,I692712,I692729,I692746,I692763,I692794,I692825,I692842,I692859,I692876,I692893,I692924,I692955,I692972,I692989,I693006,I693023,I693040,I693071,I693088,I693105,I693164,I693209,I693226,I693290,I693307,I693324,I693341,I693372,I693403,I693420,I693437,I693454,I693471,I693502,I693533,I693550,I693567,I693584,I693601,I693618,I693649,I693666,I693683,I693742,I693787,I693804,I693868,I693885,I693902,I693919,I693950,I693981,I693998,I694015,I694032,I694049,I694080,I694111,I694128,I694145,I694162,I694179,I694196,I694227,I694244,I694261,I694320,I694365,I694382,I694446,I694463,I694480,I694497,I694528,I694559,I694576,I694593,I694610,I694627,I694658,I694689,I694706,I694723,I694740,I694757,I694774,I694805,I694822,I694839,I694898,I694943,I694960,I695024,I695041,I695058,I695075,I695106,I695137,I695154,I695171,I695188,I695205,I695236,I695267,I695284,I695301,I695318,I695335,I695352,I695383,I695400,I695417,I695476,I695521,I695538,I695602,I695619,I695636,I695653,I695684,I695715,I695732,I695749,I695766,I695783,I695814,I695845,I695862,I695879,I695896,I695913,I695930,I695961,I695978,I695995,I696054,I696099,I696116,I696180,I696197,I696214,I696231,I696262,I696293,I696310,I696327,I696344,I696361,I696392,I696423,I696440,I696457,I696474,I696491,I696508,I696539,I696556,I696573,I696632,I696677,I696694,I696758,I696775,I696792,I696809,I696840,I696871,I696888,I696905,I696922,I696939,I696970,I697001,I697018,I697035,I697052,I697069,I697086,I697117,I697134,I697151,I697210,I697255,I697272,I697336,I697353,I697370,I697387,I697418,I697449,I697466,I697483,I697500,I697517,I697548,I697579,I697596,I697613,I697630,I697647,I697664,I697695,I697712,I697729,I697788,I697833,I697850,I697914,I697931,I697948,I697965,I697996,I698027,I698044,I698061,I698078,I698095,I698126,I698157,I698174,I698191,I698208,I698225,I698242,I698273,I698290,I698307,I698366,I698411,I698428,I698492,I698509,I698526,I698543,I698574,I698605,I698622,I698639,I698656,I698673,I698704,I698735,I698752,I698769,I698786,I698803,I698820,I698851,I698868,I698885,I698944,I698989,I699006,I699070,I699087,I699104,I699121,I699152,I699183,I699200,I699217,I699234,I699251,I699282,I699313,I699330,I699347,I699364,I699381,I699398,I699429,I699446,I699463,I699522,I699567,I699584,I699648,I699665,I699682,I699699,I699730,I699761,I699778,I699795,I699812,I699829,I699860,I699891,I699908,I699925,I699942,I699959,I699976,I700007,I700024,I700041,I700100,I700145,I700162,I700226,I700243,I700260,I700277,I700308,I700339,I700356,I700373,I700390,I700407,I700438,I700469,I700486,I700503,I700520,I700537,I700554,I700585,I700602,I700619,I700678,I700723,I700740,I700804,I700821,I700838,I700855,I700886,I700917,I700934,I700951,I700968,I700985,I701016,I701047,I701064,I701081,I701098,I701115,I701132,I701163,I701180,I701197,I701256,I701301,I701318,I701382,I701399,I701416,I701433,I701464,I701495,I701512,I701529,I701546,I701563,I701594,I701625,I701642,I701659,I701676,I701693,I701710,I701741,I701758,I701775,I701834,I701879,I701896,I701960,I701977,I701994,I702011,I702042,I702073,I702090,I702107,I702124,I702141,I702172,I702203,I702220,I702237,I702254,I702271,I702288,I702319,I702336,I702353,I702412,I702457,I702474,I702538,I702555,I702572,I702589,I702620,I702651,I702668,I702685,I702702,I702719,I702750,I702781,I702798,I702815,I702832,I702849,I702866,I702897,I702914,I702931,I702990,I703035,I703052,I703116,I703133,I703150,I703167,I703198,I703229,I703246,I703263,I703280,I703297,I703328,I703359,I703376,I703393,I703410,I703427,I703444,I703475,I703492,I703509,I703568,I703613,I703630,I703694,I703711,I703728,I703745,I703776,I703807,I703824,I703841,I703858,I703875,I703906,I703937,I703954,I703971,I703988,I704005,I704022,I704053,I704070,I704087,I704146,I704191,I704208,I704272,I704289,I704306,I704323,I704354,I704385,I704402,I704419,I704436,I704453,I704484,I704515,I704532,I704549,I704566,I704583,I704600,I704631,I704648,I704665,I704724,I704769,I704786,I704850,I704867,I704884,I704901,I704932,I704963,I704980,I704997,I705014,I705031,I705062,I705093,I705110,I705127,I705144,I705161,I705178,I705209,I705226,I705243,I705302,I705347,I705364,I705428,I705445,I705462,I705479,I705510,I705541,I705558,I705575,I705592,I705609,I705640,I705671,I705688,I705705,I705722,I705739,I705756,I705787,I705804,I705821,I705880,I705925,I705942,I706006,I706023,I706040,I706057,I706088,I706119,I706136,I706153,I706170,I706187,I706218,I706249,I706266,I706283,I706300,I706317,I706334,I706365,I706382,I706399,I706458,I706503,I706520,I706584,I706601,I706618,I706635,I706666,I706697,I706714,I706731,I706748,I706765,I706796,I706827,I706844,I706861,I706878,I706895,I706912,I706943,I706960,I706977,I707036,I707081,I707098,I707162,I707179,I707196,I707213,I707244,I707275,I707292,I707309,I707326,I707343,I707374,I707405,I707422,I707439,I707456,I707473,I707490,I707521,I707538,I707555,I707614,I707659,I707676,I707740,I707757,I707774,I707791,I707822,I707853,I707870,I707887,I707904,I707921,I707952,I707983,I708000,I708017,I708034,I708051,I708068,I708099,I708116,I708133,I708192,I708237,I708254,I708318,I708335,I708352,I708369,I708400,I708431,I708448,I708465,I708482,I708499,I708530,I708561,I708578,I708595,I708612,I708629,I708646,I708677,I708694,I708711,I708770,I708815,I708832,I708896,I708913,I708930,I708947,I708978,I709009,I709026,I709043,I709060,I709077,I709108,I709139,I709156,I709173,I709190,I709207,I709224,I709255,I709272,I709289,I709348,I709393,I709410,I709474,I709491,I709508,I709525,I709556,I709587,I709604,I709621,I709638,I709655,I709686,I709717,I709734,I709751,I709768,I709785,I709802,I709833,I709850,I709867,I709926,I709971,I709988,I710052,I710069,I710086,I710103,I710134,I710165,I710182,I710199,I710216,I710233,I710264,I710295,I710312,I710329,I710346,I710363,I710380,I710411,I710428,I710445,I710504,I710549,I710566,I710630,I710647,I710664,I710681,I710712,I710743,I710760,I710777,I710794,I710811,I710842,I710873,I710890,I710907,I710924,I710941,I710958,I710989,I711006,I711023,I711082,I711127,I711144,I711208,I711225,I711242,I711259,I711290,I711321,I711338,I711355,I711372,I711389,I711420,I711451,I711468,I711485,I711502,I711519,I711536,I711567,I711584,I711601,I711660,I711705,I711722,I711786,I711803,I711820,I711837,I711868,I711899,I711916,I711933,I711950,I711967,I711998,I712029,I712046,I712063,I712080,I712097,I712114,I712145,I712162,I712179,I712238,I712283,I712300,I712364,I712381,I712398,I712415,I712446,I712477,I712494,I712511,I712528,I712545,I712576,I712607,I712624,I712641,I712658,I712675,I712692,I712723,I712740,I712757,I712816,I712861,I712878,I712942,I712959,I712976,I712993,I713024,I713055,I713072,I713089,I713106,I713123,I713154,I713185,I713202,I713219,I713236,I713253,I713270,I713301,I713318,I713335,I713394,I713439,I713456,I713520,I713537,I713554,I713571,I713602,I713633,I713650,I713667,I713684,I713701,I713732,I713763,I713780,I713797,I713814,I713831,I713848,I713879,I713896,I713913,I713972,I714017,I714034,I714098,I714115,I714132,I714149,I714180,I714211,I714228,I714245,I714262,I714279,I714310,I714341,I714358,I714375,I714392,I714409,I714426,I714457,I714474,I714491,I714550,I714595,I714612,I714676,I714693,I714710,I714727,I714758,I714789,I714806,I714823,I714840,I714857,I714888,I714919,I714936,I714953,I714970,I714987,I715004,I715035,I715052,I715069,I715128,I715173,I715190,I715254,I715271,I715288,I715305,I715336,I715367,I715384,I715401,I715418,I715435,I715466,I715497,I715514,I715531,I715548,I715565,I715582,I715613,I715630,I715647,I715706,I715751,I715768,I715832,I715849,I715866,I715883,I715914,I715945,I715962,I715979,I715996,I716013,I716044,I716075,I716092,I716109,I716126,I716143,I716160,I716191,I716208,I716225,I716284,I716329,I716346,I716410,I716427,I716444,I716461,I716492,I716523,I716540,I716557,I716574,I716591,I716622,I716653,I716670,I716687,I716704,I716721,I716738,I716769,I716786,I716803,I716862,I716907,I716924,I716988,I717005,I717022,I717039,I717070,I717101,I717118,I717135,I717152,I717169,I717200,I717231,I717248,I717265,I717282,I717299,I717316,I717347,I717364,I717381,I717440,I717485,I717502,I717566,I717583,I717600,I717617,I717648,I717679,I717696,I717713,I717730,I717747,I717778,I717809,I717826,I717843,I717860,I717877,I717894,I717925,I717942,I717959,I718018,I718063,I718080,I718144,I718161,I718178,I718195,I718226,I718257,I718274,I718291,I718308,I718325,I718356,I718387,I718404,I718421,I718438,I718455,I718472,I718503,I718520,I718537,I718596,I718641,I718658,I718722,I718739,I718756,I718773,I718804,I718835,I718852,I718869,I718886,I718903,I718934,I718965,I718982,I718999,I719016,I719033,I719050,I719081,I719098,I719115,I719174,I719219,I719236,I719300,I719317,I719334,I719351,I719382,I719413,I719430,I719447,I719464,I719481,I719512,I719543,I719560,I719577,I719594,I719611,I719628,I719659,I719676,I719693,I719752,I719797,I719814,I719878,I719895,I719912,I719929,I719960,I719991,I720008,I720025,I720042,I720059,I720090,I720121,I720138,I720155,I720172,I720189,I720206,I720237,I720254,I720271,I720330,I720375,I720392,I720456,I720473,I720490,I720507,I720538,I720569,I720586,I720603,I720620,I720637,I720668,I720699,I720716,I720733,I720750,I720767,I720784,I720815,I720832,I720849,I720908,I720953,I720970,I721034,I721051,I721068,I721085,I721116,I721147,I721164,I721181,I721198,I721215,I721246,I721277,I721294,I721311,I721328,I721345,I721362,I721393,I721410,I721427,I721486,I721531,I721548,I721612,I721629,I721646,I721663,I721694,I721725,I721742,I721759,I721776,I721793,I721824,I721855,I721872,I721889,I721906,I721923,I721940,I721971,I721988,I722005,I722064,I722109,I722126,I722190,I722207,I722224,I722241,I722272,I722303,I722320,I722337,I722354,I722371,I722402,I722433,I722450,I722467,I722484,I722501,I722518,I722549,I722566,I722583,I722642,I722687,I722704,I722768,I722785,I722802,I722819,I722850,I722881,I722898,I722915,I722932,I722949,I722980,I723011,I723028,I723045,I723062,I723079,I723096,I723127,I723144,I723161,I723220,I723265,I723282,I723346,I723363,I723380,I723397,I723428,I723459,I723476,I723493,I723510,I723527,I723558,I723589,I723606,I723623,I723640,I723657,I723674,I723705,I723722,I723739,I723798,I723843,I723860,I723924,I723941,I723958,I723975,I724006,I724037,I724054,I724071,I724088,I724105,I724136,I724167,I724184,I724201,I724218,I724235,I724252,I724283,I724300,I724317,I724376,I724421,I724438,I724502,I724519,I724536,I724553,I724584,I724615,I724632,I724649,I724666,I724683,I724714,I724745,I724762,I724779,I724796,I724813,I724830,I724861,I724878,I724895,I724954,I724999,I725016,I725080,I725097,I725114,I725131,I725162,I725193,I725210,I725227,I725244,I725261,I725292,I725323,I725340,I725357,I725374,I725391,I725408,I725439,I725456,I725473,I725532,I725577,I725594,I725658,I725675,I725692,I725709,I725740,I725771,I725788,I725805,I725822,I725839,I725870,I725901,I725918,I725935,I725952,I725969,I725986,I726017,I726034,I726051,I726110,I726155,I726172,I726236,I726253,I726270,I726287,I726318,I726349,I726366,I726383,I726400,I726417,I726448,I726479,I726496,I726513,I726530,I726547,I726564,I726595,I726612,I726629,I726688,I726733,I726750,I726814,I726831,I726848,I726865,I726896,I726927,I726944,I726961,I726978,I726995,I727026,I727057,I727074,I727091,I727108,I727125,I727142,I727173,I727190,I727207,I727266,I727311,I727328,I727392,I727409,I727426,I727443,I727474,I727505,I727522,I727539,I727556,I727573,I727604,I727635,I727652,I727669,I727686,I727703,I727720,I727751,I727768,I727785,I727844,I727889,I727906;
not I_0 (I2750,I2709);
nand I_1 (I2767,I109204,I109207);
and I_2 (I2784,I2767,I109189);
DFFARX1 I_3  ( .D(I2784), .CLK(I2702), .RSTB(I2750), .Q(I2801) );
not I_4 (I2818,I2801);
nor I_5 (I2835,I109186,I109207);
or I_6 (I2733,I2835,I2801);
not I_7 (I2721,I2835);
DFFARX1 I_8  ( .D(I109210), .CLK(I2702), .RSTB(I2750), .Q(I2880) );
nor I_9 (I2897,I2880,I2835);
nand I_10 (I2914,I109195,I109201);
and I_11 (I2931,I2914,I109213);
DFFARX1 I_12  ( .D(I2931), .CLK(I2702), .RSTB(I2750), .Q(I2948) );
nor I_13 (I2730,I2948,I2801);
not I_14 (I2979,I2948);
nor I_15 (I2996,I2880,I2979);
DFFARX1 I_16  ( .D(I109192), .CLK(I2702), .RSTB(I2750), .Q(I3013) );
and I_17 (I3030,I3013,I109183);
or I_18 (I2739,I3030,I2835);
nand I_19 (I2718,I3030,I2996);
DFFARX1 I_20  ( .D(I109198), .CLK(I2702), .RSTB(I2750), .Q(I3075) );
and I_21 (I3092,I3075,I2818);
nor I_22 (I2736,I3030,I3092);
nor I_23 (I3123,I3075,I2880);
DFFARX1 I_24  ( .D(I3123), .CLK(I2702), .RSTB(I2750), .Q(I2727) );
nor I_25 (I2742,I3075,I2801);
not I_26 (I3168,I3075);
nor I_27 (I3185,I2948,I3168);
and I_28 (I3202,I2835,I3185);
or I_29 (I3219,I3030,I3202);
DFFARX1 I_30  ( .D(I3219), .CLK(I2702), .RSTB(I2750), .Q(I2715) );
nand I_31 (I2724,I3075,I2897);
nand I_32 (I2712,I3075,I2979);
not I_33 (I3311,I2709);
nand I_34 (I3328,I554212,I554215);
and I_35 (I3345,I3328,I554227);
DFFARX1 I_36  ( .D(I3345), .CLK(I2702), .RSTB(I3311), .Q(I3362) );
not I_37 (I3379,I3362);
nor I_38 (I3396,I554221,I554215);
or I_39 (I3294,I3396,I3362);
not I_40 (I3282,I3396);
DFFARX1 I_41  ( .D(I554224), .CLK(I2702), .RSTB(I3311), .Q(I3441) );
nor I_42 (I3458,I3441,I3396);
nand I_43 (I3475,I554218,I554236);
and I_44 (I3492,I3475,I554239);
DFFARX1 I_45  ( .D(I3492), .CLK(I2702), .RSTB(I3311), .Q(I3509) );
nor I_46 (I3291,I3509,I3362);
not I_47 (I3540,I3509);
nor I_48 (I3557,I3441,I3540);
DFFARX1 I_49  ( .D(I554209), .CLK(I2702), .RSTB(I3311), .Q(I3574) );
and I_50 (I3591,I3574,I554230);
or I_51 (I3300,I3591,I3396);
nand I_52 (I3279,I3591,I3557);
DFFARX1 I_53  ( .D(I554233), .CLK(I2702), .RSTB(I3311), .Q(I3636) );
and I_54 (I3653,I3636,I3379);
nor I_55 (I3297,I3591,I3653);
nor I_56 (I3684,I3636,I3441);
DFFARX1 I_57  ( .D(I3684), .CLK(I2702), .RSTB(I3311), .Q(I3288) );
nor I_58 (I3303,I3636,I3362);
not I_59 (I3729,I3636);
nor I_60 (I3746,I3509,I3729);
and I_61 (I3763,I3396,I3746);
or I_62 (I3780,I3591,I3763);
DFFARX1 I_63  ( .D(I3780), .CLK(I2702), .RSTB(I3311), .Q(I3276) );
nand I_64 (I3285,I3636,I3458);
nand I_65 (I3273,I3636,I3540);
not I_66 (I3872,I2709);
nand I_67 (I3889,I484147,I484144);
and I_68 (I3906,I3889,I484138);
DFFARX1 I_69  ( .D(I3906), .CLK(I2702), .RSTB(I3872), .Q(I3923) );
not I_70 (I3940,I3923);
nor I_71 (I3957,I484150,I484144);
or I_72 (I3855,I3957,I3923);
not I_73 (I3843,I3957);
DFFARX1 I_74  ( .D(I484162), .CLK(I2702), .RSTB(I3872), .Q(I4002) );
nor I_75 (I4019,I4002,I3957);
nand I_76 (I4036,I484153,I484135);
and I_77 (I4053,I4036,I484165);
DFFARX1 I_78  ( .D(I4053), .CLK(I2702), .RSTB(I3872), .Q(I4070) );
nor I_79 (I3852,I4070,I3923);
not I_80 (I4101,I4070);
nor I_81 (I4118,I4002,I4101);
DFFARX1 I_82  ( .D(I484141), .CLK(I2702), .RSTB(I3872), .Q(I4135) );
and I_83 (I4152,I4135,I484159);
or I_84 (I3861,I4152,I3957);
nand I_85 (I3840,I4152,I4118);
DFFARX1 I_86  ( .D(I484156), .CLK(I2702), .RSTB(I3872), .Q(I4197) );
and I_87 (I4214,I4197,I3940);
nor I_88 (I3858,I4152,I4214);
nor I_89 (I4245,I4197,I4002);
DFFARX1 I_90  ( .D(I4245), .CLK(I2702), .RSTB(I3872), .Q(I3849) );
nor I_91 (I3864,I4197,I3923);
not I_92 (I4290,I4197);
nor I_93 (I4307,I4070,I4290);
and I_94 (I4324,I3957,I4307);
or I_95 (I4341,I4152,I4324);
DFFARX1 I_96  ( .D(I4341), .CLK(I2702), .RSTB(I3872), .Q(I3837) );
nand I_97 (I3846,I4197,I4019);
nand I_98 (I3834,I4197,I4101);
not I_99 (I4433,I2709);
nand I_100 (I4450,I199224,I199221);
and I_101 (I4467,I4450,I199218);
DFFARX1 I_102  ( .D(I4467), .CLK(I2702), .RSTB(I4433), .Q(I4484) );
not I_103 (I4501,I4484);
nor I_104 (I4518,I199242,I199221);
or I_105 (I4416,I4518,I4484);
not I_106 (I4404,I4518);
DFFARX1 I_107  ( .D(I199236), .CLK(I2702), .RSTB(I4433), .Q(I4563) );
nor I_108 (I4580,I4563,I4518);
nand I_109 (I4597,I199215,I199227);
and I_110 (I4614,I4597,I199230);
DFFARX1 I_111  ( .D(I4614), .CLK(I2702), .RSTB(I4433), .Q(I4631) );
nor I_112 (I4413,I4631,I4484);
not I_113 (I4662,I4631);
nor I_114 (I4679,I4563,I4662);
DFFARX1 I_115  ( .D(I199239), .CLK(I2702), .RSTB(I4433), .Q(I4696) );
and I_116 (I4713,I4696,I199245);
or I_117 (I4422,I4713,I4518);
nand I_118 (I4401,I4713,I4679);
DFFARX1 I_119  ( .D(I199233), .CLK(I2702), .RSTB(I4433), .Q(I4758) );
and I_120 (I4775,I4758,I4501);
nor I_121 (I4419,I4713,I4775);
nor I_122 (I4806,I4758,I4563);
DFFARX1 I_123  ( .D(I4806), .CLK(I2702), .RSTB(I4433), .Q(I4410) );
nor I_124 (I4425,I4758,I4484);
not I_125 (I4851,I4758);
nor I_126 (I4868,I4631,I4851);
and I_127 (I4885,I4518,I4868);
or I_128 (I4902,I4713,I4885);
DFFARX1 I_129  ( .D(I4902), .CLK(I2702), .RSTB(I4433), .Q(I4398) );
nand I_130 (I4407,I4758,I4580);
nand I_131 (I4395,I4758,I4662);
not I_132 (I4994,I2709);
nand I_133 (I5011,I386143,I386134);
and I_134 (I5028,I5011,I386137);
DFFARX1 I_135  ( .D(I5028), .CLK(I2702), .RSTB(I4994), .Q(I5045) );
not I_136 (I5062,I5045);
nor I_137 (I5079,I386113,I386134);
or I_138 (I4977,I5079,I5045);
not I_139 (I4965,I5079);
DFFARX1 I_140  ( .D(I386128), .CLK(I2702), .RSTB(I4994), .Q(I5124) );
nor I_141 (I5141,I5124,I5079);
nand I_142 (I5158,I386116,I386131);
and I_143 (I5175,I5158,I386125);
DFFARX1 I_144  ( .D(I5175), .CLK(I2702), .RSTB(I4994), .Q(I5192) );
nor I_145 (I4974,I5192,I5045);
not I_146 (I5223,I5192);
nor I_147 (I5240,I5124,I5223);
DFFARX1 I_148  ( .D(I386140), .CLK(I2702), .RSTB(I4994), .Q(I5257) );
and I_149 (I5274,I5257,I386119);
or I_150 (I4983,I5274,I5079);
nand I_151 (I4962,I5274,I5240);
DFFARX1 I_152  ( .D(I386122), .CLK(I2702), .RSTB(I4994), .Q(I5319) );
and I_153 (I5336,I5319,I5062);
nor I_154 (I4980,I5274,I5336);
nor I_155 (I5367,I5319,I5124);
DFFARX1 I_156  ( .D(I5367), .CLK(I2702), .RSTB(I4994), .Q(I4971) );
nor I_157 (I4986,I5319,I5045);
not I_158 (I5412,I5319);
nor I_159 (I5429,I5192,I5412);
and I_160 (I5446,I5079,I5429);
or I_161 (I5463,I5274,I5446);
DFFARX1 I_162  ( .D(I5463), .CLK(I2702), .RSTB(I4994), .Q(I4959) );
nand I_163 (I4968,I5319,I5141);
nand I_164 (I4956,I5319,I5223);
not I_165 (I5555,I2709);
nand I_166 (I5572,I282114,I282105);
and I_167 (I5589,I5572,I282120);
DFFARX1 I_168  ( .D(I5589), .CLK(I2702), .RSTB(I5555), .Q(I5606) );
not I_169 (I5623,I5606);
nor I_170 (I5640,I282090,I282105);
or I_171 (I5538,I5640,I5606);
not I_172 (I5526,I5640);
DFFARX1 I_173  ( .D(I282093), .CLK(I2702), .RSTB(I5555), .Q(I5685) );
nor I_174 (I5702,I5685,I5640);
nand I_175 (I5719,I282111,I282108);
and I_176 (I5736,I5719,I282096);
DFFARX1 I_177  ( .D(I5736), .CLK(I2702), .RSTB(I5555), .Q(I5753) );
nor I_178 (I5535,I5753,I5606);
not I_179 (I5784,I5753);
nor I_180 (I5801,I5685,I5784);
DFFARX1 I_181  ( .D(I282117), .CLK(I2702), .RSTB(I5555), .Q(I5818) );
and I_182 (I5835,I5818,I282102);
or I_183 (I5544,I5835,I5640);
nand I_184 (I5523,I5835,I5801);
DFFARX1 I_185  ( .D(I282099), .CLK(I2702), .RSTB(I5555), .Q(I5880) );
and I_186 (I5897,I5880,I5623);
nor I_187 (I5541,I5835,I5897);
nor I_188 (I5928,I5880,I5685);
DFFARX1 I_189  ( .D(I5928), .CLK(I2702), .RSTB(I5555), .Q(I5532) );
nor I_190 (I5547,I5880,I5606);
not I_191 (I5973,I5880);
nor I_192 (I5990,I5753,I5973);
and I_193 (I6007,I5640,I5990);
or I_194 (I6024,I5835,I6007);
DFFARX1 I_195  ( .D(I6024), .CLK(I2702), .RSTB(I5555), .Q(I5520) );
nand I_196 (I5529,I5880,I5702);
nand I_197 (I5517,I5880,I5784);
not I_198 (I6116,I2709);
nand I_199 (I6133,I74966,I74969);
and I_200 (I6150,I6133,I74951);
DFFARX1 I_201  ( .D(I6150), .CLK(I2702), .RSTB(I6116), .Q(I6167) );
not I_202 (I6184,I6167);
nor I_203 (I6201,I74948,I74969);
or I_204 (I6099,I6201,I6167);
not I_205 (I6087,I6201);
DFFARX1 I_206  ( .D(I74972), .CLK(I2702), .RSTB(I6116), .Q(I6246) );
nor I_207 (I6263,I6246,I6201);
nand I_208 (I6280,I74957,I74963);
and I_209 (I6297,I6280,I74975);
DFFARX1 I_210  ( .D(I6297), .CLK(I2702), .RSTB(I6116), .Q(I6314) );
nor I_211 (I6096,I6314,I6167);
not I_212 (I6345,I6314);
nor I_213 (I6362,I6246,I6345);
DFFARX1 I_214  ( .D(I74954), .CLK(I2702), .RSTB(I6116), .Q(I6379) );
and I_215 (I6396,I6379,I74945);
or I_216 (I6105,I6396,I6201);
nand I_217 (I6084,I6396,I6362);
DFFARX1 I_218  ( .D(I74960), .CLK(I2702), .RSTB(I6116), .Q(I6441) );
and I_219 (I6458,I6441,I6184);
nor I_220 (I6102,I6396,I6458);
nor I_221 (I6489,I6441,I6246);
DFFARX1 I_222  ( .D(I6489), .CLK(I2702), .RSTB(I6116), .Q(I6093) );
nor I_223 (I6108,I6441,I6167);
not I_224 (I6534,I6441);
nor I_225 (I6551,I6314,I6534);
and I_226 (I6568,I6201,I6551);
or I_227 (I6585,I6396,I6568);
DFFARX1 I_228  ( .D(I6585), .CLK(I2702), .RSTB(I6116), .Q(I6081) );
nand I_229 (I6090,I6441,I6263);
nand I_230 (I6078,I6441,I6345);
not I_231 (I6677,I2709);
nand I_232 (I6694,I621852,I621855);
and I_233 (I6711,I6694,I621861);
DFFARX1 I_234  ( .D(I6711), .CLK(I2702), .RSTB(I6677), .Q(I6728) );
not I_235 (I6745,I6728);
nor I_236 (I6762,I621873,I621855);
or I_237 (I6660,I6762,I6728);
not I_238 (I6648,I6762);
DFFARX1 I_239  ( .D(I621882), .CLK(I2702), .RSTB(I6677), .Q(I6807) );
nor I_240 (I6824,I6807,I6762);
nand I_241 (I6841,I621870,I621867);
and I_242 (I6858,I6841,I621879);
DFFARX1 I_243  ( .D(I6858), .CLK(I2702), .RSTB(I6677), .Q(I6875) );
nor I_244 (I6657,I6875,I6728);
not I_245 (I6906,I6875);
nor I_246 (I6923,I6807,I6906);
DFFARX1 I_247  ( .D(I621876), .CLK(I2702), .RSTB(I6677), .Q(I6940) );
and I_248 (I6957,I6940,I621864);
or I_249 (I6666,I6957,I6762);
nand I_250 (I6645,I6957,I6923);
DFFARX1 I_251  ( .D(I621858), .CLK(I2702), .RSTB(I6677), .Q(I7002) );
and I_252 (I7019,I7002,I6745);
nor I_253 (I6663,I6957,I7019);
nor I_254 (I7050,I7002,I6807);
DFFARX1 I_255  ( .D(I7050), .CLK(I2702), .RSTB(I6677), .Q(I6654) );
nor I_256 (I6669,I7002,I6728);
not I_257 (I7095,I7002);
nor I_258 (I7112,I6875,I7095);
and I_259 (I7129,I6762,I7112);
or I_260 (I7146,I6957,I7129);
DFFARX1 I_261  ( .D(I7146), .CLK(I2702), .RSTB(I6677), .Q(I6642) );
nand I_262 (I6651,I7002,I6824);
nand I_263 (I6639,I7002,I6906);
not I_264 (I7238,I2709);
nand I_265 (I7255,I432705,I432702);
and I_266 (I7272,I7255,I432696);
DFFARX1 I_267  ( .D(I7272), .CLK(I2702), .RSTB(I7238), .Q(I7289) );
not I_268 (I7306,I7289);
nor I_269 (I7323,I432708,I432702);
or I_270 (I7221,I7323,I7289);
not I_271 (I7209,I7323);
DFFARX1 I_272  ( .D(I432720), .CLK(I2702), .RSTB(I7238), .Q(I7368) );
nor I_273 (I7385,I7368,I7323);
nand I_274 (I7402,I432711,I432693);
and I_275 (I7419,I7402,I432723);
DFFARX1 I_276  ( .D(I7419), .CLK(I2702), .RSTB(I7238), .Q(I7436) );
nor I_277 (I7218,I7436,I7289);
not I_278 (I7467,I7436);
nor I_279 (I7484,I7368,I7467);
DFFARX1 I_280  ( .D(I432699), .CLK(I2702), .RSTB(I7238), .Q(I7501) );
and I_281 (I7518,I7501,I432717);
or I_282 (I7227,I7518,I7323);
nand I_283 (I7206,I7518,I7484);
DFFARX1 I_284  ( .D(I432714), .CLK(I2702), .RSTB(I7238), .Q(I7563) );
and I_285 (I7580,I7563,I7306);
nor I_286 (I7224,I7518,I7580);
nor I_287 (I7611,I7563,I7368);
DFFARX1 I_288  ( .D(I7611), .CLK(I2702), .RSTB(I7238), .Q(I7215) );
nor I_289 (I7230,I7563,I7289);
not I_290 (I7656,I7563);
nor I_291 (I7673,I7436,I7656);
and I_292 (I7690,I7323,I7673);
or I_293 (I7707,I7518,I7690);
DFFARX1 I_294  ( .D(I7707), .CLK(I2702), .RSTB(I7238), .Q(I7203) );
nand I_295 (I7212,I7563,I7385);
nand I_296 (I7200,I7563,I7467);
not I_297 (I7799,I2709);
nand I_298 (I7816,I586955,I586943);
and I_299 (I7833,I7816,I586940);
DFFARX1 I_300  ( .D(I7833), .CLK(I2702), .RSTB(I7799), .Q(I7850) );
not I_301 (I7867,I7850);
nor I_302 (I7884,I586961,I586943);
or I_303 (I7782,I7884,I7850);
not I_304 (I7770,I7884);
DFFARX1 I_305  ( .D(I586964), .CLK(I2702), .RSTB(I7799), .Q(I7929) );
nor I_306 (I7946,I7929,I7884);
nand I_307 (I7963,I586934,I586952);
and I_308 (I7980,I7963,I586949);
DFFARX1 I_309  ( .D(I7980), .CLK(I2702), .RSTB(I7799), .Q(I7997) );
nor I_310 (I7779,I7997,I7850);
not I_311 (I8028,I7997);
nor I_312 (I8045,I7929,I8028);
DFFARX1 I_313  ( .D(I586958), .CLK(I2702), .RSTB(I7799), .Q(I8062) );
and I_314 (I8079,I8062,I586946);
or I_315 (I7788,I8079,I7884);
nand I_316 (I7767,I8079,I8045);
DFFARX1 I_317  ( .D(I586937), .CLK(I2702), .RSTB(I7799), .Q(I8124) );
and I_318 (I8141,I8124,I7867);
nor I_319 (I7785,I8079,I8141);
nor I_320 (I8172,I8124,I7929);
DFFARX1 I_321  ( .D(I8172), .CLK(I2702), .RSTB(I7799), .Q(I7776) );
nor I_322 (I7791,I8124,I7850);
not I_323 (I8217,I8124);
nor I_324 (I8234,I7997,I8217);
and I_325 (I8251,I7884,I8234);
or I_326 (I8268,I8079,I8251);
DFFARX1 I_327  ( .D(I8268), .CLK(I2702), .RSTB(I7799), .Q(I7764) );
nand I_328 (I7773,I8124,I7946);
nand I_329 (I7761,I8124,I8028);
not I_330 (I8360,I2709);
nand I_331 (I8377,I624997,I625000);
and I_332 (I8394,I8377,I625006);
DFFARX1 I_333  ( .D(I8394), .CLK(I2702), .RSTB(I8360), .Q(I8411) );
not I_334 (I8428,I8411);
nor I_335 (I8445,I625018,I625000);
or I_336 (I8343,I8445,I8411);
not I_337 (I8331,I8445);
DFFARX1 I_338  ( .D(I625027), .CLK(I2702), .RSTB(I8360), .Q(I8490) );
nor I_339 (I8507,I8490,I8445);
nand I_340 (I8524,I625015,I625012);
and I_341 (I8541,I8524,I625024);
DFFARX1 I_342  ( .D(I8541), .CLK(I2702), .RSTB(I8360), .Q(I8558) );
nor I_343 (I8340,I8558,I8411);
not I_344 (I8589,I8558);
nor I_345 (I8606,I8490,I8589);
DFFARX1 I_346  ( .D(I625021), .CLK(I2702), .RSTB(I8360), .Q(I8623) );
and I_347 (I8640,I8623,I625009);
or I_348 (I8349,I8640,I8445);
nand I_349 (I8328,I8640,I8606);
DFFARX1 I_350  ( .D(I625003), .CLK(I2702), .RSTB(I8360), .Q(I8685) );
and I_351 (I8702,I8685,I8428);
nor I_352 (I8346,I8640,I8702);
nor I_353 (I8733,I8685,I8490);
DFFARX1 I_354  ( .D(I8733), .CLK(I2702), .RSTB(I8360), .Q(I8337) );
nor I_355 (I8352,I8685,I8411);
not I_356 (I8778,I8685);
nor I_357 (I8795,I8558,I8778);
and I_358 (I8812,I8445,I8795);
or I_359 (I8829,I8640,I8812);
DFFARX1 I_360  ( .D(I8829), .CLK(I2702), .RSTB(I8360), .Q(I8325) );
nand I_361 (I8334,I8685,I8507);
nand I_362 (I8322,I8685,I8589);
not I_363 (I8921,I2709);
nand I_364 (I8938,I142206,I142203);
and I_365 (I8955,I8938,I142200);
DFFARX1 I_366  ( .D(I8955), .CLK(I2702), .RSTB(I8921), .Q(I8972) );
not I_367 (I8989,I8972);
nor I_368 (I9006,I142224,I142203);
or I_369 (I8904,I9006,I8972);
not I_370 (I8892,I9006);
DFFARX1 I_371  ( .D(I142218), .CLK(I2702), .RSTB(I8921), .Q(I9051) );
nor I_372 (I9068,I9051,I9006);
nand I_373 (I9085,I142197,I142209);
and I_374 (I9102,I9085,I142212);
DFFARX1 I_375  ( .D(I9102), .CLK(I2702), .RSTB(I8921), .Q(I9119) );
nor I_376 (I8901,I9119,I8972);
not I_377 (I9150,I9119);
nor I_378 (I9167,I9051,I9150);
DFFARX1 I_379  ( .D(I142221), .CLK(I2702), .RSTB(I8921), .Q(I9184) );
and I_380 (I9201,I9184,I142227);
or I_381 (I8910,I9201,I9006);
nand I_382 (I8889,I9201,I9167);
DFFARX1 I_383  ( .D(I142215), .CLK(I2702), .RSTB(I8921), .Q(I9246) );
and I_384 (I9263,I9246,I8989);
nor I_385 (I8907,I9201,I9263);
nor I_386 (I9294,I9246,I9051);
DFFARX1 I_387  ( .D(I9294), .CLK(I2702), .RSTB(I8921), .Q(I8898) );
nor I_388 (I8913,I9246,I8972);
not I_389 (I9339,I9246);
nor I_390 (I9356,I9119,I9339);
and I_391 (I9373,I9006,I9356);
or I_392 (I9390,I9201,I9373);
DFFARX1 I_393  ( .D(I9390), .CLK(I2702), .RSTB(I8921), .Q(I8886) );
nand I_394 (I8895,I9246,I9068);
nand I_395 (I8883,I9246,I9150);
not I_396 (I9482,I2709);
nand I_397 (I9499,I54294,I54297);
and I_398 (I9516,I9499,I54279);
DFFARX1 I_399  ( .D(I9516), .CLK(I2702), .RSTB(I9482), .Q(I9533) );
not I_400 (I9550,I9533);
nor I_401 (I9567,I54276,I54297);
or I_402 (I9465,I9567,I9533);
not I_403 (I9453,I9567);
DFFARX1 I_404  ( .D(I54300), .CLK(I2702), .RSTB(I9482), .Q(I9612) );
nor I_405 (I9629,I9612,I9567);
nand I_406 (I9646,I54285,I54291);
and I_407 (I9663,I9646,I54303);
DFFARX1 I_408  ( .D(I9663), .CLK(I2702), .RSTB(I9482), .Q(I9680) );
nor I_409 (I9462,I9680,I9533);
not I_410 (I9711,I9680);
nor I_411 (I9728,I9612,I9711);
DFFARX1 I_412  ( .D(I54282), .CLK(I2702), .RSTB(I9482), .Q(I9745) );
and I_413 (I9762,I9745,I54273);
or I_414 (I9471,I9762,I9567);
nand I_415 (I9450,I9762,I9728);
DFFARX1 I_416  ( .D(I54288), .CLK(I2702), .RSTB(I9482), .Q(I9807) );
and I_417 (I9824,I9807,I9550);
nor I_418 (I9468,I9762,I9824);
nor I_419 (I9855,I9807,I9612);
DFFARX1 I_420  ( .D(I9855), .CLK(I2702), .RSTB(I9482), .Q(I9459) );
nor I_421 (I9474,I9807,I9533);
not I_422 (I9900,I9807);
nor I_423 (I9917,I9680,I9900);
and I_424 (I9934,I9567,I9917);
or I_425 (I9951,I9762,I9934);
DFFARX1 I_426  ( .D(I9951), .CLK(I2702), .RSTB(I9482), .Q(I9447) );
nand I_427 (I9456,I9807,I9629);
nand I_428 (I9444,I9807,I9711);
not I_429 (I10043,I2709);
nand I_430 (I10060,I721005,I721026);
and I_431 (I10077,I10060,I721014);
DFFARX1 I_432  ( .D(I10077), .CLK(I2702), .RSTB(I10043), .Q(I10094) );
not I_433 (I10111,I10094);
nor I_434 (I10128,I721020,I721026);
or I_435 (I10026,I10128,I10094);
not I_436 (I10014,I10128);
DFFARX1 I_437  ( .D(I721008), .CLK(I2702), .RSTB(I10043), .Q(I10173) );
nor I_438 (I10190,I10173,I10128);
nand I_439 (I10207,I720999,I721017);
and I_440 (I10224,I10207,I721011);
DFFARX1 I_441  ( .D(I10224), .CLK(I2702), .RSTB(I10043), .Q(I10241) );
nor I_442 (I10023,I10241,I10094);
not I_443 (I10272,I10241);
nor I_444 (I10289,I10173,I10272);
DFFARX1 I_445  ( .D(I721023), .CLK(I2702), .RSTB(I10043), .Q(I10306) );
and I_446 (I10323,I10306,I720996);
or I_447 (I10032,I10323,I10128);
nand I_448 (I10011,I10323,I10289);
DFFARX1 I_449  ( .D(I721002), .CLK(I2702), .RSTB(I10043), .Q(I10368) );
and I_450 (I10385,I10368,I10111);
nor I_451 (I10029,I10323,I10385);
nor I_452 (I10416,I10368,I10173);
DFFARX1 I_453  ( .D(I10416), .CLK(I2702), .RSTB(I10043), .Q(I10020) );
nor I_454 (I10035,I10368,I10094);
not I_455 (I10461,I10368);
nor I_456 (I10478,I10241,I10461);
and I_457 (I10495,I10128,I10478);
or I_458 (I10512,I10323,I10495);
DFFARX1 I_459  ( .D(I10512), .CLK(I2702), .RSTB(I10043), .Q(I10008) );
nand I_460 (I10017,I10368,I10190);
nand I_461 (I10005,I10368,I10272);
not I_462 (I10604,I2709);
nand I_463 (I10621,I497935,I497929);
and I_464 (I10638,I10621,I497920);
DFFARX1 I_465  ( .D(I10638), .CLK(I2702), .RSTB(I10604), .Q(I10655) );
not I_466 (I10672,I10655);
nor I_467 (I10689,I497911,I497929);
or I_468 (I10587,I10689,I10655);
not I_469 (I10575,I10689);
DFFARX1 I_470  ( .D(I497926), .CLK(I2702), .RSTB(I10604), .Q(I10734) );
nor I_471 (I10751,I10734,I10689);
nand I_472 (I10768,I497917,I497932);
and I_473 (I10785,I10768,I497914);
DFFARX1 I_474  ( .D(I10785), .CLK(I2702), .RSTB(I10604), .Q(I10802) );
nor I_475 (I10584,I10802,I10655);
not I_476 (I10833,I10802);
nor I_477 (I10850,I10734,I10833);
DFFARX1 I_478  ( .D(I497923), .CLK(I2702), .RSTB(I10604), .Q(I10867) );
and I_479 (I10884,I10867,I497905);
or I_480 (I10593,I10884,I10689);
nand I_481 (I10572,I10884,I10850);
DFFARX1 I_482  ( .D(I497908), .CLK(I2702), .RSTB(I10604), .Q(I10929) );
and I_483 (I10946,I10929,I10672);
nor I_484 (I10590,I10884,I10946);
nor I_485 (I10977,I10929,I10734);
DFFARX1 I_486  ( .D(I10977), .CLK(I2702), .RSTB(I10604), .Q(I10581) );
nor I_487 (I10596,I10929,I10655);
not I_488 (I11022,I10929);
nor I_489 (I11039,I10802,I11022);
and I_490 (I11056,I10689,I11039);
or I_491 (I11073,I10884,I11056);
DFFARX1 I_492  ( .D(I11073), .CLK(I2702), .RSTB(I10604), .Q(I10569) );
nand I_493 (I10578,I10929,I10751);
nand I_494 (I10566,I10929,I10833);
not I_495 (I11165,I2709);
nand I_496 (I11182,I321894,I321885);
and I_497 (I11199,I11182,I321900);
DFFARX1 I_498  ( .D(I11199), .CLK(I2702), .RSTB(I11165), .Q(I11216) );
not I_499 (I11233,I11216);
nor I_500 (I11250,I321870,I321885);
or I_501 (I11148,I11250,I11216);
not I_502 (I11136,I11250);
DFFARX1 I_503  ( .D(I321873), .CLK(I2702), .RSTB(I11165), .Q(I11295) );
nor I_504 (I11312,I11295,I11250);
nand I_505 (I11329,I321891,I321888);
and I_506 (I11346,I11329,I321876);
DFFARX1 I_507  ( .D(I11346), .CLK(I2702), .RSTB(I11165), .Q(I11363) );
nor I_508 (I11145,I11363,I11216);
not I_509 (I11394,I11363);
nor I_510 (I11411,I11295,I11394);
DFFARX1 I_511  ( .D(I321897), .CLK(I2702), .RSTB(I11165), .Q(I11428) );
and I_512 (I11445,I11428,I321882);
or I_513 (I11154,I11445,I11250);
nand I_514 (I11133,I11445,I11411);
DFFARX1 I_515  ( .D(I321879), .CLK(I2702), .RSTB(I11165), .Q(I11490) );
and I_516 (I11507,I11490,I11233);
nor I_517 (I11151,I11445,I11507);
nor I_518 (I11538,I11490,I11295);
DFFARX1 I_519  ( .D(I11538), .CLK(I2702), .RSTB(I11165), .Q(I11142) );
nor I_520 (I11157,I11490,I11216);
not I_521 (I11583,I11490);
nor I_522 (I11600,I11363,I11583);
and I_523 (I11617,I11250,I11600);
or I_524 (I11634,I11445,I11617);
DFFARX1 I_525  ( .D(I11634), .CLK(I2702), .RSTB(I11165), .Q(I11130) );
nand I_526 (I11139,I11490,I11312);
nand I_527 (I11127,I11490,I11394);
not I_528 (I11726,I2709);
nand I_529 (I11743,I689793,I689814);
and I_530 (I11760,I11743,I689802);
DFFARX1 I_531  ( .D(I11760), .CLK(I2702), .RSTB(I11726), .Q(I11777) );
not I_532 (I11794,I11777);
nor I_533 (I11811,I689808,I689814);
or I_534 (I11709,I11811,I11777);
not I_535 (I11697,I11811);
DFFARX1 I_536  ( .D(I689796), .CLK(I2702), .RSTB(I11726), .Q(I11856) );
nor I_537 (I11873,I11856,I11811);
nand I_538 (I11890,I689787,I689805);
and I_539 (I11907,I11890,I689799);
DFFARX1 I_540  ( .D(I11907), .CLK(I2702), .RSTB(I11726), .Q(I11924) );
nor I_541 (I11706,I11924,I11777);
not I_542 (I11955,I11924);
nor I_543 (I11972,I11856,I11955);
DFFARX1 I_544  ( .D(I689811), .CLK(I2702), .RSTB(I11726), .Q(I11989) );
and I_545 (I12006,I11989,I689784);
or I_546 (I11715,I12006,I11811);
nand I_547 (I11694,I12006,I11972);
DFFARX1 I_548  ( .D(I689790), .CLK(I2702), .RSTB(I11726), .Q(I12051) );
and I_549 (I12068,I12051,I11794);
nor I_550 (I11712,I12006,I12068);
nor I_551 (I12099,I12051,I11856);
DFFARX1 I_552  ( .D(I12099), .CLK(I2702), .RSTB(I11726), .Q(I11703) );
nor I_553 (I11718,I12051,I11777);
not I_554 (I12144,I12051);
nor I_555 (I12161,I11924,I12144);
and I_556 (I12178,I11811,I12161);
or I_557 (I12195,I12006,I12178);
DFFARX1 I_558  ( .D(I12195), .CLK(I2702), .RSTB(I11726), .Q(I11691) );
nand I_559 (I11700,I12051,I11873);
nand I_560 (I11688,I12051,I11955);
not I_561 (I12287,I2709);
nand I_562 (I12304,I227855,I227849);
and I_563 (I12321,I12304,I227843);
DFFARX1 I_564  ( .D(I12321), .CLK(I2702), .RSTB(I12287), .Q(I12338) );
not I_565 (I12355,I12338);
nor I_566 (I12372,I227870,I227849);
or I_567 (I12270,I12372,I12338);
not I_568 (I12258,I12372);
DFFARX1 I_569  ( .D(I227867), .CLK(I2702), .RSTB(I12287), .Q(I12417) );
nor I_570 (I12434,I12417,I12372);
nand I_571 (I12451,I227873,I227861);
and I_572 (I12468,I12451,I227858);
DFFARX1 I_573  ( .D(I12468), .CLK(I2702), .RSTB(I12287), .Q(I12485) );
nor I_574 (I12267,I12485,I12338);
not I_575 (I12516,I12485);
nor I_576 (I12533,I12417,I12516);
DFFARX1 I_577  ( .D(I227846), .CLK(I2702), .RSTB(I12287), .Q(I12550) );
and I_578 (I12567,I12550,I227864);
or I_579 (I12276,I12567,I12372);
nand I_580 (I12255,I12567,I12533);
DFFARX1 I_581  ( .D(I227852), .CLK(I2702), .RSTB(I12287), .Q(I12612) );
and I_582 (I12629,I12612,I12355);
nor I_583 (I12273,I12567,I12629);
nor I_584 (I12660,I12612,I12417);
DFFARX1 I_585  ( .D(I12660), .CLK(I2702), .RSTB(I12287), .Q(I12264) );
nor I_586 (I12279,I12612,I12338);
not I_587 (I12705,I12612);
nor I_588 (I12722,I12485,I12705);
and I_589 (I12739,I12372,I12722);
or I_590 (I12756,I12567,I12739);
DFFARX1 I_591  ( .D(I12756), .CLK(I2702), .RSTB(I12287), .Q(I12252) );
nand I_592 (I12261,I12612,I12434);
nand I_593 (I12249,I12612,I12516);
not I_594 (I12848,I2709);
nand I_595 (I12865,I374515,I374506);
and I_596 (I12882,I12865,I374509);
DFFARX1 I_597  ( .D(I12882), .CLK(I2702), .RSTB(I12848), .Q(I12899) );
not I_598 (I12916,I12899);
nor I_599 (I12933,I374485,I374506);
or I_600 (I12831,I12933,I12899);
not I_601 (I12819,I12933);
DFFARX1 I_602  ( .D(I374500), .CLK(I2702), .RSTB(I12848), .Q(I12978) );
nor I_603 (I12995,I12978,I12933);
nand I_604 (I13012,I374488,I374503);
and I_605 (I13029,I13012,I374497);
DFFARX1 I_606  ( .D(I13029), .CLK(I2702), .RSTB(I12848), .Q(I13046) );
nor I_607 (I12828,I13046,I12899);
not I_608 (I13077,I13046);
nor I_609 (I13094,I12978,I13077);
DFFARX1 I_610  ( .D(I374512), .CLK(I2702), .RSTB(I12848), .Q(I13111) );
and I_611 (I13128,I13111,I374491);
or I_612 (I12837,I13128,I12933);
nand I_613 (I12816,I13128,I13094);
DFFARX1 I_614  ( .D(I374494), .CLK(I2702), .RSTB(I12848), .Q(I13173) );
and I_615 (I13190,I13173,I12916);
nor I_616 (I12834,I13128,I13190);
nor I_617 (I13221,I13173,I12978);
DFFARX1 I_618  ( .D(I13221), .CLK(I2702), .RSTB(I12848), .Q(I12825) );
nor I_619 (I12840,I13173,I12899);
not I_620 (I13266,I13173);
nor I_621 (I13283,I13046,I13266);
and I_622 (I13300,I12933,I13283);
or I_623 (I13317,I13128,I13300);
DFFARX1 I_624  ( .D(I13317), .CLK(I2702), .RSTB(I12848), .Q(I12813) );
nand I_625 (I12822,I13173,I12995);
nand I_626 (I12810,I13173,I13077);
not I_627 (I13409,I2709);
nand I_628 (I13426,I523867,I523870);
and I_629 (I13443,I13426,I523882);
DFFARX1 I_630  ( .D(I13443), .CLK(I2702), .RSTB(I13409), .Q(I13460) );
not I_631 (I13477,I13460);
nor I_632 (I13494,I523876,I523870);
or I_633 (I13392,I13494,I13460);
not I_634 (I13380,I13494);
DFFARX1 I_635  ( .D(I523879), .CLK(I2702), .RSTB(I13409), .Q(I13539) );
nor I_636 (I13556,I13539,I13494);
nand I_637 (I13573,I523873,I523891);
and I_638 (I13590,I13573,I523894);
DFFARX1 I_639  ( .D(I13590), .CLK(I2702), .RSTB(I13409), .Q(I13607) );
nor I_640 (I13389,I13607,I13460);
not I_641 (I13638,I13607);
nor I_642 (I13655,I13539,I13638);
DFFARX1 I_643  ( .D(I523864), .CLK(I2702), .RSTB(I13409), .Q(I13672) );
and I_644 (I13689,I13672,I523885);
or I_645 (I13398,I13689,I13494);
nand I_646 (I13377,I13689,I13655);
DFFARX1 I_647  ( .D(I523888), .CLK(I2702), .RSTB(I13409), .Q(I13734) );
and I_648 (I13751,I13734,I13477);
nor I_649 (I13395,I13689,I13751);
nor I_650 (I13782,I13734,I13539);
DFFARX1 I_651  ( .D(I13782), .CLK(I2702), .RSTB(I13409), .Q(I13386) );
nor I_652 (I13401,I13734,I13460);
not I_653 (I13827,I13734);
nor I_654 (I13844,I13607,I13827);
and I_655 (I13861,I13494,I13844);
or I_656 (I13878,I13689,I13861);
DFFARX1 I_657  ( .D(I13878), .CLK(I2702), .RSTB(I13409), .Q(I13374) );
nand I_658 (I13383,I13734,I13556);
nand I_659 (I13371,I13734,I13638);
not I_660 (I13970,I2709);
nand I_661 (I13987,I408753,I408744);
and I_662 (I14004,I13987,I408747);
DFFARX1 I_663  ( .D(I14004), .CLK(I2702), .RSTB(I13970), .Q(I14021) );
not I_664 (I14038,I14021);
nor I_665 (I14055,I408723,I408744);
or I_666 (I13953,I14055,I14021);
not I_667 (I13941,I14055);
DFFARX1 I_668  ( .D(I408738), .CLK(I2702), .RSTB(I13970), .Q(I14100) );
nor I_669 (I14117,I14100,I14055);
nand I_670 (I14134,I408726,I408741);
and I_671 (I14151,I14134,I408735);
DFFARX1 I_672  ( .D(I14151), .CLK(I2702), .RSTB(I13970), .Q(I14168) );
nor I_673 (I13950,I14168,I14021);
not I_674 (I14199,I14168);
nor I_675 (I14216,I14100,I14199);
DFFARX1 I_676  ( .D(I408750), .CLK(I2702), .RSTB(I13970), .Q(I14233) );
and I_677 (I14250,I14233,I408729);
or I_678 (I13959,I14250,I14055);
nand I_679 (I13938,I14250,I14216);
DFFARX1 I_680  ( .D(I408732), .CLK(I2702), .RSTB(I13970), .Q(I14295) );
and I_681 (I14312,I14295,I14038);
nor I_682 (I13956,I14250,I14312);
nor I_683 (I14343,I14295,I14100);
DFFARX1 I_684  ( .D(I14343), .CLK(I2702), .RSTB(I13970), .Q(I13947) );
nor I_685 (I13962,I14295,I14021);
not I_686 (I14388,I14295);
nor I_687 (I14405,I14168,I14388);
and I_688 (I14422,I14055,I14405);
or I_689 (I14439,I14250,I14422);
DFFARX1 I_690  ( .D(I14439), .CLK(I2702), .RSTB(I13970), .Q(I13935) );
nand I_691 (I13944,I14295,I14117);
nand I_692 (I13932,I14295,I14199);
not I_693 (I14531,I2709);
nand I_694 (I14548,I538147,I538150);
and I_695 (I14565,I14548,I538162);
DFFARX1 I_696  ( .D(I14565), .CLK(I2702), .RSTB(I14531), .Q(I14582) );
not I_697 (I14599,I14582);
nor I_698 (I14616,I538156,I538150);
or I_699 (I14514,I14616,I14582);
not I_700 (I14502,I14616);
DFFARX1 I_701  ( .D(I538159), .CLK(I2702), .RSTB(I14531), .Q(I14661) );
nor I_702 (I14678,I14661,I14616);
nand I_703 (I14695,I538153,I538171);
and I_704 (I14712,I14695,I538174);
DFFARX1 I_705  ( .D(I14712), .CLK(I2702), .RSTB(I14531), .Q(I14729) );
nor I_706 (I14511,I14729,I14582);
not I_707 (I14760,I14729);
nor I_708 (I14777,I14661,I14760);
DFFARX1 I_709  ( .D(I538144), .CLK(I2702), .RSTB(I14531), .Q(I14794) );
and I_710 (I14811,I14794,I538165);
or I_711 (I14520,I14811,I14616);
nand I_712 (I14499,I14811,I14777);
DFFARX1 I_713  ( .D(I538168), .CLK(I2702), .RSTB(I14531), .Q(I14856) );
and I_714 (I14873,I14856,I14599);
nor I_715 (I14517,I14811,I14873);
nor I_716 (I14904,I14856,I14661);
DFFARX1 I_717  ( .D(I14904), .CLK(I2702), .RSTB(I14531), .Q(I14508) );
nor I_718 (I14523,I14856,I14582);
not I_719 (I14949,I14856);
nor I_720 (I14966,I14729,I14949);
and I_721 (I14983,I14616,I14966);
or I_722 (I15000,I14811,I14983);
DFFARX1 I_723  ( .D(I15000), .CLK(I2702), .RSTB(I14531), .Q(I14496) );
nand I_724 (I14505,I14856,I14678);
nand I_725 (I14493,I14856,I14760);
not I_726 (I15092,I2709);
nand I_727 (I15109,I404877,I404868);
and I_728 (I15126,I15109,I404871);
DFFARX1 I_729  ( .D(I15126), .CLK(I2702), .RSTB(I15092), .Q(I15143) );
not I_730 (I15160,I15143);
nor I_731 (I15177,I404847,I404868);
or I_732 (I15075,I15177,I15143);
not I_733 (I15063,I15177);
DFFARX1 I_734  ( .D(I404862), .CLK(I2702), .RSTB(I15092), .Q(I15222) );
nor I_735 (I15239,I15222,I15177);
nand I_736 (I15256,I404850,I404865);
and I_737 (I15273,I15256,I404859);
DFFARX1 I_738  ( .D(I15273), .CLK(I2702), .RSTB(I15092), .Q(I15290) );
nor I_739 (I15072,I15290,I15143);
not I_740 (I15321,I15290);
nor I_741 (I15338,I15222,I15321);
DFFARX1 I_742  ( .D(I404874), .CLK(I2702), .RSTB(I15092), .Q(I15355) );
and I_743 (I15372,I15355,I404853);
or I_744 (I15081,I15372,I15177);
nand I_745 (I15060,I15372,I15338);
DFFARX1 I_746  ( .D(I404856), .CLK(I2702), .RSTB(I15092), .Q(I15417) );
and I_747 (I15434,I15417,I15160);
nor I_748 (I15078,I15372,I15434);
nor I_749 (I15465,I15417,I15222);
DFFARX1 I_750  ( .D(I15465), .CLK(I2702), .RSTB(I15092), .Q(I15069) );
nor I_751 (I15084,I15417,I15143);
not I_752 (I15510,I15417);
nor I_753 (I15527,I15290,I15510);
and I_754 (I15544,I15177,I15527);
or I_755 (I15561,I15372,I15544);
DFFARX1 I_756  ( .D(I15561), .CLK(I2702), .RSTB(I15092), .Q(I15057) );
nand I_757 (I15066,I15417,I15239);
nand I_758 (I15054,I15417,I15321);
not I_759 (I15653,I2709);
nand I_760 (I15670,I1447,I1207);
and I_761 (I15687,I15670,I2631);
DFFARX1 I_762  ( .D(I15687), .CLK(I2702), .RSTB(I15653), .Q(I15704) );
not I_763 (I15721,I15704);
nor I_764 (I15738,I1863,I1207);
or I_765 (I15636,I15738,I15704);
not I_766 (I15624,I15738);
DFFARX1 I_767  ( .D(I1679), .CLK(I2702), .RSTB(I15653), .Q(I15783) );
nor I_768 (I15800,I15783,I15738);
nand I_769 (I15817,I1463,I1535);
and I_770 (I15834,I15817,I2511);
DFFARX1 I_771  ( .D(I15834), .CLK(I2702), .RSTB(I15653), .Q(I15851) );
nor I_772 (I15633,I15851,I15704);
not I_773 (I15882,I15851);
nor I_774 (I15899,I15783,I15882);
DFFARX1 I_775  ( .D(I2039), .CLK(I2702), .RSTB(I15653), .Q(I15916) );
and I_776 (I15933,I15916,I1631);
or I_777 (I15642,I15933,I15738);
nand I_778 (I15621,I15933,I15899);
DFFARX1 I_779  ( .D(I2207), .CLK(I2702), .RSTB(I15653), .Q(I15978) );
and I_780 (I15995,I15978,I15721);
nor I_781 (I15639,I15933,I15995);
nor I_782 (I16026,I15978,I15783);
DFFARX1 I_783  ( .D(I16026), .CLK(I2702), .RSTB(I15653), .Q(I15630) );
nor I_784 (I15645,I15978,I15704);
not I_785 (I16071,I15978);
nor I_786 (I16088,I15851,I16071);
and I_787 (I16105,I15738,I16088);
or I_788 (I16122,I15933,I16105);
DFFARX1 I_789  ( .D(I16122), .CLK(I2702), .RSTB(I15653), .Q(I15618) );
nand I_790 (I15627,I15978,I15800);
nand I_791 (I15615,I15978,I15882);
not I_792 (I16214,I2709);
nand I_793 (I16231,I264213,I264204);
and I_794 (I16248,I16231,I264219);
DFFARX1 I_795  ( .D(I16248), .CLK(I2702), .RSTB(I16214), .Q(I16265) );
not I_796 (I16282,I16265);
nor I_797 (I16299,I264189,I264204);
or I_798 (I16197,I16299,I16265);
not I_799 (I16185,I16299);
DFFARX1 I_800  ( .D(I264192), .CLK(I2702), .RSTB(I16214), .Q(I16344) );
nor I_801 (I16361,I16344,I16299);
nand I_802 (I16378,I264210,I264207);
and I_803 (I16395,I16378,I264195);
DFFARX1 I_804  ( .D(I16395), .CLK(I2702), .RSTB(I16214), .Q(I16412) );
nor I_805 (I16194,I16412,I16265);
not I_806 (I16443,I16412);
nor I_807 (I16460,I16344,I16443);
DFFARX1 I_808  ( .D(I264216), .CLK(I2702), .RSTB(I16214), .Q(I16477) );
and I_809 (I16494,I16477,I264201);
or I_810 (I16203,I16494,I16299);
nand I_811 (I16182,I16494,I16460);
DFFARX1 I_812  ( .D(I264198), .CLK(I2702), .RSTB(I16214), .Q(I16539) );
and I_813 (I16556,I16539,I16282);
nor I_814 (I16200,I16494,I16556);
nor I_815 (I16587,I16539,I16344);
DFFARX1 I_816  ( .D(I16587), .CLK(I2702), .RSTB(I16214), .Q(I16191) );
nor I_817 (I16206,I16539,I16265);
not I_818 (I16632,I16539);
nor I_819 (I16649,I16412,I16632);
and I_820 (I16666,I16299,I16649);
or I_821 (I16683,I16494,I16666);
DFFARX1 I_822  ( .D(I16683), .CLK(I2702), .RSTB(I16214), .Q(I16179) );
nand I_823 (I16188,I16539,I16361);
nand I_824 (I16176,I16539,I16443);
not I_825 (I16775,I2709);
nand I_826 (I16792,I382267,I382258);
and I_827 (I16809,I16792,I382261);
DFFARX1 I_828  ( .D(I16809), .CLK(I2702), .RSTB(I16775), .Q(I16826) );
not I_829 (I16843,I16826);
nor I_830 (I16860,I382237,I382258);
or I_831 (I16758,I16860,I16826);
not I_832 (I16746,I16860);
DFFARX1 I_833  ( .D(I382252), .CLK(I2702), .RSTB(I16775), .Q(I16905) );
nor I_834 (I16922,I16905,I16860);
nand I_835 (I16939,I382240,I382255);
and I_836 (I16956,I16939,I382249);
DFFARX1 I_837  ( .D(I16956), .CLK(I2702), .RSTB(I16775), .Q(I16973) );
nor I_838 (I16755,I16973,I16826);
not I_839 (I17004,I16973);
nor I_840 (I17021,I16905,I17004);
DFFARX1 I_841  ( .D(I382264), .CLK(I2702), .RSTB(I16775), .Q(I17038) );
and I_842 (I17055,I17038,I382243);
or I_843 (I16764,I17055,I16860);
nand I_844 (I16743,I17055,I17021);
DFFARX1 I_845  ( .D(I382246), .CLK(I2702), .RSTB(I16775), .Q(I17100) );
and I_846 (I17117,I17100,I16843);
nor I_847 (I16761,I17055,I17117);
nor I_848 (I17148,I17100,I16905);
DFFARX1 I_849  ( .D(I17148), .CLK(I2702), .RSTB(I16775), .Q(I16752) );
nor I_850 (I16767,I17100,I16826);
not I_851 (I17193,I17100);
nor I_852 (I17210,I16973,I17193);
and I_853 (I17227,I16860,I17210);
or I_854 (I17244,I17055,I17227);
DFFARX1 I_855  ( .D(I17244), .CLK(I2702), .RSTB(I16775), .Q(I16740) );
nand I_856 (I16749,I17100,I16922);
nand I_857 (I16737,I17100,I17004);
not I_858 (I17336,I2709);
nand I_859 (I17353,I156792,I156789);
and I_860 (I17370,I17353,I156786);
DFFARX1 I_861  ( .D(I17370), .CLK(I2702), .RSTB(I17336), .Q(I17387) );
not I_862 (I17404,I17387);
nor I_863 (I17421,I156810,I156789);
or I_864 (I17319,I17421,I17387);
not I_865 (I17307,I17421);
DFFARX1 I_866  ( .D(I156804), .CLK(I2702), .RSTB(I17336), .Q(I17466) );
nor I_867 (I17483,I17466,I17421);
nand I_868 (I17500,I156783,I156795);
and I_869 (I17517,I17500,I156798);
DFFARX1 I_870  ( .D(I17517), .CLK(I2702), .RSTB(I17336), .Q(I17534) );
nor I_871 (I17316,I17534,I17387);
not I_872 (I17565,I17534);
nor I_873 (I17582,I17466,I17565);
DFFARX1 I_874  ( .D(I156807), .CLK(I2702), .RSTB(I17336), .Q(I17599) );
and I_875 (I17616,I17599,I156813);
or I_876 (I17325,I17616,I17421);
nand I_877 (I17304,I17616,I17582);
DFFARX1 I_878  ( .D(I156801), .CLK(I2702), .RSTB(I17336), .Q(I17661) );
and I_879 (I17678,I17661,I17404);
nor I_880 (I17322,I17616,I17678);
nor I_881 (I17709,I17661,I17466);
DFFARX1 I_882  ( .D(I17709), .CLK(I2702), .RSTB(I17336), .Q(I17313) );
nor I_883 (I17328,I17661,I17387);
not I_884 (I17754,I17661);
nor I_885 (I17771,I17534,I17754);
and I_886 (I17788,I17421,I17771);
or I_887 (I17805,I17616,I17788);
DFFARX1 I_888  ( .D(I17805), .CLK(I2702), .RSTB(I17336), .Q(I17301) );
nand I_889 (I17310,I17661,I17483);
nand I_890 (I17298,I17661,I17565);
not I_891 (I17897,I2709);
nand I_892 (I17914,I454091,I454088);
and I_893 (I17931,I17914,I454082);
DFFARX1 I_894  ( .D(I17931), .CLK(I2702), .RSTB(I17897), .Q(I17948) );
not I_895 (I17965,I17948);
nor I_896 (I17982,I454094,I454088);
or I_897 (I17880,I17982,I17948);
not I_898 (I17868,I17982);
DFFARX1 I_899  ( .D(I454106), .CLK(I2702), .RSTB(I17897), .Q(I18027) );
nor I_900 (I18044,I18027,I17982);
nand I_901 (I18061,I454097,I454079);
and I_902 (I18078,I18061,I454109);
DFFARX1 I_903  ( .D(I18078), .CLK(I2702), .RSTB(I17897), .Q(I18095) );
nor I_904 (I17877,I18095,I17948);
not I_905 (I18126,I18095);
nor I_906 (I18143,I18027,I18126);
DFFARX1 I_907  ( .D(I454085), .CLK(I2702), .RSTB(I17897), .Q(I18160) );
and I_908 (I18177,I18160,I454103);
or I_909 (I17886,I18177,I17982);
nand I_910 (I17865,I18177,I18143);
DFFARX1 I_911  ( .D(I454100), .CLK(I2702), .RSTB(I17897), .Q(I18222) );
and I_912 (I18239,I18222,I17965);
nor I_913 (I17883,I18177,I18239);
nor I_914 (I18270,I18222,I18027);
DFFARX1 I_915  ( .D(I18270), .CLK(I2702), .RSTB(I17897), .Q(I17874) );
nor I_916 (I17889,I18222,I17948);
not I_917 (I18315,I18222);
nor I_918 (I18332,I18095,I18315);
and I_919 (I18349,I17982,I18332);
or I_920 (I18366,I18177,I18349);
DFFARX1 I_921  ( .D(I18366), .CLK(I2702), .RSTB(I17897), .Q(I17862) );
nand I_922 (I17871,I18222,I18044);
nand I_923 (I17859,I18222,I18126);
not I_924 (I18458,I2709);
nand I_925 (I18475,I212397,I212400);
and I_926 (I18492,I18475,I212394);
DFFARX1 I_927  ( .D(I18492), .CLK(I2702), .RSTB(I18458), .Q(I18509) );
not I_928 (I18526,I18509);
nor I_929 (I18543,I212385,I212400);
or I_930 (I18441,I18543,I18509);
not I_931 (I18429,I18543);
DFFARX1 I_932  ( .D(I212373), .CLK(I2702), .RSTB(I18458), .Q(I18588) );
nor I_933 (I18605,I18588,I18543);
nand I_934 (I18622,I212382,I212376);
and I_935 (I18639,I18622,I212388);
DFFARX1 I_936  ( .D(I18639), .CLK(I2702), .RSTB(I18458), .Q(I18656) );
nor I_937 (I18438,I18656,I18509);
not I_938 (I18687,I18656);
nor I_939 (I18704,I18588,I18687);
DFFARX1 I_940  ( .D(I212403), .CLK(I2702), .RSTB(I18458), .Q(I18721) );
and I_941 (I18738,I18721,I212391);
or I_942 (I18447,I18738,I18543);
nand I_943 (I18426,I18738,I18704);
DFFARX1 I_944  ( .D(I212379), .CLK(I2702), .RSTB(I18458), .Q(I18783) );
and I_945 (I18800,I18783,I18526);
nor I_946 (I18444,I18738,I18800);
nor I_947 (I18831,I18783,I18588);
DFFARX1 I_948  ( .D(I18831), .CLK(I2702), .RSTB(I18458), .Q(I18435) );
nor I_949 (I18450,I18783,I18509);
not I_950 (I18876,I18783);
nor I_951 (I18893,I18656,I18876);
and I_952 (I18910,I18543,I18893);
or I_953 (I18927,I18738,I18910);
DFFARX1 I_954  ( .D(I18927), .CLK(I2702), .RSTB(I18458), .Q(I18423) );
nand I_955 (I18432,I18783,I18605);
nand I_956 (I18420,I18783,I18687);
not I_957 (I19019,I2709);
nand I_958 (I19036,I470275,I470272);
and I_959 (I19053,I19036,I470266);
DFFARX1 I_960  ( .D(I19053), .CLK(I2702), .RSTB(I19019), .Q(I19070) );
not I_961 (I19087,I19070);
nor I_962 (I19104,I470278,I470272);
or I_963 (I19002,I19104,I19070);
not I_964 (I18990,I19104);
DFFARX1 I_965  ( .D(I470290), .CLK(I2702), .RSTB(I19019), .Q(I19149) );
nor I_966 (I19166,I19149,I19104);
nand I_967 (I19183,I470281,I470263);
and I_968 (I19200,I19183,I470293);
DFFARX1 I_969  ( .D(I19200), .CLK(I2702), .RSTB(I19019), .Q(I19217) );
nor I_970 (I18999,I19217,I19070);
not I_971 (I19248,I19217);
nor I_972 (I19265,I19149,I19248);
DFFARX1 I_973  ( .D(I470269), .CLK(I2702), .RSTB(I19019), .Q(I19282) );
and I_974 (I19299,I19282,I470287);
or I_975 (I19008,I19299,I19104);
nand I_976 (I18987,I19299,I19265);
DFFARX1 I_977  ( .D(I470284), .CLK(I2702), .RSTB(I19019), .Q(I19344) );
and I_978 (I19361,I19344,I19087);
nor I_979 (I19005,I19299,I19361);
nor I_980 (I19392,I19344,I19149);
DFFARX1 I_981  ( .D(I19392), .CLK(I2702), .RSTB(I19019), .Q(I18996) );
nor I_982 (I19011,I19344,I19070);
not I_983 (I19437,I19344);
nor I_984 (I19454,I19217,I19437);
and I_985 (I19471,I19104,I19454);
or I_986 (I19488,I19299,I19471);
DFFARX1 I_987  ( .D(I19488), .CLK(I2702), .RSTB(I19019), .Q(I18984) );
nand I_988 (I18993,I19344,I19166);
nand I_989 (I18981,I19344,I19248);
not I_990 (I19580,I2709);
nand I_991 (I19597,I692683,I692704);
and I_992 (I19614,I19597,I692692);
DFFARX1 I_993  ( .D(I19614), .CLK(I2702), .RSTB(I19580), .Q(I19631) );
not I_994 (I19648,I19631);
nor I_995 (I19665,I692698,I692704);
or I_996 (I19563,I19665,I19631);
not I_997 (I19551,I19665);
DFFARX1 I_998  ( .D(I692686), .CLK(I2702), .RSTB(I19580), .Q(I19710) );
nor I_999 (I19727,I19710,I19665);
nand I_1000 (I19744,I692677,I692695);
and I_1001 (I19761,I19744,I692689);
DFFARX1 I_1002  ( .D(I19761), .CLK(I2702), .RSTB(I19580), .Q(I19778) );
nor I_1003 (I19560,I19778,I19631);
not I_1004 (I19809,I19778);
nor I_1005 (I19826,I19710,I19809);
DFFARX1 I_1006  ( .D(I692701), .CLK(I2702), .RSTB(I19580), .Q(I19843) );
and I_1007 (I19860,I19843,I692674);
or I_1008 (I19569,I19860,I19665);
nand I_1009 (I19548,I19860,I19826);
DFFARX1 I_1010  ( .D(I692680), .CLK(I2702), .RSTB(I19580), .Q(I19905) );
and I_1011 (I19922,I19905,I19648);
nor I_1012 (I19566,I19860,I19922);
nor I_1013 (I19953,I19905,I19710);
DFFARX1 I_1014  ( .D(I19953), .CLK(I2702), .RSTB(I19580), .Q(I19557) );
nor I_1015 (I19572,I19905,I19631);
not I_1016 (I19998,I19905);
nor I_1017 (I20015,I19778,I19998);
and I_1018 (I20032,I19665,I20015);
or I_1019 (I20049,I19860,I20032);
DFFARX1 I_1020  ( .D(I20049), .CLK(I2702), .RSTB(I19580), .Q(I19545) );
nand I_1021 (I19554,I19905,I19727);
nand I_1022 (I19542,I19905,I19809);
not I_1023 (I20141,I2709);
nand I_1024 (I20158,I227272,I227275);
and I_1025 (I20175,I20158,I227269);
DFFARX1 I_1026  ( .D(I20175), .CLK(I2702), .RSTB(I20141), .Q(I20192) );
not I_1027 (I20209,I20192);
nor I_1028 (I20226,I227260,I227275);
or I_1029 (I20124,I20226,I20192);
not I_1030 (I20112,I20226);
DFFARX1 I_1031  ( .D(I227248), .CLK(I2702), .RSTB(I20141), .Q(I20271) );
nor I_1032 (I20288,I20271,I20226);
nand I_1033 (I20305,I227257,I227251);
and I_1034 (I20322,I20305,I227263);
DFFARX1 I_1035  ( .D(I20322), .CLK(I2702), .RSTB(I20141), .Q(I20339) );
nor I_1036 (I20121,I20339,I20192);
not I_1037 (I20370,I20339);
nor I_1038 (I20387,I20271,I20370);
DFFARX1 I_1039  ( .D(I227278), .CLK(I2702), .RSTB(I20141), .Q(I20404) );
and I_1040 (I20421,I20404,I227266);
or I_1041 (I20130,I20421,I20226);
nand I_1042 (I20109,I20421,I20387);
DFFARX1 I_1043  ( .D(I227254), .CLK(I2702), .RSTB(I20141), .Q(I20466) );
and I_1044 (I20483,I20466,I20209);
nor I_1045 (I20127,I20421,I20483);
nor I_1046 (I20514,I20466,I20271);
DFFARX1 I_1047  ( .D(I20514), .CLK(I2702), .RSTB(I20141), .Q(I20118) );
nor I_1048 (I20133,I20466,I20192);
not I_1049 (I20559,I20466);
nor I_1050 (I20576,I20339,I20559);
and I_1051 (I20593,I20226,I20576);
or I_1052 (I20610,I20421,I20593);
DFFARX1 I_1053  ( .D(I20610), .CLK(I2702), .RSTB(I20141), .Q(I20106) );
nand I_1054 (I20115,I20466,I20288);
nand I_1055 (I20103,I20466,I20370);
not I_1056 (I20702,I2709);
nand I_1057 (I20719,I719271,I719292);
and I_1058 (I20736,I20719,I719280);
DFFARX1 I_1059  ( .D(I20736), .CLK(I2702), .RSTB(I20702), .Q(I20753) );
not I_1060 (I20770,I20753);
nor I_1061 (I20787,I719286,I719292);
or I_1062 (I20685,I20787,I20753);
not I_1063 (I20673,I20787);
DFFARX1 I_1064  ( .D(I719274), .CLK(I2702), .RSTB(I20702), .Q(I20832) );
nor I_1065 (I20849,I20832,I20787);
nand I_1066 (I20866,I719265,I719283);
and I_1067 (I20883,I20866,I719277);
DFFARX1 I_1068  ( .D(I20883), .CLK(I2702), .RSTB(I20702), .Q(I20900) );
nor I_1069 (I20682,I20900,I20753);
not I_1070 (I20931,I20900);
nor I_1071 (I20948,I20832,I20931);
DFFARX1 I_1072  ( .D(I719289), .CLK(I2702), .RSTB(I20702), .Q(I20965) );
and I_1073 (I20982,I20965,I719262);
or I_1074 (I20691,I20982,I20787);
nand I_1075 (I20670,I20982,I20948);
DFFARX1 I_1076  ( .D(I719268), .CLK(I2702), .RSTB(I20702), .Q(I21027) );
and I_1077 (I21044,I21027,I20770);
nor I_1078 (I20688,I20982,I21044);
nor I_1079 (I21075,I21027,I20832);
DFFARX1 I_1080  ( .D(I21075), .CLK(I2702), .RSTB(I20702), .Q(I20679) );
nor I_1081 (I20694,I21027,I20753);
not I_1082 (I21120,I21027);
nor I_1083 (I21137,I20900,I21120);
and I_1084 (I21154,I20787,I21137);
or I_1085 (I21171,I20982,I21154);
DFFARX1 I_1086  ( .D(I21171), .CLK(I2702), .RSTB(I20702), .Q(I20667) );
nand I_1087 (I20676,I21027,I20849);
nand I_1088 (I20664,I21027,I20931);
not I_1089 (I21263,I2709);
nand I_1090 (I21280,I288744,I288735);
and I_1091 (I21297,I21280,I288750);
DFFARX1 I_1092  ( .D(I21297), .CLK(I2702), .RSTB(I21263), .Q(I21314) );
not I_1093 (I21331,I21314);
nor I_1094 (I21348,I288720,I288735);
or I_1095 (I21246,I21348,I21314);
not I_1096 (I21234,I21348);
DFFARX1 I_1097  ( .D(I288723), .CLK(I2702), .RSTB(I21263), .Q(I21393) );
nor I_1098 (I21410,I21393,I21348);
nand I_1099 (I21427,I288741,I288738);
and I_1100 (I21444,I21427,I288726);
DFFARX1 I_1101  ( .D(I21444), .CLK(I2702), .RSTB(I21263), .Q(I21461) );
nor I_1102 (I21243,I21461,I21314);
not I_1103 (I21492,I21461);
nor I_1104 (I21509,I21393,I21492);
DFFARX1 I_1105  ( .D(I288747), .CLK(I2702), .RSTB(I21263), .Q(I21526) );
and I_1106 (I21543,I21526,I288732);
or I_1107 (I21252,I21543,I21348);
nand I_1108 (I21231,I21543,I21509);
DFFARX1 I_1109  ( .D(I288729), .CLK(I2702), .RSTB(I21263), .Q(I21588) );
and I_1110 (I21605,I21588,I21331);
nor I_1111 (I21249,I21543,I21605);
nor I_1112 (I21636,I21588,I21393);
DFFARX1 I_1113  ( .D(I21636), .CLK(I2702), .RSTB(I21263), .Q(I21240) );
nor I_1114 (I21255,I21588,I21314);
not I_1115 (I21681,I21588);
nor I_1116 (I21698,I21461,I21681);
and I_1117 (I21715,I21348,I21698);
or I_1118 (I21732,I21543,I21715);
DFFARX1 I_1119  ( .D(I21732), .CLK(I2702), .RSTB(I21263), .Q(I21228) );
nand I_1120 (I21237,I21588,I21410);
nand I_1121 (I21225,I21588,I21492);
not I_1122 (I21824,I2709);
nand I_1123 (I21841,I591715,I591703);
and I_1124 (I21858,I21841,I591700);
DFFARX1 I_1125  ( .D(I21858), .CLK(I2702), .RSTB(I21824), .Q(I21875) );
not I_1126 (I21892,I21875);
nor I_1127 (I21909,I591721,I591703);
or I_1128 (I21807,I21909,I21875);
not I_1129 (I21795,I21909);
DFFARX1 I_1130  ( .D(I591724), .CLK(I2702), .RSTB(I21824), .Q(I21954) );
nor I_1131 (I21971,I21954,I21909);
nand I_1132 (I21988,I591694,I591712);
and I_1133 (I22005,I21988,I591709);
DFFARX1 I_1134  ( .D(I22005), .CLK(I2702), .RSTB(I21824), .Q(I22022) );
nor I_1135 (I21804,I22022,I21875);
not I_1136 (I22053,I22022);
nor I_1137 (I22070,I21954,I22053);
DFFARX1 I_1138  ( .D(I591718), .CLK(I2702), .RSTB(I21824), .Q(I22087) );
and I_1139 (I22104,I22087,I591706);
or I_1140 (I21813,I22104,I21909);
nand I_1141 (I21792,I22104,I22070);
DFFARX1 I_1142  ( .D(I591697), .CLK(I2702), .RSTB(I21824), .Q(I22149) );
and I_1143 (I22166,I22149,I21892);
nor I_1144 (I21810,I22104,I22166);
nor I_1145 (I22197,I22149,I21954);
DFFARX1 I_1146  ( .D(I22197), .CLK(I2702), .RSTB(I21824), .Q(I21801) );
nor I_1147 (I21816,I22149,I21875);
not I_1148 (I22242,I22149);
nor I_1149 (I22259,I22022,I22242);
and I_1150 (I22276,I21909,I22259);
or I_1151 (I22293,I22104,I22276);
DFFARX1 I_1152  ( .D(I22293), .CLK(I2702), .RSTB(I21824), .Q(I21789) );
nand I_1153 (I21798,I22149,I21971);
nand I_1154 (I21786,I22149,I22053);
not I_1155 (I22385,I2709);
nand I_1156 (I22402,I525057,I525060);
and I_1157 (I22419,I22402,I525072);
DFFARX1 I_1158  ( .D(I22419), .CLK(I2702), .RSTB(I22385), .Q(I22436) );
not I_1159 (I22453,I22436);
nor I_1160 (I22470,I525066,I525060);
or I_1161 (I22368,I22470,I22436);
not I_1162 (I22356,I22470);
DFFARX1 I_1163  ( .D(I525069), .CLK(I2702), .RSTB(I22385), .Q(I22515) );
nor I_1164 (I22532,I22515,I22470);
nand I_1165 (I22549,I525063,I525081);
and I_1166 (I22566,I22549,I525084);
DFFARX1 I_1167  ( .D(I22566), .CLK(I2702), .RSTB(I22385), .Q(I22583) );
nor I_1168 (I22365,I22583,I22436);
not I_1169 (I22614,I22583);
nor I_1170 (I22631,I22515,I22614);
DFFARX1 I_1171  ( .D(I525054), .CLK(I2702), .RSTB(I22385), .Q(I22648) );
and I_1172 (I22665,I22648,I525075);
or I_1173 (I22374,I22665,I22470);
nand I_1174 (I22353,I22665,I22631);
DFFARX1 I_1175  ( .D(I525078), .CLK(I2702), .RSTB(I22385), .Q(I22710) );
and I_1176 (I22727,I22710,I22453);
nor I_1177 (I22371,I22665,I22727);
nor I_1178 (I22758,I22710,I22515);
DFFARX1 I_1179  ( .D(I22758), .CLK(I2702), .RSTB(I22385), .Q(I22362) );
nor I_1180 (I22377,I22710,I22436);
not I_1181 (I22803,I22710);
nor I_1182 (I22820,I22583,I22803);
and I_1183 (I22837,I22470,I22820);
or I_1184 (I22854,I22665,I22837);
DFFARX1 I_1185  ( .D(I22854), .CLK(I2702), .RSTB(I22385), .Q(I22350) );
nand I_1186 (I22359,I22710,I22532);
nand I_1187 (I22347,I22710,I22614);
not I_1188 (I22946,I2709);
nand I_1189 (I22963,I303330,I303321);
and I_1190 (I22980,I22963,I303336);
DFFARX1 I_1191  ( .D(I22980), .CLK(I2702), .RSTB(I22946), .Q(I22997) );
not I_1192 (I23014,I22997);
nor I_1193 (I23031,I303306,I303321);
or I_1194 (I22929,I23031,I22997);
not I_1195 (I22917,I23031);
DFFARX1 I_1196  ( .D(I303309), .CLK(I2702), .RSTB(I22946), .Q(I23076) );
nor I_1197 (I23093,I23076,I23031);
nand I_1198 (I23110,I303327,I303324);
and I_1199 (I23127,I23110,I303312);
DFFARX1 I_1200  ( .D(I23127), .CLK(I2702), .RSTB(I22946), .Q(I23144) );
nor I_1201 (I22926,I23144,I22997);
not I_1202 (I23175,I23144);
nor I_1203 (I23192,I23076,I23175);
DFFARX1 I_1204  ( .D(I303333), .CLK(I2702), .RSTB(I22946), .Q(I23209) );
and I_1205 (I23226,I23209,I303318);
or I_1206 (I22935,I23226,I23031);
nand I_1207 (I22914,I23226,I23192);
DFFARX1 I_1208  ( .D(I303315), .CLK(I2702), .RSTB(I22946), .Q(I23271) );
and I_1209 (I23288,I23271,I23014);
nor I_1210 (I22932,I23226,I23288);
nor I_1211 (I23319,I23271,I23076);
DFFARX1 I_1212  ( .D(I23319), .CLK(I2702), .RSTB(I22946), .Q(I22923) );
nor I_1213 (I22938,I23271,I22997);
not I_1214 (I23364,I23271);
nor I_1215 (I23381,I23144,I23364);
and I_1216 (I23398,I23031,I23381);
or I_1217 (I23415,I23226,I23398);
DFFARX1 I_1218  ( .D(I23415), .CLK(I2702), .RSTB(I22946), .Q(I22911) );
nand I_1219 (I22920,I23271,I23093);
nand I_1220 (I22908,I23271,I23175);
not I_1221 (I23507,I2709);
nand I_1222 (I23524,I517322,I517325);
and I_1223 (I23541,I23524,I517337);
DFFARX1 I_1224  ( .D(I23541), .CLK(I2702), .RSTB(I23507), .Q(I23558) );
not I_1225 (I23575,I23558);
nor I_1226 (I23592,I517331,I517325);
or I_1227 (I23490,I23592,I23558);
not I_1228 (I23478,I23592);
DFFARX1 I_1229  ( .D(I517334), .CLK(I2702), .RSTB(I23507), .Q(I23637) );
nor I_1230 (I23654,I23637,I23592);
nand I_1231 (I23671,I517328,I517346);
and I_1232 (I23688,I23671,I517349);
DFFARX1 I_1233  ( .D(I23688), .CLK(I2702), .RSTB(I23507), .Q(I23705) );
nor I_1234 (I23487,I23705,I23558);
not I_1235 (I23736,I23705);
nor I_1236 (I23753,I23637,I23736);
DFFARX1 I_1237  ( .D(I517319), .CLK(I2702), .RSTB(I23507), .Q(I23770) );
and I_1238 (I23787,I23770,I517340);
or I_1239 (I23496,I23787,I23592);
nand I_1240 (I23475,I23787,I23753);
DFFARX1 I_1241  ( .D(I517343), .CLK(I2702), .RSTB(I23507), .Q(I23832) );
and I_1242 (I23849,I23832,I23575);
nor I_1243 (I23493,I23787,I23849);
nor I_1244 (I23880,I23832,I23637);
DFFARX1 I_1245  ( .D(I23880), .CLK(I2702), .RSTB(I23507), .Q(I23484) );
nor I_1246 (I23499,I23832,I23558);
not I_1247 (I23925,I23832);
nor I_1248 (I23942,I23705,I23925);
and I_1249 (I23959,I23592,I23942);
or I_1250 (I23976,I23787,I23959);
DFFARX1 I_1251  ( .D(I23976), .CLK(I2702), .RSTB(I23507), .Q(I23472) );
nand I_1252 (I23481,I23832,I23654);
nand I_1253 (I23469,I23832,I23736);
not I_1254 (I24068,I2709);
nand I_1255 (I24085,I377745,I377736);
and I_1256 (I24102,I24085,I377739);
DFFARX1 I_1257  ( .D(I24102), .CLK(I2702), .RSTB(I24068), .Q(I24119) );
not I_1258 (I24136,I24119);
nor I_1259 (I24153,I377715,I377736);
or I_1260 (I24051,I24153,I24119);
not I_1261 (I24039,I24153);
DFFARX1 I_1262  ( .D(I377730), .CLK(I2702), .RSTB(I24068), .Q(I24198) );
nor I_1263 (I24215,I24198,I24153);
nand I_1264 (I24232,I377718,I377733);
and I_1265 (I24249,I24232,I377727);
DFFARX1 I_1266  ( .D(I24249), .CLK(I2702), .RSTB(I24068), .Q(I24266) );
nor I_1267 (I24048,I24266,I24119);
not I_1268 (I24297,I24266);
nor I_1269 (I24314,I24198,I24297);
DFFARX1 I_1270  ( .D(I377742), .CLK(I2702), .RSTB(I24068), .Q(I24331) );
and I_1271 (I24348,I24331,I377721);
or I_1272 (I24057,I24348,I24153);
nand I_1273 (I24036,I24348,I24314);
DFFARX1 I_1274  ( .D(I377724), .CLK(I2702), .RSTB(I24068), .Q(I24393) );
and I_1275 (I24410,I24393,I24136);
nor I_1276 (I24054,I24348,I24410);
nor I_1277 (I24441,I24393,I24198);
DFFARX1 I_1278  ( .D(I24441), .CLK(I2702), .RSTB(I24068), .Q(I24045) );
nor I_1279 (I24060,I24393,I24119);
not I_1280 (I24486,I24393);
nor I_1281 (I24503,I24266,I24486);
and I_1282 (I24520,I24153,I24503);
or I_1283 (I24537,I24348,I24520);
DFFARX1 I_1284  ( .D(I24537), .CLK(I2702), .RSTB(I24068), .Q(I24033) );
nand I_1285 (I24042,I24393,I24215);
nand I_1286 (I24030,I24393,I24297);
not I_1287 (I24629,I2709);
nand I_1288 (I24646,I131168,I131171);
and I_1289 (I24663,I24646,I131153);
DFFARX1 I_1290  ( .D(I24663), .CLK(I2702), .RSTB(I24629), .Q(I24680) );
not I_1291 (I24697,I24680);
nor I_1292 (I24714,I131150,I131171);
or I_1293 (I24612,I24714,I24680);
not I_1294 (I24600,I24714);
DFFARX1 I_1295  ( .D(I131174), .CLK(I2702), .RSTB(I24629), .Q(I24759) );
nor I_1296 (I24776,I24759,I24714);
nand I_1297 (I24793,I131159,I131165);
and I_1298 (I24810,I24793,I131177);
DFFARX1 I_1299  ( .D(I24810), .CLK(I2702), .RSTB(I24629), .Q(I24827) );
nor I_1300 (I24609,I24827,I24680);
not I_1301 (I24858,I24827);
nor I_1302 (I24875,I24759,I24858);
DFFARX1 I_1303  ( .D(I131156), .CLK(I2702), .RSTB(I24629), .Q(I24892) );
and I_1304 (I24909,I24892,I131147);
or I_1305 (I24618,I24909,I24714);
nand I_1306 (I24597,I24909,I24875);
DFFARX1 I_1307  ( .D(I131162), .CLK(I2702), .RSTB(I24629), .Q(I24954) );
and I_1308 (I24971,I24954,I24697);
nor I_1309 (I24615,I24909,I24971);
nor I_1310 (I25002,I24954,I24759);
DFFARX1 I_1311  ( .D(I25002), .CLK(I2702), .RSTB(I24629), .Q(I24606) );
nor I_1312 (I24621,I24954,I24680);
not I_1313 (I25047,I24954);
nor I_1314 (I25064,I24827,I25047);
and I_1315 (I25081,I24714,I25064);
or I_1316 (I25098,I24909,I25081);
DFFARX1 I_1317  ( .D(I25098), .CLK(I2702), .RSTB(I24629), .Q(I24594) );
nand I_1318 (I24603,I24954,I24776);
nand I_1319 (I24591,I24954,I24858);
not I_1320 (I25190,I2709);
nand I_1321 (I25207,I146847,I146844);
and I_1322 (I25224,I25207,I146841);
DFFARX1 I_1323  ( .D(I25224), .CLK(I2702), .RSTB(I25190), .Q(I25241) );
not I_1324 (I25258,I25241);
nor I_1325 (I25275,I146865,I146844);
or I_1326 (I25173,I25275,I25241);
not I_1327 (I25161,I25275);
DFFARX1 I_1328  ( .D(I146859), .CLK(I2702), .RSTB(I25190), .Q(I25320) );
nor I_1329 (I25337,I25320,I25275);
nand I_1330 (I25354,I146838,I146850);
and I_1331 (I25371,I25354,I146853);
DFFARX1 I_1332  ( .D(I25371), .CLK(I2702), .RSTB(I25190), .Q(I25388) );
nor I_1333 (I25170,I25388,I25241);
not I_1334 (I25419,I25388);
nor I_1335 (I25436,I25320,I25419);
DFFARX1 I_1336  ( .D(I146862), .CLK(I2702), .RSTB(I25190), .Q(I25453) );
and I_1337 (I25470,I25453,I146868);
or I_1338 (I25179,I25470,I25275);
nand I_1339 (I25158,I25470,I25436);
DFFARX1 I_1340  ( .D(I146856), .CLK(I2702), .RSTB(I25190), .Q(I25515) );
and I_1341 (I25532,I25515,I25258);
nor I_1342 (I25176,I25470,I25532);
nor I_1343 (I25563,I25515,I25320);
DFFARX1 I_1344  ( .D(I25563), .CLK(I2702), .RSTB(I25190), .Q(I25167) );
nor I_1345 (I25182,I25515,I25241);
not I_1346 (I25608,I25515);
nor I_1347 (I25625,I25388,I25608);
and I_1348 (I25642,I25275,I25625);
or I_1349 (I25659,I25470,I25642);
DFFARX1 I_1350  ( .D(I25659), .CLK(I2702), .RSTB(I25190), .Q(I25155) );
nand I_1351 (I25164,I25515,I25337);
nand I_1352 (I25152,I25515,I25419);
not I_1353 (I25751,I2709);
nand I_1354 (I25768,I694417,I694438);
and I_1355 (I25785,I25768,I694426);
DFFARX1 I_1356  ( .D(I25785), .CLK(I2702), .RSTB(I25751), .Q(I25802) );
not I_1357 (I25819,I25802);
nor I_1358 (I25836,I694432,I694438);
or I_1359 (I25734,I25836,I25802);
not I_1360 (I25722,I25836);
DFFARX1 I_1361  ( .D(I694420), .CLK(I2702), .RSTB(I25751), .Q(I25881) );
nor I_1362 (I25898,I25881,I25836);
nand I_1363 (I25915,I694411,I694429);
and I_1364 (I25932,I25915,I694423);
DFFARX1 I_1365  ( .D(I25932), .CLK(I2702), .RSTB(I25751), .Q(I25949) );
nor I_1366 (I25731,I25949,I25802);
not I_1367 (I25980,I25949);
nor I_1368 (I25997,I25881,I25980);
DFFARX1 I_1369  ( .D(I694435), .CLK(I2702), .RSTB(I25751), .Q(I26014) );
and I_1370 (I26031,I26014,I694408);
or I_1371 (I25740,I26031,I25836);
nand I_1372 (I25719,I26031,I25997);
DFFARX1 I_1373  ( .D(I694414), .CLK(I2702), .RSTB(I25751), .Q(I26076) );
and I_1374 (I26093,I26076,I25819);
nor I_1375 (I25737,I26031,I26093);
nor I_1376 (I26124,I26076,I25881);
DFFARX1 I_1377  ( .D(I26124), .CLK(I2702), .RSTB(I25751), .Q(I25728) );
nor I_1378 (I25743,I26076,I25802);
not I_1379 (I26169,I26076);
nor I_1380 (I26186,I25949,I26169);
and I_1381 (I26203,I25836,I26186);
or I_1382 (I26220,I26031,I26203);
DFFARX1 I_1383  ( .D(I26220), .CLK(I2702), .RSTB(I25751), .Q(I25716) );
nand I_1384 (I25725,I26076,I25898);
nand I_1385 (I25713,I26076,I25980);
not I_1386 (I26312,I2709);
nand I_1387 (I26329,I205257,I205260);
and I_1388 (I26346,I26329,I205254);
DFFARX1 I_1389  ( .D(I26346), .CLK(I2702), .RSTB(I26312), .Q(I26363) );
not I_1390 (I26380,I26363);
nor I_1391 (I26397,I205245,I205260);
or I_1392 (I26295,I26397,I26363);
not I_1393 (I26283,I26397);
DFFARX1 I_1394  ( .D(I205233), .CLK(I2702), .RSTB(I26312), .Q(I26442) );
nor I_1395 (I26459,I26442,I26397);
nand I_1396 (I26476,I205242,I205236);
and I_1397 (I26493,I26476,I205248);
DFFARX1 I_1398  ( .D(I26493), .CLK(I2702), .RSTB(I26312), .Q(I26510) );
nor I_1399 (I26292,I26510,I26363);
not I_1400 (I26541,I26510);
nor I_1401 (I26558,I26442,I26541);
DFFARX1 I_1402  ( .D(I205263), .CLK(I2702), .RSTB(I26312), .Q(I26575) );
and I_1403 (I26592,I26575,I205251);
or I_1404 (I26301,I26592,I26397);
nand I_1405 (I26280,I26592,I26558);
DFFARX1 I_1406  ( .D(I205239), .CLK(I2702), .RSTB(I26312), .Q(I26637) );
and I_1407 (I26654,I26637,I26380);
nor I_1408 (I26298,I26592,I26654);
nor I_1409 (I26685,I26637,I26442);
DFFARX1 I_1410  ( .D(I26685), .CLK(I2702), .RSTB(I26312), .Q(I26289) );
nor I_1411 (I26304,I26637,I26363);
not I_1412 (I26730,I26637);
nor I_1413 (I26747,I26510,I26730);
and I_1414 (I26764,I26397,I26747);
or I_1415 (I26781,I26592,I26764);
DFFARX1 I_1416  ( .D(I26781), .CLK(I2702), .RSTB(I26312), .Q(I26277) );
nand I_1417 (I26286,I26637,I26459);
nand I_1418 (I26274,I26637,I26541);
not I_1419 (I26873,I2709);
nand I_1420 (I26890,I350613,I350604);
and I_1421 (I26907,I26890,I350607);
DFFARX1 I_1422  ( .D(I26907), .CLK(I2702), .RSTB(I26873), .Q(I26924) );
not I_1423 (I26941,I26924);
nor I_1424 (I26958,I350583,I350604);
or I_1425 (I26856,I26958,I26924);
not I_1426 (I26844,I26958);
DFFARX1 I_1427  ( .D(I350598), .CLK(I2702), .RSTB(I26873), .Q(I27003) );
nor I_1428 (I27020,I27003,I26958);
nand I_1429 (I27037,I350586,I350601);
and I_1430 (I27054,I27037,I350595);
DFFARX1 I_1431  ( .D(I27054), .CLK(I2702), .RSTB(I26873), .Q(I27071) );
nor I_1432 (I26853,I27071,I26924);
not I_1433 (I27102,I27071);
nor I_1434 (I27119,I27003,I27102);
DFFARX1 I_1435  ( .D(I350610), .CLK(I2702), .RSTB(I26873), .Q(I27136) );
and I_1436 (I27153,I27136,I350589);
or I_1437 (I26862,I27153,I26958);
nand I_1438 (I26841,I27153,I27119);
DFFARX1 I_1439  ( .D(I350592), .CLK(I2702), .RSTB(I26873), .Q(I27198) );
and I_1440 (I27215,I27198,I26941);
nor I_1441 (I26859,I27153,I27215);
nor I_1442 (I27246,I27198,I27003);
DFFARX1 I_1443  ( .D(I27246), .CLK(I2702), .RSTB(I26873), .Q(I26850) );
nor I_1444 (I26865,I27198,I26924);
not I_1445 (I27291,I27198);
nor I_1446 (I27308,I27071,I27291);
and I_1447 (I27325,I26958,I27308);
or I_1448 (I27342,I27153,I27325);
DFFARX1 I_1449  ( .D(I27342), .CLK(I2702), .RSTB(I26873), .Q(I26838) );
nand I_1450 (I26847,I27198,I27020);
nand I_1451 (I26835,I27198,I27102);
not I_1452 (I27434,I2709);
nand I_1453 (I27451,I635690,I635693);
and I_1454 (I27468,I27451,I635699);
DFFARX1 I_1455  ( .D(I27468), .CLK(I2702), .RSTB(I27434), .Q(I27485) );
not I_1456 (I27502,I27485);
nor I_1457 (I27519,I635711,I635693);
or I_1458 (I27417,I27519,I27485);
not I_1459 (I27405,I27519);
DFFARX1 I_1460  ( .D(I635720), .CLK(I2702), .RSTB(I27434), .Q(I27564) );
nor I_1461 (I27581,I27564,I27519);
nand I_1462 (I27598,I635708,I635705);
and I_1463 (I27615,I27598,I635717);
DFFARX1 I_1464  ( .D(I27615), .CLK(I2702), .RSTB(I27434), .Q(I27632) );
nor I_1465 (I27414,I27632,I27485);
not I_1466 (I27663,I27632);
nor I_1467 (I27680,I27564,I27663);
DFFARX1 I_1468  ( .D(I635714), .CLK(I2702), .RSTB(I27434), .Q(I27697) );
and I_1469 (I27714,I27697,I635702);
or I_1470 (I27423,I27714,I27519);
nand I_1471 (I27402,I27714,I27680);
DFFARX1 I_1472  ( .D(I635696), .CLK(I2702), .RSTB(I27434), .Q(I27759) );
and I_1473 (I27776,I27759,I27502);
nor I_1474 (I27420,I27714,I27776);
nor I_1475 (I27807,I27759,I27564);
DFFARX1 I_1476  ( .D(I27807), .CLK(I2702), .RSTB(I27434), .Q(I27411) );
nor I_1477 (I27426,I27759,I27485);
not I_1478 (I27852,I27759);
nor I_1479 (I27869,I27632,I27852);
and I_1480 (I27886,I27519,I27869);
or I_1481 (I27903,I27714,I27886);
DFFARX1 I_1482  ( .D(I27903), .CLK(I2702), .RSTB(I27434), .Q(I27399) );
nand I_1483 (I27408,I27759,I27581);
nand I_1484 (I27396,I27759,I27663);
not I_1485 (I27995,I2709);
nand I_1486 (I28012,I422990,I422984);
and I_1487 (I28029,I28012,I422996);
DFFARX1 I_1488  ( .D(I28029), .CLK(I2702), .RSTB(I27995), .Q(I28046) );
not I_1489 (I28063,I28046);
nor I_1490 (I28080,I422993,I422984);
or I_1491 (I27978,I28080,I28046);
not I_1492 (I27966,I28080);
DFFARX1 I_1493  ( .D(I422972), .CLK(I2702), .RSTB(I27995), .Q(I28125) );
nor I_1494 (I28142,I28125,I28080);
nand I_1495 (I28159,I422978,I422987);
and I_1496 (I28176,I28159,I422975);
DFFARX1 I_1497  ( .D(I28176), .CLK(I2702), .RSTB(I27995), .Q(I28193) );
nor I_1498 (I27975,I28193,I28046);
not I_1499 (I28224,I28193);
nor I_1500 (I28241,I28125,I28224);
DFFARX1 I_1501  ( .D(I422999), .CLK(I2702), .RSTB(I27995), .Q(I28258) );
and I_1502 (I28275,I28258,I422969);
or I_1503 (I27984,I28275,I28080);
nand I_1504 (I27963,I28275,I28241);
DFFARX1 I_1505  ( .D(I422981), .CLK(I2702), .RSTB(I27995), .Q(I28320) );
and I_1506 (I28337,I28320,I28063);
nor I_1507 (I27981,I28275,I28337);
nor I_1508 (I28368,I28320,I28125);
DFFARX1 I_1509  ( .D(I28368), .CLK(I2702), .RSTB(I27995), .Q(I27972) );
nor I_1510 (I27987,I28320,I28046);
not I_1511 (I28413,I28320);
nor I_1512 (I28430,I28193,I28413);
and I_1513 (I28447,I28080,I28430);
or I_1514 (I28464,I28275,I28447);
DFFARX1 I_1515  ( .D(I28464), .CLK(I2702), .RSTB(I27995), .Q(I27960) );
nand I_1516 (I27969,I28320,I28142);
nand I_1517 (I27957,I28320,I28224);
not I_1518 (I28556,I2709);
nand I_1519 (I28573,I316590,I316581);
and I_1520 (I28590,I28573,I316596);
DFFARX1 I_1521  ( .D(I28590), .CLK(I2702), .RSTB(I28556), .Q(I28607) );
not I_1522 (I28624,I28607);
nor I_1523 (I28641,I316566,I316581);
or I_1524 (I28539,I28641,I28607);
not I_1525 (I28527,I28641);
DFFARX1 I_1526  ( .D(I316569), .CLK(I2702), .RSTB(I28556), .Q(I28686) );
nor I_1527 (I28703,I28686,I28641);
nand I_1528 (I28720,I316587,I316584);
and I_1529 (I28737,I28720,I316572);
DFFARX1 I_1530  ( .D(I28737), .CLK(I2702), .RSTB(I28556), .Q(I28754) );
nor I_1531 (I28536,I28754,I28607);
not I_1532 (I28785,I28754);
nor I_1533 (I28802,I28686,I28785);
DFFARX1 I_1534  ( .D(I316593), .CLK(I2702), .RSTB(I28556), .Q(I28819) );
and I_1535 (I28836,I28819,I316578);
or I_1536 (I28545,I28836,I28641);
nand I_1537 (I28524,I28836,I28802);
DFFARX1 I_1538  ( .D(I316575), .CLK(I2702), .RSTB(I28556), .Q(I28881) );
and I_1539 (I28898,I28881,I28624);
nor I_1540 (I28542,I28836,I28898);
nor I_1541 (I28929,I28881,I28686);
DFFARX1 I_1542  ( .D(I28929), .CLK(I2702), .RSTB(I28556), .Q(I28533) );
nor I_1543 (I28548,I28881,I28607);
not I_1544 (I28974,I28881);
nor I_1545 (I28991,I28754,I28974);
and I_1546 (I29008,I28641,I28991);
or I_1547 (I29025,I28836,I29008);
DFFARX1 I_1548  ( .D(I29025), .CLK(I2702), .RSTB(I28556), .Q(I28521) );
nand I_1549 (I28530,I28881,I28703);
nand I_1550 (I28518,I28881,I28785);
not I_1551 (I29117,I2709);
nand I_1552 (I29134,I700197,I700218);
and I_1553 (I29151,I29134,I700206);
DFFARX1 I_1554  ( .D(I29151), .CLK(I2702), .RSTB(I29117), .Q(I29168) );
not I_1555 (I29185,I29168);
nor I_1556 (I29202,I700212,I700218);
or I_1557 (I29100,I29202,I29168);
not I_1558 (I29088,I29202);
DFFARX1 I_1559  ( .D(I700200), .CLK(I2702), .RSTB(I29117), .Q(I29247) );
nor I_1560 (I29264,I29247,I29202);
nand I_1561 (I29281,I700191,I700209);
and I_1562 (I29298,I29281,I700203);
DFFARX1 I_1563  ( .D(I29298), .CLK(I2702), .RSTB(I29117), .Q(I29315) );
nor I_1564 (I29097,I29315,I29168);
not I_1565 (I29346,I29315);
nor I_1566 (I29363,I29247,I29346);
DFFARX1 I_1567  ( .D(I700215), .CLK(I2702), .RSTB(I29117), .Q(I29380) );
and I_1568 (I29397,I29380,I700188);
or I_1569 (I29106,I29397,I29202);
nand I_1570 (I29085,I29397,I29363);
DFFARX1 I_1571  ( .D(I700194), .CLK(I2702), .RSTB(I29117), .Q(I29442) );
and I_1572 (I29459,I29442,I29185);
nor I_1573 (I29103,I29397,I29459);
nor I_1574 (I29490,I29442,I29247);
DFFARX1 I_1575  ( .D(I29490), .CLK(I2702), .RSTB(I29117), .Q(I29094) );
nor I_1576 (I29109,I29442,I29168);
not I_1577 (I29535,I29442);
nor I_1578 (I29552,I29315,I29535);
and I_1579 (I29569,I29202,I29552);
or I_1580 (I29586,I29397,I29569);
DFFARX1 I_1581  ( .D(I29586), .CLK(I2702), .RSTB(I29117), .Q(I29082) );
nand I_1582 (I29091,I29442,I29264);
nand I_1583 (I29079,I29442,I29346);
not I_1584 (I29678,I2709);
nand I_1585 (I29695,I230235,I230229);
and I_1586 (I29712,I29695,I230223);
DFFARX1 I_1587  ( .D(I29712), .CLK(I2702), .RSTB(I29678), .Q(I29729) );
not I_1588 (I29746,I29729);
nor I_1589 (I29763,I230250,I230229);
or I_1590 (I29661,I29763,I29729);
not I_1591 (I29649,I29763);
DFFARX1 I_1592  ( .D(I230247), .CLK(I2702), .RSTB(I29678), .Q(I29808) );
nor I_1593 (I29825,I29808,I29763);
nand I_1594 (I29842,I230253,I230241);
and I_1595 (I29859,I29842,I230238);
DFFARX1 I_1596  ( .D(I29859), .CLK(I2702), .RSTB(I29678), .Q(I29876) );
nor I_1597 (I29658,I29876,I29729);
not I_1598 (I29907,I29876);
nor I_1599 (I29924,I29808,I29907);
DFFARX1 I_1600  ( .D(I230226), .CLK(I2702), .RSTB(I29678), .Q(I29941) );
and I_1601 (I29958,I29941,I230244);
or I_1602 (I29667,I29958,I29763);
nand I_1603 (I29646,I29958,I29924);
DFFARX1 I_1604  ( .D(I230232), .CLK(I2702), .RSTB(I29678), .Q(I30003) );
and I_1605 (I30020,I30003,I29746);
nor I_1606 (I29664,I29958,I30020);
nor I_1607 (I30051,I30003,I29808);
DFFARX1 I_1608  ( .D(I30051), .CLK(I2702), .RSTB(I29678), .Q(I29655) );
nor I_1609 (I29670,I30003,I29729);
not I_1610 (I30096,I30003);
nor I_1611 (I30113,I29876,I30096);
and I_1612 (I30130,I29763,I30113);
or I_1613 (I30147,I29958,I30130);
DFFARX1 I_1614  ( .D(I30147), .CLK(I2702), .RSTB(I29678), .Q(I29643) );
nand I_1615 (I29652,I30003,I29825);
nand I_1616 (I29640,I30003,I29907);
not I_1617 (I30239,I2709);
nand I_1618 (I30256,I448311,I448308);
and I_1619 (I30273,I30256,I448302);
DFFARX1 I_1620  ( .D(I30273), .CLK(I2702), .RSTB(I30239), .Q(I30290) );
not I_1621 (I30307,I30290);
nor I_1622 (I30324,I448314,I448308);
or I_1623 (I30222,I30324,I30290);
not I_1624 (I30210,I30324);
DFFARX1 I_1625  ( .D(I448326), .CLK(I2702), .RSTB(I30239), .Q(I30369) );
nor I_1626 (I30386,I30369,I30324);
nand I_1627 (I30403,I448317,I448299);
and I_1628 (I30420,I30403,I448329);
DFFARX1 I_1629  ( .D(I30420), .CLK(I2702), .RSTB(I30239), .Q(I30437) );
nor I_1630 (I30219,I30437,I30290);
not I_1631 (I30468,I30437);
nor I_1632 (I30485,I30369,I30468);
DFFARX1 I_1633  ( .D(I448305), .CLK(I2702), .RSTB(I30239), .Q(I30502) );
and I_1634 (I30519,I30502,I448323);
or I_1635 (I30228,I30519,I30324);
nand I_1636 (I30207,I30519,I30485);
DFFARX1 I_1637  ( .D(I448320), .CLK(I2702), .RSTB(I30239), .Q(I30564) );
and I_1638 (I30581,I30564,I30307);
nor I_1639 (I30225,I30519,I30581);
nor I_1640 (I30612,I30564,I30369);
DFFARX1 I_1641  ( .D(I30612), .CLK(I2702), .RSTB(I30239), .Q(I30216) );
nor I_1642 (I30231,I30564,I30290);
not I_1643 (I30657,I30564);
nor I_1644 (I30674,I30437,I30657);
and I_1645 (I30691,I30324,I30674);
or I_1646 (I30708,I30519,I30691);
DFFARX1 I_1647  ( .D(I30708), .CLK(I2702), .RSTB(I30239), .Q(I30204) );
nand I_1648 (I30213,I30564,I30386);
nand I_1649 (I30201,I30564,I30468);
not I_1650 (I30800,I2709);
nand I_1651 (I30817,I94992,I94995);
and I_1652 (I30834,I30817,I94977);
DFFARX1 I_1653  ( .D(I30834), .CLK(I2702), .RSTB(I30800), .Q(I30851) );
not I_1654 (I30868,I30851);
nor I_1655 (I30885,I94974,I94995);
or I_1656 (I30783,I30885,I30851);
not I_1657 (I30771,I30885);
DFFARX1 I_1658  ( .D(I94998), .CLK(I2702), .RSTB(I30800), .Q(I30930) );
nor I_1659 (I30947,I30930,I30885);
nand I_1660 (I30964,I94983,I94989);
and I_1661 (I30981,I30964,I95001);
DFFARX1 I_1662  ( .D(I30981), .CLK(I2702), .RSTB(I30800), .Q(I30998) );
nor I_1663 (I30780,I30998,I30851);
not I_1664 (I31029,I30998);
nor I_1665 (I31046,I30930,I31029);
DFFARX1 I_1666  ( .D(I94980), .CLK(I2702), .RSTB(I30800), .Q(I31063) );
and I_1667 (I31080,I31063,I94971);
or I_1668 (I30789,I31080,I30885);
nand I_1669 (I30768,I31080,I31046);
DFFARX1 I_1670  ( .D(I94986), .CLK(I2702), .RSTB(I30800), .Q(I31125) );
and I_1671 (I31142,I31125,I30868);
nor I_1672 (I30786,I31080,I31142);
nor I_1673 (I31173,I31125,I30930);
DFFARX1 I_1674  ( .D(I31173), .CLK(I2702), .RSTB(I30800), .Q(I30777) );
nor I_1675 (I30792,I31125,I30851);
not I_1676 (I31218,I31125);
nor I_1677 (I31235,I30998,I31218);
and I_1678 (I31252,I30885,I31235);
or I_1679 (I31269,I31080,I31252);
DFFARX1 I_1680  ( .D(I31269), .CLK(I2702), .RSTB(I30800), .Q(I30765) );
nand I_1681 (I30774,I31125,I30947);
nand I_1682 (I30762,I31125,I31029);
not I_1683 (I31361,I2709);
nand I_1684 (I31378,I598855,I598843);
and I_1685 (I31395,I31378,I598840);
DFFARX1 I_1686  ( .D(I31395), .CLK(I2702), .RSTB(I31361), .Q(I31412) );
not I_1687 (I31429,I31412);
nor I_1688 (I31446,I598861,I598843);
or I_1689 (I31344,I31446,I31412);
not I_1690 (I31332,I31446);
DFFARX1 I_1691  ( .D(I598864), .CLK(I2702), .RSTB(I31361), .Q(I31491) );
nor I_1692 (I31508,I31491,I31446);
nand I_1693 (I31525,I598834,I598852);
and I_1694 (I31542,I31525,I598849);
DFFARX1 I_1695  ( .D(I31542), .CLK(I2702), .RSTB(I31361), .Q(I31559) );
nor I_1696 (I31341,I31559,I31412);
not I_1697 (I31590,I31559);
nor I_1698 (I31607,I31491,I31590);
DFFARX1 I_1699  ( .D(I598858), .CLK(I2702), .RSTB(I31361), .Q(I31624) );
and I_1700 (I31641,I31624,I598846);
or I_1701 (I31350,I31641,I31446);
nand I_1702 (I31329,I31641,I31607);
DFFARX1 I_1703  ( .D(I598837), .CLK(I2702), .RSTB(I31361), .Q(I31686) );
and I_1704 (I31703,I31686,I31429);
nor I_1705 (I31347,I31641,I31703);
nor I_1706 (I31734,I31686,I31491);
DFFARX1 I_1707  ( .D(I31734), .CLK(I2702), .RSTB(I31361), .Q(I31338) );
nor I_1708 (I31353,I31686,I31412);
not I_1709 (I31779,I31686);
nor I_1710 (I31796,I31559,I31779);
and I_1711 (I31813,I31446,I31796);
or I_1712 (I31830,I31641,I31813);
DFFARX1 I_1713  ( .D(I31830), .CLK(I2702), .RSTB(I31361), .Q(I31326) );
nand I_1714 (I31335,I31686,I31508);
nand I_1715 (I31323,I31686,I31590);
not I_1716 (I31922,I2709);
nand I_1717 (I31939,I108558,I108561);
and I_1718 (I31956,I31939,I108543);
DFFARX1 I_1719  ( .D(I31956), .CLK(I2702), .RSTB(I31922), .Q(I31973) );
not I_1720 (I31990,I31973);
nor I_1721 (I32007,I108540,I108561);
or I_1722 (I31905,I32007,I31973);
not I_1723 (I31893,I32007);
DFFARX1 I_1724  ( .D(I108564), .CLK(I2702), .RSTB(I31922), .Q(I32052) );
nor I_1725 (I32069,I32052,I32007);
nand I_1726 (I32086,I108549,I108555);
and I_1727 (I32103,I32086,I108567);
DFFARX1 I_1728  ( .D(I32103), .CLK(I2702), .RSTB(I31922), .Q(I32120) );
nor I_1729 (I31902,I32120,I31973);
not I_1730 (I32151,I32120);
nor I_1731 (I32168,I32052,I32151);
DFFARX1 I_1732  ( .D(I108546), .CLK(I2702), .RSTB(I31922), .Q(I32185) );
and I_1733 (I32202,I32185,I108537);
or I_1734 (I31911,I32202,I32007);
nand I_1735 (I31890,I32202,I32168);
DFFARX1 I_1736  ( .D(I108552), .CLK(I2702), .RSTB(I31922), .Q(I32247) );
and I_1737 (I32264,I32247,I31990);
nor I_1738 (I31908,I32202,I32264);
nor I_1739 (I32295,I32247,I32052);
DFFARX1 I_1740  ( .D(I32295), .CLK(I2702), .RSTB(I31922), .Q(I31899) );
nor I_1741 (I31914,I32247,I31973);
not I_1742 (I32340,I32247);
nor I_1743 (I32357,I32120,I32340);
and I_1744 (I32374,I32007,I32357);
or I_1745 (I32391,I32202,I32374);
DFFARX1 I_1746  ( .D(I32391), .CLK(I2702), .RSTB(I31922), .Q(I31887) );
nand I_1747 (I31896,I32247,I32069);
nand I_1748 (I31884,I32247,I32151);
not I_1749 (I32483,I2709);
nand I_1750 (I32500,I612540,I612528);
and I_1751 (I32517,I32500,I612525);
DFFARX1 I_1752  ( .D(I32517), .CLK(I2702), .RSTB(I32483), .Q(I32534) );
not I_1753 (I32551,I32534);
nor I_1754 (I32568,I612546,I612528);
or I_1755 (I32466,I32568,I32534);
not I_1756 (I32454,I32568);
DFFARX1 I_1757  ( .D(I612549), .CLK(I2702), .RSTB(I32483), .Q(I32613) );
nor I_1758 (I32630,I32613,I32568);
nand I_1759 (I32647,I612519,I612537);
and I_1760 (I32664,I32647,I612534);
DFFARX1 I_1761  ( .D(I32664), .CLK(I2702), .RSTB(I32483), .Q(I32681) );
nor I_1762 (I32463,I32681,I32534);
not I_1763 (I32712,I32681);
nor I_1764 (I32729,I32613,I32712);
DFFARX1 I_1765  ( .D(I612543), .CLK(I2702), .RSTB(I32483), .Q(I32746) );
and I_1766 (I32763,I32746,I612531);
or I_1767 (I32472,I32763,I32568);
nand I_1768 (I32451,I32763,I32729);
DFFARX1 I_1769  ( .D(I612522), .CLK(I2702), .RSTB(I32483), .Q(I32808) );
and I_1770 (I32825,I32808,I32551);
nor I_1771 (I32469,I32763,I32825);
nor I_1772 (I32856,I32808,I32613);
DFFARX1 I_1773  ( .D(I32856), .CLK(I2702), .RSTB(I32483), .Q(I32460) );
nor I_1774 (I32475,I32808,I32534);
not I_1775 (I32901,I32808);
nor I_1776 (I32918,I32681,I32901);
and I_1777 (I32935,I32568,I32918);
or I_1778 (I32952,I32763,I32935);
DFFARX1 I_1779  ( .D(I32952), .CLK(I2702), .RSTB(I32483), .Q(I32448) );
nand I_1780 (I32457,I32808,I32630);
nand I_1781 (I32445,I32808,I32712);
not I_1782 (I33044,I2709);
nand I_1783 (I33061,I314601,I314592);
and I_1784 (I33078,I33061,I314607);
DFFARX1 I_1785  ( .D(I33078), .CLK(I2702), .RSTB(I33044), .Q(I33095) );
not I_1786 (I33112,I33095);
nor I_1787 (I33129,I314577,I314592);
or I_1788 (I33027,I33129,I33095);
not I_1789 (I33015,I33129);
DFFARX1 I_1790  ( .D(I314580), .CLK(I2702), .RSTB(I33044), .Q(I33174) );
nor I_1791 (I33191,I33174,I33129);
nand I_1792 (I33208,I314598,I314595);
and I_1793 (I33225,I33208,I314583);
DFFARX1 I_1794  ( .D(I33225), .CLK(I2702), .RSTB(I33044), .Q(I33242) );
nor I_1795 (I33024,I33242,I33095);
not I_1796 (I33273,I33242);
nor I_1797 (I33290,I33174,I33273);
DFFARX1 I_1798  ( .D(I314604), .CLK(I2702), .RSTB(I33044), .Q(I33307) );
and I_1799 (I33324,I33307,I314589);
or I_1800 (I33033,I33324,I33129);
nand I_1801 (I33012,I33324,I33290);
DFFARX1 I_1802  ( .D(I314586), .CLK(I2702), .RSTB(I33044), .Q(I33369) );
and I_1803 (I33386,I33369,I33112);
nor I_1804 (I33030,I33324,I33386);
nor I_1805 (I33417,I33369,I33174);
DFFARX1 I_1806  ( .D(I33417), .CLK(I2702), .RSTB(I33044), .Q(I33021) );
nor I_1807 (I33036,I33369,I33095);
not I_1808 (I33462,I33369);
nor I_1809 (I33479,I33242,I33462);
and I_1810 (I33496,I33129,I33479);
or I_1811 (I33513,I33324,I33496);
DFFARX1 I_1812  ( .D(I33513), .CLK(I2702), .RSTB(I33044), .Q(I33009) );
nand I_1813 (I33018,I33369,I33191);
nand I_1814 (I33006,I33369,I33273);
not I_1815 (I33605,I2709);
nand I_1816 (I33622,I718693,I718714);
and I_1817 (I33639,I33622,I718702);
DFFARX1 I_1818  ( .D(I33639), .CLK(I2702), .RSTB(I33605), .Q(I33656) );
not I_1819 (I33673,I33656);
nor I_1820 (I33690,I718708,I718714);
or I_1821 (I33588,I33690,I33656);
not I_1822 (I33576,I33690);
DFFARX1 I_1823  ( .D(I718696), .CLK(I2702), .RSTB(I33605), .Q(I33735) );
nor I_1824 (I33752,I33735,I33690);
nand I_1825 (I33769,I718687,I718705);
and I_1826 (I33786,I33769,I718699);
DFFARX1 I_1827  ( .D(I33786), .CLK(I2702), .RSTB(I33605), .Q(I33803) );
nor I_1828 (I33585,I33803,I33656);
not I_1829 (I33834,I33803);
nor I_1830 (I33851,I33735,I33834);
DFFARX1 I_1831  ( .D(I718711), .CLK(I2702), .RSTB(I33605), .Q(I33868) );
and I_1832 (I33885,I33868,I718684);
or I_1833 (I33594,I33885,I33690);
nand I_1834 (I33573,I33885,I33851);
DFFARX1 I_1835  ( .D(I718690), .CLK(I2702), .RSTB(I33605), .Q(I33930) );
and I_1836 (I33947,I33930,I33673);
nor I_1837 (I33591,I33885,I33947);
nor I_1838 (I33978,I33930,I33735);
DFFARX1 I_1839  ( .D(I33978), .CLK(I2702), .RSTB(I33605), .Q(I33582) );
nor I_1840 (I33597,I33930,I33656);
not I_1841 (I34023,I33930);
nor I_1842 (I34040,I33803,I34023);
and I_1843 (I34057,I33690,I34040);
or I_1844 (I34074,I33885,I34057);
DFFARX1 I_1845  ( .D(I34074), .CLK(I2702), .RSTB(I33605), .Q(I33570) );
nand I_1846 (I33579,I33930,I33752);
nand I_1847 (I33567,I33930,I33834);
not I_1848 (I34166,I2709);
nand I_1849 (I34183,I679091,I679094);
and I_1850 (I34200,I34183,I679100);
DFFARX1 I_1851  ( .D(I34200), .CLK(I2702), .RSTB(I34166), .Q(I34217) );
not I_1852 (I34234,I34217);
nor I_1853 (I34251,I679112,I679094);
or I_1854 (I34149,I34251,I34217);
not I_1855 (I34137,I34251);
DFFARX1 I_1856  ( .D(I679121), .CLK(I2702), .RSTB(I34166), .Q(I34296) );
nor I_1857 (I34313,I34296,I34251);
nand I_1858 (I34330,I679109,I679106);
and I_1859 (I34347,I34330,I679118);
DFFARX1 I_1860  ( .D(I34347), .CLK(I2702), .RSTB(I34166), .Q(I34364) );
nor I_1861 (I34146,I34364,I34217);
not I_1862 (I34395,I34364);
nor I_1863 (I34412,I34296,I34395);
DFFARX1 I_1864  ( .D(I679115), .CLK(I2702), .RSTB(I34166), .Q(I34429) );
and I_1865 (I34446,I34429,I679103);
or I_1866 (I34155,I34446,I34251);
nand I_1867 (I34134,I34446,I34412);
DFFARX1 I_1868  ( .D(I679097), .CLK(I2702), .RSTB(I34166), .Q(I34491) );
and I_1869 (I34508,I34491,I34234);
nor I_1870 (I34152,I34446,I34508);
nor I_1871 (I34539,I34491,I34296);
DFFARX1 I_1872  ( .D(I34539), .CLK(I2702), .RSTB(I34166), .Q(I34143) );
nor I_1873 (I34158,I34491,I34217);
not I_1874 (I34584,I34491);
nor I_1875 (I34601,I34364,I34584);
and I_1876 (I34618,I34251,I34601);
or I_1877 (I34635,I34446,I34618);
DFFARX1 I_1878  ( .D(I34635), .CLK(I2702), .RSTB(I34166), .Q(I34131) );
nand I_1879 (I34140,I34491,I34313);
nand I_1880 (I34128,I34491,I34395);
not I_1881 (I34727,I2709);
nand I_1882 (I34744,I583385,I583373);
and I_1883 (I34761,I34744,I583370);
DFFARX1 I_1884  ( .D(I34761), .CLK(I2702), .RSTB(I34727), .Q(I34778) );
not I_1885 (I34795,I34778);
nor I_1886 (I34812,I583391,I583373);
or I_1887 (I34710,I34812,I34778);
not I_1888 (I34698,I34812);
DFFARX1 I_1889  ( .D(I583394), .CLK(I2702), .RSTB(I34727), .Q(I34857) );
nor I_1890 (I34874,I34857,I34812);
nand I_1891 (I34891,I583364,I583382);
and I_1892 (I34908,I34891,I583379);
DFFARX1 I_1893  ( .D(I34908), .CLK(I2702), .RSTB(I34727), .Q(I34925) );
nor I_1894 (I34707,I34925,I34778);
not I_1895 (I34956,I34925);
nor I_1896 (I34973,I34857,I34956);
DFFARX1 I_1897  ( .D(I583388), .CLK(I2702), .RSTB(I34727), .Q(I34990) );
and I_1898 (I35007,I34990,I583376);
or I_1899 (I34716,I35007,I34812);
nand I_1900 (I34695,I35007,I34973);
DFFARX1 I_1901  ( .D(I583367), .CLK(I2702), .RSTB(I34727), .Q(I35052) );
and I_1902 (I35069,I35052,I34795);
nor I_1903 (I34713,I35007,I35069);
nor I_1904 (I35100,I35052,I34857);
DFFARX1 I_1905  ( .D(I35100), .CLK(I2702), .RSTB(I34727), .Q(I34704) );
nor I_1906 (I34719,I35052,I34778);
not I_1907 (I35145,I35052);
nor I_1908 (I35162,I34925,I35145);
and I_1909 (I35179,I34812,I35162);
or I_1910 (I35196,I35007,I35179);
DFFARX1 I_1911  ( .D(I35196), .CLK(I2702), .RSTB(I34727), .Q(I34692) );
nand I_1912 (I34701,I35052,I34874);
nand I_1913 (I34689,I35052,I34956);
not I_1914 (I35288,I2709);
nand I_1915 (I35305,I596475,I596463);
and I_1916 (I35322,I35305,I596460);
DFFARX1 I_1917  ( .D(I35322), .CLK(I2702), .RSTB(I35288), .Q(I35339) );
not I_1918 (I35356,I35339);
nor I_1919 (I35373,I596481,I596463);
or I_1920 (I35271,I35373,I35339);
not I_1921 (I35259,I35373);
DFFARX1 I_1922  ( .D(I596484), .CLK(I2702), .RSTB(I35288), .Q(I35418) );
nor I_1923 (I35435,I35418,I35373);
nand I_1924 (I35452,I596454,I596472);
and I_1925 (I35469,I35452,I596469);
DFFARX1 I_1926  ( .D(I35469), .CLK(I2702), .RSTB(I35288), .Q(I35486) );
nor I_1927 (I35268,I35486,I35339);
not I_1928 (I35517,I35486);
nor I_1929 (I35534,I35418,I35517);
DFFARX1 I_1930  ( .D(I596478), .CLK(I2702), .RSTB(I35288), .Q(I35551) );
and I_1931 (I35568,I35551,I596466);
or I_1932 (I35277,I35568,I35373);
nand I_1933 (I35256,I35568,I35534);
DFFARX1 I_1934  ( .D(I596457), .CLK(I2702), .RSTB(I35288), .Q(I35613) );
and I_1935 (I35630,I35613,I35356);
nor I_1936 (I35274,I35568,I35630);
nor I_1937 (I35661,I35613,I35418);
DFFARX1 I_1938  ( .D(I35661), .CLK(I2702), .RSTB(I35288), .Q(I35265) );
nor I_1939 (I35280,I35613,I35339);
not I_1940 (I35706,I35613);
nor I_1941 (I35723,I35486,I35706);
and I_1942 (I35740,I35373,I35723);
or I_1943 (I35757,I35568,I35740);
DFFARX1 I_1944  ( .D(I35757), .CLK(I2702), .RSTB(I35288), .Q(I35253) );
nand I_1945 (I35262,I35613,I35435);
nand I_1946 (I35250,I35613,I35517);
not I_1947 (I35849,I2709);
nand I_1948 (I35866,I491951,I491933);
and I_1949 (I35883,I35866,I491942);
DFFARX1 I_1950  ( .D(I35883), .CLK(I2702), .RSTB(I35849), .Q(I35900) );
not I_1951 (I35917,I35900);
nor I_1952 (I35934,I491927,I491933);
or I_1953 (I35832,I35934,I35900);
not I_1954 (I35820,I35934);
DFFARX1 I_1955  ( .D(I491936), .CLK(I2702), .RSTB(I35849), .Q(I35979) );
nor I_1956 (I35996,I35979,I35934);
nand I_1957 (I36013,I491924,I491930);
and I_1958 (I36030,I36013,I491939);
DFFARX1 I_1959  ( .D(I36030), .CLK(I2702), .RSTB(I35849), .Q(I36047) );
nor I_1960 (I35829,I36047,I35900);
not I_1961 (I36078,I36047);
nor I_1962 (I36095,I35979,I36078);
DFFARX1 I_1963  ( .D(I491948), .CLK(I2702), .RSTB(I35849), .Q(I36112) );
and I_1964 (I36129,I36112,I491921);
or I_1965 (I35838,I36129,I35934);
nand I_1966 (I35817,I36129,I36095);
DFFARX1 I_1967  ( .D(I491945), .CLK(I2702), .RSTB(I35849), .Q(I36174) );
and I_1968 (I36191,I36174,I35917);
nor I_1969 (I35835,I36129,I36191);
nor I_1970 (I36222,I36174,I35979);
DFFARX1 I_1971  ( .D(I36222), .CLK(I2702), .RSTB(I35849), .Q(I35826) );
nor I_1972 (I35841,I36174,I35900);
not I_1973 (I36267,I36174);
nor I_1974 (I36284,I36047,I36267);
and I_1975 (I36301,I35934,I36284);
or I_1976 (I36318,I36129,I36301);
DFFARX1 I_1977  ( .D(I36318), .CLK(I2702), .RSTB(I35849), .Q(I35814) );
nand I_1978 (I35823,I36174,I35996);
nand I_1979 (I35811,I36174,I36078);
not I_1980 (I36410,I2709);
nand I_1981 (I36427,I197235,I197232);
and I_1982 (I36444,I36427,I197229);
DFFARX1 I_1983  ( .D(I36444), .CLK(I2702), .RSTB(I36410), .Q(I36461) );
not I_1984 (I36478,I36461);
nor I_1985 (I36495,I197253,I197232);
or I_1986 (I36393,I36495,I36461);
not I_1987 (I36381,I36495);
DFFARX1 I_1988  ( .D(I197247), .CLK(I2702), .RSTB(I36410), .Q(I36540) );
nor I_1989 (I36557,I36540,I36495);
nand I_1990 (I36574,I197226,I197238);
and I_1991 (I36591,I36574,I197241);
DFFARX1 I_1992  ( .D(I36591), .CLK(I2702), .RSTB(I36410), .Q(I36608) );
nor I_1993 (I36390,I36608,I36461);
not I_1994 (I36639,I36608);
nor I_1995 (I36656,I36540,I36639);
DFFARX1 I_1996  ( .D(I197250), .CLK(I2702), .RSTB(I36410), .Q(I36673) );
and I_1997 (I36690,I36673,I197256);
or I_1998 (I36399,I36690,I36495);
nand I_1999 (I36378,I36690,I36656);
DFFARX1 I_2000  ( .D(I197244), .CLK(I2702), .RSTB(I36410), .Q(I36735) );
and I_2001 (I36752,I36735,I36478);
nor I_2002 (I36396,I36690,I36752);
nor I_2003 (I36783,I36735,I36540);
DFFARX1 I_2004  ( .D(I36783), .CLK(I2702), .RSTB(I36410), .Q(I36387) );
nor I_2005 (I36402,I36735,I36461);
not I_2006 (I36828,I36735);
nor I_2007 (I36845,I36608,I36828);
and I_2008 (I36862,I36495,I36845);
or I_2009 (I36879,I36690,I36862);
DFFARX1 I_2010  ( .D(I36879), .CLK(I2702), .RSTB(I36410), .Q(I36375) );
nand I_2011 (I36384,I36735,I36557);
nand I_2012 (I36372,I36735,I36639);
not I_2013 (I36971,I2709);
nand I_2014 (I36988,I467385,I467382);
and I_2015 (I37005,I36988,I467376);
DFFARX1 I_2016  ( .D(I37005), .CLK(I2702), .RSTB(I36971), .Q(I37022) );
not I_2017 (I37039,I37022);
nor I_2018 (I37056,I467388,I467382);
or I_2019 (I36954,I37056,I37022);
not I_2020 (I36942,I37056);
DFFARX1 I_2021  ( .D(I467400), .CLK(I2702), .RSTB(I36971), .Q(I37101) );
nor I_2022 (I37118,I37101,I37056);
nand I_2023 (I37135,I467391,I467373);
and I_2024 (I37152,I37135,I467403);
DFFARX1 I_2025  ( .D(I37152), .CLK(I2702), .RSTB(I36971), .Q(I37169) );
nor I_2026 (I36951,I37169,I37022);
not I_2027 (I37200,I37169);
nor I_2028 (I37217,I37101,I37200);
DFFARX1 I_2029  ( .D(I467379), .CLK(I2702), .RSTB(I36971), .Q(I37234) );
and I_2030 (I37251,I37234,I467397);
or I_2031 (I36960,I37251,I37056);
nand I_2032 (I36939,I37251,I37217);
DFFARX1 I_2033  ( .D(I467394), .CLK(I2702), .RSTB(I36971), .Q(I37296) );
and I_2034 (I37313,I37296,I37039);
nor I_2035 (I36957,I37251,I37313);
nor I_2036 (I37344,I37296,I37101);
DFFARX1 I_2037  ( .D(I37344), .CLK(I2702), .RSTB(I36971), .Q(I36948) );
nor I_2038 (I36963,I37296,I37022);
not I_2039 (I37389,I37296);
nor I_2040 (I37406,I37169,I37389);
and I_2041 (I37423,I37056,I37406);
or I_2042 (I37440,I37251,I37423);
DFFARX1 I_2043  ( .D(I37440), .CLK(I2702), .RSTB(I36971), .Q(I36936) );
nand I_2044 (I36945,I37296,I37118);
nand I_2045 (I36933,I37296,I37200);
not I_2046 (I37532,I2709);
nand I_2047 (I37549,I457559,I457556);
and I_2048 (I37566,I37549,I457550);
DFFARX1 I_2049  ( .D(I37566), .CLK(I2702), .RSTB(I37532), .Q(I37583) );
not I_2050 (I37600,I37583);
nor I_2051 (I37617,I457562,I457556);
or I_2052 (I37515,I37617,I37583);
not I_2053 (I37503,I37617);
DFFARX1 I_2054  ( .D(I457574), .CLK(I2702), .RSTB(I37532), .Q(I37662) );
nor I_2055 (I37679,I37662,I37617);
nand I_2056 (I37696,I457565,I457547);
and I_2057 (I37713,I37696,I457577);
DFFARX1 I_2058  ( .D(I37713), .CLK(I2702), .RSTB(I37532), .Q(I37730) );
nor I_2059 (I37512,I37730,I37583);
not I_2060 (I37761,I37730);
nor I_2061 (I37778,I37662,I37761);
DFFARX1 I_2062  ( .D(I457553), .CLK(I2702), .RSTB(I37532), .Q(I37795) );
and I_2063 (I37812,I37795,I457571);
or I_2064 (I37521,I37812,I37617);
nand I_2065 (I37500,I37812,I37778);
DFFARX1 I_2066  ( .D(I457568), .CLK(I2702), .RSTB(I37532), .Q(I37857) );
and I_2067 (I37874,I37857,I37600);
nor I_2068 (I37518,I37812,I37874);
nor I_2069 (I37905,I37857,I37662);
DFFARX1 I_2070  ( .D(I37905), .CLK(I2702), .RSTB(I37532), .Q(I37509) );
nor I_2071 (I37524,I37857,I37583);
not I_2072 (I37950,I37857);
nor I_2073 (I37967,I37730,I37950);
and I_2074 (I37984,I37617,I37967);
or I_2075 (I38001,I37812,I37984);
DFFARX1 I_2076  ( .D(I38001), .CLK(I2702), .RSTB(I37532), .Q(I37497) );
nand I_2077 (I37506,I37857,I37679);
nand I_2078 (I37494,I37857,I37761);
not I_2079 (I38093,I2709);
nand I_2080 (I38110,I415646,I415640);
and I_2081 (I38127,I38110,I415652);
DFFARX1 I_2082  ( .D(I38127), .CLK(I2702), .RSTB(I38093), .Q(I38144) );
not I_2083 (I38161,I38144);
nor I_2084 (I38178,I415649,I415640);
or I_2085 (I38076,I38178,I38144);
not I_2086 (I38064,I38178);
DFFARX1 I_2087  ( .D(I415628), .CLK(I2702), .RSTB(I38093), .Q(I38223) );
nor I_2088 (I38240,I38223,I38178);
nand I_2089 (I38257,I415634,I415643);
and I_2090 (I38274,I38257,I415631);
DFFARX1 I_2091  ( .D(I38274), .CLK(I2702), .RSTB(I38093), .Q(I38291) );
nor I_2092 (I38073,I38291,I38144);
not I_2093 (I38322,I38291);
nor I_2094 (I38339,I38223,I38322);
DFFARX1 I_2095  ( .D(I415655), .CLK(I2702), .RSTB(I38093), .Q(I38356) );
and I_2096 (I38373,I38356,I415625);
or I_2097 (I38082,I38373,I38178);
nand I_2098 (I38061,I38373,I38339);
DFFARX1 I_2099  ( .D(I415637), .CLK(I2702), .RSTB(I38093), .Q(I38418) );
and I_2100 (I38435,I38418,I38161);
nor I_2101 (I38079,I38373,I38435);
nor I_2102 (I38466,I38418,I38223);
DFFARX1 I_2103  ( .D(I38466), .CLK(I2702), .RSTB(I38093), .Q(I38070) );
nor I_2104 (I38085,I38418,I38144);
not I_2105 (I38511,I38418);
nor I_2106 (I38528,I38291,I38511);
and I_2107 (I38545,I38178,I38528);
or I_2108 (I38562,I38373,I38545);
DFFARX1 I_2109  ( .D(I38562), .CLK(I2702), .RSTB(I38093), .Q(I38058) );
nand I_2110 (I38067,I38418,I38240);
nand I_2111 (I38055,I38418,I38322);
not I_2112 (I38654,I2709);
nand I_2113 (I38671,I167400,I167397);
and I_2114 (I38688,I38671,I167394);
DFFARX1 I_2115  ( .D(I38688), .CLK(I2702), .RSTB(I38654), .Q(I38705) );
not I_2116 (I38722,I38705);
nor I_2117 (I38739,I167418,I167397);
or I_2118 (I38637,I38739,I38705);
not I_2119 (I38625,I38739);
DFFARX1 I_2120  ( .D(I167412), .CLK(I2702), .RSTB(I38654), .Q(I38784) );
nor I_2121 (I38801,I38784,I38739);
nand I_2122 (I38818,I167391,I167403);
and I_2123 (I38835,I38818,I167406);
DFFARX1 I_2124  ( .D(I38835), .CLK(I2702), .RSTB(I38654), .Q(I38852) );
nor I_2125 (I38634,I38852,I38705);
not I_2126 (I38883,I38852);
nor I_2127 (I38900,I38784,I38883);
DFFARX1 I_2128  ( .D(I167415), .CLK(I2702), .RSTB(I38654), .Q(I38917) );
and I_2129 (I38934,I38917,I167421);
or I_2130 (I38643,I38934,I38739);
nand I_2131 (I38622,I38934,I38900);
DFFARX1 I_2132  ( .D(I167409), .CLK(I2702), .RSTB(I38654), .Q(I38979) );
and I_2133 (I38996,I38979,I38722);
nor I_2134 (I38640,I38934,I38996);
nor I_2135 (I39027,I38979,I38784);
DFFARX1 I_2136  ( .D(I39027), .CLK(I2702), .RSTB(I38654), .Q(I38631) );
nor I_2137 (I38646,I38979,I38705);
not I_2138 (I39072,I38979);
nor I_2139 (I39089,I38852,I39072);
and I_2140 (I39106,I38739,I39089);
or I_2141 (I39123,I38934,I39106);
DFFARX1 I_2142  ( .D(I39123), .CLK(I2702), .RSTB(I38654), .Q(I38619) );
nand I_2143 (I38628,I38979,I38801);
nand I_2144 (I38616,I38979,I38883);
not I_2145 (I39215,I2709);
nand I_2146 (I39232,I203472,I203475);
and I_2147 (I39249,I39232,I203469);
DFFARX1 I_2148  ( .D(I39249), .CLK(I2702), .RSTB(I39215), .Q(I39266) );
not I_2149 (I39283,I39266);
nor I_2150 (I39300,I203460,I203475);
or I_2151 (I39198,I39300,I39266);
not I_2152 (I39186,I39300);
DFFARX1 I_2153  ( .D(I203448), .CLK(I2702), .RSTB(I39215), .Q(I39345) );
nor I_2154 (I39362,I39345,I39300);
nand I_2155 (I39379,I203457,I203451);
and I_2156 (I39396,I39379,I203463);
DFFARX1 I_2157  ( .D(I39396), .CLK(I2702), .RSTB(I39215), .Q(I39413) );
nor I_2158 (I39195,I39413,I39266);
not I_2159 (I39444,I39413);
nor I_2160 (I39461,I39345,I39444);
DFFARX1 I_2161  ( .D(I203478), .CLK(I2702), .RSTB(I39215), .Q(I39478) );
and I_2162 (I39495,I39478,I203466);
or I_2163 (I39204,I39495,I39300);
nand I_2164 (I39183,I39495,I39461);
DFFARX1 I_2165  ( .D(I203454), .CLK(I2702), .RSTB(I39215), .Q(I39540) );
and I_2166 (I39557,I39540,I39283);
nor I_2167 (I39201,I39495,I39557);
nor I_2168 (I39588,I39540,I39345);
DFFARX1 I_2169  ( .D(I39588), .CLK(I2702), .RSTB(I39215), .Q(I39192) );
nor I_2170 (I39207,I39540,I39266);
not I_2171 (I39633,I39540);
nor I_2172 (I39650,I39413,I39633);
and I_2173 (I39667,I39300,I39650);
or I_2174 (I39684,I39495,I39667);
DFFARX1 I_2175  ( .D(I39684), .CLK(I2702), .RSTB(I39215), .Q(I39180) );
nand I_2176 (I39189,I39540,I39362);
nand I_2177 (I39177,I39540,I39444);
not I_2178 (I39776,I2709);
nand I_2179 (I39793,I518512,I518515);
and I_2180 (I39810,I39793,I518527);
DFFARX1 I_2181  ( .D(I39810), .CLK(I2702), .RSTB(I39776), .Q(I39827) );
not I_2182 (I39844,I39827);
nor I_2183 (I39861,I518521,I518515);
or I_2184 (I39759,I39861,I39827);
not I_2185 (I39747,I39861);
DFFARX1 I_2186  ( .D(I518524), .CLK(I2702), .RSTB(I39776), .Q(I39906) );
nor I_2187 (I39923,I39906,I39861);
nand I_2188 (I39940,I518518,I518536);
and I_2189 (I39957,I39940,I518539);
DFFARX1 I_2190  ( .D(I39957), .CLK(I2702), .RSTB(I39776), .Q(I39974) );
nor I_2191 (I39756,I39974,I39827);
not I_2192 (I40005,I39974);
nor I_2193 (I40022,I39906,I40005);
DFFARX1 I_2194  ( .D(I518509), .CLK(I2702), .RSTB(I39776), .Q(I40039) );
and I_2195 (I40056,I40039,I518530);
or I_2196 (I39765,I40056,I39861);
nand I_2197 (I39744,I40056,I40022);
DFFARX1 I_2198  ( .D(I518533), .CLK(I2702), .RSTB(I39776), .Q(I40101) );
and I_2199 (I40118,I40101,I39844);
nor I_2200 (I39762,I40056,I40118);
nor I_2201 (I40149,I40101,I39906);
DFFARX1 I_2202  ( .D(I40149), .CLK(I2702), .RSTB(I39776), .Q(I39753) );
nor I_2203 (I39768,I40101,I39827);
not I_2204 (I40194,I40101);
nor I_2205 (I40211,I39974,I40194);
and I_2206 (I40228,I39861,I40211);
or I_2207 (I40245,I40056,I40228);
DFFARX1 I_2208  ( .D(I40245), .CLK(I2702), .RSTB(I39776), .Q(I39741) );
nand I_2209 (I39750,I40101,I39923);
nand I_2210 (I39738,I40101,I40005);
not I_2211 (I40337,I2709);
nand I_2212 (I40354,I324546,I324537);
and I_2213 (I40371,I40354,I324552);
DFFARX1 I_2214  ( .D(I40371), .CLK(I2702), .RSTB(I40337), .Q(I40388) );
not I_2215 (I40405,I40388);
nor I_2216 (I40422,I324522,I324537);
or I_2217 (I40320,I40422,I40388);
not I_2218 (I40308,I40422);
DFFARX1 I_2219  ( .D(I324525), .CLK(I2702), .RSTB(I40337), .Q(I40467) );
nor I_2220 (I40484,I40467,I40422);
nand I_2221 (I40501,I324543,I324540);
and I_2222 (I40518,I40501,I324528);
DFFARX1 I_2223  ( .D(I40518), .CLK(I2702), .RSTB(I40337), .Q(I40535) );
nor I_2224 (I40317,I40535,I40388);
not I_2225 (I40566,I40535);
nor I_2226 (I40583,I40467,I40566);
DFFARX1 I_2227  ( .D(I324549), .CLK(I2702), .RSTB(I40337), .Q(I40600) );
and I_2228 (I40617,I40600,I324534);
or I_2229 (I40326,I40617,I40422);
nand I_2230 (I40305,I40617,I40583);
DFFARX1 I_2231  ( .D(I324531), .CLK(I2702), .RSTB(I40337), .Q(I40662) );
and I_2232 (I40679,I40662,I40405);
nor I_2233 (I40323,I40617,I40679);
nor I_2234 (I40710,I40662,I40467);
DFFARX1 I_2235  ( .D(I40710), .CLK(I2702), .RSTB(I40337), .Q(I40314) );
nor I_2236 (I40329,I40662,I40388);
not I_2237 (I40755,I40662);
nor I_2238 (I40772,I40535,I40755);
and I_2239 (I40789,I40422,I40772);
or I_2240 (I40806,I40617,I40789);
DFFARX1 I_2241  ( .D(I40806), .CLK(I2702), .RSTB(I40337), .Q(I40302) );
nand I_2242 (I40311,I40662,I40484);
nand I_2243 (I40299,I40662,I40566);
not I_2244 (I40898,I2709);
nand I_2245 (I40915,I243920,I243914);
and I_2246 (I40932,I40915,I243908);
DFFARX1 I_2247  ( .D(I40932), .CLK(I2702), .RSTB(I40898), .Q(I40949) );
not I_2248 (I40966,I40949);
nor I_2249 (I40983,I243935,I243914);
or I_2250 (I40881,I40983,I40949);
not I_2251 (I40869,I40983);
DFFARX1 I_2252  ( .D(I243932), .CLK(I2702), .RSTB(I40898), .Q(I41028) );
nor I_2253 (I41045,I41028,I40983);
nand I_2254 (I41062,I243938,I243926);
and I_2255 (I41079,I41062,I243923);
DFFARX1 I_2256  ( .D(I41079), .CLK(I2702), .RSTB(I40898), .Q(I41096) );
nor I_2257 (I40878,I41096,I40949);
not I_2258 (I41127,I41096);
nor I_2259 (I41144,I41028,I41127);
DFFARX1 I_2260  ( .D(I243911), .CLK(I2702), .RSTB(I40898), .Q(I41161) );
and I_2261 (I41178,I41161,I243929);
or I_2262 (I40887,I41178,I40983);
nand I_2263 (I40866,I41178,I41144);
DFFARX1 I_2264  ( .D(I243917), .CLK(I2702), .RSTB(I40898), .Q(I41223) );
and I_2265 (I41240,I41223,I40966);
nor I_2266 (I40884,I41178,I41240);
nor I_2267 (I41271,I41223,I41028);
DFFARX1 I_2268  ( .D(I41271), .CLK(I2702), .RSTB(I40898), .Q(I40875) );
nor I_2269 (I40890,I41223,I40949);
not I_2270 (I41316,I41223);
nor I_2271 (I41333,I41096,I41316);
and I_2272 (I41350,I40983,I41333);
or I_2273 (I41367,I41178,I41350);
DFFARX1 I_2274  ( .D(I41367), .CLK(I2702), .RSTB(I40898), .Q(I40863) );
nand I_2275 (I40872,I41223,I41045);
nand I_2276 (I40860,I41223,I41127);
not I_2277 (I41459,I2709);
nand I_2278 (I41476,I501981,I501975);
and I_2279 (I41493,I41476,I501966);
DFFARX1 I_2280  ( .D(I41493), .CLK(I2702), .RSTB(I41459), .Q(I41510) );
not I_2281 (I41527,I41510);
nor I_2282 (I41544,I501957,I501975);
or I_2283 (I41442,I41544,I41510);
not I_2284 (I41430,I41544);
DFFARX1 I_2285  ( .D(I501972), .CLK(I2702), .RSTB(I41459), .Q(I41589) );
nor I_2286 (I41606,I41589,I41544);
nand I_2287 (I41623,I501963,I501978);
and I_2288 (I41640,I41623,I501960);
DFFARX1 I_2289  ( .D(I41640), .CLK(I2702), .RSTB(I41459), .Q(I41657) );
nor I_2290 (I41439,I41657,I41510);
not I_2291 (I41688,I41657);
nor I_2292 (I41705,I41589,I41688);
DFFARX1 I_2293  ( .D(I501969), .CLK(I2702), .RSTB(I41459), .Q(I41722) );
and I_2294 (I41739,I41722,I501951);
or I_2295 (I41448,I41739,I41544);
nand I_2296 (I41427,I41739,I41705);
DFFARX1 I_2297  ( .D(I501954), .CLK(I2702), .RSTB(I41459), .Q(I41784) );
and I_2298 (I41801,I41784,I41527);
nor I_2299 (I41445,I41739,I41801);
nor I_2300 (I41832,I41784,I41589);
DFFARX1 I_2301  ( .D(I41832), .CLK(I2702), .RSTB(I41459), .Q(I41436) );
nor I_2302 (I41451,I41784,I41510);
not I_2303 (I41877,I41784);
nor I_2304 (I41894,I41657,I41877);
and I_2305 (I41911,I41544,I41894);
or I_2306 (I41928,I41739,I41911);
DFFARX1 I_2307  ( .D(I41928), .CLK(I2702), .RSTB(I41459), .Q(I41424) );
nand I_2308 (I41433,I41784,I41606);
nand I_2309 (I41421,I41784,I41688);
not I_2310 (I42020,I2709);
nand I_2311 (I42037,I589930,I589918);
and I_2312 (I42054,I42037,I589915);
DFFARX1 I_2313  ( .D(I42054), .CLK(I2702), .RSTB(I42020), .Q(I42071) );
not I_2314 (I42088,I42071);
nor I_2315 (I42105,I589936,I589918);
or I_2316 (I42003,I42105,I42071);
not I_2317 (I41991,I42105);
DFFARX1 I_2318  ( .D(I589939), .CLK(I2702), .RSTB(I42020), .Q(I42150) );
nor I_2319 (I42167,I42150,I42105);
nand I_2320 (I42184,I589909,I589927);
and I_2321 (I42201,I42184,I589924);
DFFARX1 I_2322  ( .D(I42201), .CLK(I2702), .RSTB(I42020), .Q(I42218) );
nor I_2323 (I42000,I42218,I42071);
not I_2324 (I42249,I42218);
nor I_2325 (I42266,I42150,I42249);
DFFARX1 I_2326  ( .D(I589933), .CLK(I2702), .RSTB(I42020), .Q(I42283) );
and I_2327 (I42300,I42283,I589921);
or I_2328 (I42009,I42300,I42105);
nand I_2329 (I41988,I42300,I42266);
DFFARX1 I_2330  ( .D(I589912), .CLK(I2702), .RSTB(I42020), .Q(I42345) );
and I_2331 (I42362,I42345,I42088);
nor I_2332 (I42006,I42300,I42362);
nor I_2333 (I42393,I42345,I42150);
DFFARX1 I_2334  ( .D(I42393), .CLK(I2702), .RSTB(I42020), .Q(I41997) );
nor I_2335 (I42012,I42345,I42071);
not I_2336 (I42438,I42345);
nor I_2337 (I42455,I42218,I42438);
and I_2338 (I42472,I42105,I42455);
or I_2339 (I42489,I42300,I42472);
DFFARX1 I_2340  ( .D(I42489), .CLK(I2702), .RSTB(I42020), .Q(I41985) );
nand I_2341 (I41994,I42345,I42167);
nand I_2342 (I41982,I42345,I42249);
not I_2343 (I42581,I2709);
nand I_2344 (I42598,I698463,I698484);
and I_2345 (I42615,I42598,I698472);
DFFARX1 I_2346  ( .D(I42615), .CLK(I2702), .RSTB(I42581), .Q(I42632) );
not I_2347 (I42649,I42632);
nor I_2348 (I42666,I698478,I698484);
or I_2349 (I42564,I42666,I42632);
not I_2350 (I42552,I42666);
DFFARX1 I_2351  ( .D(I698466), .CLK(I2702), .RSTB(I42581), .Q(I42711) );
nor I_2352 (I42728,I42711,I42666);
nand I_2353 (I42745,I698457,I698475);
and I_2354 (I42762,I42745,I698469);
DFFARX1 I_2355  ( .D(I42762), .CLK(I2702), .RSTB(I42581), .Q(I42779) );
nor I_2356 (I42561,I42779,I42632);
not I_2357 (I42810,I42779);
nor I_2358 (I42827,I42711,I42810);
DFFARX1 I_2359  ( .D(I698481), .CLK(I2702), .RSTB(I42581), .Q(I42844) );
and I_2360 (I42861,I42844,I698454);
or I_2361 (I42570,I42861,I42666);
nand I_2362 (I42549,I42861,I42827);
DFFARX1 I_2363  ( .D(I698460), .CLK(I2702), .RSTB(I42581), .Q(I42906) );
and I_2364 (I42923,I42906,I42649);
nor I_2365 (I42567,I42861,I42923);
nor I_2366 (I42954,I42906,I42711);
DFFARX1 I_2367  ( .D(I42954), .CLK(I2702), .RSTB(I42581), .Q(I42558) );
nor I_2368 (I42573,I42906,I42632);
not I_2369 (I42999,I42906);
nor I_2370 (I43016,I42779,I42999);
and I_2371 (I43033,I42666,I43016);
or I_2372 (I43050,I42861,I43033);
DFFARX1 I_2373  ( .D(I43050), .CLK(I2702), .RSTB(I42581), .Q(I42546) );
nand I_2374 (I42555,I42906,I42728);
nand I_2375 (I42543,I42906,I42810);
not I_2376 (I43142,I2709);
nand I_2377 (I43159,I666511,I666514);
and I_2378 (I43176,I43159,I666520);
DFFARX1 I_2379  ( .D(I43176), .CLK(I2702), .RSTB(I43142), .Q(I43193) );
not I_2380 (I43210,I43193);
nor I_2381 (I43227,I666532,I666514);
or I_2382 (I43125,I43227,I43193);
not I_2383 (I43113,I43227);
DFFARX1 I_2384  ( .D(I666541), .CLK(I2702), .RSTB(I43142), .Q(I43272) );
nor I_2385 (I43289,I43272,I43227);
nand I_2386 (I43306,I666529,I666526);
and I_2387 (I43323,I43306,I666538);
DFFARX1 I_2388  ( .D(I43323), .CLK(I2702), .RSTB(I43142), .Q(I43340) );
nor I_2389 (I43122,I43340,I43193);
not I_2390 (I43371,I43340);
nor I_2391 (I43388,I43272,I43371);
DFFARX1 I_2392  ( .D(I666535), .CLK(I2702), .RSTB(I43142), .Q(I43405) );
and I_2393 (I43422,I43405,I666523);
or I_2394 (I43131,I43422,I43227);
nand I_2395 (I43110,I43422,I43388);
DFFARX1 I_2396  ( .D(I666517), .CLK(I2702), .RSTB(I43142), .Q(I43467) );
and I_2397 (I43484,I43467,I43210);
nor I_2398 (I43128,I43422,I43484);
nor I_2399 (I43515,I43467,I43272);
DFFARX1 I_2400  ( .D(I43515), .CLK(I2702), .RSTB(I43142), .Q(I43119) );
nor I_2401 (I43134,I43467,I43193);
not I_2402 (I43560,I43467);
nor I_2403 (I43577,I43340,I43560);
and I_2404 (I43594,I43227,I43577);
or I_2405 (I43611,I43422,I43594);
DFFARX1 I_2406  ( .D(I43611), .CLK(I2702), .RSTB(I43142), .Q(I43107) );
nand I_2407 (I43116,I43467,I43289);
nand I_2408 (I43104,I43467,I43371);
not I_2409 (I43703,I2709);
nand I_2410 (I43720,I159444,I159441);
and I_2411 (I43737,I43720,I159438);
DFFARX1 I_2412  ( .D(I43737), .CLK(I2702), .RSTB(I43703), .Q(I43754) );
not I_2413 (I43771,I43754);
nor I_2414 (I43788,I159462,I159441);
or I_2415 (I43686,I43788,I43754);
not I_2416 (I43674,I43788);
DFFARX1 I_2417  ( .D(I159456), .CLK(I2702), .RSTB(I43703), .Q(I43833) );
nor I_2418 (I43850,I43833,I43788);
nand I_2419 (I43867,I159435,I159447);
and I_2420 (I43884,I43867,I159450);
DFFARX1 I_2421  ( .D(I43884), .CLK(I2702), .RSTB(I43703), .Q(I43901) );
nor I_2422 (I43683,I43901,I43754);
not I_2423 (I43932,I43901);
nor I_2424 (I43949,I43833,I43932);
DFFARX1 I_2425  ( .D(I159459), .CLK(I2702), .RSTB(I43703), .Q(I43966) );
and I_2426 (I43983,I43966,I159465);
or I_2427 (I43692,I43983,I43788);
nand I_2428 (I43671,I43983,I43949);
DFFARX1 I_2429  ( .D(I159453), .CLK(I2702), .RSTB(I43703), .Q(I44028) );
and I_2430 (I44045,I44028,I43771);
nor I_2431 (I43689,I43983,I44045);
nor I_2432 (I44076,I44028,I43833);
DFFARX1 I_2433  ( .D(I44076), .CLK(I2702), .RSTB(I43703), .Q(I43680) );
nor I_2434 (I43695,I44028,I43754);
not I_2435 (I44121,I44028);
nor I_2436 (I44138,I43901,I44121);
and I_2437 (I44155,I43788,I44138);
or I_2438 (I44172,I43983,I44155);
DFFARX1 I_2439  ( .D(I44172), .CLK(I2702), .RSTB(I43703), .Q(I43668) );
nand I_2440 (I43677,I44028,I43850);
nand I_2441 (I43665,I44028,I43932);
not I_2442 (I44264,I2709);
nand I_2443 (I44281,I424826,I424820);
and I_2444 (I44298,I44281,I424832);
DFFARX1 I_2445  ( .D(I44298), .CLK(I2702), .RSTB(I44264), .Q(I44315) );
not I_2446 (I44332,I44315);
nor I_2447 (I44349,I424829,I424820);
or I_2448 (I44247,I44349,I44315);
not I_2449 (I44235,I44349);
DFFARX1 I_2450  ( .D(I424808), .CLK(I2702), .RSTB(I44264), .Q(I44394) );
nor I_2451 (I44411,I44394,I44349);
nand I_2452 (I44428,I424814,I424823);
and I_2453 (I44445,I44428,I424811);
DFFARX1 I_2454  ( .D(I44445), .CLK(I2702), .RSTB(I44264), .Q(I44462) );
nor I_2455 (I44244,I44462,I44315);
not I_2456 (I44493,I44462);
nor I_2457 (I44510,I44394,I44493);
DFFARX1 I_2458  ( .D(I424835), .CLK(I2702), .RSTB(I44264), .Q(I44527) );
and I_2459 (I44544,I44527,I424805);
or I_2460 (I44253,I44544,I44349);
nand I_2461 (I44232,I44544,I44510);
DFFARX1 I_2462  ( .D(I424817), .CLK(I2702), .RSTB(I44264), .Q(I44589) );
and I_2463 (I44606,I44589,I44332);
nor I_2464 (I44250,I44544,I44606);
nor I_2465 (I44637,I44589,I44394);
DFFARX1 I_2466  ( .D(I44637), .CLK(I2702), .RSTB(I44264), .Q(I44241) );
nor I_2467 (I44256,I44589,I44315);
not I_2468 (I44682,I44589);
nor I_2469 (I44699,I44462,I44682);
and I_2470 (I44716,I44349,I44699);
or I_2471 (I44733,I44544,I44716);
DFFARX1 I_2472  ( .D(I44733), .CLK(I2702), .RSTB(I44264), .Q(I44229) );
nand I_2473 (I44238,I44589,I44411);
nand I_2474 (I44226,I44589,I44493);
not I_2475 (I44825,I2709);
nand I_2476 (I44842,I331839,I331830);
and I_2477 (I44859,I44842,I331845);
DFFARX1 I_2478  ( .D(I44859), .CLK(I2702), .RSTB(I44825), .Q(I44876) );
not I_2479 (I44893,I44876);
nor I_2480 (I44910,I331815,I331830);
or I_2481 (I44808,I44910,I44876);
not I_2482 (I44796,I44910);
DFFARX1 I_2483  ( .D(I331818), .CLK(I2702), .RSTB(I44825), .Q(I44955) );
nor I_2484 (I44972,I44955,I44910);
nand I_2485 (I44989,I331836,I331833);
and I_2486 (I45006,I44989,I331821);
DFFARX1 I_2487  ( .D(I45006), .CLK(I2702), .RSTB(I44825), .Q(I45023) );
nor I_2488 (I44805,I45023,I44876);
not I_2489 (I45054,I45023);
nor I_2490 (I45071,I44955,I45054);
DFFARX1 I_2491  ( .D(I331842), .CLK(I2702), .RSTB(I44825), .Q(I45088) );
and I_2492 (I45105,I45088,I331827);
or I_2493 (I44814,I45105,I44910);
nand I_2494 (I44793,I45105,I45071);
DFFARX1 I_2495  ( .D(I331824), .CLK(I2702), .RSTB(I44825), .Q(I45150) );
and I_2496 (I45167,I45150,I44893);
nor I_2497 (I44811,I45105,I45167);
nor I_2498 (I45198,I45150,I44955);
DFFARX1 I_2499  ( .D(I45198), .CLK(I2702), .RSTB(I44825), .Q(I44802) );
nor I_2500 (I44817,I45150,I44876);
not I_2501 (I45243,I45150);
nor I_2502 (I45260,I45023,I45243);
and I_2503 (I45277,I44910,I45260);
or I_2504 (I45294,I45105,I45277);
DFFARX1 I_2505  ( .D(I45294), .CLK(I2702), .RSTB(I44825), .Q(I44790) );
nand I_2506 (I44799,I45150,I44972);
nand I_2507 (I44787,I45150,I45054);
not I_2508 (I45386,I2709);
nand I_2509 (I45403,I587550,I587538);
and I_2510 (I45420,I45403,I587535);
DFFARX1 I_2511  ( .D(I45420), .CLK(I2702), .RSTB(I45386), .Q(I45437) );
not I_2512 (I45454,I45437);
nor I_2513 (I45471,I587556,I587538);
or I_2514 (I45369,I45471,I45437);
not I_2515 (I45357,I45471);
DFFARX1 I_2516  ( .D(I587559), .CLK(I2702), .RSTB(I45386), .Q(I45516) );
nor I_2517 (I45533,I45516,I45471);
nand I_2518 (I45550,I587529,I587547);
and I_2519 (I45567,I45550,I587544);
DFFARX1 I_2520  ( .D(I45567), .CLK(I2702), .RSTB(I45386), .Q(I45584) );
nor I_2521 (I45366,I45584,I45437);
not I_2522 (I45615,I45584);
nor I_2523 (I45632,I45516,I45615);
DFFARX1 I_2524  ( .D(I587553), .CLK(I2702), .RSTB(I45386), .Q(I45649) );
and I_2525 (I45666,I45649,I587541);
or I_2526 (I45375,I45666,I45471);
nand I_2527 (I45354,I45666,I45632);
DFFARX1 I_2528  ( .D(I587532), .CLK(I2702), .RSTB(I45386), .Q(I45711) );
and I_2529 (I45728,I45711,I45454);
nor I_2530 (I45372,I45666,I45728);
nor I_2531 (I45759,I45711,I45516);
DFFARX1 I_2532  ( .D(I45759), .CLK(I2702), .RSTB(I45386), .Q(I45363) );
nor I_2533 (I45378,I45711,I45437);
not I_2534 (I45804,I45711);
nor I_2535 (I45821,I45584,I45804);
and I_2536 (I45838,I45471,I45821);
or I_2537 (I45855,I45666,I45838);
DFFARX1 I_2538  ( .D(I45855), .CLK(I2702), .RSTB(I45386), .Q(I45351) );
nand I_2539 (I45360,I45711,I45533);
nand I_2540 (I45348,I45711,I45615);
not I_2541 (I45947,I2709);
nand I_2542 (I45964,I499669,I499663);
and I_2543 (I45981,I45964,I499654);
DFFARX1 I_2544  ( .D(I45981), .CLK(I2702), .RSTB(I45947), .Q(I45998) );
not I_2545 (I46015,I45998);
nor I_2546 (I46032,I499645,I499663);
or I_2547 (I45930,I46032,I45998);
not I_2548 (I45918,I46032);
DFFARX1 I_2549  ( .D(I499660), .CLK(I2702), .RSTB(I45947), .Q(I46077) );
nor I_2550 (I46094,I46077,I46032);
nand I_2551 (I46111,I499651,I499666);
and I_2552 (I46128,I46111,I499648);
DFFARX1 I_2553  ( .D(I46128), .CLK(I2702), .RSTB(I45947), .Q(I46145) );
nor I_2554 (I45927,I46145,I45998);
not I_2555 (I46176,I46145);
nor I_2556 (I46193,I46077,I46176);
DFFARX1 I_2557  ( .D(I499657), .CLK(I2702), .RSTB(I45947), .Q(I46210) );
and I_2558 (I46227,I46210,I499639);
or I_2559 (I45936,I46227,I46032);
nand I_2560 (I45915,I46227,I46193);
DFFARX1 I_2561  ( .D(I499642), .CLK(I2702), .RSTB(I45947), .Q(I46272) );
and I_2562 (I46289,I46272,I46015);
nor I_2563 (I45933,I46227,I46289);
nor I_2564 (I46320,I46272,I46077);
DFFARX1 I_2565  ( .D(I46320), .CLK(I2702), .RSTB(I45947), .Q(I45924) );
nor I_2566 (I45939,I46272,I45998);
not I_2567 (I46365,I46272);
nor I_2568 (I46382,I46145,I46365);
and I_2569 (I46399,I46032,I46382);
or I_2570 (I46416,I46227,I46399);
DFFARX1 I_2571  ( .D(I46416), .CLK(I2702), .RSTB(I45947), .Q(I45912) );
nand I_2572 (I45921,I46272,I46094);
nand I_2573 (I45909,I46272,I46176);
not I_2574 (I46508,I2709);
nand I_2575 (I46525,I515537,I515540);
and I_2576 (I46542,I46525,I515552);
DFFARX1 I_2577  ( .D(I46542), .CLK(I2702), .RSTB(I46508), .Q(I46559) );
not I_2578 (I46576,I46559);
nor I_2579 (I46593,I515546,I515540);
or I_2580 (I46491,I46593,I46559);
not I_2581 (I46479,I46593);
DFFARX1 I_2582  ( .D(I515549), .CLK(I2702), .RSTB(I46508), .Q(I46638) );
nor I_2583 (I46655,I46638,I46593);
nand I_2584 (I46672,I515543,I515561);
and I_2585 (I46689,I46672,I515564);
DFFARX1 I_2586  ( .D(I46689), .CLK(I2702), .RSTB(I46508), .Q(I46706) );
nor I_2587 (I46488,I46706,I46559);
not I_2588 (I46737,I46706);
nor I_2589 (I46754,I46638,I46737);
DFFARX1 I_2590  ( .D(I515534), .CLK(I2702), .RSTB(I46508), .Q(I46771) );
and I_2591 (I46788,I46771,I515555);
or I_2592 (I46497,I46788,I46593);
nand I_2593 (I46476,I46788,I46754);
DFFARX1 I_2594  ( .D(I515558), .CLK(I2702), .RSTB(I46508), .Q(I46833) );
and I_2595 (I46850,I46833,I46576);
nor I_2596 (I46494,I46788,I46850);
nor I_2597 (I46881,I46833,I46638);
DFFARX1 I_2598  ( .D(I46881), .CLK(I2702), .RSTB(I46508), .Q(I46485) );
nor I_2599 (I46500,I46833,I46559);
not I_2600 (I46926,I46833);
nor I_2601 (I46943,I46706,I46926);
and I_2602 (I46960,I46593,I46943);
or I_2603 (I46977,I46788,I46960);
DFFARX1 I_2604  ( .D(I46977), .CLK(I2702), .RSTB(I46508), .Q(I46473) );
nand I_2605 (I46482,I46833,I46655);
nand I_2606 (I46470,I46833,I46737);
not I_2607 (I47069,I2709);
nand I_2608 (I47086,I201092,I201095);
and I_2609 (I47103,I47086,I201089);
DFFARX1 I_2610  ( .D(I47103), .CLK(I2702), .RSTB(I47069), .Q(I47120) );
not I_2611 (I47137,I47120);
nor I_2612 (I47154,I201080,I201095);
or I_2613 (I47052,I47154,I47120);
not I_2614 (I47040,I47154);
DFFARX1 I_2615  ( .D(I201068), .CLK(I2702), .RSTB(I47069), .Q(I47199) );
nor I_2616 (I47216,I47199,I47154);
nand I_2617 (I47233,I201077,I201071);
and I_2618 (I47250,I47233,I201083);
DFFARX1 I_2619  ( .D(I47250), .CLK(I2702), .RSTB(I47069), .Q(I47267) );
nor I_2620 (I47049,I47267,I47120);
not I_2621 (I47298,I47267);
nor I_2622 (I47315,I47199,I47298);
DFFARX1 I_2623  ( .D(I201098), .CLK(I2702), .RSTB(I47069), .Q(I47332) );
and I_2624 (I47349,I47332,I201086);
or I_2625 (I47058,I47349,I47154);
nand I_2626 (I47037,I47349,I47315);
DFFARX1 I_2627  ( .D(I201074), .CLK(I2702), .RSTB(I47069), .Q(I47394) );
and I_2628 (I47411,I47394,I47137);
nor I_2629 (I47055,I47349,I47411);
nor I_2630 (I47442,I47394,I47199);
DFFARX1 I_2631  ( .D(I47442), .CLK(I2702), .RSTB(I47069), .Q(I47046) );
nor I_2632 (I47061,I47394,I47120);
not I_2633 (I47487,I47394);
nor I_2634 (I47504,I47267,I47487);
and I_2635 (I47521,I47154,I47504);
or I_2636 (I47538,I47349,I47521);
DFFARX1 I_2637  ( .D(I47538), .CLK(I2702), .RSTB(I47069), .Q(I47034) );
nand I_2638 (I47043,I47394,I47216);
nand I_2639 (I47031,I47394,I47298);
not I_2640 (I47630,I2709);
nand I_2641 (I47647,I614304,I614307);
and I_2642 (I47664,I47647,I614313);
DFFARX1 I_2643  ( .D(I47664), .CLK(I2702), .RSTB(I47630), .Q(I47681) );
not I_2644 (I47698,I47681);
nor I_2645 (I47715,I614325,I614307);
or I_2646 (I47613,I47715,I47681);
not I_2647 (I47601,I47715);
DFFARX1 I_2648  ( .D(I614334), .CLK(I2702), .RSTB(I47630), .Q(I47760) );
nor I_2649 (I47777,I47760,I47715);
nand I_2650 (I47794,I614322,I614319);
and I_2651 (I47811,I47794,I614331);
DFFARX1 I_2652  ( .D(I47811), .CLK(I2702), .RSTB(I47630), .Q(I47828) );
nor I_2653 (I47610,I47828,I47681);
not I_2654 (I47859,I47828);
nor I_2655 (I47876,I47760,I47859);
DFFARX1 I_2656  ( .D(I614328), .CLK(I2702), .RSTB(I47630), .Q(I47893) );
and I_2657 (I47910,I47893,I614316);
or I_2658 (I47619,I47910,I47715);
nand I_2659 (I47598,I47910,I47876);
DFFARX1 I_2660  ( .D(I614310), .CLK(I2702), .RSTB(I47630), .Q(I47955) );
and I_2661 (I47972,I47955,I47698);
nor I_2662 (I47616,I47910,I47972);
nor I_2663 (I48003,I47955,I47760);
DFFARX1 I_2664  ( .D(I48003), .CLK(I2702), .RSTB(I47630), .Q(I47607) );
nor I_2665 (I47622,I47955,I47681);
not I_2666 (I48048,I47955);
nor I_2667 (I48065,I47828,I48048);
and I_2668 (I48082,I47715,I48065);
or I_2669 (I48099,I47910,I48082);
DFFARX1 I_2670  ( .D(I48099), .CLK(I2702), .RSTB(I47630), .Q(I47595) );
nand I_2671 (I47604,I47955,I47777);
nand I_2672 (I47592,I47955,I47859);
not I_2673 (I48191,I2709);
nand I_2674 (I48208,I426662,I426656);
and I_2675 (I48225,I48208,I426668);
DFFARX1 I_2676  ( .D(I48225), .CLK(I2702), .RSTB(I48191), .Q(I48242) );
not I_2677 (I48259,I48242);
nor I_2678 (I48276,I426665,I426656);
or I_2679 (I48174,I48276,I48242);
not I_2680 (I48162,I48276);
DFFARX1 I_2681  ( .D(I426644), .CLK(I2702), .RSTB(I48191), .Q(I48321) );
nor I_2682 (I48338,I48321,I48276);
nand I_2683 (I48355,I426650,I426659);
and I_2684 (I48372,I48355,I426647);
DFFARX1 I_2685  ( .D(I48372), .CLK(I2702), .RSTB(I48191), .Q(I48389) );
nor I_2686 (I48171,I48389,I48242);
not I_2687 (I48420,I48389);
nor I_2688 (I48437,I48321,I48420);
DFFARX1 I_2689  ( .D(I426671), .CLK(I2702), .RSTB(I48191), .Q(I48454) );
and I_2690 (I48471,I48454,I426641);
or I_2691 (I48180,I48471,I48276);
nand I_2692 (I48159,I48471,I48437);
DFFARX1 I_2693  ( .D(I426653), .CLK(I2702), .RSTB(I48191), .Q(I48516) );
and I_2694 (I48533,I48516,I48259);
nor I_2695 (I48177,I48471,I48533);
nor I_2696 (I48564,I48516,I48321);
DFFARX1 I_2697  ( .D(I48564), .CLK(I2702), .RSTB(I48191), .Q(I48168) );
nor I_2698 (I48183,I48516,I48242);
not I_2699 (I48609,I48516);
nor I_2700 (I48626,I48389,I48609);
and I_2701 (I48643,I48276,I48626);
or I_2702 (I48660,I48471,I48643);
DFFARX1 I_2703  ( .D(I48660), .CLK(I2702), .RSTB(I48191), .Q(I48156) );
nand I_2704 (I48165,I48516,I48338);
nand I_2705 (I48153,I48516,I48420);
not I_2706 (I48752,I2709);
nand I_2707 (I48769,I434439,I434436);
and I_2708 (I48786,I48769,I434430);
DFFARX1 I_2709  ( .D(I48786), .CLK(I2702), .RSTB(I48752), .Q(I48803) );
not I_2710 (I48820,I48803);
nor I_2711 (I48837,I434442,I434436);
or I_2712 (I48735,I48837,I48803);
not I_2713 (I48723,I48837);
DFFARX1 I_2714  ( .D(I434454), .CLK(I2702), .RSTB(I48752), .Q(I48882) );
nor I_2715 (I48899,I48882,I48837);
nand I_2716 (I48916,I434445,I434427);
and I_2717 (I48933,I48916,I434457);
DFFARX1 I_2718  ( .D(I48933), .CLK(I2702), .RSTB(I48752), .Q(I48950) );
nor I_2719 (I48732,I48950,I48803);
not I_2720 (I48981,I48950);
nor I_2721 (I48998,I48882,I48981);
DFFARX1 I_2722  ( .D(I434433), .CLK(I2702), .RSTB(I48752), .Q(I49015) );
and I_2723 (I49032,I49015,I434451);
or I_2724 (I48741,I49032,I48837);
nand I_2725 (I48720,I49032,I48998);
DFFARX1 I_2726  ( .D(I434448), .CLK(I2702), .RSTB(I48752), .Q(I49077) );
and I_2727 (I49094,I49077,I48820);
nor I_2728 (I48738,I49032,I49094);
nor I_2729 (I49125,I49077,I48882);
DFFARX1 I_2730  ( .D(I49125), .CLK(I2702), .RSTB(I48752), .Q(I48729) );
nor I_2731 (I48744,I49077,I48803);
not I_2732 (I49170,I49077);
nor I_2733 (I49187,I48950,I49170);
and I_2734 (I49204,I48837,I49187);
or I_2735 (I49221,I49032,I49204);
DFFARX1 I_2736  ( .D(I49221), .CLK(I2702), .RSTB(I48752), .Q(I48717) );
nand I_2737 (I48726,I49077,I48899);
nand I_2738 (I48714,I49077,I48981);
not I_2739 (I49313,I2709);
nand I_2740 (I49330,I190605,I190602);
and I_2741 (I49347,I49330,I190599);
DFFARX1 I_2742  ( .D(I49347), .CLK(I2702), .RSTB(I49313), .Q(I49364) );
not I_2743 (I49381,I49364);
nor I_2744 (I49398,I190623,I190602);
or I_2745 (I49296,I49398,I49364);
not I_2746 (I49284,I49398);
DFFARX1 I_2747  ( .D(I190617), .CLK(I2702), .RSTB(I49313), .Q(I49443) );
nor I_2748 (I49460,I49443,I49398);
nand I_2749 (I49477,I190596,I190608);
and I_2750 (I49494,I49477,I190611);
DFFARX1 I_2751  ( .D(I49494), .CLK(I2702), .RSTB(I49313), .Q(I49511) );
nor I_2752 (I49293,I49511,I49364);
not I_2753 (I49542,I49511);
nor I_2754 (I49559,I49443,I49542);
DFFARX1 I_2755  ( .D(I190620), .CLK(I2702), .RSTB(I49313), .Q(I49576) );
and I_2756 (I49593,I49576,I190626);
or I_2757 (I49302,I49593,I49398);
nand I_2758 (I49281,I49593,I49559);
DFFARX1 I_2759  ( .D(I190614), .CLK(I2702), .RSTB(I49313), .Q(I49638) );
and I_2760 (I49655,I49638,I49381);
nor I_2761 (I49299,I49593,I49655);
nor I_2762 (I49686,I49638,I49443);
DFFARX1 I_2763  ( .D(I49686), .CLK(I2702), .RSTB(I49313), .Q(I49290) );
nor I_2764 (I49305,I49638,I49364);
not I_2765 (I49731,I49638);
nor I_2766 (I49748,I49511,I49731);
and I_2767 (I49765,I49398,I49748);
or I_2768 (I49782,I49593,I49765);
DFFARX1 I_2769  ( .D(I49782), .CLK(I2702), .RSTB(I49313), .Q(I49278) );
nand I_2770 (I49287,I49638,I49460);
nand I_2771 (I49275,I49638,I49542);
not I_2772 (I49874,I2709);
nand I_2773 (I49891,I711757,I711778);
and I_2774 (I49908,I49891,I711766);
DFFARX1 I_2775  ( .D(I49908), .CLK(I2702), .RSTB(I49874), .Q(I49925) );
not I_2776 (I49942,I49925);
nor I_2777 (I49959,I711772,I711778);
or I_2778 (I49857,I49959,I49925);
not I_2779 (I49845,I49959);
DFFARX1 I_2780  ( .D(I711760), .CLK(I2702), .RSTB(I49874), .Q(I50004) );
nor I_2781 (I50021,I50004,I49959);
nand I_2782 (I50038,I711751,I711769);
and I_2783 (I50055,I50038,I711763);
DFFARX1 I_2784  ( .D(I50055), .CLK(I2702), .RSTB(I49874), .Q(I50072) );
nor I_2785 (I49854,I50072,I49925);
not I_2786 (I50103,I50072);
nor I_2787 (I50120,I50004,I50103);
DFFARX1 I_2788  ( .D(I711775), .CLK(I2702), .RSTB(I49874), .Q(I50137) );
and I_2789 (I50154,I50137,I711748);
or I_2790 (I49863,I50154,I49959);
nand I_2791 (I49842,I50154,I50120);
DFFARX1 I_2792  ( .D(I711754), .CLK(I2702), .RSTB(I49874), .Q(I50199) );
and I_2793 (I50216,I50199,I49942);
nor I_2794 (I49860,I50154,I50216);
nor I_2795 (I50247,I50199,I50004);
DFFARX1 I_2796  ( .D(I50247), .CLK(I2702), .RSTB(I49874), .Q(I49851) );
nor I_2797 (I49866,I50199,I49925);
not I_2798 (I50292,I50199);
nor I_2799 (I50309,I50072,I50292);
and I_2800 (I50326,I49959,I50309);
or I_2801 (I50343,I50154,I50326);
DFFARX1 I_2802  ( .D(I50343), .CLK(I2702), .RSTB(I49874), .Q(I49839) );
nand I_2803 (I49848,I50199,I50021);
nand I_2804 (I49836,I50199,I50103);
not I_2805 (I50435,I2709);
not I_2806 (I50452,I707133);
nor I_2807 (I50469,I707130,I707127);
nand I_2808 (I50486,I50469,I707148);
DFFARX1 I_2809  ( .D(I50486), .CLK(I2702), .RSTB(I50435), .Q(I50409) );
nor I_2810 (I50517,I50452,I707130);
nand I_2811 (I50534,I50517,I707151);
not I_2812 (I50424,I50534);
DFFARX1 I_2813  ( .D(I50534), .CLK(I2702), .RSTB(I50435), .Q(I50406) );
not I_2814 (I50579,I707130);
not I_2815 (I50596,I50579);
not I_2816 (I50613,I707124);
nor I_2817 (I50630,I50613,I707136);
and I_2818 (I50647,I50630,I707145);
or I_2819 (I50664,I50647,I707139);
DFFARX1 I_2820  ( .D(I50664), .CLK(I2702), .RSTB(I50435), .Q(I50681) );
nor I_2821 (I50698,I50681,I50534);
nor I_2822 (I50715,I50681,I50596);
nand I_2823 (I50421,I50486,I50715);
nand I_2824 (I50746,I50452,I707124);
nand I_2825 (I50763,I50746,I50681);
and I_2826 (I50780,I50746,I50763);
DFFARX1 I_2827  ( .D(I50780), .CLK(I2702), .RSTB(I50435), .Q(I50403) );
DFFARX1 I_2828  ( .D(I50746), .CLK(I2702), .RSTB(I50435), .Q(I50811) );
and I_2829 (I50400,I50579,I50811);
DFFARX1 I_2830  ( .D(I707154), .CLK(I2702), .RSTB(I50435), .Q(I50842) );
not I_2831 (I50859,I50842);
nor I_2832 (I50876,I50534,I50859);
and I_2833 (I50893,I50842,I50876);
nand I_2834 (I50415,I50842,I50596);
DFFARX1 I_2835  ( .D(I50842), .CLK(I2702), .RSTB(I50435), .Q(I50924) );
not I_2836 (I50412,I50924);
DFFARX1 I_2837  ( .D(I707142), .CLK(I2702), .RSTB(I50435), .Q(I50955) );
not I_2838 (I50972,I50955);
or I_2839 (I50989,I50972,I50893);
DFFARX1 I_2840  ( .D(I50989), .CLK(I2702), .RSTB(I50435), .Q(I50418) );
nand I_2841 (I50427,I50972,I50698);
DFFARX1 I_2842  ( .D(I50972), .CLK(I2702), .RSTB(I50435), .Q(I50397) );
not I_2843 (I51081,I2709);
not I_2844 (I51098,I418091);
nor I_2845 (I51115,I418073,I418088);
nand I_2846 (I51132,I51115,I418097);
DFFARX1 I_2847  ( .D(I51132), .CLK(I2702), .RSTB(I51081), .Q(I51055) );
nor I_2848 (I51163,I51098,I418073);
nand I_2849 (I51180,I51163,I418100);
not I_2850 (I51070,I51180);
DFFARX1 I_2851  ( .D(I51180), .CLK(I2702), .RSTB(I51081), .Q(I51052) );
not I_2852 (I51225,I418073);
not I_2853 (I51242,I51225);
not I_2854 (I51259,I418103);
nor I_2855 (I51276,I51259,I418079);
and I_2856 (I51293,I51276,I418082);
or I_2857 (I51310,I51293,I418076);
DFFARX1 I_2858  ( .D(I51310), .CLK(I2702), .RSTB(I51081), .Q(I51327) );
nor I_2859 (I51344,I51327,I51180);
nor I_2860 (I51361,I51327,I51242);
nand I_2861 (I51067,I51132,I51361);
nand I_2862 (I51392,I51098,I418103);
nand I_2863 (I51409,I51392,I51327);
and I_2864 (I51426,I51392,I51409);
DFFARX1 I_2865  ( .D(I51426), .CLK(I2702), .RSTB(I51081), .Q(I51049) );
DFFARX1 I_2866  ( .D(I51392), .CLK(I2702), .RSTB(I51081), .Q(I51457) );
and I_2867 (I51046,I51225,I51457);
DFFARX1 I_2868  ( .D(I418085), .CLK(I2702), .RSTB(I51081), .Q(I51488) );
not I_2869 (I51505,I51488);
nor I_2870 (I51522,I51180,I51505);
and I_2871 (I51539,I51488,I51522);
nand I_2872 (I51061,I51488,I51242);
DFFARX1 I_2873  ( .D(I51488), .CLK(I2702), .RSTB(I51081), .Q(I51570) );
not I_2874 (I51058,I51570);
DFFARX1 I_2875  ( .D(I418094), .CLK(I2702), .RSTB(I51081), .Q(I51601) );
not I_2876 (I51618,I51601);
or I_2877 (I51635,I51618,I51539);
DFFARX1 I_2878  ( .D(I51635), .CLK(I2702), .RSTB(I51081), .Q(I51064) );
nand I_2879 (I51073,I51618,I51344);
DFFARX1 I_2880  ( .D(I51618), .CLK(I2702), .RSTB(I51081), .Q(I51043) );
not I_2881 (I51727,I2709);
not I_2882 (I51744,I379025);
nor I_2883 (I51761,I379037,I379019);
nand I_2884 (I51778,I51761,I379034);
DFFARX1 I_2885  ( .D(I51778), .CLK(I2702), .RSTB(I51727), .Q(I51701) );
nor I_2886 (I51809,I51744,I379037);
nand I_2887 (I51826,I51809,I379022);
not I_2888 (I51716,I51826);
DFFARX1 I_2889  ( .D(I51826), .CLK(I2702), .RSTB(I51727), .Q(I51698) );
not I_2890 (I51871,I379037);
not I_2891 (I51888,I51871);
not I_2892 (I51905,I379031);
nor I_2893 (I51922,I51905,I379010);
and I_2894 (I51939,I51922,I379013);
or I_2895 (I51956,I51939,I379016);
DFFARX1 I_2896  ( .D(I51956), .CLK(I2702), .RSTB(I51727), .Q(I51973) );
nor I_2897 (I51990,I51973,I51826);
nor I_2898 (I52007,I51973,I51888);
nand I_2899 (I51713,I51778,I52007);
nand I_2900 (I52038,I51744,I379031);
nand I_2901 (I52055,I52038,I51973);
and I_2902 (I52072,I52038,I52055);
DFFARX1 I_2903  ( .D(I52072), .CLK(I2702), .RSTB(I51727), .Q(I51695) );
DFFARX1 I_2904  ( .D(I52038), .CLK(I2702), .RSTB(I51727), .Q(I52103) );
and I_2905 (I51692,I51871,I52103);
DFFARX1 I_2906  ( .D(I379007), .CLK(I2702), .RSTB(I51727), .Q(I52134) );
not I_2907 (I52151,I52134);
nor I_2908 (I52168,I51826,I52151);
and I_2909 (I52185,I52134,I52168);
nand I_2910 (I51707,I52134,I51888);
DFFARX1 I_2911  ( .D(I52134), .CLK(I2702), .RSTB(I51727), .Q(I52216) );
not I_2912 (I51704,I52216);
DFFARX1 I_2913  ( .D(I379028), .CLK(I2702), .RSTB(I51727), .Q(I52247) );
not I_2914 (I52264,I52247);
or I_2915 (I52281,I52264,I52185);
DFFARX1 I_2916  ( .D(I52281), .CLK(I2702), .RSTB(I51727), .Q(I51710) );
nand I_2917 (I51719,I52264,I51990);
DFFARX1 I_2918  ( .D(I52264), .CLK(I2702), .RSTB(I51727), .Q(I51689) );
not I_2919 (I52373,I2709);
not I_2920 (I52390,I8886);
nor I_2921 (I52407,I8898,I8883);
nand I_2922 (I52424,I52407,I8895);
DFFARX1 I_2923  ( .D(I52424), .CLK(I2702), .RSTB(I52373), .Q(I52347) );
nor I_2924 (I52455,I52390,I8898);
nand I_2925 (I52472,I52455,I8913);
not I_2926 (I52362,I52472);
DFFARX1 I_2927  ( .D(I52472), .CLK(I2702), .RSTB(I52373), .Q(I52344) );
not I_2928 (I52517,I8898);
not I_2929 (I52534,I52517);
not I_2930 (I52551,I8889);
nor I_2931 (I52568,I52551,I8901);
and I_2932 (I52585,I52568,I8892);
or I_2933 (I52602,I52585,I8907);
DFFARX1 I_2934  ( .D(I52602), .CLK(I2702), .RSTB(I52373), .Q(I52619) );
nor I_2935 (I52636,I52619,I52472);
nor I_2936 (I52653,I52619,I52534);
nand I_2937 (I52359,I52424,I52653);
nand I_2938 (I52684,I52390,I8889);
nand I_2939 (I52701,I52684,I52619);
and I_2940 (I52718,I52684,I52701);
DFFARX1 I_2941  ( .D(I52718), .CLK(I2702), .RSTB(I52373), .Q(I52341) );
DFFARX1 I_2942  ( .D(I52684), .CLK(I2702), .RSTB(I52373), .Q(I52749) );
and I_2943 (I52338,I52517,I52749);
DFFARX1 I_2944  ( .D(I8910), .CLK(I2702), .RSTB(I52373), .Q(I52780) );
not I_2945 (I52797,I52780);
nor I_2946 (I52814,I52472,I52797);
and I_2947 (I52831,I52780,I52814);
nand I_2948 (I52353,I52780,I52534);
DFFARX1 I_2949  ( .D(I52780), .CLK(I2702), .RSTB(I52373), .Q(I52862) );
not I_2950 (I52350,I52862);
DFFARX1 I_2951  ( .D(I8904), .CLK(I2702), .RSTB(I52373), .Q(I52893) );
not I_2952 (I52910,I52893);
or I_2953 (I52927,I52910,I52831);
DFFARX1 I_2954  ( .D(I52927), .CLK(I2702), .RSTB(I52373), .Q(I52356) );
nand I_2955 (I52365,I52910,I52636);
DFFARX1 I_2956  ( .D(I52910), .CLK(I2702), .RSTB(I52373), .Q(I52335) );
not I_2957 (I53019,I2709);
not I_2958 (I53036,I361583);
nor I_2959 (I53053,I361595,I361577);
nand I_2960 (I53070,I53053,I361592);
DFFARX1 I_2961  ( .D(I53070), .CLK(I2702), .RSTB(I53019), .Q(I52993) );
nor I_2962 (I53101,I53036,I361595);
nand I_2963 (I53118,I53101,I361580);
not I_2964 (I53008,I53118);
DFFARX1 I_2965  ( .D(I53118), .CLK(I2702), .RSTB(I53019), .Q(I52990) );
not I_2966 (I53163,I361595);
not I_2967 (I53180,I53163);
not I_2968 (I53197,I361589);
nor I_2969 (I53214,I53197,I361568);
and I_2970 (I53231,I53214,I361571);
or I_2971 (I53248,I53231,I361574);
DFFARX1 I_2972  ( .D(I53248), .CLK(I2702), .RSTB(I53019), .Q(I53265) );
nor I_2973 (I53282,I53265,I53118);
nor I_2974 (I53299,I53265,I53180);
nand I_2975 (I53005,I53070,I53299);
nand I_2976 (I53330,I53036,I361589);
nand I_2977 (I53347,I53330,I53265);
and I_2978 (I53364,I53330,I53347);
DFFARX1 I_2979  ( .D(I53364), .CLK(I2702), .RSTB(I53019), .Q(I52987) );
DFFARX1 I_2980  ( .D(I53330), .CLK(I2702), .RSTB(I53019), .Q(I53395) );
and I_2981 (I52984,I53163,I53395);
DFFARX1 I_2982  ( .D(I361565), .CLK(I2702), .RSTB(I53019), .Q(I53426) );
not I_2983 (I53443,I53426);
nor I_2984 (I53460,I53118,I53443);
and I_2985 (I53477,I53426,I53460);
nand I_2986 (I52999,I53426,I53180);
DFFARX1 I_2987  ( .D(I53426), .CLK(I2702), .RSTB(I53019), .Q(I53508) );
not I_2988 (I52996,I53508);
DFFARX1 I_2989  ( .D(I361586), .CLK(I2702), .RSTB(I53019), .Q(I53539) );
not I_2990 (I53556,I53539);
or I_2991 (I53573,I53556,I53477);
DFFARX1 I_2992  ( .D(I53573), .CLK(I2702), .RSTB(I53019), .Q(I53002) );
nand I_2993 (I53011,I53556,I53282);
DFFARX1 I_2994  ( .D(I53556), .CLK(I2702), .RSTB(I53019), .Q(I52981) );
not I_2995 (I53665,I2709);
not I_2996 (I53682,I455828);
nor I_2997 (I53699,I455816,I455822);
nand I_2998 (I53716,I53699,I455813);
DFFARX1 I_2999  ( .D(I53716), .CLK(I2702), .RSTB(I53665), .Q(I53639) );
nor I_3000 (I53747,I53682,I455816);
nand I_3001 (I53764,I53747,I455819);
not I_3002 (I53654,I53764);
DFFARX1 I_3003  ( .D(I53764), .CLK(I2702), .RSTB(I53665), .Q(I53636) );
not I_3004 (I53809,I455816);
not I_3005 (I53826,I53809);
not I_3006 (I53843,I455831);
nor I_3007 (I53860,I53843,I455843);
and I_3008 (I53877,I53860,I455825);
or I_3009 (I53894,I53877,I455840);
DFFARX1 I_3010  ( .D(I53894), .CLK(I2702), .RSTB(I53665), .Q(I53911) );
nor I_3011 (I53928,I53911,I53764);
nor I_3012 (I53945,I53911,I53826);
nand I_3013 (I53651,I53716,I53945);
nand I_3014 (I53976,I53682,I455831);
nand I_3015 (I53993,I53976,I53911);
and I_3016 (I54010,I53976,I53993);
DFFARX1 I_3017  ( .D(I54010), .CLK(I2702), .RSTB(I53665), .Q(I53633) );
DFFARX1 I_3018  ( .D(I53976), .CLK(I2702), .RSTB(I53665), .Q(I54041) );
and I_3019 (I53630,I53809,I54041);
DFFARX1 I_3020  ( .D(I455834), .CLK(I2702), .RSTB(I53665), .Q(I54072) );
not I_3021 (I54089,I54072);
nor I_3022 (I54106,I53764,I54089);
and I_3023 (I54123,I54072,I54106);
nand I_3024 (I53645,I54072,I53826);
DFFARX1 I_3025  ( .D(I54072), .CLK(I2702), .RSTB(I53665), .Q(I54154) );
not I_3026 (I53642,I54154);
DFFARX1 I_3027  ( .D(I455837), .CLK(I2702), .RSTB(I53665), .Q(I54185) );
not I_3028 (I54202,I54185);
or I_3029 (I54219,I54202,I54123);
DFFARX1 I_3030  ( .D(I54219), .CLK(I2702), .RSTB(I53665), .Q(I53648) );
nand I_3031 (I53657,I54202,I53928);
DFFARX1 I_3032  ( .D(I54202), .CLK(I2702), .RSTB(I53665), .Q(I53627) );
not I_3033 (I54311,I2709);
not I_3034 (I54328,I646383);
nor I_3035 (I54345,I646398,I646413);
nand I_3036 (I54362,I54345,I646401);
DFFARX1 I_3037  ( .D(I54362), .CLK(I2702), .RSTB(I54311), .Q(I54285) );
nor I_3038 (I54393,I54328,I646398);
nand I_3039 (I54410,I54393,I646404);
not I_3040 (I54300,I54410);
DFFARX1 I_3041  ( .D(I54410), .CLK(I2702), .RSTB(I54311), .Q(I54282) );
not I_3042 (I54455,I646398);
not I_3043 (I54472,I54455);
not I_3044 (I54489,I646410);
nor I_3045 (I54506,I54489,I646407);
and I_3046 (I54523,I54506,I646386);
or I_3047 (I54540,I54523,I646395);
DFFARX1 I_3048  ( .D(I54540), .CLK(I2702), .RSTB(I54311), .Q(I54557) );
nor I_3049 (I54574,I54557,I54410);
nor I_3050 (I54591,I54557,I54472);
nand I_3051 (I54297,I54362,I54591);
nand I_3052 (I54622,I54328,I646410);
nand I_3053 (I54639,I54622,I54557);
and I_3054 (I54656,I54622,I54639);
DFFARX1 I_3055  ( .D(I54656), .CLK(I2702), .RSTB(I54311), .Q(I54279) );
DFFARX1 I_3056  ( .D(I54622), .CLK(I2702), .RSTB(I54311), .Q(I54687) );
and I_3057 (I54276,I54455,I54687);
DFFARX1 I_3058  ( .D(I646392), .CLK(I2702), .RSTB(I54311), .Q(I54718) );
not I_3059 (I54735,I54718);
nor I_3060 (I54752,I54410,I54735);
and I_3061 (I54769,I54718,I54752);
nand I_3062 (I54291,I54718,I54472);
DFFARX1 I_3063  ( .D(I54718), .CLK(I2702), .RSTB(I54311), .Q(I54800) );
not I_3064 (I54288,I54800);
DFFARX1 I_3065  ( .D(I646389), .CLK(I2702), .RSTB(I54311), .Q(I54831) );
not I_3066 (I54848,I54831);
or I_3067 (I54865,I54848,I54769);
DFFARX1 I_3068  ( .D(I54865), .CLK(I2702), .RSTB(I54311), .Q(I54294) );
nand I_3069 (I54303,I54848,I54574);
DFFARX1 I_3070  ( .D(I54848), .CLK(I2702), .RSTB(I54311), .Q(I54273) );
not I_3071 (I54957,I2709);
not I_3072 (I54974,I238559);
nor I_3073 (I54991,I238580,I238553);
nand I_3074 (I55008,I54991,I238568);
DFFARX1 I_3075  ( .D(I55008), .CLK(I2702), .RSTB(I54957), .Q(I54931) );
nor I_3076 (I55039,I54974,I238580);
nand I_3077 (I55056,I55039,I238583);
not I_3078 (I54946,I55056);
DFFARX1 I_3079  ( .D(I55056), .CLK(I2702), .RSTB(I54957), .Q(I54928) );
not I_3080 (I55101,I238580);
not I_3081 (I55118,I55101);
not I_3082 (I55135,I238556);
nor I_3083 (I55152,I55135,I238574);
and I_3084 (I55169,I55152,I238562);
or I_3085 (I55186,I55169,I238565);
DFFARX1 I_3086  ( .D(I55186), .CLK(I2702), .RSTB(I54957), .Q(I55203) );
nor I_3087 (I55220,I55203,I55056);
nor I_3088 (I55237,I55203,I55118);
nand I_3089 (I54943,I55008,I55237);
nand I_3090 (I55268,I54974,I238556);
nand I_3091 (I55285,I55268,I55203);
and I_3092 (I55302,I55268,I55285);
DFFARX1 I_3093  ( .D(I55302), .CLK(I2702), .RSTB(I54957), .Q(I54925) );
DFFARX1 I_3094  ( .D(I55268), .CLK(I2702), .RSTB(I54957), .Q(I55333) );
and I_3095 (I54922,I55101,I55333);
DFFARX1 I_3096  ( .D(I238577), .CLK(I2702), .RSTB(I54957), .Q(I55364) );
not I_3097 (I55381,I55364);
nor I_3098 (I55398,I55056,I55381);
and I_3099 (I55415,I55364,I55398);
nand I_3100 (I54937,I55364,I55118);
DFFARX1 I_3101  ( .D(I55364), .CLK(I2702), .RSTB(I54957), .Q(I55446) );
not I_3102 (I54934,I55446);
DFFARX1 I_3103  ( .D(I238571), .CLK(I2702), .RSTB(I54957), .Q(I55477) );
not I_3104 (I55494,I55477);
or I_3105 (I55511,I55494,I55415);
DFFARX1 I_3106  ( .D(I55511), .CLK(I2702), .RSTB(I54957), .Q(I54940) );
nand I_3107 (I54949,I55494,I55220);
DFFARX1 I_3108  ( .D(I55494), .CLK(I2702), .RSTB(I54957), .Q(I54919) );
not I_3109 (I55603,I2709);
not I_3110 (I55620,I675317);
nor I_3111 (I55637,I675332,I675347);
nand I_3112 (I55654,I55637,I675335);
DFFARX1 I_3113  ( .D(I55654), .CLK(I2702), .RSTB(I55603), .Q(I55577) );
nor I_3114 (I55685,I55620,I675332);
nand I_3115 (I55702,I55685,I675338);
not I_3116 (I55592,I55702);
DFFARX1 I_3117  ( .D(I55702), .CLK(I2702), .RSTB(I55603), .Q(I55574) );
not I_3118 (I55747,I675332);
not I_3119 (I55764,I55747);
not I_3120 (I55781,I675344);
nor I_3121 (I55798,I55781,I675341);
and I_3122 (I55815,I55798,I675320);
or I_3123 (I55832,I55815,I675329);
DFFARX1 I_3124  ( .D(I55832), .CLK(I2702), .RSTB(I55603), .Q(I55849) );
nor I_3125 (I55866,I55849,I55702);
nor I_3126 (I55883,I55849,I55764);
nand I_3127 (I55589,I55654,I55883);
nand I_3128 (I55914,I55620,I675344);
nand I_3129 (I55931,I55914,I55849);
and I_3130 (I55948,I55914,I55931);
DFFARX1 I_3131  ( .D(I55948), .CLK(I2702), .RSTB(I55603), .Q(I55571) );
DFFARX1 I_3132  ( .D(I55914), .CLK(I2702), .RSTB(I55603), .Q(I55979) );
and I_3133 (I55568,I55747,I55979);
DFFARX1 I_3134  ( .D(I675326), .CLK(I2702), .RSTB(I55603), .Q(I56010) );
not I_3135 (I56027,I56010);
nor I_3136 (I56044,I55702,I56027);
and I_3137 (I56061,I56010,I56044);
nand I_3138 (I55583,I56010,I55764);
DFFARX1 I_3139  ( .D(I56010), .CLK(I2702), .RSTB(I55603), .Q(I56092) );
not I_3140 (I55580,I56092);
DFFARX1 I_3141  ( .D(I675323), .CLK(I2702), .RSTB(I55603), .Q(I56123) );
not I_3142 (I56140,I56123);
or I_3143 (I56157,I56140,I56061);
DFFARX1 I_3144  ( .D(I56157), .CLK(I2702), .RSTB(I55603), .Q(I55586) );
nand I_3145 (I55595,I56140,I55866);
DFFARX1 I_3146  ( .D(I56140), .CLK(I2702), .RSTB(I55603), .Q(I55565) );
not I_3147 (I56249,I2709);
not I_3148 (I56266,I556021);
nor I_3149 (I56283,I555997,I556003);
nand I_3150 (I56300,I56283,I556006);
DFFARX1 I_3151  ( .D(I56300), .CLK(I2702), .RSTB(I56249), .Q(I56223) );
nor I_3152 (I56331,I56266,I555997);
nand I_3153 (I56348,I56331,I556015);
not I_3154 (I56238,I56348);
DFFARX1 I_3155  ( .D(I56348), .CLK(I2702), .RSTB(I56249), .Q(I56220) );
not I_3156 (I56393,I555997);
not I_3157 (I56410,I56393);
not I_3158 (I56427,I555994);
nor I_3159 (I56444,I56427,I556009);
and I_3160 (I56461,I56444,I556000);
or I_3161 (I56478,I56461,I556012);
DFFARX1 I_3162  ( .D(I56478), .CLK(I2702), .RSTB(I56249), .Q(I56495) );
nor I_3163 (I56512,I56495,I56348);
nor I_3164 (I56529,I56495,I56410);
nand I_3165 (I56235,I56300,I56529);
nand I_3166 (I56560,I56266,I555994);
nand I_3167 (I56577,I56560,I56495);
and I_3168 (I56594,I56560,I56577);
DFFARX1 I_3169  ( .D(I56594), .CLK(I2702), .RSTB(I56249), .Q(I56217) );
DFFARX1 I_3170  ( .D(I56560), .CLK(I2702), .RSTB(I56249), .Q(I56625) );
and I_3171 (I56214,I56393,I56625);
DFFARX1 I_3172  ( .D(I556024), .CLK(I2702), .RSTB(I56249), .Q(I56656) );
not I_3173 (I56673,I56656);
nor I_3174 (I56690,I56348,I56673);
and I_3175 (I56707,I56656,I56690);
nand I_3176 (I56229,I56656,I56410);
DFFARX1 I_3177  ( .D(I56656), .CLK(I2702), .RSTB(I56249), .Q(I56738) );
not I_3178 (I56226,I56738);
DFFARX1 I_3179  ( .D(I556018), .CLK(I2702), .RSTB(I56249), .Q(I56769) );
not I_3180 (I56786,I56769);
or I_3181 (I56803,I56786,I56707);
DFFARX1 I_3182  ( .D(I56803), .CLK(I2702), .RSTB(I56249), .Q(I56232) );
nand I_3183 (I56241,I56786,I56512);
DFFARX1 I_3184  ( .D(I56786), .CLK(I2702), .RSTB(I56249), .Q(I56211) );
not I_3185 (I56895,I2709);
not I_3186 (I56912,I570896);
nor I_3187 (I56929,I570872,I570878);
nand I_3188 (I56946,I56929,I570881);
DFFARX1 I_3189  ( .D(I56946), .CLK(I2702), .RSTB(I56895), .Q(I56869) );
nor I_3190 (I56977,I56912,I570872);
nand I_3191 (I56994,I56977,I570890);
not I_3192 (I56884,I56994);
DFFARX1 I_3193  ( .D(I56994), .CLK(I2702), .RSTB(I56895), .Q(I56866) );
not I_3194 (I57039,I570872);
not I_3195 (I57056,I57039);
not I_3196 (I57073,I570869);
nor I_3197 (I57090,I57073,I570884);
and I_3198 (I57107,I57090,I570875);
or I_3199 (I57124,I57107,I570887);
DFFARX1 I_3200  ( .D(I57124), .CLK(I2702), .RSTB(I56895), .Q(I57141) );
nor I_3201 (I57158,I57141,I56994);
nor I_3202 (I57175,I57141,I57056);
nand I_3203 (I56881,I56946,I57175);
nand I_3204 (I57206,I56912,I570869);
nand I_3205 (I57223,I57206,I57141);
and I_3206 (I57240,I57206,I57223);
DFFARX1 I_3207  ( .D(I57240), .CLK(I2702), .RSTB(I56895), .Q(I56863) );
DFFARX1 I_3208  ( .D(I57206), .CLK(I2702), .RSTB(I56895), .Q(I57271) );
and I_3209 (I56860,I57039,I57271);
DFFARX1 I_3210  ( .D(I570899), .CLK(I2702), .RSTB(I56895), .Q(I57302) );
not I_3211 (I57319,I57302);
nor I_3212 (I57336,I56994,I57319);
and I_3213 (I57353,I57302,I57336);
nand I_3214 (I56875,I57302,I57056);
DFFARX1 I_3215  ( .D(I57302), .CLK(I2702), .RSTB(I56895), .Q(I57384) );
not I_3216 (I56872,I57384);
DFFARX1 I_3217  ( .D(I570893), .CLK(I2702), .RSTB(I56895), .Q(I57415) );
not I_3218 (I57432,I57415);
or I_3219 (I57449,I57432,I57353);
DFFARX1 I_3220  ( .D(I57449), .CLK(I2702), .RSTB(I56895), .Q(I56878) );
nand I_3221 (I56887,I57432,I57158);
DFFARX1 I_3222  ( .D(I57432), .CLK(I2702), .RSTB(I56895), .Q(I56857) );
not I_3223 (I57541,I2709);
not I_3224 (I57558,I505446);
nor I_3225 (I57575,I505422,I505428);
nand I_3226 (I57592,I57575,I505431);
DFFARX1 I_3227  ( .D(I57592), .CLK(I2702), .RSTB(I57541), .Q(I57515) );
nor I_3228 (I57623,I57558,I505422);
nand I_3229 (I57640,I57623,I505440);
not I_3230 (I57530,I57640);
DFFARX1 I_3231  ( .D(I57640), .CLK(I2702), .RSTB(I57541), .Q(I57512) );
not I_3232 (I57685,I505422);
not I_3233 (I57702,I57685);
not I_3234 (I57719,I505419);
nor I_3235 (I57736,I57719,I505434);
and I_3236 (I57753,I57736,I505425);
or I_3237 (I57770,I57753,I505437);
DFFARX1 I_3238  ( .D(I57770), .CLK(I2702), .RSTB(I57541), .Q(I57787) );
nor I_3239 (I57804,I57787,I57640);
nor I_3240 (I57821,I57787,I57702);
nand I_3241 (I57527,I57592,I57821);
nand I_3242 (I57852,I57558,I505419);
nand I_3243 (I57869,I57852,I57787);
and I_3244 (I57886,I57852,I57869);
DFFARX1 I_3245  ( .D(I57886), .CLK(I2702), .RSTB(I57541), .Q(I57509) );
DFFARX1 I_3246  ( .D(I57852), .CLK(I2702), .RSTB(I57541), .Q(I57917) );
and I_3247 (I57506,I57685,I57917);
DFFARX1 I_3248  ( .D(I505449), .CLK(I2702), .RSTB(I57541), .Q(I57948) );
not I_3249 (I57965,I57948);
nor I_3250 (I57982,I57640,I57965);
and I_3251 (I57999,I57948,I57982);
nand I_3252 (I57521,I57948,I57702);
DFFARX1 I_3253  ( .D(I57948), .CLK(I2702), .RSTB(I57541), .Q(I58030) );
not I_3254 (I57518,I58030);
DFFARX1 I_3255  ( .D(I505443), .CLK(I2702), .RSTB(I57541), .Q(I58061) );
not I_3256 (I58078,I58061);
or I_3257 (I58095,I58078,I57999);
DFFARX1 I_3258  ( .D(I58095), .CLK(I2702), .RSTB(I57541), .Q(I57524) );
nand I_3259 (I57533,I58078,I57804);
DFFARX1 I_3260  ( .D(I58078), .CLK(I2702), .RSTB(I57541), .Q(I57503) );
not I_3261 (I58187,I2709);
not I_3262 (I58204,I424211);
nor I_3263 (I58221,I424193,I424208);
nand I_3264 (I58238,I58221,I424217);
DFFARX1 I_3265  ( .D(I58238), .CLK(I2702), .RSTB(I58187), .Q(I58161) );
nor I_3266 (I58269,I58204,I424193);
nand I_3267 (I58286,I58269,I424220);
not I_3268 (I58176,I58286);
DFFARX1 I_3269  ( .D(I58286), .CLK(I2702), .RSTB(I58187), .Q(I58158) );
not I_3270 (I58331,I424193);
not I_3271 (I58348,I58331);
not I_3272 (I58365,I424223);
nor I_3273 (I58382,I58365,I424199);
and I_3274 (I58399,I58382,I424202);
or I_3275 (I58416,I58399,I424196);
DFFARX1 I_3276  ( .D(I58416), .CLK(I2702), .RSTB(I58187), .Q(I58433) );
nor I_3277 (I58450,I58433,I58286);
nor I_3278 (I58467,I58433,I58348);
nand I_3279 (I58173,I58238,I58467);
nand I_3280 (I58498,I58204,I424223);
nand I_3281 (I58515,I58498,I58433);
and I_3282 (I58532,I58498,I58515);
DFFARX1 I_3283  ( .D(I58532), .CLK(I2702), .RSTB(I58187), .Q(I58155) );
DFFARX1 I_3284  ( .D(I58498), .CLK(I2702), .RSTB(I58187), .Q(I58563) );
and I_3285 (I58152,I58331,I58563);
DFFARX1 I_3286  ( .D(I424205), .CLK(I2702), .RSTB(I58187), .Q(I58594) );
not I_3287 (I58611,I58594);
nor I_3288 (I58628,I58286,I58611);
and I_3289 (I58645,I58594,I58628);
nand I_3290 (I58167,I58594,I58348);
DFFARX1 I_3291  ( .D(I58594), .CLK(I2702), .RSTB(I58187), .Q(I58676) );
not I_3292 (I58164,I58676);
DFFARX1 I_3293  ( .D(I424214), .CLK(I2702), .RSTB(I58187), .Q(I58707) );
not I_3294 (I58724,I58707);
or I_3295 (I58741,I58724,I58645);
DFFARX1 I_3296  ( .D(I58741), .CLK(I2702), .RSTB(I58187), .Q(I58170) );
nand I_3297 (I58179,I58724,I58450);
DFFARX1 I_3298  ( .D(I58724), .CLK(I2702), .RSTB(I58187), .Q(I58149) );
not I_3299 (I58833,I2709);
not I_3300 (I58850,I504859);
nor I_3301 (I58867,I504871,I504853);
nand I_3302 (I58884,I58867,I504862);
DFFARX1 I_3303  ( .D(I58884), .CLK(I2702), .RSTB(I58833), .Q(I58807) );
nor I_3304 (I58915,I58850,I504871);
nand I_3305 (I58932,I58915,I504868);
not I_3306 (I58822,I58932);
DFFARX1 I_3307  ( .D(I58932), .CLK(I2702), .RSTB(I58833), .Q(I58804) );
not I_3308 (I58977,I504871);
not I_3309 (I58994,I58977);
not I_3310 (I59011,I504841);
nor I_3311 (I59028,I59011,I504844);
and I_3312 (I59045,I59028,I504850);
or I_3313 (I59062,I59045,I504865);
DFFARX1 I_3314  ( .D(I59062), .CLK(I2702), .RSTB(I58833), .Q(I59079) );
nor I_3315 (I59096,I59079,I58932);
nor I_3316 (I59113,I59079,I58994);
nand I_3317 (I58819,I58884,I59113);
nand I_3318 (I59144,I58850,I504841);
nand I_3319 (I59161,I59144,I59079);
and I_3320 (I59178,I59144,I59161);
DFFARX1 I_3321  ( .D(I59178), .CLK(I2702), .RSTB(I58833), .Q(I58801) );
DFFARX1 I_3322  ( .D(I59144), .CLK(I2702), .RSTB(I58833), .Q(I59209) );
and I_3323 (I58798,I58977,I59209);
DFFARX1 I_3324  ( .D(I504847), .CLK(I2702), .RSTB(I58833), .Q(I59240) );
not I_3325 (I59257,I59240);
nor I_3326 (I59274,I58932,I59257);
and I_3327 (I59291,I59240,I59274);
nand I_3328 (I58813,I59240,I58994);
DFFARX1 I_3329  ( .D(I59240), .CLK(I2702), .RSTB(I58833), .Q(I59322) );
not I_3330 (I58810,I59322);
DFFARX1 I_3331  ( .D(I504856), .CLK(I2702), .RSTB(I58833), .Q(I59353) );
not I_3332 (I59370,I59353);
or I_3333 (I59387,I59370,I59291);
DFFARX1 I_3334  ( .D(I59387), .CLK(I2702), .RSTB(I58833), .Q(I58816) );
nand I_3335 (I58825,I59370,I59096);
DFFARX1 I_3336  ( .D(I59370), .CLK(I2702), .RSTB(I58833), .Q(I58795) );
not I_3337 (I59479,I2709);
not I_3338 (I59496,I244509);
nor I_3339 (I59513,I244530,I244503);
nand I_3340 (I59530,I59513,I244518);
DFFARX1 I_3341  ( .D(I59530), .CLK(I2702), .RSTB(I59479), .Q(I59453) );
nor I_3342 (I59561,I59496,I244530);
nand I_3343 (I59578,I59561,I244533);
not I_3344 (I59468,I59578);
DFFARX1 I_3345  ( .D(I59578), .CLK(I2702), .RSTB(I59479), .Q(I59450) );
not I_3346 (I59623,I244530);
not I_3347 (I59640,I59623);
not I_3348 (I59657,I244506);
nor I_3349 (I59674,I59657,I244524);
and I_3350 (I59691,I59674,I244512);
or I_3351 (I59708,I59691,I244515);
DFFARX1 I_3352  ( .D(I59708), .CLK(I2702), .RSTB(I59479), .Q(I59725) );
nor I_3353 (I59742,I59725,I59578);
nor I_3354 (I59759,I59725,I59640);
nand I_3355 (I59465,I59530,I59759);
nand I_3356 (I59790,I59496,I244506);
nand I_3357 (I59807,I59790,I59725);
and I_3358 (I59824,I59790,I59807);
DFFARX1 I_3359  ( .D(I59824), .CLK(I2702), .RSTB(I59479), .Q(I59447) );
DFFARX1 I_3360  ( .D(I59790), .CLK(I2702), .RSTB(I59479), .Q(I59855) );
and I_3361 (I59444,I59623,I59855);
DFFARX1 I_3362  ( .D(I244527), .CLK(I2702), .RSTB(I59479), .Q(I59886) );
not I_3363 (I59903,I59886);
nor I_3364 (I59920,I59578,I59903);
and I_3365 (I59937,I59886,I59920);
nand I_3366 (I59459,I59886,I59640);
DFFARX1 I_3367  ( .D(I59886), .CLK(I2702), .RSTB(I59479), .Q(I59968) );
not I_3368 (I59456,I59968);
DFFARX1 I_3369  ( .D(I244521), .CLK(I2702), .RSTB(I59479), .Q(I59999) );
not I_3370 (I60016,I59999);
or I_3371 (I60033,I60016,I59937);
DFFARX1 I_3372  ( .D(I60033), .CLK(I2702), .RSTB(I59479), .Q(I59462) );
nand I_3373 (I59471,I60016,I59742);
DFFARX1 I_3374  ( .D(I60016), .CLK(I2702), .RSTB(I59479), .Q(I59441) );
not I_3375 (I60125,I2709);
not I_3376 (I60142,I14496);
nor I_3377 (I60159,I14508,I14493);
nand I_3378 (I60176,I60159,I14505);
DFFARX1 I_3379  ( .D(I60176), .CLK(I2702), .RSTB(I60125), .Q(I60099) );
nor I_3380 (I60207,I60142,I14508);
nand I_3381 (I60224,I60207,I14523);
not I_3382 (I60114,I60224);
DFFARX1 I_3383  ( .D(I60224), .CLK(I2702), .RSTB(I60125), .Q(I60096) );
not I_3384 (I60269,I14508);
not I_3385 (I60286,I60269);
not I_3386 (I60303,I14499);
nor I_3387 (I60320,I60303,I14511);
and I_3388 (I60337,I60320,I14502);
or I_3389 (I60354,I60337,I14517);
DFFARX1 I_3390  ( .D(I60354), .CLK(I2702), .RSTB(I60125), .Q(I60371) );
nor I_3391 (I60388,I60371,I60224);
nor I_3392 (I60405,I60371,I60286);
nand I_3393 (I60111,I60176,I60405);
nand I_3394 (I60436,I60142,I14499);
nand I_3395 (I60453,I60436,I60371);
and I_3396 (I60470,I60436,I60453);
DFFARX1 I_3397  ( .D(I60470), .CLK(I2702), .RSTB(I60125), .Q(I60093) );
DFFARX1 I_3398  ( .D(I60436), .CLK(I2702), .RSTB(I60125), .Q(I60501) );
and I_3399 (I60090,I60269,I60501);
DFFARX1 I_3400  ( .D(I14520), .CLK(I2702), .RSTB(I60125), .Q(I60532) );
not I_3401 (I60549,I60532);
nor I_3402 (I60566,I60224,I60549);
and I_3403 (I60583,I60532,I60566);
nand I_3404 (I60105,I60532,I60286);
DFFARX1 I_3405  ( .D(I60532), .CLK(I2702), .RSTB(I60125), .Q(I60614) );
not I_3406 (I60102,I60614);
DFFARX1 I_3407  ( .D(I14514), .CLK(I2702), .RSTB(I60125), .Q(I60645) );
not I_3408 (I60662,I60645);
or I_3409 (I60679,I60662,I60583);
DFFARX1 I_3410  ( .D(I60679), .CLK(I2702), .RSTB(I60125), .Q(I60108) );
nand I_3411 (I60117,I60662,I60388);
DFFARX1 I_3412  ( .D(I60662), .CLK(I2702), .RSTB(I60125), .Q(I60087) );
not I_3413 (I60771,I2709);
not I_3414 (I60788,I340265);
nor I_3415 (I60805,I340277,I340259);
nand I_3416 (I60822,I60805,I340274);
DFFARX1 I_3417  ( .D(I60822), .CLK(I2702), .RSTB(I60771), .Q(I60745) );
nor I_3418 (I60853,I60788,I340277);
nand I_3419 (I60870,I60853,I340262);
not I_3420 (I60760,I60870);
DFFARX1 I_3421  ( .D(I60870), .CLK(I2702), .RSTB(I60771), .Q(I60742) );
not I_3422 (I60915,I340277);
not I_3423 (I60932,I60915);
not I_3424 (I60949,I340271);
nor I_3425 (I60966,I60949,I340250);
and I_3426 (I60983,I60966,I340253);
or I_3427 (I61000,I60983,I340256);
DFFARX1 I_3428  ( .D(I61000), .CLK(I2702), .RSTB(I60771), .Q(I61017) );
nor I_3429 (I61034,I61017,I60870);
nor I_3430 (I61051,I61017,I60932);
nand I_3431 (I60757,I60822,I61051);
nand I_3432 (I61082,I60788,I340271);
nand I_3433 (I61099,I61082,I61017);
and I_3434 (I61116,I61082,I61099);
DFFARX1 I_3435  ( .D(I61116), .CLK(I2702), .RSTB(I60771), .Q(I60739) );
DFFARX1 I_3436  ( .D(I61082), .CLK(I2702), .RSTB(I60771), .Q(I61147) );
and I_3437 (I60736,I60915,I61147);
DFFARX1 I_3438  ( .D(I340247), .CLK(I2702), .RSTB(I60771), .Q(I61178) );
not I_3439 (I61195,I61178);
nor I_3440 (I61212,I60870,I61195);
and I_3441 (I61229,I61178,I61212);
nand I_3442 (I60751,I61178,I60932);
DFFARX1 I_3443  ( .D(I61178), .CLK(I2702), .RSTB(I60771), .Q(I61260) );
not I_3444 (I60748,I61260);
DFFARX1 I_3445  ( .D(I340268), .CLK(I2702), .RSTB(I60771), .Q(I61291) );
not I_3446 (I61308,I61291);
or I_3447 (I61325,I61308,I61229);
DFFARX1 I_3448  ( .D(I61325), .CLK(I2702), .RSTB(I60771), .Q(I60754) );
nand I_3449 (I60763,I61308,I61034);
DFFARX1 I_3450  ( .D(I61308), .CLK(I2702), .RSTB(I60771), .Q(I60733) );
not I_3451 (I61417,I2709);
not I_3452 (I61434,I204638);
nor I_3453 (I61451,I204668,I204647);
nand I_3454 (I61468,I61451,I204659);
DFFARX1 I_3455  ( .D(I61468), .CLK(I2702), .RSTB(I61417), .Q(I61391) );
nor I_3456 (I61499,I61434,I204668);
nand I_3457 (I61516,I61499,I204641);
not I_3458 (I61406,I61516);
DFFARX1 I_3459  ( .D(I61516), .CLK(I2702), .RSTB(I61417), .Q(I61388) );
not I_3460 (I61561,I204668);
not I_3461 (I61578,I61561);
not I_3462 (I61595,I204644);
nor I_3463 (I61612,I61595,I204662);
and I_3464 (I61629,I61612,I204653);
or I_3465 (I61646,I61629,I204650);
DFFARX1 I_3466  ( .D(I61646), .CLK(I2702), .RSTB(I61417), .Q(I61663) );
nor I_3467 (I61680,I61663,I61516);
nor I_3468 (I61697,I61663,I61578);
nand I_3469 (I61403,I61468,I61697);
nand I_3470 (I61728,I61434,I204644);
nand I_3471 (I61745,I61728,I61663);
and I_3472 (I61762,I61728,I61745);
DFFARX1 I_3473  ( .D(I61762), .CLK(I2702), .RSTB(I61417), .Q(I61385) );
DFFARX1 I_3474  ( .D(I61728), .CLK(I2702), .RSTB(I61417), .Q(I61793) );
and I_3475 (I61382,I61561,I61793);
DFFARX1 I_3476  ( .D(I204656), .CLK(I2702), .RSTB(I61417), .Q(I61824) );
not I_3477 (I61841,I61824);
nor I_3478 (I61858,I61516,I61841);
and I_3479 (I61875,I61824,I61858);
nand I_3480 (I61397,I61824,I61578);
DFFARX1 I_3481  ( .D(I61824), .CLK(I2702), .RSTB(I61417), .Q(I61906) );
not I_3482 (I61394,I61906);
DFFARX1 I_3483  ( .D(I204665), .CLK(I2702), .RSTB(I61417), .Q(I61937) );
not I_3484 (I61954,I61937);
or I_3485 (I61971,I61954,I61875);
DFFARX1 I_3486  ( .D(I61971), .CLK(I2702), .RSTB(I61417), .Q(I61400) );
nand I_3487 (I61409,I61954,I61680);
DFFARX1 I_3488  ( .D(I61954), .CLK(I2702), .RSTB(I61417), .Q(I61379) );
not I_3489 (I62063,I2709);
not I_3490 (I62080,I709445);
nor I_3491 (I62097,I709442,I709439);
nand I_3492 (I62114,I62097,I709460);
DFFARX1 I_3493  ( .D(I62114), .CLK(I2702), .RSTB(I62063), .Q(I62037) );
nor I_3494 (I62145,I62080,I709442);
nand I_3495 (I62162,I62145,I709463);
not I_3496 (I62052,I62162);
DFFARX1 I_3497  ( .D(I62162), .CLK(I2702), .RSTB(I62063), .Q(I62034) );
not I_3498 (I62207,I709442);
not I_3499 (I62224,I62207);
not I_3500 (I62241,I709436);
nor I_3501 (I62258,I62241,I709448);
and I_3502 (I62275,I62258,I709457);
or I_3503 (I62292,I62275,I709451);
DFFARX1 I_3504  ( .D(I62292), .CLK(I2702), .RSTB(I62063), .Q(I62309) );
nor I_3505 (I62326,I62309,I62162);
nor I_3506 (I62343,I62309,I62224);
nand I_3507 (I62049,I62114,I62343);
nand I_3508 (I62374,I62080,I709436);
nand I_3509 (I62391,I62374,I62309);
and I_3510 (I62408,I62374,I62391);
DFFARX1 I_3511  ( .D(I62408), .CLK(I2702), .RSTB(I62063), .Q(I62031) );
DFFARX1 I_3512  ( .D(I62374), .CLK(I2702), .RSTB(I62063), .Q(I62439) );
and I_3513 (I62028,I62207,I62439);
DFFARX1 I_3514  ( .D(I709466), .CLK(I2702), .RSTB(I62063), .Q(I62470) );
not I_3515 (I62487,I62470);
nor I_3516 (I62504,I62162,I62487);
and I_3517 (I62521,I62470,I62504);
nand I_3518 (I62043,I62470,I62224);
DFFARX1 I_3519  ( .D(I62470), .CLK(I2702), .RSTB(I62063), .Q(I62552) );
not I_3520 (I62040,I62552);
DFFARX1 I_3521  ( .D(I709454), .CLK(I2702), .RSTB(I62063), .Q(I62583) );
not I_3522 (I62600,I62583);
or I_3523 (I62617,I62600,I62521);
DFFARX1 I_3524  ( .D(I62617), .CLK(I2702), .RSTB(I62063), .Q(I62046) );
nand I_3525 (I62055,I62600,I62326);
DFFARX1 I_3526  ( .D(I62600), .CLK(I2702), .RSTB(I62063), .Q(I62025) );
not I_3527 (I62709,I2709);
not I_3528 (I62726,I444268);
nor I_3529 (I62743,I444256,I444262);
nand I_3530 (I62760,I62743,I444253);
DFFARX1 I_3531  ( .D(I62760), .CLK(I2702), .RSTB(I62709), .Q(I62683) );
nor I_3532 (I62791,I62726,I444256);
nand I_3533 (I62808,I62791,I444259);
not I_3534 (I62698,I62808);
DFFARX1 I_3535  ( .D(I62808), .CLK(I2702), .RSTB(I62709), .Q(I62680) );
not I_3536 (I62853,I444256);
not I_3537 (I62870,I62853);
not I_3538 (I62887,I444271);
nor I_3539 (I62904,I62887,I444283);
and I_3540 (I62921,I62904,I444265);
or I_3541 (I62938,I62921,I444280);
DFFARX1 I_3542  ( .D(I62938), .CLK(I2702), .RSTB(I62709), .Q(I62955) );
nor I_3543 (I62972,I62955,I62808);
nor I_3544 (I62989,I62955,I62870);
nand I_3545 (I62695,I62760,I62989);
nand I_3546 (I63020,I62726,I444271);
nand I_3547 (I63037,I63020,I62955);
and I_3548 (I63054,I63020,I63037);
DFFARX1 I_3549  ( .D(I63054), .CLK(I2702), .RSTB(I62709), .Q(I62677) );
DFFARX1 I_3550  ( .D(I63020), .CLK(I2702), .RSTB(I62709), .Q(I63085) );
and I_3551 (I62674,I62853,I63085);
DFFARX1 I_3552  ( .D(I444274), .CLK(I2702), .RSTB(I62709), .Q(I63116) );
not I_3553 (I63133,I63116);
nor I_3554 (I63150,I62808,I63133);
and I_3555 (I63167,I63116,I63150);
nand I_3556 (I62689,I63116,I62870);
DFFARX1 I_3557  ( .D(I63116), .CLK(I2702), .RSTB(I62709), .Q(I63198) );
not I_3558 (I62686,I63198);
DFFARX1 I_3559  ( .D(I444277), .CLK(I2702), .RSTB(I62709), .Q(I63229) );
not I_3560 (I63246,I63229);
or I_3561 (I63263,I63246,I63167);
DFFARX1 I_3562  ( .D(I63263), .CLK(I2702), .RSTB(I62709), .Q(I62692) );
nand I_3563 (I62701,I63246,I62972);
DFFARX1 I_3564  ( .D(I63246), .CLK(I2702), .RSTB(I62709), .Q(I62671) );
not I_3565 (I63355,I2709);
not I_3566 (I63372,I668398);
nor I_3567 (I63389,I668413,I668428);
nand I_3568 (I63406,I63389,I668416);
DFFARX1 I_3569  ( .D(I63406), .CLK(I2702), .RSTB(I63355), .Q(I63329) );
nor I_3570 (I63437,I63372,I668413);
nand I_3571 (I63454,I63437,I668419);
not I_3572 (I63344,I63454);
DFFARX1 I_3573  ( .D(I63454), .CLK(I2702), .RSTB(I63355), .Q(I63326) );
not I_3574 (I63499,I668413);
not I_3575 (I63516,I63499);
not I_3576 (I63533,I668425);
nor I_3577 (I63550,I63533,I668422);
and I_3578 (I63567,I63550,I668401);
or I_3579 (I63584,I63567,I668410);
DFFARX1 I_3580  ( .D(I63584), .CLK(I2702), .RSTB(I63355), .Q(I63601) );
nor I_3581 (I63618,I63601,I63454);
nor I_3582 (I63635,I63601,I63516);
nand I_3583 (I63341,I63406,I63635);
nand I_3584 (I63666,I63372,I668425);
nand I_3585 (I63683,I63666,I63601);
and I_3586 (I63700,I63666,I63683);
DFFARX1 I_3587  ( .D(I63700), .CLK(I2702), .RSTB(I63355), .Q(I63323) );
DFFARX1 I_3588  ( .D(I63666), .CLK(I2702), .RSTB(I63355), .Q(I63731) );
and I_3589 (I63320,I63499,I63731);
DFFARX1 I_3590  ( .D(I668407), .CLK(I2702), .RSTB(I63355), .Q(I63762) );
not I_3591 (I63779,I63762);
nor I_3592 (I63796,I63454,I63779);
and I_3593 (I63813,I63762,I63796);
nand I_3594 (I63335,I63762,I63516);
DFFARX1 I_3595  ( .D(I63762), .CLK(I2702), .RSTB(I63355), .Q(I63844) );
not I_3596 (I63332,I63844);
DFFARX1 I_3597  ( .D(I668404), .CLK(I2702), .RSTB(I63355), .Q(I63875) );
not I_3598 (I63892,I63875);
or I_3599 (I63909,I63892,I63813);
DFFARX1 I_3600  ( .D(I63909), .CLK(I2702), .RSTB(I63355), .Q(I63338) );
nand I_3601 (I63347,I63892,I63618);
DFFARX1 I_3602  ( .D(I63892), .CLK(I2702), .RSTB(I63355), .Q(I63317) );
not I_3603 (I64001,I2709);
not I_3604 (I64018,I357707);
nor I_3605 (I64035,I357719,I357701);
nand I_3606 (I64052,I64035,I357716);
DFFARX1 I_3607  ( .D(I64052), .CLK(I2702), .RSTB(I64001), .Q(I63975) );
nor I_3608 (I64083,I64018,I357719);
nand I_3609 (I64100,I64083,I357704);
not I_3610 (I63990,I64100);
DFFARX1 I_3611  ( .D(I64100), .CLK(I2702), .RSTB(I64001), .Q(I63972) );
not I_3612 (I64145,I357719);
not I_3613 (I64162,I64145);
not I_3614 (I64179,I357713);
nor I_3615 (I64196,I64179,I357692);
and I_3616 (I64213,I64196,I357695);
or I_3617 (I64230,I64213,I357698);
DFFARX1 I_3618  ( .D(I64230), .CLK(I2702), .RSTB(I64001), .Q(I64247) );
nor I_3619 (I64264,I64247,I64100);
nor I_3620 (I64281,I64247,I64162);
nand I_3621 (I63987,I64052,I64281);
nand I_3622 (I64312,I64018,I357713);
nand I_3623 (I64329,I64312,I64247);
and I_3624 (I64346,I64312,I64329);
DFFARX1 I_3625  ( .D(I64346), .CLK(I2702), .RSTB(I64001), .Q(I63969) );
DFFARX1 I_3626  ( .D(I64312), .CLK(I2702), .RSTB(I64001), .Q(I64377) );
and I_3627 (I63966,I64145,I64377);
DFFARX1 I_3628  ( .D(I357689), .CLK(I2702), .RSTB(I64001), .Q(I64408) );
not I_3629 (I64425,I64408);
nor I_3630 (I64442,I64100,I64425);
and I_3631 (I64459,I64408,I64442);
nand I_3632 (I63981,I64408,I64162);
DFFARX1 I_3633  ( .D(I64408), .CLK(I2702), .RSTB(I64001), .Q(I64490) );
not I_3634 (I63978,I64490);
DFFARX1 I_3635  ( .D(I357710), .CLK(I2702), .RSTB(I64001), .Q(I64521) );
not I_3636 (I64538,I64521);
or I_3637 (I64555,I64538,I64459);
DFFARX1 I_3638  ( .D(I64555), .CLK(I2702), .RSTB(I64001), .Q(I63984) );
nand I_3639 (I63993,I64538,I64264);
DFFARX1 I_3640  ( .D(I64538), .CLK(I2702), .RSTB(I64001), .Q(I63963) );
not I_3641 (I64647,I2709);
not I_3642 (I64664,I266196);
nor I_3643 (I64681,I266193,I266181);
nand I_3644 (I64698,I64681,I266184);
DFFARX1 I_3645  ( .D(I64698), .CLK(I2702), .RSTB(I64647), .Q(I64621) );
nor I_3646 (I64729,I64664,I266193);
nand I_3647 (I64746,I64729,I266190);
not I_3648 (I64636,I64746);
DFFARX1 I_3649  ( .D(I64746), .CLK(I2702), .RSTB(I64647), .Q(I64618) );
not I_3650 (I64791,I266193);
not I_3651 (I64808,I64791);
not I_3652 (I64825,I266202);
nor I_3653 (I64842,I64825,I266178);
and I_3654 (I64859,I64842,I266199);
or I_3655 (I64876,I64859,I266187);
DFFARX1 I_3656  ( .D(I64876), .CLK(I2702), .RSTB(I64647), .Q(I64893) );
nor I_3657 (I64910,I64893,I64746);
nor I_3658 (I64927,I64893,I64808);
nand I_3659 (I64633,I64698,I64927);
nand I_3660 (I64958,I64664,I266202);
nand I_3661 (I64975,I64958,I64893);
and I_3662 (I64992,I64958,I64975);
DFFARX1 I_3663  ( .D(I64992), .CLK(I2702), .RSTB(I64647), .Q(I64615) );
DFFARX1 I_3664  ( .D(I64958), .CLK(I2702), .RSTB(I64647), .Q(I65023) );
and I_3665 (I64612,I64791,I65023);
DFFARX1 I_3666  ( .D(I266208), .CLK(I2702), .RSTB(I64647), .Q(I65054) );
not I_3667 (I65071,I65054);
nor I_3668 (I65088,I64746,I65071);
and I_3669 (I65105,I65054,I65088);
nand I_3670 (I64627,I65054,I64808);
DFFARX1 I_3671  ( .D(I65054), .CLK(I2702), .RSTB(I64647), .Q(I65136) );
not I_3672 (I64624,I65136);
DFFARX1 I_3673  ( .D(I266205), .CLK(I2702), .RSTB(I64647), .Q(I65167) );
not I_3674 (I65184,I65167);
or I_3675 (I65201,I65184,I65105);
DFFARX1 I_3676  ( .D(I65201), .CLK(I2702), .RSTB(I64647), .Q(I64630) );
nand I_3677 (I64639,I65184,I64910);
DFFARX1 I_3678  ( .D(I65184), .CLK(I2702), .RSTB(I64647), .Q(I64609) );
not I_3679 (I65293,I2709);
not I_3680 (I65310,I409387);
nor I_3681 (I65327,I409399,I409381);
nand I_3682 (I65344,I65327,I409396);
DFFARX1 I_3683  ( .D(I65344), .CLK(I2702), .RSTB(I65293), .Q(I65267) );
nor I_3684 (I65375,I65310,I409399);
nand I_3685 (I65392,I65375,I409384);
not I_3686 (I65282,I65392);
DFFARX1 I_3687  ( .D(I65392), .CLK(I2702), .RSTB(I65293), .Q(I65264) );
not I_3688 (I65437,I409399);
not I_3689 (I65454,I65437);
not I_3690 (I65471,I409393);
nor I_3691 (I65488,I65471,I409372);
and I_3692 (I65505,I65488,I409375);
or I_3693 (I65522,I65505,I409378);
DFFARX1 I_3694  ( .D(I65522), .CLK(I2702), .RSTB(I65293), .Q(I65539) );
nor I_3695 (I65556,I65539,I65392);
nor I_3696 (I65573,I65539,I65454);
nand I_3697 (I65279,I65344,I65573);
nand I_3698 (I65604,I65310,I409393);
nand I_3699 (I65621,I65604,I65539);
and I_3700 (I65638,I65604,I65621);
DFFARX1 I_3701  ( .D(I65638), .CLK(I2702), .RSTB(I65293), .Q(I65261) );
DFFARX1 I_3702  ( .D(I65604), .CLK(I2702), .RSTB(I65293), .Q(I65669) );
and I_3703 (I65258,I65437,I65669);
DFFARX1 I_3704  ( .D(I409369), .CLK(I2702), .RSTB(I65293), .Q(I65700) );
not I_3705 (I65717,I65700);
nor I_3706 (I65734,I65392,I65717);
and I_3707 (I65751,I65700,I65734);
nand I_3708 (I65273,I65700,I65454);
DFFARX1 I_3709  ( .D(I65700), .CLK(I2702), .RSTB(I65293), .Q(I65782) );
not I_3710 (I65270,I65782);
DFFARX1 I_3711  ( .D(I409390), .CLK(I2702), .RSTB(I65293), .Q(I65813) );
not I_3712 (I65830,I65813);
or I_3713 (I65847,I65830,I65751);
DFFARX1 I_3714  ( .D(I65847), .CLK(I2702), .RSTB(I65293), .Q(I65276) );
nand I_3715 (I65285,I65830,I65556);
DFFARX1 I_3716  ( .D(I65830), .CLK(I2702), .RSTB(I65293), .Q(I65255) );
not I_3717 (I65939,I2709);
not I_3718 (I65956,I708867);
nor I_3719 (I65973,I708864,I708861);
nand I_3720 (I65990,I65973,I708882);
DFFARX1 I_3721  ( .D(I65990), .CLK(I2702), .RSTB(I65939), .Q(I65913) );
nor I_3722 (I66021,I65956,I708864);
nand I_3723 (I66038,I66021,I708885);
not I_3724 (I65928,I66038);
DFFARX1 I_3725  ( .D(I66038), .CLK(I2702), .RSTB(I65939), .Q(I65910) );
not I_3726 (I66083,I708864);
not I_3727 (I66100,I66083);
not I_3728 (I66117,I708858);
nor I_3729 (I66134,I66117,I708870);
and I_3730 (I66151,I66134,I708879);
or I_3731 (I66168,I66151,I708873);
DFFARX1 I_3732  ( .D(I66168), .CLK(I2702), .RSTB(I65939), .Q(I66185) );
nor I_3733 (I66202,I66185,I66038);
nor I_3734 (I66219,I66185,I66100);
nand I_3735 (I65925,I65990,I66219);
nand I_3736 (I66250,I65956,I708858);
nand I_3737 (I66267,I66250,I66185);
and I_3738 (I66284,I66250,I66267);
DFFARX1 I_3739  ( .D(I66284), .CLK(I2702), .RSTB(I65939), .Q(I65907) );
DFFARX1 I_3740  ( .D(I66250), .CLK(I2702), .RSTB(I65939), .Q(I66315) );
and I_3741 (I65904,I66083,I66315);
DFFARX1 I_3742  ( .D(I708888), .CLK(I2702), .RSTB(I65939), .Q(I66346) );
not I_3743 (I66363,I66346);
nor I_3744 (I66380,I66038,I66363);
and I_3745 (I66397,I66346,I66380);
nand I_3746 (I65919,I66346,I66100);
DFFARX1 I_3747  ( .D(I66346), .CLK(I2702), .RSTB(I65939), .Q(I66428) );
not I_3748 (I65916,I66428);
DFFARX1 I_3749  ( .D(I708876), .CLK(I2702), .RSTB(I65939), .Q(I66459) );
not I_3750 (I66476,I66459);
or I_3751 (I66493,I66476,I66397);
DFFARX1 I_3752  ( .D(I66493), .CLK(I2702), .RSTB(I65939), .Q(I65922) );
nand I_3753 (I65931,I66476,I66202);
DFFARX1 I_3754  ( .D(I66476), .CLK(I2702), .RSTB(I65939), .Q(I65901) );
not I_3755 (I66585,I2709);
not I_3756 (I66602,I613129);
nor I_3757 (I66619,I613114,I613141);
nand I_3758 (I66636,I66619,I613117);
DFFARX1 I_3759  ( .D(I66636), .CLK(I2702), .RSTB(I66585), .Q(I66559) );
nor I_3760 (I66667,I66602,I613114);
nand I_3761 (I66684,I66667,I613132);
not I_3762 (I66574,I66684);
DFFARX1 I_3763  ( .D(I66684), .CLK(I2702), .RSTB(I66585), .Q(I66556) );
not I_3764 (I66729,I613114);
not I_3765 (I66746,I66729);
not I_3766 (I66763,I613144);
nor I_3767 (I66780,I66763,I613126);
and I_3768 (I66797,I66780,I613135);
or I_3769 (I66814,I66797,I613120);
DFFARX1 I_3770  ( .D(I66814), .CLK(I2702), .RSTB(I66585), .Q(I66831) );
nor I_3771 (I66848,I66831,I66684);
nor I_3772 (I66865,I66831,I66746);
nand I_3773 (I66571,I66636,I66865);
nand I_3774 (I66896,I66602,I613144);
nand I_3775 (I66913,I66896,I66831);
and I_3776 (I66930,I66896,I66913);
DFFARX1 I_3777  ( .D(I66930), .CLK(I2702), .RSTB(I66585), .Q(I66553) );
DFFARX1 I_3778  ( .D(I66896), .CLK(I2702), .RSTB(I66585), .Q(I66961) );
and I_3779 (I66550,I66729,I66961);
DFFARX1 I_3780  ( .D(I613123), .CLK(I2702), .RSTB(I66585), .Q(I66992) );
not I_3781 (I67009,I66992);
nor I_3782 (I67026,I66684,I67009);
and I_3783 (I67043,I66992,I67026);
nand I_3784 (I66565,I66992,I66746);
DFFARX1 I_3785  ( .D(I66992), .CLK(I2702), .RSTB(I66585), .Q(I67074) );
not I_3786 (I66562,I67074);
DFFARX1 I_3787  ( .D(I613138), .CLK(I2702), .RSTB(I66585), .Q(I67105) );
not I_3788 (I67122,I67105);
or I_3789 (I67139,I67122,I67043);
DFFARX1 I_3790  ( .D(I67139), .CLK(I2702), .RSTB(I66585), .Q(I66568) );
nand I_3791 (I66577,I67122,I66848);
DFFARX1 I_3792  ( .D(I67122), .CLK(I2702), .RSTB(I66585), .Q(I66547) );
not I_3793 (I67231,I2709);
not I_3794 (I67248,I289401);
nor I_3795 (I67265,I289398,I289386);
nand I_3796 (I67282,I67265,I289389);
DFFARX1 I_3797  ( .D(I67282), .CLK(I2702), .RSTB(I67231), .Q(I67205) );
nor I_3798 (I67313,I67248,I289398);
nand I_3799 (I67330,I67313,I289395);
not I_3800 (I67220,I67330);
DFFARX1 I_3801  ( .D(I67330), .CLK(I2702), .RSTB(I67231), .Q(I67202) );
not I_3802 (I67375,I289398);
not I_3803 (I67392,I67375);
not I_3804 (I67409,I289407);
nor I_3805 (I67426,I67409,I289383);
and I_3806 (I67443,I67426,I289404);
or I_3807 (I67460,I67443,I289392);
DFFARX1 I_3808  ( .D(I67460), .CLK(I2702), .RSTB(I67231), .Q(I67477) );
nor I_3809 (I67494,I67477,I67330);
nor I_3810 (I67511,I67477,I67392);
nand I_3811 (I67217,I67282,I67511);
nand I_3812 (I67542,I67248,I289407);
nand I_3813 (I67559,I67542,I67477);
and I_3814 (I67576,I67542,I67559);
DFFARX1 I_3815  ( .D(I67576), .CLK(I2702), .RSTB(I67231), .Q(I67199) );
DFFARX1 I_3816  ( .D(I67542), .CLK(I2702), .RSTB(I67231), .Q(I67607) );
and I_3817 (I67196,I67375,I67607);
DFFARX1 I_3818  ( .D(I289413), .CLK(I2702), .RSTB(I67231), .Q(I67638) );
not I_3819 (I67655,I67638);
nor I_3820 (I67672,I67330,I67655);
and I_3821 (I67689,I67638,I67672);
nand I_3822 (I67211,I67638,I67392);
DFFARX1 I_3823  ( .D(I67638), .CLK(I2702), .RSTB(I67231), .Q(I67720) );
not I_3824 (I67208,I67720);
DFFARX1 I_3825  ( .D(I289410), .CLK(I2702), .RSTB(I67231), .Q(I67751) );
not I_3826 (I67768,I67751);
or I_3827 (I67785,I67768,I67689);
DFFARX1 I_3828  ( .D(I67785), .CLK(I2702), .RSTB(I67231), .Q(I67214) );
nand I_3829 (I67223,I67768,I67494);
DFFARX1 I_3830  ( .D(I67768), .CLK(I2702), .RSTB(I67231), .Q(I67193) );
not I_3831 (I67877,I2709);
not I_3832 (I67894,I503703);
nor I_3833 (I67911,I503715,I503697);
nand I_3834 (I67928,I67911,I503706);
DFFARX1 I_3835  ( .D(I67928), .CLK(I2702), .RSTB(I67877), .Q(I67851) );
nor I_3836 (I67959,I67894,I503715);
nand I_3837 (I67976,I67959,I503712);
not I_3838 (I67866,I67976);
DFFARX1 I_3839  ( .D(I67976), .CLK(I2702), .RSTB(I67877), .Q(I67848) );
not I_3840 (I68021,I503715);
not I_3841 (I68038,I68021);
not I_3842 (I68055,I503685);
nor I_3843 (I68072,I68055,I503688);
and I_3844 (I68089,I68072,I503694);
or I_3845 (I68106,I68089,I503709);
DFFARX1 I_3846  ( .D(I68106), .CLK(I2702), .RSTB(I67877), .Q(I68123) );
nor I_3847 (I68140,I68123,I67976);
nor I_3848 (I68157,I68123,I68038);
nand I_3849 (I67863,I67928,I68157);
nand I_3850 (I68188,I67894,I503685);
nand I_3851 (I68205,I68188,I68123);
and I_3852 (I68222,I68188,I68205);
DFFARX1 I_3853  ( .D(I68222), .CLK(I2702), .RSTB(I67877), .Q(I67845) );
DFFARX1 I_3854  ( .D(I68188), .CLK(I2702), .RSTB(I67877), .Q(I68253) );
and I_3855 (I67842,I68021,I68253);
DFFARX1 I_3856  ( .D(I503691), .CLK(I2702), .RSTB(I67877), .Q(I68284) );
not I_3857 (I68301,I68284);
nor I_3858 (I68318,I67976,I68301);
and I_3859 (I68335,I68284,I68318);
nand I_3860 (I67857,I68284,I68038);
DFFARX1 I_3861  ( .D(I68284), .CLK(I2702), .RSTB(I67877), .Q(I68366) );
not I_3862 (I67854,I68366);
DFFARX1 I_3863  ( .D(I503700), .CLK(I2702), .RSTB(I67877), .Q(I68397) );
not I_3864 (I68414,I68397);
or I_3865 (I68431,I68414,I68335);
DFFARX1 I_3866  ( .D(I68431), .CLK(I2702), .RSTB(I67877), .Q(I67860) );
nand I_3867 (I67869,I68414,I68140);
DFFARX1 I_3868  ( .D(I68414), .CLK(I2702), .RSTB(I67877), .Q(I67839) );
not I_3869 (I68523,I2709);
not I_3870 (I68540,I397759);
nor I_3871 (I68557,I397771,I397753);
nand I_3872 (I68574,I68557,I397768);
DFFARX1 I_3873  ( .D(I68574), .CLK(I2702), .RSTB(I68523), .Q(I68497) );
nor I_3874 (I68605,I68540,I397771);
nand I_3875 (I68622,I68605,I397756);
not I_3876 (I68512,I68622);
DFFARX1 I_3877  ( .D(I68622), .CLK(I2702), .RSTB(I68523), .Q(I68494) );
not I_3878 (I68667,I397771);
not I_3879 (I68684,I68667);
not I_3880 (I68701,I397765);
nor I_3881 (I68718,I68701,I397744);
and I_3882 (I68735,I68718,I397747);
or I_3883 (I68752,I68735,I397750);
DFFARX1 I_3884  ( .D(I68752), .CLK(I2702), .RSTB(I68523), .Q(I68769) );
nor I_3885 (I68786,I68769,I68622);
nor I_3886 (I68803,I68769,I68684);
nand I_3887 (I68509,I68574,I68803);
nand I_3888 (I68834,I68540,I397765);
nand I_3889 (I68851,I68834,I68769);
and I_3890 (I68868,I68834,I68851);
DFFARX1 I_3891  ( .D(I68868), .CLK(I2702), .RSTB(I68523), .Q(I68491) );
DFFARX1 I_3892  ( .D(I68834), .CLK(I2702), .RSTB(I68523), .Q(I68899) );
and I_3893 (I68488,I68667,I68899);
DFFARX1 I_3894  ( .D(I397741), .CLK(I2702), .RSTB(I68523), .Q(I68930) );
not I_3895 (I68947,I68930);
nor I_3896 (I68964,I68622,I68947);
and I_3897 (I68981,I68930,I68964);
nand I_3898 (I68503,I68930,I68684);
DFFARX1 I_3899  ( .D(I68930), .CLK(I2702), .RSTB(I68523), .Q(I69012) );
not I_3900 (I68500,I69012);
DFFARX1 I_3901  ( .D(I397762), .CLK(I2702), .RSTB(I68523), .Q(I69043) );
not I_3902 (I69060,I69043);
or I_3903 (I69077,I69060,I68981);
DFFARX1 I_3904  ( .D(I69077), .CLK(I2702), .RSTB(I68523), .Q(I68506) );
nand I_3905 (I68515,I69060,I68786);
DFFARX1 I_3906  ( .D(I69060), .CLK(I2702), .RSTB(I68523), .Q(I68485) );
not I_3907 (I69169,I2709);
not I_3908 (I69186,I693261);
nor I_3909 (I69203,I693258,I693255);
nand I_3910 (I69220,I69203,I693276);
DFFARX1 I_3911  ( .D(I69220), .CLK(I2702), .RSTB(I69169), .Q(I69143) );
nor I_3912 (I69251,I69186,I693258);
nand I_3913 (I69268,I69251,I693279);
not I_3914 (I69158,I69268);
DFFARX1 I_3915  ( .D(I69268), .CLK(I2702), .RSTB(I69169), .Q(I69140) );
not I_3916 (I69313,I693258);
not I_3917 (I69330,I69313);
not I_3918 (I69347,I693252);
nor I_3919 (I69364,I69347,I693264);
and I_3920 (I69381,I69364,I693273);
or I_3921 (I69398,I69381,I693267);
DFFARX1 I_3922  ( .D(I69398), .CLK(I2702), .RSTB(I69169), .Q(I69415) );
nor I_3923 (I69432,I69415,I69268);
nor I_3924 (I69449,I69415,I69330);
nand I_3925 (I69155,I69220,I69449);
nand I_3926 (I69480,I69186,I693252);
nand I_3927 (I69497,I69480,I69415);
and I_3928 (I69514,I69480,I69497);
DFFARX1 I_3929  ( .D(I69514), .CLK(I2702), .RSTB(I69169), .Q(I69137) );
DFFARX1 I_3930  ( .D(I69480), .CLK(I2702), .RSTB(I69169), .Q(I69545) );
and I_3931 (I69134,I69313,I69545);
DFFARX1 I_3932  ( .D(I693282), .CLK(I2702), .RSTB(I69169), .Q(I69576) );
not I_3933 (I69593,I69576);
nor I_3934 (I69610,I69268,I69593);
and I_3935 (I69627,I69576,I69610);
nand I_3936 (I69149,I69576,I69330);
DFFARX1 I_3937  ( .D(I69576), .CLK(I2702), .RSTB(I69169), .Q(I69658) );
not I_3938 (I69146,I69658);
DFFARX1 I_3939  ( .D(I693270), .CLK(I2702), .RSTB(I69169), .Q(I69689) );
not I_3940 (I69706,I69689);
or I_3941 (I69723,I69706,I69627);
DFFARX1 I_3942  ( .D(I69723), .CLK(I2702), .RSTB(I69169), .Q(I69152) );
nand I_3943 (I69161,I69706,I69432);
DFFARX1 I_3944  ( .D(I69706), .CLK(I2702), .RSTB(I69169), .Q(I69131) );
not I_3945 (I69815,I2709);
not I_3946 (I69832,I1399);
nor I_3947 (I69849,I1423,I2223);
nand I_3948 (I69866,I69849,I2295);
DFFARX1 I_3949  ( .D(I69866), .CLK(I2702), .RSTB(I69815), .Q(I69789) );
nor I_3950 (I69897,I69832,I1423);
nand I_3951 (I69914,I69897,I1303);
not I_3952 (I69804,I69914);
DFFARX1 I_3953  ( .D(I69914), .CLK(I2702), .RSTB(I69815), .Q(I69786) );
not I_3954 (I69959,I1423);
not I_3955 (I69976,I69959);
not I_3956 (I69993,I1375);
nor I_3957 (I70010,I69993,I2535);
and I_3958 (I70027,I70010,I2007);
or I_3959 (I70044,I70027,I1351);
DFFARX1 I_3960  ( .D(I70044), .CLK(I2702), .RSTB(I69815), .Q(I70061) );
nor I_3961 (I70078,I70061,I69914);
nor I_3962 (I70095,I70061,I69976);
nand I_3963 (I69801,I69866,I70095);
nand I_3964 (I70126,I69832,I1375);
nand I_3965 (I70143,I70126,I70061);
and I_3966 (I70160,I70126,I70143);
DFFARX1 I_3967  ( .D(I70160), .CLK(I2702), .RSTB(I69815), .Q(I69783) );
DFFARX1 I_3968  ( .D(I70126), .CLK(I2702), .RSTB(I69815), .Q(I70191) );
and I_3969 (I69780,I69959,I70191);
DFFARX1 I_3970  ( .D(I1527), .CLK(I2702), .RSTB(I69815), .Q(I70222) );
not I_3971 (I70239,I70222);
nor I_3972 (I70256,I69914,I70239);
and I_3973 (I70273,I70222,I70256);
nand I_3974 (I69795,I70222,I69976);
DFFARX1 I_3975  ( .D(I70222), .CLK(I2702), .RSTB(I69815), .Q(I70304) );
not I_3976 (I69792,I70304);
DFFARX1 I_3977  ( .D(I1879), .CLK(I2702), .RSTB(I69815), .Q(I70335) );
not I_3978 (I70352,I70335);
or I_3979 (I70369,I70352,I70273);
DFFARX1 I_3980  ( .D(I70369), .CLK(I2702), .RSTB(I69815), .Q(I69798) );
nand I_3981 (I69807,I70352,I70078);
DFFARX1 I_3982  ( .D(I70352), .CLK(I2702), .RSTB(I69815), .Q(I69777) );
not I_3983 (I70461,I2709);
not I_3984 (I70478,I465654);
nor I_3985 (I70495,I465642,I465648);
nand I_3986 (I70512,I70495,I465639);
DFFARX1 I_3987  ( .D(I70512), .CLK(I2702), .RSTB(I70461), .Q(I70435) );
nor I_3988 (I70543,I70478,I465642);
nand I_3989 (I70560,I70543,I465645);
not I_3990 (I70450,I70560);
DFFARX1 I_3991  ( .D(I70560), .CLK(I2702), .RSTB(I70461), .Q(I70432) );
not I_3992 (I70605,I465642);
not I_3993 (I70622,I70605);
not I_3994 (I70639,I465657);
nor I_3995 (I70656,I70639,I465669);
and I_3996 (I70673,I70656,I465651);
or I_3997 (I70690,I70673,I465666);
DFFARX1 I_3998  ( .D(I70690), .CLK(I2702), .RSTB(I70461), .Q(I70707) );
nor I_3999 (I70724,I70707,I70560);
nor I_4000 (I70741,I70707,I70622);
nand I_4001 (I70447,I70512,I70741);
nand I_4002 (I70772,I70478,I465657);
nand I_4003 (I70789,I70772,I70707);
and I_4004 (I70806,I70772,I70789);
DFFARX1 I_4005  ( .D(I70806), .CLK(I2702), .RSTB(I70461), .Q(I70429) );
DFFARX1 I_4006  ( .D(I70772), .CLK(I2702), .RSTB(I70461), .Q(I70837) );
and I_4007 (I70426,I70605,I70837);
DFFARX1 I_4008  ( .D(I465660), .CLK(I2702), .RSTB(I70461), .Q(I70868) );
not I_4009 (I70885,I70868);
nor I_4010 (I70902,I70560,I70885);
and I_4011 (I70919,I70868,I70902);
nand I_4012 (I70441,I70868,I70622);
DFFARX1 I_4013  ( .D(I70868), .CLK(I2702), .RSTB(I70461), .Q(I70950) );
not I_4014 (I70438,I70950);
DFFARX1 I_4015  ( .D(I465663), .CLK(I2702), .RSTB(I70461), .Q(I70981) );
not I_4016 (I70998,I70981);
or I_4017 (I71015,I70998,I70919);
DFFARX1 I_4018  ( .D(I71015), .CLK(I2702), .RSTB(I70461), .Q(I70444) );
nand I_4019 (I70453,I70998,I70724);
DFFARX1 I_4020  ( .D(I70998), .CLK(I2702), .RSTB(I70461), .Q(I70423) );
not I_4021 (I71107,I2709);
not I_4022 (I71124,I365459);
nor I_4023 (I71141,I365471,I365453);
nand I_4024 (I71158,I71141,I365468);
DFFARX1 I_4025  ( .D(I71158), .CLK(I2702), .RSTB(I71107), .Q(I71081) );
nor I_4026 (I71189,I71124,I365471);
nand I_4027 (I71206,I71189,I365456);
not I_4028 (I71096,I71206);
DFFARX1 I_4029  ( .D(I71206), .CLK(I2702), .RSTB(I71107), .Q(I71078) );
not I_4030 (I71251,I365471);
not I_4031 (I71268,I71251);
not I_4032 (I71285,I365465);
nor I_4033 (I71302,I71285,I365444);
and I_4034 (I71319,I71302,I365447);
or I_4035 (I71336,I71319,I365450);
DFFARX1 I_4036  ( .D(I71336), .CLK(I2702), .RSTB(I71107), .Q(I71353) );
nor I_4037 (I71370,I71353,I71206);
nor I_4038 (I71387,I71353,I71268);
nand I_4039 (I71093,I71158,I71387);
nand I_4040 (I71418,I71124,I365465);
nand I_4041 (I71435,I71418,I71353);
and I_4042 (I71452,I71418,I71435);
DFFARX1 I_4043  ( .D(I71452), .CLK(I2702), .RSTB(I71107), .Q(I71075) );
DFFARX1 I_4044  ( .D(I71418), .CLK(I2702), .RSTB(I71107), .Q(I71483) );
and I_4045 (I71072,I71251,I71483);
DFFARX1 I_4046  ( .D(I365441), .CLK(I2702), .RSTB(I71107), .Q(I71514) );
not I_4047 (I71531,I71514);
nor I_4048 (I71548,I71206,I71531);
and I_4049 (I71565,I71514,I71548);
nand I_4050 (I71087,I71514,I71268);
DFFARX1 I_4051  ( .D(I71514), .CLK(I2702), .RSTB(I71107), .Q(I71596) );
not I_4052 (I71084,I71596);
DFFARX1 I_4053  ( .D(I365462), .CLK(I2702), .RSTB(I71107), .Q(I71627) );
not I_4054 (I71644,I71627);
or I_4055 (I71661,I71644,I71565);
DFFARX1 I_4056  ( .D(I71661), .CLK(I2702), .RSTB(I71107), .Q(I71090) );
nand I_4057 (I71099,I71644,I71370);
DFFARX1 I_4058  ( .D(I71644), .CLK(I2702), .RSTB(I71107), .Q(I71069) );
not I_4059 (I71753,I2709);
not I_4060 (I71770,I466232);
nor I_4061 (I71787,I466220,I466226);
nand I_4062 (I71804,I71787,I466217);
DFFARX1 I_4063  ( .D(I71804), .CLK(I2702), .RSTB(I71753), .Q(I71727) );
nor I_4064 (I71835,I71770,I466220);
nand I_4065 (I71852,I71835,I466223);
not I_4066 (I71742,I71852);
DFFARX1 I_4067  ( .D(I71852), .CLK(I2702), .RSTB(I71753), .Q(I71724) );
not I_4068 (I71897,I466220);
not I_4069 (I71914,I71897);
not I_4070 (I71931,I466235);
nor I_4071 (I71948,I71931,I466247);
and I_4072 (I71965,I71948,I466229);
or I_4073 (I71982,I71965,I466244);
DFFARX1 I_4074  ( .D(I71982), .CLK(I2702), .RSTB(I71753), .Q(I71999) );
nor I_4075 (I72016,I71999,I71852);
nor I_4076 (I72033,I71999,I71914);
nand I_4077 (I71739,I71804,I72033);
nand I_4078 (I72064,I71770,I466235);
nand I_4079 (I72081,I72064,I71999);
and I_4080 (I72098,I72064,I72081);
DFFARX1 I_4081  ( .D(I72098), .CLK(I2702), .RSTB(I71753), .Q(I71721) );
DFFARX1 I_4082  ( .D(I72064), .CLK(I2702), .RSTB(I71753), .Q(I72129) );
and I_4083 (I71718,I71897,I72129);
DFFARX1 I_4084  ( .D(I466238), .CLK(I2702), .RSTB(I71753), .Q(I72160) );
not I_4085 (I72177,I72160);
nor I_4086 (I72194,I71852,I72177);
and I_4087 (I72211,I72160,I72194);
nand I_4088 (I71733,I72160,I71914);
DFFARX1 I_4089  ( .D(I72160), .CLK(I2702), .RSTB(I71753), .Q(I72242) );
not I_4090 (I71730,I72242);
DFFARX1 I_4091  ( .D(I466241), .CLK(I2702), .RSTB(I71753), .Q(I72273) );
not I_4092 (I72290,I72273);
or I_4093 (I72307,I72290,I72211);
DFFARX1 I_4094  ( .D(I72307), .CLK(I2702), .RSTB(I71753), .Q(I71736) );
nand I_4095 (I71745,I72290,I72016);
DFFARX1 I_4096  ( .D(I72290), .CLK(I2702), .RSTB(I71753), .Q(I71715) );
not I_4097 (I72399,I2709);
not I_4098 (I72416,I610154);
nor I_4099 (I72433,I610139,I610166);
nand I_4100 (I72450,I72433,I610142);
DFFARX1 I_4101  ( .D(I72450), .CLK(I2702), .RSTB(I72399), .Q(I72373) );
nor I_4102 (I72481,I72416,I610139);
nand I_4103 (I72498,I72481,I610157);
not I_4104 (I72388,I72498);
DFFARX1 I_4105  ( .D(I72498), .CLK(I2702), .RSTB(I72399), .Q(I72370) );
not I_4106 (I72543,I610139);
not I_4107 (I72560,I72543);
not I_4108 (I72577,I610169);
nor I_4109 (I72594,I72577,I610151);
and I_4110 (I72611,I72594,I610160);
or I_4111 (I72628,I72611,I610145);
DFFARX1 I_4112  ( .D(I72628), .CLK(I2702), .RSTB(I72399), .Q(I72645) );
nor I_4113 (I72662,I72645,I72498);
nor I_4114 (I72679,I72645,I72560);
nand I_4115 (I72385,I72450,I72679);
nand I_4116 (I72710,I72416,I610169);
nand I_4117 (I72727,I72710,I72645);
and I_4118 (I72744,I72710,I72727);
DFFARX1 I_4119  ( .D(I72744), .CLK(I2702), .RSTB(I72399), .Q(I72367) );
DFFARX1 I_4120  ( .D(I72710), .CLK(I2702), .RSTB(I72399), .Q(I72775) );
and I_4121 (I72364,I72543,I72775);
DFFARX1 I_4122  ( .D(I610148), .CLK(I2702), .RSTB(I72399), .Q(I72806) );
not I_4123 (I72823,I72806);
nor I_4124 (I72840,I72498,I72823);
and I_4125 (I72857,I72806,I72840);
nand I_4126 (I72379,I72806,I72560);
DFFARX1 I_4127  ( .D(I72806), .CLK(I2702), .RSTB(I72399), .Q(I72888) );
not I_4128 (I72376,I72888);
DFFARX1 I_4129  ( .D(I610163), .CLK(I2702), .RSTB(I72399), .Q(I72919) );
not I_4130 (I72936,I72919);
or I_4131 (I72953,I72936,I72857);
DFFARX1 I_4132  ( .D(I72953), .CLK(I2702), .RSTB(I72399), .Q(I72382) );
nand I_4133 (I72391,I72936,I72662);
DFFARX1 I_4134  ( .D(I72936), .CLK(I2702), .RSTB(I72399), .Q(I72361) );
not I_4135 (I73045,I2709);
not I_4136 (I73062,I22911);
nor I_4137 (I73079,I22923,I22908);
nand I_4138 (I73096,I73079,I22920);
DFFARX1 I_4139  ( .D(I73096), .CLK(I2702), .RSTB(I73045), .Q(I73019) );
nor I_4140 (I73127,I73062,I22923);
nand I_4141 (I73144,I73127,I22938);
not I_4142 (I73034,I73144);
DFFARX1 I_4143  ( .D(I73144), .CLK(I2702), .RSTB(I73045), .Q(I73016) );
not I_4144 (I73189,I22923);
not I_4145 (I73206,I73189);
not I_4146 (I73223,I22914);
nor I_4147 (I73240,I73223,I22926);
and I_4148 (I73257,I73240,I22917);
or I_4149 (I73274,I73257,I22932);
DFFARX1 I_4150  ( .D(I73274), .CLK(I2702), .RSTB(I73045), .Q(I73291) );
nor I_4151 (I73308,I73291,I73144);
nor I_4152 (I73325,I73291,I73206);
nand I_4153 (I73031,I73096,I73325);
nand I_4154 (I73356,I73062,I22914);
nand I_4155 (I73373,I73356,I73291);
and I_4156 (I73390,I73356,I73373);
DFFARX1 I_4157  ( .D(I73390), .CLK(I2702), .RSTB(I73045), .Q(I73013) );
DFFARX1 I_4158  ( .D(I73356), .CLK(I2702), .RSTB(I73045), .Q(I73421) );
and I_4159 (I73010,I73189,I73421);
DFFARX1 I_4160  ( .D(I22935), .CLK(I2702), .RSTB(I73045), .Q(I73452) );
not I_4161 (I73469,I73452);
nor I_4162 (I73486,I73144,I73469);
and I_4163 (I73503,I73452,I73486);
nand I_4164 (I73025,I73452,I73206);
DFFARX1 I_4165  ( .D(I73452), .CLK(I2702), .RSTB(I73045), .Q(I73534) );
not I_4166 (I73022,I73534);
DFFARX1 I_4167  ( .D(I22929), .CLK(I2702), .RSTB(I73045), .Q(I73565) );
not I_4168 (I73582,I73565);
or I_4169 (I73599,I73582,I73503);
DFFARX1 I_4170  ( .D(I73599), .CLK(I2702), .RSTB(I73045), .Q(I73028) );
nand I_4171 (I73037,I73582,I73308);
DFFARX1 I_4172  ( .D(I73582), .CLK(I2702), .RSTB(I73045), .Q(I73007) );
not I_4173 (I73691,I2709);
not I_4174 (I73708,I497345);
nor I_4175 (I73725,I497357,I497339);
nand I_4176 (I73742,I73725,I497348);
DFFARX1 I_4177  ( .D(I73742), .CLK(I2702), .RSTB(I73691), .Q(I73665) );
nor I_4178 (I73773,I73708,I497357);
nand I_4179 (I73790,I73773,I497354);
not I_4180 (I73680,I73790);
DFFARX1 I_4181  ( .D(I73790), .CLK(I2702), .RSTB(I73691), .Q(I73662) );
not I_4182 (I73835,I497357);
not I_4183 (I73852,I73835);
not I_4184 (I73869,I497327);
nor I_4185 (I73886,I73869,I497330);
and I_4186 (I73903,I73886,I497336);
or I_4187 (I73920,I73903,I497351);
DFFARX1 I_4188  ( .D(I73920), .CLK(I2702), .RSTB(I73691), .Q(I73937) );
nor I_4189 (I73954,I73937,I73790);
nor I_4190 (I73971,I73937,I73852);
nand I_4191 (I73677,I73742,I73971);
nand I_4192 (I74002,I73708,I497327);
nand I_4193 (I74019,I74002,I73937);
and I_4194 (I74036,I74002,I74019);
DFFARX1 I_4195  ( .D(I74036), .CLK(I2702), .RSTB(I73691), .Q(I73659) );
DFFARX1 I_4196  ( .D(I74002), .CLK(I2702), .RSTB(I73691), .Q(I74067) );
and I_4197 (I73656,I73835,I74067);
DFFARX1 I_4198  ( .D(I497333), .CLK(I2702), .RSTB(I73691), .Q(I74098) );
not I_4199 (I74115,I74098);
nor I_4200 (I74132,I73790,I74115);
and I_4201 (I74149,I74098,I74132);
nand I_4202 (I73671,I74098,I73852);
DFFARX1 I_4203  ( .D(I74098), .CLK(I2702), .RSTB(I73691), .Q(I74180) );
not I_4204 (I73668,I74180);
DFFARX1 I_4205  ( .D(I497342), .CLK(I2702), .RSTB(I73691), .Q(I74211) );
not I_4206 (I74228,I74211);
or I_4207 (I74245,I74228,I74149);
DFFARX1 I_4208  ( .D(I74245), .CLK(I2702), .RSTB(I73691), .Q(I73674) );
nand I_4209 (I73683,I74228,I73954);
DFFARX1 I_4210  ( .D(I74228), .CLK(I2702), .RSTB(I73691), .Q(I73653) );
not I_4211 (I74337,I2709);
not I_4212 (I74354,I309291);
nor I_4213 (I74371,I309288,I309276);
nand I_4214 (I74388,I74371,I309279);
DFFARX1 I_4215  ( .D(I74388), .CLK(I2702), .RSTB(I74337), .Q(I74311) );
nor I_4216 (I74419,I74354,I309288);
nand I_4217 (I74436,I74419,I309285);
not I_4218 (I74326,I74436);
DFFARX1 I_4219  ( .D(I74436), .CLK(I2702), .RSTB(I74337), .Q(I74308) );
not I_4220 (I74481,I309288);
not I_4221 (I74498,I74481);
not I_4222 (I74515,I309297);
nor I_4223 (I74532,I74515,I309273);
and I_4224 (I74549,I74532,I309294);
or I_4225 (I74566,I74549,I309282);
DFFARX1 I_4226  ( .D(I74566), .CLK(I2702), .RSTB(I74337), .Q(I74583) );
nor I_4227 (I74600,I74583,I74436);
nor I_4228 (I74617,I74583,I74498);
nand I_4229 (I74323,I74388,I74617);
nand I_4230 (I74648,I74354,I309297);
nand I_4231 (I74665,I74648,I74583);
and I_4232 (I74682,I74648,I74665);
DFFARX1 I_4233  ( .D(I74682), .CLK(I2702), .RSTB(I74337), .Q(I74305) );
DFFARX1 I_4234  ( .D(I74648), .CLK(I2702), .RSTB(I74337), .Q(I74713) );
and I_4235 (I74302,I74481,I74713);
DFFARX1 I_4236  ( .D(I309303), .CLK(I2702), .RSTB(I74337), .Q(I74744) );
not I_4237 (I74761,I74744);
nor I_4238 (I74778,I74436,I74761);
and I_4239 (I74795,I74744,I74778);
nand I_4240 (I74317,I74744,I74498);
DFFARX1 I_4241  ( .D(I74744), .CLK(I2702), .RSTB(I74337), .Q(I74826) );
not I_4242 (I74314,I74826);
DFFARX1 I_4243  ( .D(I309300), .CLK(I2702), .RSTB(I74337), .Q(I74857) );
not I_4244 (I74874,I74857);
or I_4245 (I74891,I74874,I74795);
DFFARX1 I_4246  ( .D(I74891), .CLK(I2702), .RSTB(I74337), .Q(I74320) );
nand I_4247 (I74329,I74874,I74600);
DFFARX1 I_4248  ( .D(I74874), .CLK(I2702), .RSTB(I74337), .Q(I74299) );
not I_4249 (I74983,I2709);
not I_4250 (I75000,I3276);
nor I_4251 (I75017,I3288,I3273);
nand I_4252 (I75034,I75017,I3285);
DFFARX1 I_4253  ( .D(I75034), .CLK(I2702), .RSTB(I74983), .Q(I74957) );
nor I_4254 (I75065,I75000,I3288);
nand I_4255 (I75082,I75065,I3303);
not I_4256 (I74972,I75082);
DFFARX1 I_4257  ( .D(I75082), .CLK(I2702), .RSTB(I74983), .Q(I74954) );
not I_4258 (I75127,I3288);
not I_4259 (I75144,I75127);
not I_4260 (I75161,I3279);
nor I_4261 (I75178,I75161,I3291);
and I_4262 (I75195,I75178,I3282);
or I_4263 (I75212,I75195,I3297);
DFFARX1 I_4264  ( .D(I75212), .CLK(I2702), .RSTB(I74983), .Q(I75229) );
nor I_4265 (I75246,I75229,I75082);
nor I_4266 (I75263,I75229,I75144);
nand I_4267 (I74969,I75034,I75263);
nand I_4268 (I75294,I75000,I3279);
nand I_4269 (I75311,I75294,I75229);
and I_4270 (I75328,I75294,I75311);
DFFARX1 I_4271  ( .D(I75328), .CLK(I2702), .RSTB(I74983), .Q(I74951) );
DFFARX1 I_4272  ( .D(I75294), .CLK(I2702), .RSTB(I74983), .Q(I75359) );
and I_4273 (I74948,I75127,I75359);
DFFARX1 I_4274  ( .D(I3300), .CLK(I2702), .RSTB(I74983), .Q(I75390) );
not I_4275 (I75407,I75390);
nor I_4276 (I75424,I75082,I75407);
and I_4277 (I75441,I75390,I75424);
nand I_4278 (I74963,I75390,I75144);
DFFARX1 I_4279  ( .D(I75390), .CLK(I2702), .RSTB(I74983), .Q(I75472) );
not I_4280 (I74960,I75472);
DFFARX1 I_4281  ( .D(I3294), .CLK(I2702), .RSTB(I74983), .Q(I75503) );
not I_4282 (I75520,I75503);
or I_4283 (I75537,I75520,I75441);
DFFARX1 I_4284  ( .D(I75537), .CLK(I2702), .RSTB(I74983), .Q(I74966) );
nand I_4285 (I74975,I75520,I75246);
DFFARX1 I_4286  ( .D(I75520), .CLK(I2702), .RSTB(I74983), .Q(I74945) );
not I_4287 (I75629,I2709);
not I_4288 (I75646,I213563);
nor I_4289 (I75663,I213593,I213572);
nand I_4290 (I75680,I75663,I213584);
DFFARX1 I_4291  ( .D(I75680), .CLK(I2702), .RSTB(I75629), .Q(I75603) );
nor I_4292 (I75711,I75646,I213593);
nand I_4293 (I75728,I75711,I213566);
not I_4294 (I75618,I75728);
DFFARX1 I_4295  ( .D(I75728), .CLK(I2702), .RSTB(I75629), .Q(I75600) );
not I_4296 (I75773,I213593);
not I_4297 (I75790,I75773);
not I_4298 (I75807,I213569);
nor I_4299 (I75824,I75807,I213587);
and I_4300 (I75841,I75824,I213578);
or I_4301 (I75858,I75841,I213575);
DFFARX1 I_4302  ( .D(I75858), .CLK(I2702), .RSTB(I75629), .Q(I75875) );
nor I_4303 (I75892,I75875,I75728);
nor I_4304 (I75909,I75875,I75790);
nand I_4305 (I75615,I75680,I75909);
nand I_4306 (I75940,I75646,I213569);
nand I_4307 (I75957,I75940,I75875);
and I_4308 (I75974,I75940,I75957);
DFFARX1 I_4309  ( .D(I75974), .CLK(I2702), .RSTB(I75629), .Q(I75597) );
DFFARX1 I_4310  ( .D(I75940), .CLK(I2702), .RSTB(I75629), .Q(I76005) );
and I_4311 (I75594,I75773,I76005);
DFFARX1 I_4312  ( .D(I213581), .CLK(I2702), .RSTB(I75629), .Q(I76036) );
not I_4313 (I76053,I76036);
nor I_4314 (I76070,I75728,I76053);
and I_4315 (I76087,I76036,I76070);
nand I_4316 (I75609,I76036,I75790);
DFFARX1 I_4317  ( .D(I76036), .CLK(I2702), .RSTB(I75629), .Q(I76118) );
not I_4318 (I75606,I76118);
DFFARX1 I_4319  ( .D(I213590), .CLK(I2702), .RSTB(I75629), .Q(I76149) );
not I_4320 (I76166,I76149);
or I_4321 (I76183,I76166,I76087);
DFFARX1 I_4322  ( .D(I76183), .CLK(I2702), .RSTB(I75629), .Q(I75612) );
nand I_4323 (I75621,I76166,I75892);
DFFARX1 I_4324  ( .D(I76166), .CLK(I2702), .RSTB(I75629), .Q(I75591) );
not I_4325 (I76275,I2709);
not I_4326 (I76292,I362875);
nor I_4327 (I76309,I362887,I362869);
nand I_4328 (I76326,I76309,I362884);
DFFARX1 I_4329  ( .D(I76326), .CLK(I2702), .RSTB(I76275), .Q(I76249) );
nor I_4330 (I76357,I76292,I362887);
nand I_4331 (I76374,I76357,I362872);
not I_4332 (I76264,I76374);
DFFARX1 I_4333  ( .D(I76374), .CLK(I2702), .RSTB(I76275), .Q(I76246) );
not I_4334 (I76419,I362887);
not I_4335 (I76436,I76419);
not I_4336 (I76453,I362881);
nor I_4337 (I76470,I76453,I362860);
and I_4338 (I76487,I76470,I362863);
or I_4339 (I76504,I76487,I362866);
DFFARX1 I_4340  ( .D(I76504), .CLK(I2702), .RSTB(I76275), .Q(I76521) );
nor I_4341 (I76538,I76521,I76374);
nor I_4342 (I76555,I76521,I76436);
nand I_4343 (I76261,I76326,I76555);
nand I_4344 (I76586,I76292,I362881);
nand I_4345 (I76603,I76586,I76521);
and I_4346 (I76620,I76586,I76603);
DFFARX1 I_4347  ( .D(I76620), .CLK(I2702), .RSTB(I76275), .Q(I76243) );
DFFARX1 I_4348  ( .D(I76586), .CLK(I2702), .RSTB(I76275), .Q(I76651) );
and I_4349 (I76240,I76419,I76651);
DFFARX1 I_4350  ( .D(I362857), .CLK(I2702), .RSTB(I76275), .Q(I76682) );
not I_4351 (I76699,I76682);
nor I_4352 (I76716,I76374,I76699);
and I_4353 (I76733,I76682,I76716);
nand I_4354 (I76255,I76682,I76436);
DFFARX1 I_4355  ( .D(I76682), .CLK(I2702), .RSTB(I76275), .Q(I76764) );
not I_4356 (I76252,I76764);
DFFARX1 I_4357  ( .D(I362878), .CLK(I2702), .RSTB(I76275), .Q(I76795) );
not I_4358 (I76812,I76795);
or I_4359 (I76829,I76812,I76733);
DFFARX1 I_4360  ( .D(I76829), .CLK(I2702), .RSTB(I76275), .Q(I76258) );
nand I_4361 (I76267,I76812,I76538);
DFFARX1 I_4362  ( .D(I76812), .CLK(I2702), .RSTB(I76275), .Q(I76237) );
not I_4363 (I76921,I2709);
not I_4364 (I76938,I270837);
nor I_4365 (I76955,I270834,I270822);
nand I_4366 (I76972,I76955,I270825);
DFFARX1 I_4367  ( .D(I76972), .CLK(I2702), .RSTB(I76921), .Q(I76895) );
nor I_4368 (I77003,I76938,I270834);
nand I_4369 (I77020,I77003,I270831);
not I_4370 (I76910,I77020);
DFFARX1 I_4371  ( .D(I77020), .CLK(I2702), .RSTB(I76921), .Q(I76892) );
not I_4372 (I77065,I270834);
not I_4373 (I77082,I77065);
not I_4374 (I77099,I270843);
nor I_4375 (I77116,I77099,I270819);
and I_4376 (I77133,I77116,I270840);
or I_4377 (I77150,I77133,I270828);
DFFARX1 I_4378  ( .D(I77150), .CLK(I2702), .RSTB(I76921), .Q(I77167) );
nor I_4379 (I77184,I77167,I77020);
nor I_4380 (I77201,I77167,I77082);
nand I_4381 (I76907,I76972,I77201);
nand I_4382 (I77232,I76938,I270843);
nand I_4383 (I77249,I77232,I77167);
and I_4384 (I77266,I77232,I77249);
DFFARX1 I_4385  ( .D(I77266), .CLK(I2702), .RSTB(I76921), .Q(I76889) );
DFFARX1 I_4386  ( .D(I77232), .CLK(I2702), .RSTB(I76921), .Q(I77297) );
and I_4387 (I76886,I77065,I77297);
DFFARX1 I_4388  ( .D(I270849), .CLK(I2702), .RSTB(I76921), .Q(I77328) );
not I_4389 (I77345,I77328);
nor I_4390 (I77362,I77020,I77345);
and I_4391 (I77379,I77328,I77362);
nand I_4392 (I76901,I77328,I77082);
DFFARX1 I_4393  ( .D(I77328), .CLK(I2702), .RSTB(I76921), .Q(I77410) );
not I_4394 (I76898,I77410);
DFFARX1 I_4395  ( .D(I270846), .CLK(I2702), .RSTB(I76921), .Q(I77441) );
not I_4396 (I77458,I77441);
or I_4397 (I77475,I77458,I77379);
DFFARX1 I_4398  ( .D(I77475), .CLK(I2702), .RSTB(I76921), .Q(I76904) );
nand I_4399 (I76913,I77458,I77184);
DFFARX1 I_4400  ( .D(I77458), .CLK(I2702), .RSTB(I76921), .Q(I76883) );
not I_4401 (I77567,I2709);
not I_4402 (I77584,I622481);
nor I_4403 (I77601,I622496,I622511);
nand I_4404 (I77618,I77601,I622499);
DFFARX1 I_4405  ( .D(I77618), .CLK(I2702), .RSTB(I77567), .Q(I77541) );
nor I_4406 (I77649,I77584,I622496);
nand I_4407 (I77666,I77649,I622502);
not I_4408 (I77556,I77666);
DFFARX1 I_4409  ( .D(I77666), .CLK(I2702), .RSTB(I77567), .Q(I77538) );
not I_4410 (I77711,I622496);
not I_4411 (I77728,I77711);
not I_4412 (I77745,I622508);
nor I_4413 (I77762,I77745,I622505);
and I_4414 (I77779,I77762,I622484);
or I_4415 (I77796,I77779,I622493);
DFFARX1 I_4416  ( .D(I77796), .CLK(I2702), .RSTB(I77567), .Q(I77813) );
nor I_4417 (I77830,I77813,I77666);
nor I_4418 (I77847,I77813,I77728);
nand I_4419 (I77553,I77618,I77847);
nand I_4420 (I77878,I77584,I622508);
nand I_4421 (I77895,I77878,I77813);
and I_4422 (I77912,I77878,I77895);
DFFARX1 I_4423  ( .D(I77912), .CLK(I2702), .RSTB(I77567), .Q(I77535) );
DFFARX1 I_4424  ( .D(I77878), .CLK(I2702), .RSTB(I77567), .Q(I77943) );
and I_4425 (I77532,I77711,I77943);
DFFARX1 I_4426  ( .D(I622490), .CLK(I2702), .RSTB(I77567), .Q(I77974) );
not I_4427 (I77991,I77974);
nor I_4428 (I78008,I77666,I77991);
and I_4429 (I78025,I77974,I78008);
nand I_4430 (I77547,I77974,I77728);
DFFARX1 I_4431  ( .D(I77974), .CLK(I2702), .RSTB(I77567), .Q(I78056) );
not I_4432 (I77544,I78056);
DFFARX1 I_4433  ( .D(I622487), .CLK(I2702), .RSTB(I77567), .Q(I78087) );
not I_4434 (I78104,I78087);
or I_4435 (I78121,I78104,I78025);
DFFARX1 I_4436  ( .D(I78121), .CLK(I2702), .RSTB(I77567), .Q(I77550) );
nand I_4437 (I77559,I78104,I77830);
DFFARX1 I_4438  ( .D(I78104), .CLK(I2702), .RSTB(I77567), .Q(I77529) );
not I_4439 (I78213,I2709);
not I_4440 (I78230,I473746);
nor I_4441 (I78247,I473734,I473740);
nand I_4442 (I78264,I78247,I473731);
DFFARX1 I_4443  ( .D(I78264), .CLK(I2702), .RSTB(I78213), .Q(I78187) );
nor I_4444 (I78295,I78230,I473734);
nand I_4445 (I78312,I78295,I473737);
not I_4446 (I78202,I78312);
DFFARX1 I_4447  ( .D(I78312), .CLK(I2702), .RSTB(I78213), .Q(I78184) );
not I_4448 (I78357,I473734);
not I_4449 (I78374,I78357);
not I_4450 (I78391,I473749);
nor I_4451 (I78408,I78391,I473761);
and I_4452 (I78425,I78408,I473743);
or I_4453 (I78442,I78425,I473758);
DFFARX1 I_4454  ( .D(I78442), .CLK(I2702), .RSTB(I78213), .Q(I78459) );
nor I_4455 (I78476,I78459,I78312);
nor I_4456 (I78493,I78459,I78374);
nand I_4457 (I78199,I78264,I78493);
nand I_4458 (I78524,I78230,I473749);
nand I_4459 (I78541,I78524,I78459);
and I_4460 (I78558,I78524,I78541);
DFFARX1 I_4461  ( .D(I78558), .CLK(I2702), .RSTB(I78213), .Q(I78181) );
DFFARX1 I_4462  ( .D(I78524), .CLK(I2702), .RSTB(I78213), .Q(I78589) );
and I_4463 (I78178,I78357,I78589);
DFFARX1 I_4464  ( .D(I473752), .CLK(I2702), .RSTB(I78213), .Q(I78620) );
not I_4465 (I78637,I78620);
nor I_4466 (I78654,I78312,I78637);
and I_4467 (I78671,I78620,I78654);
nand I_4468 (I78193,I78620,I78374);
DFFARX1 I_4469  ( .D(I78620), .CLK(I2702), .RSTB(I78213), .Q(I78702) );
not I_4470 (I78190,I78702);
DFFARX1 I_4471  ( .D(I473755), .CLK(I2702), .RSTB(I78213), .Q(I78733) );
not I_4472 (I78750,I78733);
or I_4473 (I78767,I78750,I78671);
DFFARX1 I_4474  ( .D(I78767), .CLK(I2702), .RSTB(I78213), .Q(I78196) );
nand I_4475 (I78205,I78750,I78476);
DFFARX1 I_4476  ( .D(I78750), .CLK(I2702), .RSTB(I78213), .Q(I78175) );
not I_4477 (I78859,I2709);
not I_4478 (I78876,I504281);
nor I_4479 (I78893,I504293,I504275);
nand I_4480 (I78910,I78893,I504284);
DFFARX1 I_4481  ( .D(I78910), .CLK(I2702), .RSTB(I78859), .Q(I78833) );
nor I_4482 (I78941,I78876,I504293);
nand I_4483 (I78958,I78941,I504290);
not I_4484 (I78848,I78958);
DFFARX1 I_4485  ( .D(I78958), .CLK(I2702), .RSTB(I78859), .Q(I78830) );
not I_4486 (I79003,I504293);
not I_4487 (I79020,I79003);
not I_4488 (I79037,I504263);
nor I_4489 (I79054,I79037,I504266);
and I_4490 (I79071,I79054,I504272);
or I_4491 (I79088,I79071,I504287);
DFFARX1 I_4492  ( .D(I79088), .CLK(I2702), .RSTB(I78859), .Q(I79105) );
nor I_4493 (I79122,I79105,I78958);
nor I_4494 (I79139,I79105,I79020);
nand I_4495 (I78845,I78910,I79139);
nand I_4496 (I79170,I78876,I504263);
nand I_4497 (I79187,I79170,I79105);
and I_4498 (I79204,I79170,I79187);
DFFARX1 I_4499  ( .D(I79204), .CLK(I2702), .RSTB(I78859), .Q(I78827) );
DFFARX1 I_4500  ( .D(I79170), .CLK(I2702), .RSTB(I78859), .Q(I79235) );
and I_4501 (I78824,I79003,I79235);
DFFARX1 I_4502  ( .D(I504269), .CLK(I2702), .RSTB(I78859), .Q(I79266) );
not I_4503 (I79283,I79266);
nor I_4504 (I79300,I78958,I79283);
and I_4505 (I79317,I79266,I79300);
nand I_4506 (I78839,I79266,I79020);
DFFARX1 I_4507  ( .D(I79266), .CLK(I2702), .RSTB(I78859), .Q(I79348) );
not I_4508 (I78836,I79348);
DFFARX1 I_4509  ( .D(I504278), .CLK(I2702), .RSTB(I78859), .Q(I79379) );
not I_4510 (I79396,I79379);
or I_4511 (I79413,I79396,I79317);
DFFARX1 I_4512  ( .D(I79413), .CLK(I2702), .RSTB(I78859), .Q(I78842) );
nand I_4513 (I78851,I79396,I79122);
DFFARX1 I_4514  ( .D(I79396), .CLK(I2702), .RSTB(I78859), .Q(I78821) );
not I_4515 (I79505,I2709);
not I_4516 (I79522,I262881);
nor I_4517 (I79539,I262878,I262866);
nand I_4518 (I79556,I79539,I262869);
DFFARX1 I_4519  ( .D(I79556), .CLK(I2702), .RSTB(I79505), .Q(I79479) );
nor I_4520 (I79587,I79522,I262878);
nand I_4521 (I79604,I79587,I262875);
not I_4522 (I79494,I79604);
DFFARX1 I_4523  ( .D(I79604), .CLK(I2702), .RSTB(I79505), .Q(I79476) );
not I_4524 (I79649,I262878);
not I_4525 (I79666,I79649);
not I_4526 (I79683,I262887);
nor I_4527 (I79700,I79683,I262863);
and I_4528 (I79717,I79700,I262884);
or I_4529 (I79734,I79717,I262872);
DFFARX1 I_4530  ( .D(I79734), .CLK(I2702), .RSTB(I79505), .Q(I79751) );
nor I_4531 (I79768,I79751,I79604);
nor I_4532 (I79785,I79751,I79666);
nand I_4533 (I79491,I79556,I79785);
nand I_4534 (I79816,I79522,I262887);
nand I_4535 (I79833,I79816,I79751);
and I_4536 (I79850,I79816,I79833);
DFFARX1 I_4537  ( .D(I79850), .CLK(I2702), .RSTB(I79505), .Q(I79473) );
DFFARX1 I_4538  ( .D(I79816), .CLK(I2702), .RSTB(I79505), .Q(I79881) );
and I_4539 (I79470,I79649,I79881);
DFFARX1 I_4540  ( .D(I262893), .CLK(I2702), .RSTB(I79505), .Q(I79912) );
not I_4541 (I79929,I79912);
nor I_4542 (I79946,I79604,I79929);
and I_4543 (I79963,I79912,I79946);
nand I_4544 (I79485,I79912,I79666);
DFFARX1 I_4545  ( .D(I79912), .CLK(I2702), .RSTB(I79505), .Q(I79994) );
not I_4546 (I79482,I79994);
DFFARX1 I_4547  ( .D(I262890), .CLK(I2702), .RSTB(I79505), .Q(I80025) );
not I_4548 (I80042,I80025);
or I_4549 (I80059,I80042,I79963);
DFFARX1 I_4550  ( .D(I80059), .CLK(I2702), .RSTB(I79505), .Q(I79488) );
nand I_4551 (I79497,I80042,I79768);
DFFARX1 I_4552  ( .D(I80042), .CLK(I2702), .RSTB(I79505), .Q(I79467) );
not I_4553 (I80151,I2709);
not I_4554 (I80168,I547096);
nor I_4555 (I80185,I547072,I547078);
nand I_4556 (I80202,I80185,I547081);
DFFARX1 I_4557  ( .D(I80202), .CLK(I2702), .RSTB(I80151), .Q(I80125) );
nor I_4558 (I80233,I80168,I547072);
nand I_4559 (I80250,I80233,I547090);
not I_4560 (I80140,I80250);
DFFARX1 I_4561  ( .D(I80250), .CLK(I2702), .RSTB(I80151), .Q(I80122) );
not I_4562 (I80295,I547072);
not I_4563 (I80312,I80295);
not I_4564 (I80329,I547069);
nor I_4565 (I80346,I80329,I547084);
and I_4566 (I80363,I80346,I547075);
or I_4567 (I80380,I80363,I547087);
DFFARX1 I_4568  ( .D(I80380), .CLK(I2702), .RSTB(I80151), .Q(I80397) );
nor I_4569 (I80414,I80397,I80250);
nor I_4570 (I80431,I80397,I80312);
nand I_4571 (I80137,I80202,I80431);
nand I_4572 (I80462,I80168,I547069);
nand I_4573 (I80479,I80462,I80397);
and I_4574 (I80496,I80462,I80479);
DFFARX1 I_4575  ( .D(I80496), .CLK(I2702), .RSTB(I80151), .Q(I80119) );
DFFARX1 I_4576  ( .D(I80462), .CLK(I2702), .RSTB(I80151), .Q(I80527) );
and I_4577 (I80116,I80295,I80527);
DFFARX1 I_4578  ( .D(I547099), .CLK(I2702), .RSTB(I80151), .Q(I80558) );
not I_4579 (I80575,I80558);
nor I_4580 (I80592,I80250,I80575);
and I_4581 (I80609,I80558,I80592);
nand I_4582 (I80131,I80558,I80312);
DFFARX1 I_4583  ( .D(I80558), .CLK(I2702), .RSTB(I80151), .Q(I80640) );
not I_4584 (I80128,I80640);
DFFARX1 I_4585  ( .D(I547093), .CLK(I2702), .RSTB(I80151), .Q(I80671) );
not I_4586 (I80688,I80671);
or I_4587 (I80705,I80688,I80609);
DFFARX1 I_4588  ( .D(I80705), .CLK(I2702), .RSTB(I80151), .Q(I80134) );
nand I_4589 (I80143,I80688,I80414);
DFFARX1 I_4590  ( .D(I80688), .CLK(I2702), .RSTB(I80151), .Q(I80113) );
not I_4591 (I80797,I2709);
not I_4592 (I80814,I151497);
nor I_4593 (I80831,I151485,I151491);
nand I_4594 (I80848,I80831,I151500);
DFFARX1 I_4595  ( .D(I80848), .CLK(I2702), .RSTB(I80797), .Q(I80771) );
nor I_4596 (I80879,I80814,I151485);
nand I_4597 (I80896,I80879,I151488);
not I_4598 (I80786,I80896);
DFFARX1 I_4599  ( .D(I80896), .CLK(I2702), .RSTB(I80797), .Q(I80768) );
not I_4600 (I80941,I151485);
not I_4601 (I80958,I80941);
not I_4602 (I80975,I151509);
nor I_4603 (I80992,I80975,I151482);
and I_4604 (I81009,I80992,I151503);
or I_4605 (I81026,I81009,I151494);
DFFARX1 I_4606  ( .D(I81026), .CLK(I2702), .RSTB(I80797), .Q(I81043) );
nor I_4607 (I81060,I81043,I80896);
nor I_4608 (I81077,I81043,I80958);
nand I_4609 (I80783,I80848,I81077);
nand I_4610 (I81108,I80814,I151509);
nand I_4611 (I81125,I81108,I81043);
and I_4612 (I81142,I81108,I81125);
DFFARX1 I_4613  ( .D(I81142), .CLK(I2702), .RSTB(I80797), .Q(I80765) );
DFFARX1 I_4614  ( .D(I81108), .CLK(I2702), .RSTB(I80797), .Q(I81173) );
and I_4615 (I80762,I80941,I81173);
DFFARX1 I_4616  ( .D(I151479), .CLK(I2702), .RSTB(I80797), .Q(I81204) );
not I_4617 (I81221,I81204);
nor I_4618 (I81238,I80896,I81221);
and I_4619 (I81255,I81204,I81238);
nand I_4620 (I80777,I81204,I80958);
DFFARX1 I_4621  ( .D(I81204), .CLK(I2702), .RSTB(I80797), .Q(I81286) );
not I_4622 (I80774,I81286);
DFFARX1 I_4623  ( .D(I151506), .CLK(I2702), .RSTB(I80797), .Q(I81317) );
not I_4624 (I81334,I81317);
or I_4625 (I81351,I81334,I81255);
DFFARX1 I_4626  ( .D(I81351), .CLK(I2702), .RSTB(I80797), .Q(I80780) );
nand I_4627 (I80789,I81334,I81060);
DFFARX1 I_4628  ( .D(I81334), .CLK(I2702), .RSTB(I80797), .Q(I80759) );
not I_4629 (I81443,I2709);
not I_4630 (I81460,I433286);
nor I_4631 (I81477,I433274,I433280);
nand I_4632 (I81494,I81477,I433271);
DFFARX1 I_4633  ( .D(I81494), .CLK(I2702), .RSTB(I81443), .Q(I81417) );
nor I_4634 (I81525,I81460,I433274);
nand I_4635 (I81542,I81525,I433277);
not I_4636 (I81432,I81542);
DFFARX1 I_4637  ( .D(I81542), .CLK(I2702), .RSTB(I81443), .Q(I81414) );
not I_4638 (I81587,I433274);
not I_4639 (I81604,I81587);
not I_4640 (I81621,I433289);
nor I_4641 (I81638,I81621,I433301);
and I_4642 (I81655,I81638,I433283);
or I_4643 (I81672,I81655,I433298);
DFFARX1 I_4644  ( .D(I81672), .CLK(I2702), .RSTB(I81443), .Q(I81689) );
nor I_4645 (I81706,I81689,I81542);
nor I_4646 (I81723,I81689,I81604);
nand I_4647 (I81429,I81494,I81723);
nand I_4648 (I81754,I81460,I433289);
nand I_4649 (I81771,I81754,I81689);
and I_4650 (I81788,I81754,I81771);
DFFARX1 I_4651  ( .D(I81788), .CLK(I2702), .RSTB(I81443), .Q(I81411) );
DFFARX1 I_4652  ( .D(I81754), .CLK(I2702), .RSTB(I81443), .Q(I81819) );
and I_4653 (I81408,I81587,I81819);
DFFARX1 I_4654  ( .D(I433292), .CLK(I2702), .RSTB(I81443), .Q(I81850) );
not I_4655 (I81867,I81850);
nor I_4656 (I81884,I81542,I81867);
and I_4657 (I81901,I81850,I81884);
nand I_4658 (I81423,I81850,I81604);
DFFARX1 I_4659  ( .D(I81850), .CLK(I2702), .RSTB(I81443), .Q(I81932) );
not I_4660 (I81420,I81932);
DFFARX1 I_4661  ( .D(I433295), .CLK(I2702), .RSTB(I81443), .Q(I81963) );
not I_4662 (I81980,I81963);
or I_4663 (I81997,I81980,I81901);
DFFARX1 I_4664  ( .D(I81997), .CLK(I2702), .RSTB(I81443), .Q(I81426) );
nand I_4665 (I81435,I81980,I81706);
DFFARX1 I_4666  ( .D(I81980), .CLK(I2702), .RSTB(I81443), .Q(I81405) );
not I_4667 (I82089,I2709);
not I_4668 (I82106,I280782);
nor I_4669 (I82123,I280779,I280767);
nand I_4670 (I82140,I82123,I280770);
DFFARX1 I_4671  ( .D(I82140), .CLK(I2702), .RSTB(I82089), .Q(I82063) );
nor I_4672 (I82171,I82106,I280779);
nand I_4673 (I82188,I82171,I280776);
not I_4674 (I82078,I82188);
DFFARX1 I_4675  ( .D(I82188), .CLK(I2702), .RSTB(I82089), .Q(I82060) );
not I_4676 (I82233,I280779);
not I_4677 (I82250,I82233);
not I_4678 (I82267,I280788);
nor I_4679 (I82284,I82267,I280764);
and I_4680 (I82301,I82284,I280785);
or I_4681 (I82318,I82301,I280773);
DFFARX1 I_4682  ( .D(I82318), .CLK(I2702), .RSTB(I82089), .Q(I82335) );
nor I_4683 (I82352,I82335,I82188);
nor I_4684 (I82369,I82335,I82250);
nand I_4685 (I82075,I82140,I82369);
nand I_4686 (I82400,I82106,I280788);
nand I_4687 (I82417,I82400,I82335);
and I_4688 (I82434,I82400,I82417);
DFFARX1 I_4689  ( .D(I82434), .CLK(I2702), .RSTB(I82089), .Q(I82057) );
DFFARX1 I_4690  ( .D(I82400), .CLK(I2702), .RSTB(I82089), .Q(I82465) );
and I_4691 (I82054,I82233,I82465);
DFFARX1 I_4692  ( .D(I280794), .CLK(I2702), .RSTB(I82089), .Q(I82496) );
not I_4693 (I82513,I82496);
nor I_4694 (I82530,I82188,I82513);
and I_4695 (I82547,I82496,I82530);
nand I_4696 (I82069,I82496,I82250);
DFFARX1 I_4697  ( .D(I82496), .CLK(I2702), .RSTB(I82089), .Q(I82578) );
not I_4698 (I82066,I82578);
DFFARX1 I_4699  ( .D(I280791), .CLK(I2702), .RSTB(I82089), .Q(I82609) );
not I_4700 (I82626,I82609);
or I_4701 (I82643,I82626,I82547);
DFFARX1 I_4702  ( .D(I82643), .CLK(I2702), .RSTB(I82089), .Q(I82072) );
nand I_4703 (I82081,I82626,I82352);
DFFARX1 I_4704  ( .D(I82626), .CLK(I2702), .RSTB(I82089), .Q(I82051) );
not I_4705 (I82735,I2709);
not I_4706 (I82752,I352539);
nor I_4707 (I82769,I352551,I352533);
nand I_4708 (I82786,I82769,I352548);
DFFARX1 I_4709  ( .D(I82786), .CLK(I2702), .RSTB(I82735), .Q(I82709) );
nor I_4710 (I82817,I82752,I352551);
nand I_4711 (I82834,I82817,I352536);
not I_4712 (I82724,I82834);
DFFARX1 I_4713  ( .D(I82834), .CLK(I2702), .RSTB(I82735), .Q(I82706) );
not I_4714 (I82879,I352551);
not I_4715 (I82896,I82879);
not I_4716 (I82913,I352545);
nor I_4717 (I82930,I82913,I352524);
and I_4718 (I82947,I82930,I352527);
or I_4719 (I82964,I82947,I352530);
DFFARX1 I_4720  ( .D(I82964), .CLK(I2702), .RSTB(I82735), .Q(I82981) );
nor I_4721 (I82998,I82981,I82834);
nor I_4722 (I83015,I82981,I82896);
nand I_4723 (I82721,I82786,I83015);
nand I_4724 (I83046,I82752,I352545);
nand I_4725 (I83063,I83046,I82981);
and I_4726 (I83080,I83046,I83063);
DFFARX1 I_4727  ( .D(I83080), .CLK(I2702), .RSTB(I82735), .Q(I82703) );
DFFARX1 I_4728  ( .D(I83046), .CLK(I2702), .RSTB(I82735), .Q(I83111) );
and I_4729 (I82700,I82879,I83111);
DFFARX1 I_4730  ( .D(I352521), .CLK(I2702), .RSTB(I82735), .Q(I83142) );
not I_4731 (I83159,I83142);
nor I_4732 (I83176,I82834,I83159);
and I_4733 (I83193,I83142,I83176);
nand I_4734 (I82715,I83142,I82896);
DFFARX1 I_4735  ( .D(I83142), .CLK(I2702), .RSTB(I82735), .Q(I83224) );
not I_4736 (I82712,I83224);
DFFARX1 I_4737  ( .D(I352542), .CLK(I2702), .RSTB(I82735), .Q(I83255) );
not I_4738 (I83272,I83255);
or I_4739 (I83289,I83272,I83193);
DFFARX1 I_4740  ( .D(I83289), .CLK(I2702), .RSTB(I82735), .Q(I82718) );
nand I_4741 (I82727,I83272,I82998);
DFFARX1 I_4742  ( .D(I83272), .CLK(I2702), .RSTB(I82735), .Q(I82697) );
not I_4743 (I83381,I2709);
not I_4744 (I83398,I148845);
nor I_4745 (I83415,I148833,I148839);
nand I_4746 (I83432,I83415,I148848);
DFFARX1 I_4747  ( .D(I83432), .CLK(I2702), .RSTB(I83381), .Q(I83355) );
nor I_4748 (I83463,I83398,I148833);
nand I_4749 (I83480,I83463,I148836);
not I_4750 (I83370,I83480);
DFFARX1 I_4751  ( .D(I83480), .CLK(I2702), .RSTB(I83381), .Q(I83352) );
not I_4752 (I83525,I148833);
not I_4753 (I83542,I83525);
not I_4754 (I83559,I148857);
nor I_4755 (I83576,I83559,I148830);
and I_4756 (I83593,I83576,I148851);
or I_4757 (I83610,I83593,I148842);
DFFARX1 I_4758  ( .D(I83610), .CLK(I2702), .RSTB(I83381), .Q(I83627) );
nor I_4759 (I83644,I83627,I83480);
nor I_4760 (I83661,I83627,I83542);
nand I_4761 (I83367,I83432,I83661);
nand I_4762 (I83692,I83398,I148857);
nand I_4763 (I83709,I83692,I83627);
and I_4764 (I83726,I83692,I83709);
DFFARX1 I_4765  ( .D(I83726), .CLK(I2702), .RSTB(I83381), .Q(I83349) );
DFFARX1 I_4766  ( .D(I83692), .CLK(I2702), .RSTB(I83381), .Q(I83757) );
and I_4767 (I83346,I83525,I83757);
DFFARX1 I_4768  ( .D(I148827), .CLK(I2702), .RSTB(I83381), .Q(I83788) );
not I_4769 (I83805,I83788);
nor I_4770 (I83822,I83480,I83805);
and I_4771 (I83839,I83788,I83822);
nand I_4772 (I83361,I83788,I83542);
DFFARX1 I_4773  ( .D(I83788), .CLK(I2702), .RSTB(I83381), .Q(I83870) );
not I_4774 (I83358,I83870);
DFFARX1 I_4775  ( .D(I148854), .CLK(I2702), .RSTB(I83381), .Q(I83901) );
not I_4776 (I83918,I83901);
or I_4777 (I83935,I83918,I83839);
DFFARX1 I_4778  ( .D(I83935), .CLK(I2702), .RSTB(I83381), .Q(I83364) );
nand I_4779 (I83373,I83918,I83644);
DFFARX1 I_4780  ( .D(I83918), .CLK(I2702), .RSTB(I83381), .Q(I83343) );
not I_4781 (I84027,I2709);
not I_4782 (I84044,I1495);
nor I_4783 (I84061,I2127,I1607);
nand I_4784 (I84078,I84061,I1615);
DFFARX1 I_4785  ( .D(I84078), .CLK(I2702), .RSTB(I84027), .Q(I84001) );
nor I_4786 (I84109,I84044,I2127);
nand I_4787 (I84126,I84109,I1855);
not I_4788 (I84016,I84126);
DFFARX1 I_4789  ( .D(I84126), .CLK(I2702), .RSTB(I84027), .Q(I83998) );
not I_4790 (I84171,I2127);
not I_4791 (I84188,I84171);
not I_4792 (I84205,I2287);
nor I_4793 (I84222,I84205,I1255);
and I_4794 (I84239,I84222,I2079);
or I_4795 (I84256,I84239,I1599);
DFFARX1 I_4796  ( .D(I84256), .CLK(I2702), .RSTB(I84027), .Q(I84273) );
nor I_4797 (I84290,I84273,I84126);
nor I_4798 (I84307,I84273,I84188);
nand I_4799 (I84013,I84078,I84307);
nand I_4800 (I84338,I84044,I2287);
nand I_4801 (I84355,I84338,I84273);
and I_4802 (I84372,I84338,I84355);
DFFARX1 I_4803  ( .D(I84372), .CLK(I2702), .RSTB(I84027), .Q(I83995) );
DFFARX1 I_4804  ( .D(I84338), .CLK(I2702), .RSTB(I84027), .Q(I84403) );
and I_4805 (I83992,I84171,I84403);
DFFARX1 I_4806  ( .D(I2231), .CLK(I2702), .RSTB(I84027), .Q(I84434) );
not I_4807 (I84451,I84434);
nor I_4808 (I84468,I84126,I84451);
and I_4809 (I84485,I84434,I84468);
nand I_4810 (I84007,I84434,I84188);
DFFARX1 I_4811  ( .D(I84434), .CLK(I2702), .RSTB(I84027), .Q(I84516) );
not I_4812 (I84004,I84516);
DFFARX1 I_4813  ( .D(I2415), .CLK(I2702), .RSTB(I84027), .Q(I84547) );
not I_4814 (I84564,I84547);
or I_4815 (I84581,I84564,I84485);
DFFARX1 I_4816  ( .D(I84581), .CLK(I2702), .RSTB(I84027), .Q(I84010) );
nand I_4817 (I84019,I84564,I84290);
DFFARX1 I_4818  ( .D(I84564), .CLK(I2702), .RSTB(I84027), .Q(I83989) );
not I_4819 (I84673,I2709);
not I_4820 (I84690,I608964);
nor I_4821 (I84707,I608949,I608976);
nand I_4822 (I84724,I84707,I608952);
DFFARX1 I_4823  ( .D(I84724), .CLK(I2702), .RSTB(I84673), .Q(I84647) );
nor I_4824 (I84755,I84690,I608949);
nand I_4825 (I84772,I84755,I608967);
not I_4826 (I84662,I84772);
DFFARX1 I_4827  ( .D(I84772), .CLK(I2702), .RSTB(I84673), .Q(I84644) );
not I_4828 (I84817,I608949);
not I_4829 (I84834,I84817);
not I_4830 (I84851,I608979);
nor I_4831 (I84868,I84851,I608961);
and I_4832 (I84885,I84868,I608970);
or I_4833 (I84902,I84885,I608955);
DFFARX1 I_4834  ( .D(I84902), .CLK(I2702), .RSTB(I84673), .Q(I84919) );
nor I_4835 (I84936,I84919,I84772);
nor I_4836 (I84953,I84919,I84834);
nand I_4837 (I84659,I84724,I84953);
nand I_4838 (I84984,I84690,I608979);
nand I_4839 (I85001,I84984,I84919);
and I_4840 (I85018,I84984,I85001);
DFFARX1 I_4841  ( .D(I85018), .CLK(I2702), .RSTB(I84673), .Q(I84641) );
DFFARX1 I_4842  ( .D(I84984), .CLK(I2702), .RSTB(I84673), .Q(I85049) );
and I_4843 (I84638,I84817,I85049);
DFFARX1 I_4844  ( .D(I608958), .CLK(I2702), .RSTB(I84673), .Q(I85080) );
not I_4845 (I85097,I85080);
nor I_4846 (I85114,I84772,I85097);
and I_4847 (I85131,I85080,I85114);
nand I_4848 (I84653,I85080,I84834);
DFFARX1 I_4849  ( .D(I85080), .CLK(I2702), .RSTB(I84673), .Q(I85162) );
not I_4850 (I84650,I85162);
DFFARX1 I_4851  ( .D(I608973), .CLK(I2702), .RSTB(I84673), .Q(I85193) );
not I_4852 (I85210,I85193);
or I_4853 (I85227,I85210,I85131);
DFFARX1 I_4854  ( .D(I85227), .CLK(I2702), .RSTB(I84673), .Q(I84656) );
nand I_4855 (I84665,I85210,I84936);
DFFARX1 I_4856  ( .D(I85210), .CLK(I2702), .RSTB(I84673), .Q(I84635) );
not I_4857 (I85319,I2709);
not I_4858 (I85336,I689155);
nor I_4859 (I85353,I689170,I689185);
nand I_4860 (I85370,I85353,I689173);
DFFARX1 I_4861  ( .D(I85370), .CLK(I2702), .RSTB(I85319), .Q(I85293) );
nor I_4862 (I85401,I85336,I689170);
nand I_4863 (I85418,I85401,I689176);
not I_4864 (I85308,I85418);
DFFARX1 I_4865  ( .D(I85418), .CLK(I2702), .RSTB(I85319), .Q(I85290) );
not I_4866 (I85463,I689170);
not I_4867 (I85480,I85463);
not I_4868 (I85497,I689182);
nor I_4869 (I85514,I85497,I689179);
and I_4870 (I85531,I85514,I689158);
or I_4871 (I85548,I85531,I689167);
DFFARX1 I_4872  ( .D(I85548), .CLK(I2702), .RSTB(I85319), .Q(I85565) );
nor I_4873 (I85582,I85565,I85418);
nor I_4874 (I85599,I85565,I85480);
nand I_4875 (I85305,I85370,I85599);
nand I_4876 (I85630,I85336,I689182);
nand I_4877 (I85647,I85630,I85565);
and I_4878 (I85664,I85630,I85647);
DFFARX1 I_4879  ( .D(I85664), .CLK(I2702), .RSTB(I85319), .Q(I85287) );
DFFARX1 I_4880  ( .D(I85630), .CLK(I2702), .RSTB(I85319), .Q(I85695) );
and I_4881 (I85284,I85463,I85695);
DFFARX1 I_4882  ( .D(I689164), .CLK(I2702), .RSTB(I85319), .Q(I85726) );
not I_4883 (I85743,I85726);
nor I_4884 (I85760,I85418,I85743);
and I_4885 (I85777,I85726,I85760);
nand I_4886 (I85299,I85726,I85480);
DFFARX1 I_4887  ( .D(I85726), .CLK(I2702), .RSTB(I85319), .Q(I85808) );
not I_4888 (I85296,I85808);
DFFARX1 I_4889  ( .D(I689161), .CLK(I2702), .RSTB(I85319), .Q(I85839) );
not I_4890 (I85856,I85839);
or I_4891 (I85873,I85856,I85777);
DFFARX1 I_4892  ( .D(I85873), .CLK(I2702), .RSTB(I85319), .Q(I85302) );
nand I_4893 (I85311,I85856,I85582);
DFFARX1 I_4894  ( .D(I85856), .CLK(I2702), .RSTB(I85319), .Q(I85281) );
not I_4895 (I85965,I2709);
not I_4896 (I85982,I664624);
nor I_4897 (I85999,I664639,I664654);
nand I_4898 (I86016,I85999,I664642);
DFFARX1 I_4899  ( .D(I86016), .CLK(I2702), .RSTB(I85965), .Q(I85939) );
nor I_4900 (I86047,I85982,I664639);
nand I_4901 (I86064,I86047,I664645);
not I_4902 (I85954,I86064);
DFFARX1 I_4903  ( .D(I86064), .CLK(I2702), .RSTB(I85965), .Q(I85936) );
not I_4904 (I86109,I664639);
not I_4905 (I86126,I86109);
not I_4906 (I86143,I664651);
nor I_4907 (I86160,I86143,I664648);
and I_4908 (I86177,I86160,I664627);
or I_4909 (I86194,I86177,I664636);
DFFARX1 I_4910  ( .D(I86194), .CLK(I2702), .RSTB(I85965), .Q(I86211) );
nor I_4911 (I86228,I86211,I86064);
nor I_4912 (I86245,I86211,I86126);
nand I_4913 (I85951,I86016,I86245);
nand I_4914 (I86276,I85982,I664651);
nand I_4915 (I86293,I86276,I86211);
and I_4916 (I86310,I86276,I86293);
DFFARX1 I_4917  ( .D(I86310), .CLK(I2702), .RSTB(I85965), .Q(I85933) );
DFFARX1 I_4918  ( .D(I86276), .CLK(I2702), .RSTB(I85965), .Q(I86341) );
and I_4919 (I85930,I86109,I86341);
DFFARX1 I_4920  ( .D(I664633), .CLK(I2702), .RSTB(I85965), .Q(I86372) );
not I_4921 (I86389,I86372);
nor I_4922 (I86406,I86064,I86389);
and I_4923 (I86423,I86372,I86406);
nand I_4924 (I85945,I86372,I86126);
DFFARX1 I_4925  ( .D(I86372), .CLK(I2702), .RSTB(I85965), .Q(I86454) );
not I_4926 (I85942,I86454);
DFFARX1 I_4927  ( .D(I664630), .CLK(I2702), .RSTB(I85965), .Q(I86485) );
not I_4928 (I86502,I86485);
or I_4929 (I86519,I86502,I86423);
DFFARX1 I_4930  ( .D(I86519), .CLK(I2702), .RSTB(I85965), .Q(I85948) );
nand I_4931 (I85957,I86502,I86228);
DFFARX1 I_4932  ( .D(I86502), .CLK(I2702), .RSTB(I85965), .Q(I85927) );
not I_4933 (I86611,I2709);
not I_4934 (I86628,I602419);
nor I_4935 (I86645,I602404,I602431);
nand I_4936 (I86662,I86645,I602407);
DFFARX1 I_4937  ( .D(I86662), .CLK(I2702), .RSTB(I86611), .Q(I86585) );
nor I_4938 (I86693,I86628,I602404);
nand I_4939 (I86710,I86693,I602422);
not I_4940 (I86600,I86710);
DFFARX1 I_4941  ( .D(I86710), .CLK(I2702), .RSTB(I86611), .Q(I86582) );
not I_4942 (I86755,I602404);
not I_4943 (I86772,I86755);
not I_4944 (I86789,I602434);
nor I_4945 (I86806,I86789,I602416);
and I_4946 (I86823,I86806,I602425);
or I_4947 (I86840,I86823,I602410);
DFFARX1 I_4948  ( .D(I86840), .CLK(I2702), .RSTB(I86611), .Q(I86857) );
nor I_4949 (I86874,I86857,I86710);
nor I_4950 (I86891,I86857,I86772);
nand I_4951 (I86597,I86662,I86891);
nand I_4952 (I86922,I86628,I602434);
nand I_4953 (I86939,I86922,I86857);
and I_4954 (I86956,I86922,I86939);
DFFARX1 I_4955  ( .D(I86956), .CLK(I2702), .RSTB(I86611), .Q(I86579) );
DFFARX1 I_4956  ( .D(I86922), .CLK(I2702), .RSTB(I86611), .Q(I86987) );
and I_4957 (I86576,I86755,I86987);
DFFARX1 I_4958  ( .D(I602413), .CLK(I2702), .RSTB(I86611), .Q(I87018) );
not I_4959 (I87035,I87018);
nor I_4960 (I87052,I86710,I87035);
and I_4961 (I87069,I87018,I87052);
nand I_4962 (I86591,I87018,I86772);
DFFARX1 I_4963  ( .D(I87018), .CLK(I2702), .RSTB(I86611), .Q(I87100) );
not I_4964 (I86588,I87100);
DFFARX1 I_4965  ( .D(I602428), .CLK(I2702), .RSTB(I86611), .Q(I87131) );
not I_4966 (I87148,I87131);
or I_4967 (I87165,I87148,I87069);
DFFARX1 I_4968  ( .D(I87165), .CLK(I2702), .RSTB(I86611), .Q(I86594) );
nand I_4969 (I86603,I87148,I86874);
DFFARX1 I_4970  ( .D(I87148), .CLK(I2702), .RSTB(I86611), .Q(I86573) );
not I_4971 (I87257,I2709);
not I_4972 (I87274,I388069);
nor I_4973 (I87291,I388081,I388063);
nand I_4974 (I87308,I87291,I388078);
DFFARX1 I_4975  ( .D(I87308), .CLK(I2702), .RSTB(I87257), .Q(I87231) );
nor I_4976 (I87339,I87274,I388081);
nand I_4977 (I87356,I87339,I388066);
not I_4978 (I87246,I87356);
DFFARX1 I_4979  ( .D(I87356), .CLK(I2702), .RSTB(I87257), .Q(I87228) );
not I_4980 (I87401,I388081);
not I_4981 (I87418,I87401);
not I_4982 (I87435,I388075);
nor I_4983 (I87452,I87435,I388054);
and I_4984 (I87469,I87452,I388057);
or I_4985 (I87486,I87469,I388060);
DFFARX1 I_4986  ( .D(I87486), .CLK(I2702), .RSTB(I87257), .Q(I87503) );
nor I_4987 (I87520,I87503,I87356);
nor I_4988 (I87537,I87503,I87418);
nand I_4989 (I87243,I87308,I87537);
nand I_4990 (I87568,I87274,I388075);
nand I_4991 (I87585,I87568,I87503);
and I_4992 (I87602,I87568,I87585);
DFFARX1 I_4993  ( .D(I87602), .CLK(I2702), .RSTB(I87257), .Q(I87225) );
DFFARX1 I_4994  ( .D(I87568), .CLK(I2702), .RSTB(I87257), .Q(I87633) );
and I_4995 (I87222,I87401,I87633);
DFFARX1 I_4996  ( .D(I388051), .CLK(I2702), .RSTB(I87257), .Q(I87664) );
not I_4997 (I87681,I87664);
nor I_4998 (I87698,I87356,I87681);
and I_4999 (I87715,I87664,I87698);
nand I_5000 (I87237,I87664,I87418);
DFFARX1 I_5001  ( .D(I87664), .CLK(I2702), .RSTB(I87257), .Q(I87746) );
not I_5002 (I87234,I87746);
DFFARX1 I_5003  ( .D(I388072), .CLK(I2702), .RSTB(I87257), .Q(I87777) );
not I_5004 (I87794,I87777);
or I_5005 (I87811,I87794,I87715);
DFFARX1 I_5006  ( .D(I87811), .CLK(I2702), .RSTB(I87257), .Q(I87240) );
nand I_5007 (I87249,I87794,I87520);
DFFARX1 I_5008  ( .D(I87794), .CLK(I2702), .RSTB(I87257), .Q(I87219) );
not I_5009 (I87903,I2709);
not I_5010 (I87920,I247632);
nor I_5011 (I87937,I247629,I247617);
nand I_5012 (I87954,I87937,I247620);
DFFARX1 I_5013  ( .D(I87954), .CLK(I2702), .RSTB(I87903), .Q(I87877) );
nor I_5014 (I87985,I87920,I247629);
nand I_5015 (I88002,I87985,I247626);
not I_5016 (I87892,I88002);
DFFARX1 I_5017  ( .D(I88002), .CLK(I2702), .RSTB(I87903), .Q(I87874) );
not I_5018 (I88047,I247629);
not I_5019 (I88064,I88047);
not I_5020 (I88081,I247638);
nor I_5021 (I88098,I88081,I247614);
and I_5022 (I88115,I88098,I247635);
or I_5023 (I88132,I88115,I247623);
DFFARX1 I_5024  ( .D(I88132), .CLK(I2702), .RSTB(I87903), .Q(I88149) );
nor I_5025 (I88166,I88149,I88002);
nor I_5026 (I88183,I88149,I88064);
nand I_5027 (I87889,I87954,I88183);
nand I_5028 (I88214,I87920,I247638);
nand I_5029 (I88231,I88214,I88149);
and I_5030 (I88248,I88214,I88231);
DFFARX1 I_5031  ( .D(I88248), .CLK(I2702), .RSTB(I87903), .Q(I87871) );
DFFARX1 I_5032  ( .D(I88214), .CLK(I2702), .RSTB(I87903), .Q(I88279) );
and I_5033 (I87868,I88047,I88279);
DFFARX1 I_5034  ( .D(I247644), .CLK(I2702), .RSTB(I87903), .Q(I88310) );
not I_5035 (I88327,I88310);
nor I_5036 (I88344,I88002,I88327);
and I_5037 (I88361,I88310,I88344);
nand I_5038 (I87883,I88310,I88064);
DFFARX1 I_5039  ( .D(I88310), .CLK(I2702), .RSTB(I87903), .Q(I88392) );
not I_5040 (I87880,I88392);
DFFARX1 I_5041  ( .D(I247641), .CLK(I2702), .RSTB(I87903), .Q(I88423) );
not I_5042 (I88440,I88423);
or I_5043 (I88457,I88440,I88361);
DFFARX1 I_5044  ( .D(I88457), .CLK(I2702), .RSTB(I87903), .Q(I87886) );
nand I_5045 (I87895,I88440,I88166);
DFFARX1 I_5046  ( .D(I88440), .CLK(I2702), .RSTB(I87903), .Q(I87865) );
not I_5047 (I88549,I2709);
not I_5048 (I88566,I410033);
nor I_5049 (I88583,I410045,I410027);
nand I_5050 (I88600,I88583,I410042);
DFFARX1 I_5051  ( .D(I88600), .CLK(I2702), .RSTB(I88549), .Q(I88523) );
nor I_5052 (I88631,I88566,I410045);
nand I_5053 (I88648,I88631,I410030);
not I_5054 (I88538,I88648);
DFFARX1 I_5055  ( .D(I88648), .CLK(I2702), .RSTB(I88549), .Q(I88520) );
not I_5056 (I88693,I410045);
not I_5057 (I88710,I88693);
not I_5058 (I88727,I410039);
nor I_5059 (I88744,I88727,I410018);
and I_5060 (I88761,I88744,I410021);
or I_5061 (I88778,I88761,I410024);
DFFARX1 I_5062  ( .D(I88778), .CLK(I2702), .RSTB(I88549), .Q(I88795) );
nor I_5063 (I88812,I88795,I88648);
nor I_5064 (I88829,I88795,I88710);
nand I_5065 (I88535,I88600,I88829);
nand I_5066 (I88860,I88566,I410039);
nand I_5067 (I88877,I88860,I88795);
and I_5068 (I88894,I88860,I88877);
DFFARX1 I_5069  ( .D(I88894), .CLK(I2702), .RSTB(I88549), .Q(I88517) );
DFFARX1 I_5070  ( .D(I88860), .CLK(I2702), .RSTB(I88549), .Q(I88925) );
and I_5071 (I88514,I88693,I88925);
DFFARX1 I_5072  ( .D(I410015), .CLK(I2702), .RSTB(I88549), .Q(I88956) );
not I_5073 (I88973,I88956);
nor I_5074 (I88990,I88648,I88973);
and I_5075 (I89007,I88956,I88990);
nand I_5076 (I88529,I88956,I88710);
DFFARX1 I_5077  ( .D(I88956), .CLK(I2702), .RSTB(I88549), .Q(I89038) );
not I_5078 (I88526,I89038);
DFFARX1 I_5079  ( .D(I410036), .CLK(I2702), .RSTB(I88549), .Q(I89069) );
not I_5080 (I89086,I89069);
or I_5081 (I89103,I89086,I89007);
DFFARX1 I_5082  ( .D(I89103), .CLK(I2702), .RSTB(I88549), .Q(I88532) );
nand I_5083 (I88541,I89086,I88812);
DFFARX1 I_5084  ( .D(I89086), .CLK(I2702), .RSTB(I88549), .Q(I88511) );
not I_5085 (I89195,I2709);
not I_5086 (I89212,I478370);
nor I_5087 (I89229,I478358,I478364);
nand I_5088 (I89246,I89229,I478355);
DFFARX1 I_5089  ( .D(I89246), .CLK(I2702), .RSTB(I89195), .Q(I89169) );
nor I_5090 (I89277,I89212,I478358);
nand I_5091 (I89294,I89277,I478361);
not I_5092 (I89184,I89294);
DFFARX1 I_5093  ( .D(I89294), .CLK(I2702), .RSTB(I89195), .Q(I89166) );
not I_5094 (I89339,I478358);
not I_5095 (I89356,I89339);
not I_5096 (I89373,I478373);
nor I_5097 (I89390,I89373,I478385);
and I_5098 (I89407,I89390,I478367);
or I_5099 (I89424,I89407,I478382);
DFFARX1 I_5100  ( .D(I89424), .CLK(I2702), .RSTB(I89195), .Q(I89441) );
nor I_5101 (I89458,I89441,I89294);
nor I_5102 (I89475,I89441,I89356);
nand I_5103 (I89181,I89246,I89475);
nand I_5104 (I89506,I89212,I478373);
nand I_5105 (I89523,I89506,I89441);
and I_5106 (I89540,I89506,I89523);
DFFARX1 I_5107  ( .D(I89540), .CLK(I2702), .RSTB(I89195), .Q(I89163) );
DFFARX1 I_5108  ( .D(I89506), .CLK(I2702), .RSTB(I89195), .Q(I89571) );
and I_5109 (I89160,I89339,I89571);
DFFARX1 I_5110  ( .D(I478376), .CLK(I2702), .RSTB(I89195), .Q(I89602) );
not I_5111 (I89619,I89602);
nor I_5112 (I89636,I89294,I89619);
and I_5113 (I89653,I89602,I89636);
nand I_5114 (I89175,I89602,I89356);
DFFARX1 I_5115  ( .D(I89602), .CLK(I2702), .RSTB(I89195), .Q(I89684) );
not I_5116 (I89172,I89684);
DFFARX1 I_5117  ( .D(I478379), .CLK(I2702), .RSTB(I89195), .Q(I89715) );
not I_5118 (I89732,I89715);
or I_5119 (I89749,I89732,I89653);
DFFARX1 I_5120  ( .D(I89749), .CLK(I2702), .RSTB(I89195), .Q(I89178) );
nand I_5121 (I89187,I89732,I89458);
DFFARX1 I_5122  ( .D(I89732), .CLK(I2702), .RSTB(I89195), .Q(I89157) );
not I_5123 (I89841,I2709);
not I_5124 (I89858,I139563);
nor I_5125 (I89875,I139551,I139557);
nand I_5126 (I89892,I89875,I139566);
DFFARX1 I_5127  ( .D(I89892), .CLK(I2702), .RSTB(I89841), .Q(I89815) );
nor I_5128 (I89923,I89858,I139551);
nand I_5129 (I89940,I89923,I139554);
not I_5130 (I89830,I89940);
DFFARX1 I_5131  ( .D(I89940), .CLK(I2702), .RSTB(I89841), .Q(I89812) );
not I_5132 (I89985,I139551);
not I_5133 (I90002,I89985);
not I_5134 (I90019,I139575);
nor I_5135 (I90036,I90019,I139548);
and I_5136 (I90053,I90036,I139569);
or I_5137 (I90070,I90053,I139560);
DFFARX1 I_5138  ( .D(I90070), .CLK(I2702), .RSTB(I89841), .Q(I90087) );
nor I_5139 (I90104,I90087,I89940);
nor I_5140 (I90121,I90087,I90002);
nand I_5141 (I89827,I89892,I90121);
nand I_5142 (I90152,I89858,I139575);
nand I_5143 (I90169,I90152,I90087);
and I_5144 (I90186,I90152,I90169);
DFFARX1 I_5145  ( .D(I90186), .CLK(I2702), .RSTB(I89841), .Q(I89809) );
DFFARX1 I_5146  ( .D(I90152), .CLK(I2702), .RSTB(I89841), .Q(I90217) );
and I_5147 (I89806,I89985,I90217);
DFFARX1 I_5148  ( .D(I139545), .CLK(I2702), .RSTB(I89841), .Q(I90248) );
not I_5149 (I90265,I90248);
nor I_5150 (I90282,I89940,I90265);
and I_5151 (I90299,I90248,I90282);
nand I_5152 (I89821,I90248,I90002);
DFFARX1 I_5153  ( .D(I90248), .CLK(I2702), .RSTB(I89841), .Q(I90330) );
not I_5154 (I89818,I90330);
DFFARX1 I_5155  ( .D(I139572), .CLK(I2702), .RSTB(I89841), .Q(I90361) );
not I_5156 (I90378,I90361);
or I_5157 (I90395,I90378,I90299);
DFFARX1 I_5158  ( .D(I90395), .CLK(I2702), .RSTB(I89841), .Q(I89824) );
nand I_5159 (I89833,I90378,I90104);
DFFARX1 I_5160  ( .D(I90378), .CLK(I2702), .RSTB(I89841), .Q(I89803) );
not I_5161 (I90487,I2709);
not I_5162 (I90504,I570301);
nor I_5163 (I90521,I570277,I570283);
nand I_5164 (I90538,I90521,I570286);
DFFARX1 I_5165  ( .D(I90538), .CLK(I2702), .RSTB(I90487), .Q(I90461) );
nor I_5166 (I90569,I90504,I570277);
nand I_5167 (I90586,I90569,I570295);
not I_5168 (I90476,I90586);
DFFARX1 I_5169  ( .D(I90586), .CLK(I2702), .RSTB(I90487), .Q(I90458) );
not I_5170 (I90631,I570277);
not I_5171 (I90648,I90631);
not I_5172 (I90665,I570274);
nor I_5173 (I90682,I90665,I570289);
and I_5174 (I90699,I90682,I570280);
or I_5175 (I90716,I90699,I570292);
DFFARX1 I_5176  ( .D(I90716), .CLK(I2702), .RSTB(I90487), .Q(I90733) );
nor I_5177 (I90750,I90733,I90586);
nor I_5178 (I90767,I90733,I90648);
nand I_5179 (I90473,I90538,I90767);
nand I_5180 (I90798,I90504,I570274);
nand I_5181 (I90815,I90798,I90733);
and I_5182 (I90832,I90798,I90815);
DFFARX1 I_5183  ( .D(I90832), .CLK(I2702), .RSTB(I90487), .Q(I90455) );
DFFARX1 I_5184  ( .D(I90798), .CLK(I2702), .RSTB(I90487), .Q(I90863) );
and I_5185 (I90452,I90631,I90863);
DFFARX1 I_5186  ( .D(I570304), .CLK(I2702), .RSTB(I90487), .Q(I90894) );
not I_5187 (I90911,I90894);
nor I_5188 (I90928,I90586,I90911);
and I_5189 (I90945,I90894,I90928);
nand I_5190 (I90467,I90894,I90648);
DFFARX1 I_5191  ( .D(I90894), .CLK(I2702), .RSTB(I90487), .Q(I90976) );
not I_5192 (I90464,I90976);
DFFARX1 I_5193  ( .D(I570298), .CLK(I2702), .RSTB(I90487), .Q(I91007) );
not I_5194 (I91024,I91007);
or I_5195 (I91041,I91024,I90945);
DFFARX1 I_5196  ( .D(I91041), .CLK(I2702), .RSTB(I90487), .Q(I90470) );
nand I_5197 (I90479,I91024,I90750);
DFFARX1 I_5198  ( .D(I91024), .CLK(I2702), .RSTB(I90487), .Q(I90449) );
not I_5199 (I91133,I2709);
not I_5200 (I91150,I703665);
nor I_5201 (I91167,I703662,I703659);
nand I_5202 (I91184,I91167,I703680);
DFFARX1 I_5203  ( .D(I91184), .CLK(I2702), .RSTB(I91133), .Q(I91107) );
nor I_5204 (I91215,I91150,I703662);
nand I_5205 (I91232,I91215,I703683);
not I_5206 (I91122,I91232);
DFFARX1 I_5207  ( .D(I91232), .CLK(I2702), .RSTB(I91133), .Q(I91104) );
not I_5208 (I91277,I703662);
not I_5209 (I91294,I91277);
not I_5210 (I91311,I703656);
nor I_5211 (I91328,I91311,I703668);
and I_5212 (I91345,I91328,I703677);
or I_5213 (I91362,I91345,I703671);
DFFARX1 I_5214  ( .D(I91362), .CLK(I2702), .RSTB(I91133), .Q(I91379) );
nor I_5215 (I91396,I91379,I91232);
nor I_5216 (I91413,I91379,I91294);
nand I_5217 (I91119,I91184,I91413);
nand I_5218 (I91444,I91150,I703656);
nand I_5219 (I91461,I91444,I91379);
and I_5220 (I91478,I91444,I91461);
DFFARX1 I_5221  ( .D(I91478), .CLK(I2702), .RSTB(I91133), .Q(I91101) );
DFFARX1 I_5222  ( .D(I91444), .CLK(I2702), .RSTB(I91133), .Q(I91509) );
and I_5223 (I91098,I91277,I91509);
DFFARX1 I_5224  ( .D(I703686), .CLK(I2702), .RSTB(I91133), .Q(I91540) );
not I_5225 (I91557,I91540);
nor I_5226 (I91574,I91232,I91557);
and I_5227 (I91591,I91540,I91574);
nand I_5228 (I91113,I91540,I91294);
DFFARX1 I_5229  ( .D(I91540), .CLK(I2702), .RSTB(I91133), .Q(I91622) );
not I_5230 (I91110,I91622);
DFFARX1 I_5231  ( .D(I703674), .CLK(I2702), .RSTB(I91133), .Q(I91653) );
not I_5232 (I91670,I91653);
or I_5233 (I91687,I91670,I91591);
DFFARX1 I_5234  ( .D(I91687), .CLK(I2702), .RSTB(I91133), .Q(I91116) );
nand I_5235 (I91125,I91670,I91396);
DFFARX1 I_5236  ( .D(I91670), .CLK(I2702), .RSTB(I91133), .Q(I91095) );
not I_5237 (I91779,I2709);
not I_5238 (I91796,I144867);
nor I_5239 (I91813,I144855,I144861);
nand I_5240 (I91830,I91813,I144870);
DFFARX1 I_5241  ( .D(I91830), .CLK(I2702), .RSTB(I91779), .Q(I91753) );
nor I_5242 (I91861,I91796,I144855);
nand I_5243 (I91878,I91861,I144858);
not I_5244 (I91768,I91878);
DFFARX1 I_5245  ( .D(I91878), .CLK(I2702), .RSTB(I91779), .Q(I91750) );
not I_5246 (I91923,I144855);
not I_5247 (I91940,I91923);
not I_5248 (I91957,I144879);
nor I_5249 (I91974,I91957,I144852);
and I_5250 (I91991,I91974,I144873);
or I_5251 (I92008,I91991,I144864);
DFFARX1 I_5252  ( .D(I92008), .CLK(I2702), .RSTB(I91779), .Q(I92025) );
nor I_5253 (I92042,I92025,I91878);
nor I_5254 (I92059,I92025,I91940);
nand I_5255 (I91765,I91830,I92059);
nand I_5256 (I92090,I91796,I144879);
nand I_5257 (I92107,I92090,I92025);
and I_5258 (I92124,I92090,I92107);
DFFARX1 I_5259  ( .D(I92124), .CLK(I2702), .RSTB(I91779), .Q(I91747) );
DFFARX1 I_5260  ( .D(I92090), .CLK(I2702), .RSTB(I91779), .Q(I92155) );
and I_5261 (I91744,I91923,I92155);
DFFARX1 I_5262  ( .D(I144849), .CLK(I2702), .RSTB(I91779), .Q(I92186) );
not I_5263 (I92203,I92186);
nor I_5264 (I92220,I91878,I92203);
and I_5265 (I92237,I92186,I92220);
nand I_5266 (I91759,I92186,I91940);
DFFARX1 I_5267  ( .D(I92186), .CLK(I2702), .RSTB(I91779), .Q(I92268) );
not I_5268 (I91756,I92268);
DFFARX1 I_5269  ( .D(I144876), .CLK(I2702), .RSTB(I91779), .Q(I92299) );
not I_5270 (I92316,I92299);
or I_5271 (I92333,I92316,I92237);
DFFARX1 I_5272  ( .D(I92333), .CLK(I2702), .RSTB(I91779), .Q(I91762) );
nand I_5273 (I91771,I92316,I92042);
DFFARX1 I_5274  ( .D(I92316), .CLK(I2702), .RSTB(I91779), .Q(I91741) );
not I_5275 (I92425,I2709);
not I_5276 (I92442,I717537);
nor I_5277 (I92459,I717534,I717531);
nand I_5278 (I92476,I92459,I717552);
DFFARX1 I_5279  ( .D(I92476), .CLK(I2702), .RSTB(I92425), .Q(I92399) );
nor I_5280 (I92507,I92442,I717534);
nand I_5281 (I92524,I92507,I717555);
not I_5282 (I92414,I92524);
DFFARX1 I_5283  ( .D(I92524), .CLK(I2702), .RSTB(I92425), .Q(I92396) );
not I_5284 (I92569,I717534);
not I_5285 (I92586,I92569);
not I_5286 (I92603,I717528);
nor I_5287 (I92620,I92603,I717540);
and I_5288 (I92637,I92620,I717549);
or I_5289 (I92654,I92637,I717543);
DFFARX1 I_5290  ( .D(I92654), .CLK(I2702), .RSTB(I92425), .Q(I92671) );
nor I_5291 (I92688,I92671,I92524);
nor I_5292 (I92705,I92671,I92586);
nand I_5293 (I92411,I92476,I92705);
nand I_5294 (I92736,I92442,I717528);
nand I_5295 (I92753,I92736,I92671);
and I_5296 (I92770,I92736,I92753);
DFFARX1 I_5297  ( .D(I92770), .CLK(I2702), .RSTB(I92425), .Q(I92393) );
DFFARX1 I_5298  ( .D(I92736), .CLK(I2702), .RSTB(I92425), .Q(I92801) );
and I_5299 (I92390,I92569,I92801);
DFFARX1 I_5300  ( .D(I717558), .CLK(I2702), .RSTB(I92425), .Q(I92832) );
not I_5301 (I92849,I92832);
nor I_5302 (I92866,I92524,I92849);
and I_5303 (I92883,I92832,I92866);
nand I_5304 (I92405,I92832,I92586);
DFFARX1 I_5305  ( .D(I92832), .CLK(I2702), .RSTB(I92425), .Q(I92914) );
not I_5306 (I92402,I92914);
DFFARX1 I_5307  ( .D(I717546), .CLK(I2702), .RSTB(I92425), .Q(I92945) );
not I_5308 (I92962,I92945);
or I_5309 (I92979,I92962,I92883);
DFFARX1 I_5310  ( .D(I92979), .CLK(I2702), .RSTB(I92425), .Q(I92408) );
nand I_5311 (I92417,I92962,I92688);
DFFARX1 I_5312  ( .D(I92962), .CLK(I2702), .RSTB(I92425), .Q(I92387) );
not I_5313 (I93071,I2709);
not I_5314 (I93088,I296694);
nor I_5315 (I93105,I296691,I296679);
nand I_5316 (I93122,I93105,I296682);
DFFARX1 I_5317  ( .D(I93122), .CLK(I2702), .RSTB(I93071), .Q(I93045) );
nor I_5318 (I93153,I93088,I296691);
nand I_5319 (I93170,I93153,I296688);
not I_5320 (I93060,I93170);
DFFARX1 I_5321  ( .D(I93170), .CLK(I2702), .RSTB(I93071), .Q(I93042) );
not I_5322 (I93215,I296691);
not I_5323 (I93232,I93215);
not I_5324 (I93249,I296700);
nor I_5325 (I93266,I93249,I296676);
and I_5326 (I93283,I93266,I296697);
or I_5327 (I93300,I93283,I296685);
DFFARX1 I_5328  ( .D(I93300), .CLK(I2702), .RSTB(I93071), .Q(I93317) );
nor I_5329 (I93334,I93317,I93170);
nor I_5330 (I93351,I93317,I93232);
nand I_5331 (I93057,I93122,I93351);
nand I_5332 (I93382,I93088,I296700);
nand I_5333 (I93399,I93382,I93317);
and I_5334 (I93416,I93382,I93399);
DFFARX1 I_5335  ( .D(I93416), .CLK(I2702), .RSTB(I93071), .Q(I93039) );
DFFARX1 I_5336  ( .D(I93382), .CLK(I2702), .RSTB(I93071), .Q(I93447) );
and I_5337 (I93036,I93215,I93447);
DFFARX1 I_5338  ( .D(I296706), .CLK(I2702), .RSTB(I93071), .Q(I93478) );
not I_5339 (I93495,I93478);
nor I_5340 (I93512,I93170,I93495);
and I_5341 (I93529,I93478,I93512);
nand I_5342 (I93051,I93478,I93232);
DFFARX1 I_5343  ( .D(I93478), .CLK(I2702), .RSTB(I93071), .Q(I93560) );
not I_5344 (I93048,I93560);
DFFARX1 I_5345  ( .D(I296703), .CLK(I2702), .RSTB(I93071), .Q(I93591) );
not I_5346 (I93608,I93591);
or I_5347 (I93625,I93608,I93529);
DFFARX1 I_5348  ( .D(I93625), .CLK(I2702), .RSTB(I93071), .Q(I93054) );
nand I_5349 (I93063,I93608,I93334);
DFFARX1 I_5350  ( .D(I93608), .CLK(I2702), .RSTB(I93071), .Q(I93033) );
not I_5351 (I93717,I2709);
not I_5352 (I93734,I346725);
nor I_5353 (I93751,I346737,I346719);
nand I_5354 (I93768,I93751,I346734);
DFFARX1 I_5355  ( .D(I93768), .CLK(I2702), .RSTB(I93717), .Q(I93691) );
nor I_5356 (I93799,I93734,I346737);
nand I_5357 (I93816,I93799,I346722);
not I_5358 (I93706,I93816);
DFFARX1 I_5359  ( .D(I93816), .CLK(I2702), .RSTB(I93717), .Q(I93688) );
not I_5360 (I93861,I346737);
not I_5361 (I93878,I93861);
not I_5362 (I93895,I346731);
nor I_5363 (I93912,I93895,I346710);
and I_5364 (I93929,I93912,I346713);
or I_5365 (I93946,I93929,I346716);
DFFARX1 I_5366  ( .D(I93946), .CLK(I2702), .RSTB(I93717), .Q(I93963) );
nor I_5367 (I93980,I93963,I93816);
nor I_5368 (I93997,I93963,I93878);
nand I_5369 (I93703,I93768,I93997);
nand I_5370 (I94028,I93734,I346731);
nand I_5371 (I94045,I94028,I93963);
and I_5372 (I94062,I94028,I94045);
DFFARX1 I_5373  ( .D(I94062), .CLK(I2702), .RSTB(I93717), .Q(I93685) );
DFFARX1 I_5374  ( .D(I94028), .CLK(I2702), .RSTB(I93717), .Q(I94093) );
and I_5375 (I93682,I93861,I94093);
DFFARX1 I_5376  ( .D(I346707), .CLK(I2702), .RSTB(I93717), .Q(I94124) );
not I_5377 (I94141,I94124);
nor I_5378 (I94158,I93816,I94141);
and I_5379 (I94175,I94124,I94158);
nand I_5380 (I93697,I94124,I93878);
DFFARX1 I_5381  ( .D(I94124), .CLK(I2702), .RSTB(I93717), .Q(I94206) );
not I_5382 (I93694,I94206);
DFFARX1 I_5383  ( .D(I346728), .CLK(I2702), .RSTB(I93717), .Q(I94237) );
not I_5384 (I94254,I94237);
or I_5385 (I94271,I94254,I94175);
DFFARX1 I_5386  ( .D(I94271), .CLK(I2702), .RSTB(I93717), .Q(I93700) );
nand I_5387 (I93709,I94254,I93980);
DFFARX1 I_5388  ( .D(I94254), .CLK(I2702), .RSTB(I93717), .Q(I93679) );
not I_5389 (I94363,I2709);
not I_5390 (I94380,I443112);
nor I_5391 (I94397,I443100,I443106);
nand I_5392 (I94414,I94397,I443097);
DFFARX1 I_5393  ( .D(I94414), .CLK(I2702), .RSTB(I94363), .Q(I94337) );
nor I_5394 (I94445,I94380,I443100);
nand I_5395 (I94462,I94445,I443103);
not I_5396 (I94352,I94462);
DFFARX1 I_5397  ( .D(I94462), .CLK(I2702), .RSTB(I94363), .Q(I94334) );
not I_5398 (I94507,I443100);
not I_5399 (I94524,I94507);
not I_5400 (I94541,I443115);
nor I_5401 (I94558,I94541,I443127);
and I_5402 (I94575,I94558,I443109);
or I_5403 (I94592,I94575,I443124);
DFFARX1 I_5404  ( .D(I94592), .CLK(I2702), .RSTB(I94363), .Q(I94609) );
nor I_5405 (I94626,I94609,I94462);
nor I_5406 (I94643,I94609,I94524);
nand I_5407 (I94349,I94414,I94643);
nand I_5408 (I94674,I94380,I443115);
nand I_5409 (I94691,I94674,I94609);
and I_5410 (I94708,I94674,I94691);
DFFARX1 I_5411  ( .D(I94708), .CLK(I2702), .RSTB(I94363), .Q(I94331) );
DFFARX1 I_5412  ( .D(I94674), .CLK(I2702), .RSTB(I94363), .Q(I94739) );
and I_5413 (I94328,I94507,I94739);
DFFARX1 I_5414  ( .D(I443118), .CLK(I2702), .RSTB(I94363), .Q(I94770) );
not I_5415 (I94787,I94770);
nor I_5416 (I94804,I94462,I94787);
and I_5417 (I94821,I94770,I94804);
nand I_5418 (I94343,I94770,I94524);
DFFARX1 I_5419  ( .D(I94770), .CLK(I2702), .RSTB(I94363), .Q(I94852) );
not I_5420 (I94340,I94852);
DFFARX1 I_5421  ( .D(I443121), .CLK(I2702), .RSTB(I94363), .Q(I94883) );
not I_5422 (I94900,I94883);
or I_5423 (I94917,I94900,I94821);
DFFARX1 I_5424  ( .D(I94917), .CLK(I2702), .RSTB(I94363), .Q(I94346) );
nand I_5425 (I94355,I94900,I94626);
DFFARX1 I_5426  ( .D(I94900), .CLK(I2702), .RSTB(I94363), .Q(I94325) );
not I_5427 (I95009,I2709);
not I_5428 (I95026,I255588);
nor I_5429 (I95043,I255585,I255573);
nand I_5430 (I95060,I95043,I255576);
DFFARX1 I_5431  ( .D(I95060), .CLK(I2702), .RSTB(I95009), .Q(I94983) );
nor I_5432 (I95091,I95026,I255585);
nand I_5433 (I95108,I95091,I255582);
not I_5434 (I94998,I95108);
DFFARX1 I_5435  ( .D(I95108), .CLK(I2702), .RSTB(I95009), .Q(I94980) );
not I_5436 (I95153,I255585);
not I_5437 (I95170,I95153);
not I_5438 (I95187,I255594);
nor I_5439 (I95204,I95187,I255570);
and I_5440 (I95221,I95204,I255591);
or I_5441 (I95238,I95221,I255579);
DFFARX1 I_5442  ( .D(I95238), .CLK(I2702), .RSTB(I95009), .Q(I95255) );
nor I_5443 (I95272,I95255,I95108);
nor I_5444 (I95289,I95255,I95170);
nand I_5445 (I94995,I95060,I95289);
nand I_5446 (I95320,I95026,I255594);
nand I_5447 (I95337,I95320,I95255);
and I_5448 (I95354,I95320,I95337);
DFFARX1 I_5449  ( .D(I95354), .CLK(I2702), .RSTB(I95009), .Q(I94977) );
DFFARX1 I_5450  ( .D(I95320), .CLK(I2702), .RSTB(I95009), .Q(I95385) );
and I_5451 (I94974,I95153,I95385);
DFFARX1 I_5452  ( .D(I255600), .CLK(I2702), .RSTB(I95009), .Q(I95416) );
not I_5453 (I95433,I95416);
nor I_5454 (I95450,I95108,I95433);
and I_5455 (I95467,I95416,I95450);
nand I_5456 (I94989,I95416,I95170);
DFFARX1 I_5457  ( .D(I95416), .CLK(I2702), .RSTB(I95009), .Q(I95498) );
not I_5458 (I94986,I95498);
DFFARX1 I_5459  ( .D(I255597), .CLK(I2702), .RSTB(I95009), .Q(I95529) );
not I_5460 (I95546,I95529);
or I_5461 (I95563,I95546,I95467);
DFFARX1 I_5462  ( .D(I95563), .CLK(I2702), .RSTB(I95009), .Q(I94992) );
nand I_5463 (I95001,I95546,I95272);
DFFARX1 I_5464  ( .D(I95546), .CLK(I2702), .RSTB(I95009), .Q(I94971) );
not I_5465 (I95655,I2709);
not I_5466 (I95672,I2047);
nor I_5467 (I95689,I1343,I1847);
nand I_5468 (I95706,I95689,I1831);
DFFARX1 I_5469  ( .D(I95706), .CLK(I2702), .RSTB(I95655), .Q(I95629) );
nor I_5470 (I95737,I95672,I1343);
nand I_5471 (I95754,I95737,I2615);
not I_5472 (I95644,I95754);
DFFARX1 I_5473  ( .D(I95754), .CLK(I2702), .RSTB(I95655), .Q(I95626) );
not I_5474 (I95799,I1343);
not I_5475 (I95816,I95799);
not I_5476 (I95833,I2071);
nor I_5477 (I95850,I95833,I2447);
and I_5478 (I95867,I95850,I2455);
or I_5479 (I95884,I95867,I2159);
DFFARX1 I_5480  ( .D(I95884), .CLK(I2702), .RSTB(I95655), .Q(I95901) );
nor I_5481 (I95918,I95901,I95754);
nor I_5482 (I95935,I95901,I95816);
nand I_5483 (I95641,I95706,I95935);
nand I_5484 (I95966,I95672,I2071);
nand I_5485 (I95983,I95966,I95901);
and I_5486 (I96000,I95966,I95983);
DFFARX1 I_5487  ( .D(I96000), .CLK(I2702), .RSTB(I95655), .Q(I95623) );
DFFARX1 I_5488  ( .D(I95966), .CLK(I2702), .RSTB(I95655), .Q(I96031) );
and I_5489 (I95620,I95799,I96031);
DFFARX1 I_5490  ( .D(I1703), .CLK(I2702), .RSTB(I95655), .Q(I96062) );
not I_5491 (I96079,I96062);
nor I_5492 (I96096,I95754,I96079);
and I_5493 (I96113,I96062,I96096);
nand I_5494 (I95635,I96062,I95816);
DFFARX1 I_5495  ( .D(I96062), .CLK(I2702), .RSTB(I95655), .Q(I96144) );
not I_5496 (I95632,I96144);
DFFARX1 I_5497  ( .D(I2135), .CLK(I2702), .RSTB(I95655), .Q(I96175) );
not I_5498 (I96192,I96175);
or I_5499 (I96209,I96192,I96113);
DFFARX1 I_5500  ( .D(I96209), .CLK(I2702), .RSTB(I95655), .Q(I95638) );
nand I_5501 (I95647,I96192,I95918);
DFFARX1 I_5502  ( .D(I96192), .CLK(I2702), .RSTB(I95655), .Q(I95617) );
not I_5503 (I96301,I2709);
not I_5504 (I96318,I173376);
nor I_5505 (I96335,I173364,I173370);
nand I_5506 (I96352,I96335,I173379);
DFFARX1 I_5507  ( .D(I96352), .CLK(I2702), .RSTB(I96301), .Q(I96275) );
nor I_5508 (I96383,I96318,I173364);
nand I_5509 (I96400,I96383,I173367);
not I_5510 (I96290,I96400);
DFFARX1 I_5511  ( .D(I96400), .CLK(I2702), .RSTB(I96301), .Q(I96272) );
not I_5512 (I96445,I173364);
not I_5513 (I96462,I96445);
not I_5514 (I96479,I173388);
nor I_5515 (I96496,I96479,I173361);
and I_5516 (I96513,I96496,I173382);
or I_5517 (I96530,I96513,I173373);
DFFARX1 I_5518  ( .D(I96530), .CLK(I2702), .RSTB(I96301), .Q(I96547) );
nor I_5519 (I96564,I96547,I96400);
nor I_5520 (I96581,I96547,I96462);
nand I_5521 (I96287,I96352,I96581);
nand I_5522 (I96612,I96318,I173388);
nand I_5523 (I96629,I96612,I96547);
and I_5524 (I96646,I96612,I96629);
DFFARX1 I_5525  ( .D(I96646), .CLK(I2702), .RSTB(I96301), .Q(I96269) );
DFFARX1 I_5526  ( .D(I96612), .CLK(I2702), .RSTB(I96301), .Q(I96677) );
and I_5527 (I96266,I96445,I96677);
DFFARX1 I_5528  ( .D(I173358), .CLK(I2702), .RSTB(I96301), .Q(I96708) );
not I_5529 (I96725,I96708);
nor I_5530 (I96742,I96400,I96725);
and I_5531 (I96759,I96708,I96742);
nand I_5532 (I96281,I96708,I96462);
DFFARX1 I_5533  ( .D(I96708), .CLK(I2702), .RSTB(I96301), .Q(I96790) );
not I_5534 (I96278,I96790);
DFFARX1 I_5535  ( .D(I173385), .CLK(I2702), .RSTB(I96301), .Q(I96821) );
not I_5536 (I96838,I96821);
or I_5537 (I96855,I96838,I96759);
DFFARX1 I_5538  ( .D(I96855), .CLK(I2702), .RSTB(I96301), .Q(I96284) );
nand I_5539 (I96293,I96838,I96564);
DFFARX1 I_5540  ( .D(I96838), .CLK(I2702), .RSTB(I96301), .Q(I96263) );
not I_5541 (I96947,I2709);
not I_5542 (I96964,I353185);
nor I_5543 (I96981,I353197,I353179);
nand I_5544 (I96998,I96981,I353194);
DFFARX1 I_5545  ( .D(I96998), .CLK(I2702), .RSTB(I96947), .Q(I96921) );
nor I_5546 (I97029,I96964,I353197);
nand I_5547 (I97046,I97029,I353182);
not I_5548 (I96936,I97046);
DFFARX1 I_5549  ( .D(I97046), .CLK(I2702), .RSTB(I96947), .Q(I96918) );
not I_5550 (I97091,I353197);
not I_5551 (I97108,I97091);
not I_5552 (I97125,I353191);
nor I_5553 (I97142,I97125,I353170);
and I_5554 (I97159,I97142,I353173);
or I_5555 (I97176,I97159,I353176);
DFFARX1 I_5556  ( .D(I97176), .CLK(I2702), .RSTB(I96947), .Q(I97193) );
nor I_5557 (I97210,I97193,I97046);
nor I_5558 (I97227,I97193,I97108);
nand I_5559 (I96933,I96998,I97227);
nand I_5560 (I97258,I96964,I353191);
nand I_5561 (I97275,I97258,I97193);
and I_5562 (I97292,I97258,I97275);
DFFARX1 I_5563  ( .D(I97292), .CLK(I2702), .RSTB(I96947), .Q(I96915) );
DFFARX1 I_5564  ( .D(I97258), .CLK(I2702), .RSTB(I96947), .Q(I97323) );
and I_5565 (I96912,I97091,I97323);
DFFARX1 I_5566  ( .D(I353167), .CLK(I2702), .RSTB(I96947), .Q(I97354) );
not I_5567 (I97371,I97354);
nor I_5568 (I97388,I97046,I97371);
and I_5569 (I97405,I97354,I97388);
nand I_5570 (I96927,I97354,I97108);
DFFARX1 I_5571  ( .D(I97354), .CLK(I2702), .RSTB(I96947), .Q(I97436) );
not I_5572 (I96924,I97436);
DFFARX1 I_5573  ( .D(I353188), .CLK(I2702), .RSTB(I96947), .Q(I97467) );
not I_5574 (I97484,I97467);
or I_5575 (I97501,I97484,I97405);
DFFARX1 I_5576  ( .D(I97501), .CLK(I2702), .RSTB(I96947), .Q(I96930) );
nand I_5577 (I96939,I97484,I97210);
DFFARX1 I_5578  ( .D(I97484), .CLK(I2702), .RSTB(I96947), .Q(I96909) );
not I_5579 (I97593,I2709);
not I_5580 (I97610,I342203);
nor I_5581 (I97627,I342215,I342197);
nand I_5582 (I97644,I97627,I342212);
DFFARX1 I_5583  ( .D(I97644), .CLK(I2702), .RSTB(I97593), .Q(I97567) );
nor I_5584 (I97675,I97610,I342215);
nand I_5585 (I97692,I97675,I342200);
not I_5586 (I97582,I97692);
DFFARX1 I_5587  ( .D(I97692), .CLK(I2702), .RSTB(I97593), .Q(I97564) );
not I_5588 (I97737,I342215);
not I_5589 (I97754,I97737);
not I_5590 (I97771,I342209);
nor I_5591 (I97788,I97771,I342188);
and I_5592 (I97805,I97788,I342191);
or I_5593 (I97822,I97805,I342194);
DFFARX1 I_5594  ( .D(I97822), .CLK(I2702), .RSTB(I97593), .Q(I97839) );
nor I_5595 (I97856,I97839,I97692);
nor I_5596 (I97873,I97839,I97754);
nand I_5597 (I97579,I97644,I97873);
nand I_5598 (I97904,I97610,I342209);
nand I_5599 (I97921,I97904,I97839);
and I_5600 (I97938,I97904,I97921);
DFFARX1 I_5601  ( .D(I97938), .CLK(I2702), .RSTB(I97593), .Q(I97561) );
DFFARX1 I_5602  ( .D(I97904), .CLK(I2702), .RSTB(I97593), .Q(I97969) );
and I_5603 (I97558,I97737,I97969);
DFFARX1 I_5604  ( .D(I342185), .CLK(I2702), .RSTB(I97593), .Q(I98000) );
not I_5605 (I98017,I98000);
nor I_5606 (I98034,I97692,I98017);
and I_5607 (I98051,I98000,I98034);
nand I_5608 (I97573,I98000,I97754);
DFFARX1 I_5609  ( .D(I98000), .CLK(I2702), .RSTB(I97593), .Q(I98082) );
not I_5610 (I97570,I98082);
DFFARX1 I_5611  ( .D(I342206), .CLK(I2702), .RSTB(I97593), .Q(I98113) );
not I_5612 (I98130,I98113);
or I_5613 (I98147,I98130,I98051);
DFFARX1 I_5614  ( .D(I98147), .CLK(I2702), .RSTB(I97593), .Q(I97576) );
nand I_5615 (I97585,I98130,I97856);
DFFARX1 I_5616  ( .D(I98130), .CLK(I2702), .RSTB(I97593), .Q(I97555) );
not I_5617 (I98239,I2709);
not I_5618 (I98256,I315921);
nor I_5619 (I98273,I315918,I315906);
nand I_5620 (I98290,I98273,I315909);
DFFARX1 I_5621  ( .D(I98290), .CLK(I2702), .RSTB(I98239), .Q(I98213) );
nor I_5622 (I98321,I98256,I315918);
nand I_5623 (I98338,I98321,I315915);
not I_5624 (I98228,I98338);
DFFARX1 I_5625  ( .D(I98338), .CLK(I2702), .RSTB(I98239), .Q(I98210) );
not I_5626 (I98383,I315918);
not I_5627 (I98400,I98383);
not I_5628 (I98417,I315927);
nor I_5629 (I98434,I98417,I315903);
and I_5630 (I98451,I98434,I315924);
or I_5631 (I98468,I98451,I315912);
DFFARX1 I_5632  ( .D(I98468), .CLK(I2702), .RSTB(I98239), .Q(I98485) );
nor I_5633 (I98502,I98485,I98338);
nor I_5634 (I98519,I98485,I98400);
nand I_5635 (I98225,I98290,I98519);
nand I_5636 (I98550,I98256,I315927);
nand I_5637 (I98567,I98550,I98485);
and I_5638 (I98584,I98550,I98567);
DFFARX1 I_5639  ( .D(I98584), .CLK(I2702), .RSTB(I98239), .Q(I98207) );
DFFARX1 I_5640  ( .D(I98550), .CLK(I2702), .RSTB(I98239), .Q(I98615) );
and I_5641 (I98204,I98383,I98615);
DFFARX1 I_5642  ( .D(I315933), .CLK(I2702), .RSTB(I98239), .Q(I98646) );
not I_5643 (I98663,I98646);
nor I_5644 (I98680,I98338,I98663);
and I_5645 (I98697,I98646,I98680);
nand I_5646 (I98219,I98646,I98400);
DFFARX1 I_5647  ( .D(I98646), .CLK(I2702), .RSTB(I98239), .Q(I98728) );
not I_5648 (I98216,I98728);
DFFARX1 I_5649  ( .D(I315930), .CLK(I2702), .RSTB(I98239), .Q(I98759) );
not I_5650 (I98776,I98759);
or I_5651 (I98793,I98776,I98697);
DFFARX1 I_5652  ( .D(I98793), .CLK(I2702), .RSTB(I98239), .Q(I98222) );
nand I_5653 (I98231,I98776,I98502);
DFFARX1 I_5654  ( .D(I98776), .CLK(I2702), .RSTB(I98239), .Q(I98201) );
not I_5655 (I98885,I2709);
not I_5656 (I98902,I576251);
nor I_5657 (I98919,I576227,I576233);
nand I_5658 (I98936,I98919,I576236);
DFFARX1 I_5659  ( .D(I98936), .CLK(I2702), .RSTB(I98885), .Q(I98859) );
nor I_5660 (I98967,I98902,I576227);
nand I_5661 (I98984,I98967,I576245);
not I_5662 (I98874,I98984);
DFFARX1 I_5663  ( .D(I98984), .CLK(I2702), .RSTB(I98885), .Q(I98856) );
not I_5664 (I99029,I576227);
not I_5665 (I99046,I99029);
not I_5666 (I99063,I576224);
nor I_5667 (I99080,I99063,I576239);
and I_5668 (I99097,I99080,I576230);
or I_5669 (I99114,I99097,I576242);
DFFARX1 I_5670  ( .D(I99114), .CLK(I2702), .RSTB(I98885), .Q(I99131) );
nor I_5671 (I99148,I99131,I98984);
nor I_5672 (I99165,I99131,I99046);
nand I_5673 (I98871,I98936,I99165);
nand I_5674 (I99196,I98902,I576224);
nand I_5675 (I99213,I99196,I99131);
and I_5676 (I99230,I99196,I99213);
DFFARX1 I_5677  ( .D(I99230), .CLK(I2702), .RSTB(I98885), .Q(I98853) );
DFFARX1 I_5678  ( .D(I99196), .CLK(I2702), .RSTB(I98885), .Q(I99261) );
and I_5679 (I98850,I99029,I99261);
DFFARX1 I_5680  ( .D(I576254), .CLK(I2702), .RSTB(I98885), .Q(I99292) );
not I_5681 (I99309,I99292);
nor I_5682 (I99326,I98984,I99309);
and I_5683 (I99343,I99292,I99326);
nand I_5684 (I98865,I99292,I99046);
DFFARX1 I_5685  ( .D(I99292), .CLK(I2702), .RSTB(I98885), .Q(I99374) );
not I_5686 (I98862,I99374);
DFFARX1 I_5687  ( .D(I576248), .CLK(I2702), .RSTB(I98885), .Q(I99405) );
not I_5688 (I99422,I99405);
or I_5689 (I99439,I99422,I99343);
DFFARX1 I_5690  ( .D(I99439), .CLK(I2702), .RSTB(I98885), .Q(I98868) );
nand I_5691 (I98877,I99422,I99148);
DFFARX1 I_5692  ( .D(I99422), .CLK(I2702), .RSTB(I98885), .Q(I98847) );
not I_5693 (I99531,I2709);
not I_5694 (I99548,I461030);
nor I_5695 (I99565,I461018,I461024);
nand I_5696 (I99582,I99565,I461015);
DFFARX1 I_5697  ( .D(I99582), .CLK(I2702), .RSTB(I99531), .Q(I99505) );
nor I_5698 (I99613,I99548,I461018);
nand I_5699 (I99630,I99613,I461021);
not I_5700 (I99520,I99630);
DFFARX1 I_5701  ( .D(I99630), .CLK(I2702), .RSTB(I99531), .Q(I99502) );
not I_5702 (I99675,I461018);
not I_5703 (I99692,I99675);
not I_5704 (I99709,I461033);
nor I_5705 (I99726,I99709,I461045);
and I_5706 (I99743,I99726,I461027);
or I_5707 (I99760,I99743,I461042);
DFFARX1 I_5708  ( .D(I99760), .CLK(I2702), .RSTB(I99531), .Q(I99777) );
nor I_5709 (I99794,I99777,I99630);
nor I_5710 (I99811,I99777,I99692);
nand I_5711 (I99517,I99582,I99811);
nand I_5712 (I99842,I99548,I461033);
nand I_5713 (I99859,I99842,I99777);
and I_5714 (I99876,I99842,I99859);
DFFARX1 I_5715  ( .D(I99876), .CLK(I2702), .RSTB(I99531), .Q(I99499) );
DFFARX1 I_5716  ( .D(I99842), .CLK(I2702), .RSTB(I99531), .Q(I99907) );
and I_5717 (I99496,I99675,I99907);
DFFARX1 I_5718  ( .D(I461036), .CLK(I2702), .RSTB(I99531), .Q(I99938) );
not I_5719 (I99955,I99938);
nor I_5720 (I99972,I99630,I99955);
and I_5721 (I99989,I99938,I99972);
nand I_5722 (I99511,I99938,I99692);
DFFARX1 I_5723  ( .D(I99938), .CLK(I2702), .RSTB(I99531), .Q(I100020) );
not I_5724 (I99508,I100020);
DFFARX1 I_5725  ( .D(I461039), .CLK(I2702), .RSTB(I99531), .Q(I100051) );
not I_5726 (I100068,I100051);
or I_5727 (I100085,I100068,I99989);
DFFARX1 I_5728  ( .D(I100085), .CLK(I2702), .RSTB(I99531), .Q(I99514) );
nand I_5729 (I99523,I100068,I99794);
DFFARX1 I_5730  ( .D(I100068), .CLK(I2702), .RSTB(I99531), .Q(I99493) );
not I_5731 (I100177,I2709);
not I_5732 (I100194,I399697);
nor I_5733 (I100211,I399709,I399691);
nand I_5734 (I100228,I100211,I399706);
DFFARX1 I_5735  ( .D(I100228), .CLK(I2702), .RSTB(I100177), .Q(I100151) );
nor I_5736 (I100259,I100194,I399709);
nand I_5737 (I100276,I100259,I399694);
not I_5738 (I100166,I100276);
DFFARX1 I_5739  ( .D(I100276), .CLK(I2702), .RSTB(I100177), .Q(I100148) );
not I_5740 (I100321,I399709);
not I_5741 (I100338,I100321);
not I_5742 (I100355,I399703);
nor I_5743 (I100372,I100355,I399682);
and I_5744 (I100389,I100372,I399685);
or I_5745 (I100406,I100389,I399688);
DFFARX1 I_5746  ( .D(I100406), .CLK(I2702), .RSTB(I100177), .Q(I100423) );
nor I_5747 (I100440,I100423,I100276);
nor I_5748 (I100457,I100423,I100338);
nand I_5749 (I100163,I100228,I100457);
nand I_5750 (I100488,I100194,I399703);
nand I_5751 (I100505,I100488,I100423);
and I_5752 (I100522,I100488,I100505);
DFFARX1 I_5753  ( .D(I100522), .CLK(I2702), .RSTB(I100177), .Q(I100145) );
DFFARX1 I_5754  ( .D(I100488), .CLK(I2702), .RSTB(I100177), .Q(I100553) );
and I_5755 (I100142,I100321,I100553);
DFFARX1 I_5756  ( .D(I399679), .CLK(I2702), .RSTB(I100177), .Q(I100584) );
not I_5757 (I100601,I100584);
nor I_5758 (I100618,I100276,I100601);
and I_5759 (I100635,I100584,I100618);
nand I_5760 (I100157,I100584,I100338);
DFFARX1 I_5761  ( .D(I100584), .CLK(I2702), .RSTB(I100177), .Q(I100666) );
not I_5762 (I100154,I100666);
DFFARX1 I_5763  ( .D(I399700), .CLK(I2702), .RSTB(I100177), .Q(I100697) );
not I_5764 (I100714,I100697);
or I_5765 (I100731,I100714,I100635);
DFFARX1 I_5766  ( .D(I100731), .CLK(I2702), .RSTB(I100177), .Q(I100160) );
nand I_5767 (I100169,I100714,I100440);
DFFARX1 I_5768  ( .D(I100714), .CLK(I2702), .RSTB(I100177), .Q(I100139) );
not I_5769 (I100823,I2709);
not I_5770 (I100840,I419315);
nor I_5771 (I100857,I419297,I419312);
nand I_5772 (I100874,I100857,I419321);
DFFARX1 I_5773  ( .D(I100874), .CLK(I2702), .RSTB(I100823), .Q(I100797) );
nor I_5774 (I100905,I100840,I419297);
nand I_5775 (I100922,I100905,I419324);
not I_5776 (I100812,I100922);
DFFARX1 I_5777  ( .D(I100922), .CLK(I2702), .RSTB(I100823), .Q(I100794) );
not I_5778 (I100967,I419297);
not I_5779 (I100984,I100967);
not I_5780 (I101001,I419327);
nor I_5781 (I101018,I101001,I419303);
and I_5782 (I101035,I101018,I419306);
or I_5783 (I101052,I101035,I419300);
DFFARX1 I_5784  ( .D(I101052), .CLK(I2702), .RSTB(I100823), .Q(I101069) );
nor I_5785 (I101086,I101069,I100922);
nor I_5786 (I101103,I101069,I100984);
nand I_5787 (I100809,I100874,I101103);
nand I_5788 (I101134,I100840,I419327);
nand I_5789 (I101151,I101134,I101069);
and I_5790 (I101168,I101134,I101151);
DFFARX1 I_5791  ( .D(I101168), .CLK(I2702), .RSTB(I100823), .Q(I100791) );
DFFARX1 I_5792  ( .D(I101134), .CLK(I2702), .RSTB(I100823), .Q(I101199) );
and I_5793 (I100788,I100967,I101199);
DFFARX1 I_5794  ( .D(I419309), .CLK(I2702), .RSTB(I100823), .Q(I101230) );
not I_5795 (I101247,I101230);
nor I_5796 (I101264,I100922,I101247);
and I_5797 (I101281,I101230,I101264);
nand I_5798 (I100803,I101230,I100984);
DFFARX1 I_5799  ( .D(I101230), .CLK(I2702), .RSTB(I100823), .Q(I101312) );
not I_5800 (I100800,I101312);
DFFARX1 I_5801  ( .D(I419318), .CLK(I2702), .RSTB(I100823), .Q(I101343) );
not I_5802 (I101360,I101343);
or I_5803 (I101377,I101360,I101281);
DFFARX1 I_5804  ( .D(I101377), .CLK(I2702), .RSTB(I100823), .Q(I100806) );
nand I_5805 (I100815,I101360,I101086);
DFFARX1 I_5806  ( .D(I101360), .CLK(I2702), .RSTB(I100823), .Q(I100785) );
not I_5807 (I101469,I2709);
not I_5808 (I101486,I218918);
nor I_5809 (I101503,I218948,I218927);
nand I_5810 (I101520,I101503,I218939);
DFFARX1 I_5811  ( .D(I101520), .CLK(I2702), .RSTB(I101469), .Q(I101443) );
nor I_5812 (I101551,I101486,I218948);
nand I_5813 (I101568,I101551,I218921);
not I_5814 (I101458,I101568);
DFFARX1 I_5815  ( .D(I101568), .CLK(I2702), .RSTB(I101469), .Q(I101440) );
not I_5816 (I101613,I218948);
not I_5817 (I101630,I101613);
not I_5818 (I101647,I218924);
nor I_5819 (I101664,I101647,I218942);
and I_5820 (I101681,I101664,I218933);
or I_5821 (I101698,I101681,I218930);
DFFARX1 I_5822  ( .D(I101698), .CLK(I2702), .RSTB(I101469), .Q(I101715) );
nor I_5823 (I101732,I101715,I101568);
nor I_5824 (I101749,I101715,I101630);
nand I_5825 (I101455,I101520,I101749);
nand I_5826 (I101780,I101486,I218924);
nand I_5827 (I101797,I101780,I101715);
and I_5828 (I101814,I101780,I101797);
DFFARX1 I_5829  ( .D(I101814), .CLK(I2702), .RSTB(I101469), .Q(I101437) );
DFFARX1 I_5830  ( .D(I101780), .CLK(I2702), .RSTB(I101469), .Q(I101845) );
and I_5831 (I101434,I101613,I101845);
DFFARX1 I_5832  ( .D(I218936), .CLK(I2702), .RSTB(I101469), .Q(I101876) );
not I_5833 (I101893,I101876);
nor I_5834 (I101910,I101568,I101893);
and I_5835 (I101927,I101876,I101910);
nand I_5836 (I101449,I101876,I101630);
DFFARX1 I_5837  ( .D(I101876), .CLK(I2702), .RSTB(I101469), .Q(I101958) );
not I_5838 (I101446,I101958);
DFFARX1 I_5839  ( .D(I218945), .CLK(I2702), .RSTB(I101469), .Q(I101989) );
not I_5840 (I102006,I101989);
or I_5841 (I102023,I102006,I101927);
DFFARX1 I_5842  ( .D(I102023), .CLK(I2702), .RSTB(I101469), .Q(I101452) );
nand I_5843 (I101461,I102006,I101732);
DFFARX1 I_5844  ( .D(I102006), .CLK(I2702), .RSTB(I101469), .Q(I101431) );
not I_5845 (I102115,I2709);
not I_5846 (I102132,I158127);
nor I_5847 (I102149,I158115,I158121);
nand I_5848 (I102166,I102149,I158130);
DFFARX1 I_5849  ( .D(I102166), .CLK(I2702), .RSTB(I102115), .Q(I102089) );
nor I_5850 (I102197,I102132,I158115);
nand I_5851 (I102214,I102197,I158118);
not I_5852 (I102104,I102214);
DFFARX1 I_5853  ( .D(I102214), .CLK(I2702), .RSTB(I102115), .Q(I102086) );
not I_5854 (I102259,I158115);
not I_5855 (I102276,I102259);
not I_5856 (I102293,I158139);
nor I_5857 (I102310,I102293,I158112);
and I_5858 (I102327,I102310,I158133);
or I_5859 (I102344,I102327,I158124);
DFFARX1 I_5860  ( .D(I102344), .CLK(I2702), .RSTB(I102115), .Q(I102361) );
nor I_5861 (I102378,I102361,I102214);
nor I_5862 (I102395,I102361,I102276);
nand I_5863 (I102101,I102166,I102395);
nand I_5864 (I102426,I102132,I158139);
nand I_5865 (I102443,I102426,I102361);
and I_5866 (I102460,I102426,I102443);
DFFARX1 I_5867  ( .D(I102460), .CLK(I2702), .RSTB(I102115), .Q(I102083) );
DFFARX1 I_5868  ( .D(I102426), .CLK(I2702), .RSTB(I102115), .Q(I102491) );
and I_5869 (I102080,I102259,I102491);
DFFARX1 I_5870  ( .D(I158109), .CLK(I2702), .RSTB(I102115), .Q(I102522) );
not I_5871 (I102539,I102522);
nor I_5872 (I102556,I102214,I102539);
and I_5873 (I102573,I102522,I102556);
nand I_5874 (I102095,I102522,I102276);
DFFARX1 I_5875  ( .D(I102522), .CLK(I2702), .RSTB(I102115), .Q(I102604) );
not I_5876 (I102092,I102604);
DFFARX1 I_5877  ( .D(I158136), .CLK(I2702), .RSTB(I102115), .Q(I102635) );
not I_5878 (I102652,I102635);
or I_5879 (I102669,I102652,I102573);
DFFARX1 I_5880  ( .D(I102669), .CLK(I2702), .RSTB(I102115), .Q(I102098) );
nand I_5881 (I102107,I102652,I102378);
DFFARX1 I_5882  ( .D(I102652), .CLK(I2702), .RSTB(I102115), .Q(I102077) );
not I_5883 (I102761,I2709);
not I_5884 (I102778,I368043);
nor I_5885 (I102795,I368055,I368037);
nand I_5886 (I102812,I102795,I368052);
DFFARX1 I_5887  ( .D(I102812), .CLK(I2702), .RSTB(I102761), .Q(I102735) );
nor I_5888 (I102843,I102778,I368055);
nand I_5889 (I102860,I102843,I368040);
not I_5890 (I102750,I102860);
DFFARX1 I_5891  ( .D(I102860), .CLK(I2702), .RSTB(I102761), .Q(I102732) );
not I_5892 (I102905,I368055);
not I_5893 (I102922,I102905);
not I_5894 (I102939,I368049);
nor I_5895 (I102956,I102939,I368028);
and I_5896 (I102973,I102956,I368031);
or I_5897 (I102990,I102973,I368034);
DFFARX1 I_5898  ( .D(I102990), .CLK(I2702), .RSTB(I102761), .Q(I103007) );
nor I_5899 (I103024,I103007,I102860);
nor I_5900 (I103041,I103007,I102922);
nand I_5901 (I102747,I102812,I103041);
nand I_5902 (I103072,I102778,I368049);
nand I_5903 (I103089,I103072,I103007);
and I_5904 (I103106,I103072,I103089);
DFFARX1 I_5905  ( .D(I103106), .CLK(I2702), .RSTB(I102761), .Q(I102729) );
DFFARX1 I_5906  ( .D(I103072), .CLK(I2702), .RSTB(I102761), .Q(I103137) );
and I_5907 (I102726,I102905,I103137);
DFFARX1 I_5908  ( .D(I368025), .CLK(I2702), .RSTB(I102761), .Q(I103168) );
not I_5909 (I103185,I103168);
nor I_5910 (I103202,I102860,I103185);
and I_5911 (I103219,I103168,I103202);
nand I_5912 (I102741,I103168,I102922);
DFFARX1 I_5913  ( .D(I103168), .CLK(I2702), .RSTB(I102761), .Q(I103250) );
not I_5914 (I102738,I103250);
DFFARX1 I_5915  ( .D(I368046), .CLK(I2702), .RSTB(I102761), .Q(I103281) );
not I_5916 (I103298,I103281);
or I_5917 (I103315,I103298,I103219);
DFFARX1 I_5918  ( .D(I103315), .CLK(I2702), .RSTB(I102761), .Q(I102744) );
nand I_5919 (I102753,I103298,I103024);
DFFARX1 I_5920  ( .D(I103298), .CLK(I2702), .RSTB(I102761), .Q(I102723) );
not I_5921 (I103407,I2709);
not I_5922 (I103424,I7203);
nor I_5923 (I103441,I7215,I7200);
nand I_5924 (I103458,I103441,I7212);
DFFARX1 I_5925  ( .D(I103458), .CLK(I2702), .RSTB(I103407), .Q(I103381) );
nor I_5926 (I103489,I103424,I7215);
nand I_5927 (I103506,I103489,I7230);
not I_5928 (I103396,I103506);
DFFARX1 I_5929  ( .D(I103506), .CLK(I2702), .RSTB(I103407), .Q(I103378) );
not I_5930 (I103551,I7215);
not I_5931 (I103568,I103551);
not I_5932 (I103585,I7206);
nor I_5933 (I103602,I103585,I7218);
and I_5934 (I103619,I103602,I7209);
or I_5935 (I103636,I103619,I7224);
DFFARX1 I_5936  ( .D(I103636), .CLK(I2702), .RSTB(I103407), .Q(I103653) );
nor I_5937 (I103670,I103653,I103506);
nor I_5938 (I103687,I103653,I103568);
nand I_5939 (I103393,I103458,I103687);
nand I_5940 (I103718,I103424,I7206);
nand I_5941 (I103735,I103718,I103653);
and I_5942 (I103752,I103718,I103735);
DFFARX1 I_5943  ( .D(I103752), .CLK(I2702), .RSTB(I103407), .Q(I103375) );
DFFARX1 I_5944  ( .D(I103718), .CLK(I2702), .RSTB(I103407), .Q(I103783) );
and I_5945 (I103372,I103551,I103783);
DFFARX1 I_5946  ( .D(I7227), .CLK(I2702), .RSTB(I103407), .Q(I103814) );
not I_5947 (I103831,I103814);
nor I_5948 (I103848,I103506,I103831);
and I_5949 (I103865,I103814,I103848);
nand I_5950 (I103387,I103814,I103568);
DFFARX1 I_5951  ( .D(I103814), .CLK(I2702), .RSTB(I103407), .Q(I103896) );
not I_5952 (I103384,I103896);
DFFARX1 I_5953  ( .D(I7221), .CLK(I2702), .RSTB(I103407), .Q(I103927) );
not I_5954 (I103944,I103927);
or I_5955 (I103961,I103944,I103865);
DFFARX1 I_5956  ( .D(I103961), .CLK(I2702), .RSTB(I103407), .Q(I103390) );
nand I_5957 (I103399,I103944,I103670);
DFFARX1 I_5958  ( .D(I103944), .CLK(I2702), .RSTB(I103407), .Q(I103369) );
not I_5959 (I104053,I2709);
not I_5960 (I104070,I436176);
nor I_5961 (I104087,I436164,I436170);
nand I_5962 (I104104,I104087,I436161);
DFFARX1 I_5963  ( .D(I104104), .CLK(I2702), .RSTB(I104053), .Q(I104027) );
nor I_5964 (I104135,I104070,I436164);
nand I_5965 (I104152,I104135,I436167);
not I_5966 (I104042,I104152);
DFFARX1 I_5967  ( .D(I104152), .CLK(I2702), .RSTB(I104053), .Q(I104024) );
not I_5968 (I104197,I436164);
not I_5969 (I104214,I104197);
not I_5970 (I104231,I436179);
nor I_5971 (I104248,I104231,I436191);
and I_5972 (I104265,I104248,I436173);
or I_5973 (I104282,I104265,I436188);
DFFARX1 I_5974  ( .D(I104282), .CLK(I2702), .RSTB(I104053), .Q(I104299) );
nor I_5975 (I104316,I104299,I104152);
nor I_5976 (I104333,I104299,I104214);
nand I_5977 (I104039,I104104,I104333);
nand I_5978 (I104364,I104070,I436179);
nand I_5979 (I104381,I104364,I104299);
and I_5980 (I104398,I104364,I104381);
DFFARX1 I_5981  ( .D(I104398), .CLK(I2702), .RSTB(I104053), .Q(I104021) );
DFFARX1 I_5982  ( .D(I104364), .CLK(I2702), .RSTB(I104053), .Q(I104429) );
and I_5983 (I104018,I104197,I104429);
DFFARX1 I_5984  ( .D(I436182), .CLK(I2702), .RSTB(I104053), .Q(I104460) );
not I_5985 (I104477,I104460);
nor I_5986 (I104494,I104152,I104477);
and I_5987 (I104511,I104460,I104494);
nand I_5988 (I104033,I104460,I104214);
DFFARX1 I_5989  ( .D(I104460), .CLK(I2702), .RSTB(I104053), .Q(I104542) );
not I_5990 (I104030,I104542);
DFFARX1 I_5991  ( .D(I436185), .CLK(I2702), .RSTB(I104053), .Q(I104573) );
not I_5992 (I104590,I104573);
or I_5993 (I104607,I104590,I104511);
DFFARX1 I_5994  ( .D(I104607), .CLK(I2702), .RSTB(I104053), .Q(I104036) );
nand I_5995 (I104045,I104590,I104316);
DFFARX1 I_5996  ( .D(I104590), .CLK(I2702), .RSTB(I104053), .Q(I104015) );
not I_5997 (I104699,I2709);
not I_5998 (I104716,I284760);
nor I_5999 (I104733,I284757,I284745);
nand I_6000 (I104750,I104733,I284748);
DFFARX1 I_6001  ( .D(I104750), .CLK(I2702), .RSTB(I104699), .Q(I104673) );
nor I_6002 (I104781,I104716,I284757);
nand I_6003 (I104798,I104781,I284754);
not I_6004 (I104688,I104798);
DFFARX1 I_6005  ( .D(I104798), .CLK(I2702), .RSTB(I104699), .Q(I104670) );
not I_6006 (I104843,I284757);
not I_6007 (I104860,I104843);
not I_6008 (I104877,I284766);
nor I_6009 (I104894,I104877,I284742);
and I_6010 (I104911,I104894,I284763);
or I_6011 (I104928,I104911,I284751);
DFFARX1 I_6012  ( .D(I104928), .CLK(I2702), .RSTB(I104699), .Q(I104945) );
nor I_6013 (I104962,I104945,I104798);
nor I_6014 (I104979,I104945,I104860);
nand I_6015 (I104685,I104750,I104979);
nand I_6016 (I105010,I104716,I284766);
nand I_6017 (I105027,I105010,I104945);
and I_6018 (I105044,I105010,I105027);
DFFARX1 I_6019  ( .D(I105044), .CLK(I2702), .RSTB(I104699), .Q(I104667) );
DFFARX1 I_6020  ( .D(I105010), .CLK(I2702), .RSTB(I104699), .Q(I105075) );
and I_6021 (I104664,I104843,I105075);
DFFARX1 I_6022  ( .D(I284772), .CLK(I2702), .RSTB(I104699), .Q(I105106) );
not I_6023 (I105123,I105106);
nor I_6024 (I105140,I104798,I105123);
and I_6025 (I105157,I105106,I105140);
nand I_6026 (I104679,I105106,I104860);
DFFARX1 I_6027  ( .D(I105106), .CLK(I2702), .RSTB(I104699), .Q(I105188) );
not I_6028 (I104676,I105188);
DFFARX1 I_6029  ( .D(I284769), .CLK(I2702), .RSTB(I104699), .Q(I105219) );
not I_6030 (I105236,I105219);
or I_6031 (I105253,I105236,I105157);
DFFARX1 I_6032  ( .D(I105253), .CLK(I2702), .RSTB(I104699), .Q(I104682) );
nand I_6033 (I104691,I105236,I104962);
DFFARX1 I_6034  ( .D(I105236), .CLK(I2702), .RSTB(I104699), .Q(I104661) );
not I_6035 (I105345,I2709);
not I_6036 (I105362,I510801);
nor I_6037 (I105379,I510777,I510783);
nand I_6038 (I105396,I105379,I510786);
DFFARX1 I_6039  ( .D(I105396), .CLK(I2702), .RSTB(I105345), .Q(I105319) );
nor I_6040 (I105427,I105362,I510777);
nand I_6041 (I105444,I105427,I510795);
not I_6042 (I105334,I105444);
DFFARX1 I_6043  ( .D(I105444), .CLK(I2702), .RSTB(I105345), .Q(I105316) );
not I_6044 (I105489,I510777);
not I_6045 (I105506,I105489);
not I_6046 (I105523,I510774);
nor I_6047 (I105540,I105523,I510789);
and I_6048 (I105557,I105540,I510780);
or I_6049 (I105574,I105557,I510792);
DFFARX1 I_6050  ( .D(I105574), .CLK(I2702), .RSTB(I105345), .Q(I105591) );
nor I_6051 (I105608,I105591,I105444);
nor I_6052 (I105625,I105591,I105506);
nand I_6053 (I105331,I105396,I105625);
nand I_6054 (I105656,I105362,I510774);
nand I_6055 (I105673,I105656,I105591);
and I_6056 (I105690,I105656,I105673);
DFFARX1 I_6057  ( .D(I105690), .CLK(I2702), .RSTB(I105345), .Q(I105313) );
DFFARX1 I_6058  ( .D(I105656), .CLK(I2702), .RSTB(I105345), .Q(I105721) );
and I_6059 (I105310,I105489,I105721);
DFFARX1 I_6060  ( .D(I510804), .CLK(I2702), .RSTB(I105345), .Q(I105752) );
not I_6061 (I105769,I105752);
nor I_6062 (I105786,I105444,I105769);
and I_6063 (I105803,I105752,I105786);
nand I_6064 (I105325,I105752,I105506);
DFFARX1 I_6065  ( .D(I105752), .CLK(I2702), .RSTB(I105345), .Q(I105834) );
not I_6066 (I105322,I105834);
DFFARX1 I_6067  ( .D(I510798), .CLK(I2702), .RSTB(I105345), .Q(I105865) );
not I_6068 (I105882,I105865);
or I_6069 (I105899,I105882,I105803);
DFFARX1 I_6070  ( .D(I105899), .CLK(I2702), .RSTB(I105345), .Q(I105328) );
nand I_6071 (I105337,I105882,I105608);
DFFARX1 I_6072  ( .D(I105882), .CLK(I2702), .RSTB(I105345), .Q(I105307) );
not I_6073 (I105991,I2709);
not I_6074 (I106008,I575061);
nor I_6075 (I106025,I575037,I575043);
nand I_6076 (I106042,I106025,I575046);
DFFARX1 I_6077  ( .D(I106042), .CLK(I2702), .RSTB(I105991), .Q(I105965) );
nor I_6078 (I106073,I106008,I575037);
nand I_6079 (I106090,I106073,I575055);
not I_6080 (I105980,I106090);
DFFARX1 I_6081  ( .D(I106090), .CLK(I2702), .RSTB(I105991), .Q(I105962) );
not I_6082 (I106135,I575037);
not I_6083 (I106152,I106135);
not I_6084 (I106169,I575034);
nor I_6085 (I106186,I106169,I575049);
and I_6086 (I106203,I106186,I575040);
or I_6087 (I106220,I106203,I575052);
DFFARX1 I_6088  ( .D(I106220), .CLK(I2702), .RSTB(I105991), .Q(I106237) );
nor I_6089 (I106254,I106237,I106090);
nor I_6090 (I106271,I106237,I106152);
nand I_6091 (I105977,I106042,I106271);
nand I_6092 (I106302,I106008,I575034);
nand I_6093 (I106319,I106302,I106237);
and I_6094 (I106336,I106302,I106319);
DFFARX1 I_6095  ( .D(I106336), .CLK(I2702), .RSTB(I105991), .Q(I105959) );
DFFARX1 I_6096  ( .D(I106302), .CLK(I2702), .RSTB(I105991), .Q(I106367) );
and I_6097 (I105956,I106135,I106367);
DFFARX1 I_6098  ( .D(I575064), .CLK(I2702), .RSTB(I105991), .Q(I106398) );
not I_6099 (I106415,I106398);
nor I_6100 (I106432,I106090,I106415);
and I_6101 (I106449,I106398,I106432);
nand I_6102 (I105971,I106398,I106152);
DFFARX1 I_6103  ( .D(I106398), .CLK(I2702), .RSTB(I105991), .Q(I106480) );
not I_6104 (I105968,I106480);
DFFARX1 I_6105  ( .D(I575058), .CLK(I2702), .RSTB(I105991), .Q(I106511) );
not I_6106 (I106528,I106511);
or I_6107 (I106545,I106528,I106449);
DFFARX1 I_6108  ( .D(I106545), .CLK(I2702), .RSTB(I105991), .Q(I105974) );
nand I_6109 (I105983,I106528,I106254);
DFFARX1 I_6110  ( .D(I106528), .CLK(I2702), .RSTB(I105991), .Q(I105953) );
not I_6111 (I106637,I2709);
not I_6112 (I106654,I248295);
nor I_6113 (I106671,I248292,I248280);
nand I_6114 (I106688,I106671,I248283);
DFFARX1 I_6115  ( .D(I106688), .CLK(I2702), .RSTB(I106637), .Q(I106611) );
nor I_6116 (I106719,I106654,I248292);
nand I_6117 (I106736,I106719,I248289);
not I_6118 (I106626,I106736);
DFFARX1 I_6119  ( .D(I106736), .CLK(I2702), .RSTB(I106637), .Q(I106608) );
not I_6120 (I106781,I248292);
not I_6121 (I106798,I106781);
not I_6122 (I106815,I248301);
nor I_6123 (I106832,I106815,I248277);
and I_6124 (I106849,I106832,I248298);
or I_6125 (I106866,I106849,I248286);
DFFARX1 I_6126  ( .D(I106866), .CLK(I2702), .RSTB(I106637), .Q(I106883) );
nor I_6127 (I106900,I106883,I106736);
nor I_6128 (I106917,I106883,I106798);
nand I_6129 (I106623,I106688,I106917);
nand I_6130 (I106948,I106654,I248301);
nand I_6131 (I106965,I106948,I106883);
and I_6132 (I106982,I106948,I106965);
DFFARX1 I_6133  ( .D(I106982), .CLK(I2702), .RSTB(I106637), .Q(I106605) );
DFFARX1 I_6134  ( .D(I106948), .CLK(I2702), .RSTB(I106637), .Q(I107013) );
and I_6135 (I106602,I106781,I107013);
DFFARX1 I_6136  ( .D(I248307), .CLK(I2702), .RSTB(I106637), .Q(I107044) );
not I_6137 (I107061,I107044);
nor I_6138 (I107078,I106736,I107061);
and I_6139 (I107095,I107044,I107078);
nand I_6140 (I106617,I107044,I106798);
DFFARX1 I_6141  ( .D(I107044), .CLK(I2702), .RSTB(I106637), .Q(I107126) );
not I_6142 (I106614,I107126);
DFFARX1 I_6143  ( .D(I248304), .CLK(I2702), .RSTB(I106637), .Q(I107157) );
not I_6144 (I107174,I107157);
or I_6145 (I107191,I107174,I107095);
DFFARX1 I_6146  ( .D(I107191), .CLK(I2702), .RSTB(I106637), .Q(I106620) );
nand I_6147 (I106629,I107174,I106900);
DFFARX1 I_6148  ( .D(I107174), .CLK(I2702), .RSTB(I106637), .Q(I106599) );
not I_6149 (I107283,I2709);
not I_6150 (I107300,I649528);
nor I_6151 (I107317,I649543,I649558);
nand I_6152 (I107334,I107317,I649546);
DFFARX1 I_6153  ( .D(I107334), .CLK(I2702), .RSTB(I107283), .Q(I107257) );
nor I_6154 (I107365,I107300,I649543);
nand I_6155 (I107382,I107365,I649549);
not I_6156 (I107272,I107382);
DFFARX1 I_6157  ( .D(I107382), .CLK(I2702), .RSTB(I107283), .Q(I107254) );
not I_6158 (I107427,I649543);
not I_6159 (I107444,I107427);
not I_6160 (I107461,I649555);
nor I_6161 (I107478,I107461,I649552);
and I_6162 (I107495,I107478,I649531);
or I_6163 (I107512,I107495,I649540);
DFFARX1 I_6164  ( .D(I107512), .CLK(I2702), .RSTB(I107283), .Q(I107529) );
nor I_6165 (I107546,I107529,I107382);
nor I_6166 (I107563,I107529,I107444);
nand I_6167 (I107269,I107334,I107563);
nand I_6168 (I107594,I107300,I649555);
nand I_6169 (I107611,I107594,I107529);
and I_6170 (I107628,I107594,I107611);
DFFARX1 I_6171  ( .D(I107628), .CLK(I2702), .RSTB(I107283), .Q(I107251) );
DFFARX1 I_6172  ( .D(I107594), .CLK(I2702), .RSTB(I107283), .Q(I107659) );
and I_6173 (I107248,I107427,I107659);
DFFARX1 I_6174  ( .D(I649537), .CLK(I2702), .RSTB(I107283), .Q(I107690) );
not I_6175 (I107707,I107690);
nor I_6176 (I107724,I107382,I107707);
and I_6177 (I107741,I107690,I107724);
nand I_6178 (I107263,I107690,I107444);
DFFARX1 I_6179  ( .D(I107690), .CLK(I2702), .RSTB(I107283), .Q(I107772) );
not I_6180 (I107260,I107772);
DFFARX1 I_6181  ( .D(I649534), .CLK(I2702), .RSTB(I107283), .Q(I107803) );
not I_6182 (I107820,I107803);
or I_6183 (I107837,I107820,I107741);
DFFARX1 I_6184  ( .D(I107837), .CLK(I2702), .RSTB(I107283), .Q(I107266) );
nand I_6185 (I107275,I107820,I107546);
DFFARX1 I_6186  ( .D(I107820), .CLK(I2702), .RSTB(I107283), .Q(I107245) );
not I_6187 (I107929,I2709);
not I_6188 (I107946,I329181);
nor I_6189 (I107963,I329178,I329166);
nand I_6190 (I107980,I107963,I329169);
DFFARX1 I_6191  ( .D(I107980), .CLK(I2702), .RSTB(I107929), .Q(I107903) );
nor I_6192 (I108011,I107946,I329178);
nand I_6193 (I108028,I108011,I329175);
not I_6194 (I107918,I108028);
DFFARX1 I_6195  ( .D(I108028), .CLK(I2702), .RSTB(I107929), .Q(I107900) );
not I_6196 (I108073,I329178);
not I_6197 (I108090,I108073);
not I_6198 (I108107,I329187);
nor I_6199 (I108124,I108107,I329163);
and I_6200 (I108141,I108124,I329184);
or I_6201 (I108158,I108141,I329172);
DFFARX1 I_6202  ( .D(I108158), .CLK(I2702), .RSTB(I107929), .Q(I108175) );
nor I_6203 (I108192,I108175,I108028);
nor I_6204 (I108209,I108175,I108090);
nand I_6205 (I107915,I107980,I108209);
nand I_6206 (I108240,I107946,I329187);
nand I_6207 (I108257,I108240,I108175);
and I_6208 (I108274,I108240,I108257);
DFFARX1 I_6209  ( .D(I108274), .CLK(I2702), .RSTB(I107929), .Q(I107897) );
DFFARX1 I_6210  ( .D(I108240), .CLK(I2702), .RSTB(I107929), .Q(I108305) );
and I_6211 (I107894,I108073,I108305);
DFFARX1 I_6212  ( .D(I329193), .CLK(I2702), .RSTB(I107929), .Q(I108336) );
not I_6213 (I108353,I108336);
nor I_6214 (I108370,I108028,I108353);
and I_6215 (I108387,I108336,I108370);
nand I_6216 (I107909,I108336,I108090);
DFFARX1 I_6217  ( .D(I108336), .CLK(I2702), .RSTB(I107929), .Q(I108418) );
not I_6218 (I107906,I108418);
DFFARX1 I_6219  ( .D(I329190), .CLK(I2702), .RSTB(I107929), .Q(I108449) );
not I_6220 (I108466,I108449);
or I_6221 (I108483,I108466,I108387);
DFFARX1 I_6222  ( .D(I108483), .CLK(I2702), .RSTB(I107929), .Q(I107912) );
nand I_6223 (I107921,I108466,I108192);
DFFARX1 I_6224  ( .D(I108466), .CLK(I2702), .RSTB(I107929), .Q(I107891) );
not I_6225 (I108575,I2709);
not I_6226 (I108592,I181332);
nor I_6227 (I108609,I181320,I181326);
nand I_6228 (I108626,I108609,I181335);
DFFARX1 I_6229  ( .D(I108626), .CLK(I2702), .RSTB(I108575), .Q(I108549) );
nor I_6230 (I108657,I108592,I181320);
nand I_6231 (I108674,I108657,I181323);
not I_6232 (I108564,I108674);
DFFARX1 I_6233  ( .D(I108674), .CLK(I2702), .RSTB(I108575), .Q(I108546) );
not I_6234 (I108719,I181320);
not I_6235 (I108736,I108719);
not I_6236 (I108753,I181344);
nor I_6237 (I108770,I108753,I181317);
and I_6238 (I108787,I108770,I181338);
or I_6239 (I108804,I108787,I181329);
DFFARX1 I_6240  ( .D(I108804), .CLK(I2702), .RSTB(I108575), .Q(I108821) );
nor I_6241 (I108838,I108821,I108674);
nor I_6242 (I108855,I108821,I108736);
nand I_6243 (I108561,I108626,I108855);
nand I_6244 (I108886,I108592,I181344);
nand I_6245 (I108903,I108886,I108821);
and I_6246 (I108920,I108886,I108903);
DFFARX1 I_6247  ( .D(I108920), .CLK(I2702), .RSTB(I108575), .Q(I108543) );
DFFARX1 I_6248  ( .D(I108886), .CLK(I2702), .RSTB(I108575), .Q(I108951) );
and I_6249 (I108540,I108719,I108951);
DFFARX1 I_6250  ( .D(I181314), .CLK(I2702), .RSTB(I108575), .Q(I108982) );
not I_6251 (I108999,I108982);
nor I_6252 (I109016,I108674,I108999);
and I_6253 (I109033,I108982,I109016);
nand I_6254 (I108555,I108982,I108736);
DFFARX1 I_6255  ( .D(I108982), .CLK(I2702), .RSTB(I108575), .Q(I109064) );
not I_6256 (I108552,I109064);
DFFARX1 I_6257  ( .D(I181341), .CLK(I2702), .RSTB(I108575), .Q(I109095) );
not I_6258 (I109112,I109095);
or I_6259 (I109129,I109112,I109033);
DFFARX1 I_6260  ( .D(I109129), .CLK(I2702), .RSTB(I108575), .Q(I108558) );
nand I_6261 (I108567,I109112,I108838);
DFFARX1 I_6262  ( .D(I109112), .CLK(I2702), .RSTB(I108575), .Q(I108537) );
not I_6263 (I109221,I2709);
not I_6264 (I109238,I500235);
nor I_6265 (I109255,I500247,I500229);
nand I_6266 (I109272,I109255,I500238);
DFFARX1 I_6267  ( .D(I109272), .CLK(I2702), .RSTB(I109221), .Q(I109195) );
nor I_6268 (I109303,I109238,I500247);
nand I_6269 (I109320,I109303,I500244);
not I_6270 (I109210,I109320);
DFFARX1 I_6271  ( .D(I109320), .CLK(I2702), .RSTB(I109221), .Q(I109192) );
not I_6272 (I109365,I500247);
not I_6273 (I109382,I109365);
not I_6274 (I109399,I500217);
nor I_6275 (I109416,I109399,I500220);
and I_6276 (I109433,I109416,I500226);
or I_6277 (I109450,I109433,I500241);
DFFARX1 I_6278  ( .D(I109450), .CLK(I2702), .RSTB(I109221), .Q(I109467) );
nor I_6279 (I109484,I109467,I109320);
nor I_6280 (I109501,I109467,I109382);
nand I_6281 (I109207,I109272,I109501);
nand I_6282 (I109532,I109238,I500217);
nand I_6283 (I109549,I109532,I109467);
and I_6284 (I109566,I109532,I109549);
DFFARX1 I_6285  ( .D(I109566), .CLK(I2702), .RSTB(I109221), .Q(I109189) );
DFFARX1 I_6286  ( .D(I109532), .CLK(I2702), .RSTB(I109221), .Q(I109597) );
and I_6287 (I109186,I109365,I109597);
DFFARX1 I_6288  ( .D(I500223), .CLK(I2702), .RSTB(I109221), .Q(I109628) );
not I_6289 (I109645,I109628);
nor I_6290 (I109662,I109320,I109645);
and I_6291 (I109679,I109628,I109662);
nand I_6292 (I109201,I109628,I109382);
DFFARX1 I_6293  ( .D(I109628), .CLK(I2702), .RSTB(I109221), .Q(I109710) );
not I_6294 (I109198,I109710);
DFFARX1 I_6295  ( .D(I500232), .CLK(I2702), .RSTB(I109221), .Q(I109741) );
not I_6296 (I109758,I109741);
or I_6297 (I109775,I109758,I109679);
DFFARX1 I_6298  ( .D(I109775), .CLK(I2702), .RSTB(I109221), .Q(I109204) );
nand I_6299 (I109213,I109758,I109484);
DFFARX1 I_6300  ( .D(I109758), .CLK(I2702), .RSTB(I109221), .Q(I109183) );
not I_6301 (I109867,I2709);
not I_6302 (I109884,I216538);
nor I_6303 (I109901,I216568,I216547);
nand I_6304 (I109918,I109901,I216559);
DFFARX1 I_6305  ( .D(I109918), .CLK(I2702), .RSTB(I109867), .Q(I109841) );
nor I_6306 (I109949,I109884,I216568);
nand I_6307 (I109966,I109949,I216541);
not I_6308 (I109856,I109966);
DFFARX1 I_6309  ( .D(I109966), .CLK(I2702), .RSTB(I109867), .Q(I109838) );
not I_6310 (I110011,I216568);
not I_6311 (I110028,I110011);
not I_6312 (I110045,I216544);
nor I_6313 (I110062,I110045,I216562);
and I_6314 (I110079,I110062,I216553);
or I_6315 (I110096,I110079,I216550);
DFFARX1 I_6316  ( .D(I110096), .CLK(I2702), .RSTB(I109867), .Q(I110113) );
nor I_6317 (I110130,I110113,I109966);
nor I_6318 (I110147,I110113,I110028);
nand I_6319 (I109853,I109918,I110147);
nand I_6320 (I110178,I109884,I216544);
nand I_6321 (I110195,I110178,I110113);
and I_6322 (I110212,I110178,I110195);
DFFARX1 I_6323  ( .D(I110212), .CLK(I2702), .RSTB(I109867), .Q(I109835) );
DFFARX1 I_6324  ( .D(I110178), .CLK(I2702), .RSTB(I109867), .Q(I110243) );
and I_6325 (I109832,I110011,I110243);
DFFARX1 I_6326  ( .D(I216556), .CLK(I2702), .RSTB(I109867), .Q(I110274) );
not I_6327 (I110291,I110274);
nor I_6328 (I110308,I109966,I110291);
and I_6329 (I110325,I110274,I110308);
nand I_6330 (I109847,I110274,I110028);
DFFARX1 I_6331  ( .D(I110274), .CLK(I2702), .RSTB(I109867), .Q(I110356) );
not I_6332 (I109844,I110356);
DFFARX1 I_6333  ( .D(I216565), .CLK(I2702), .RSTB(I109867), .Q(I110387) );
not I_6334 (I110404,I110387);
or I_6335 (I110421,I110404,I110325);
DFFARX1 I_6336  ( .D(I110421), .CLK(I2702), .RSTB(I109867), .Q(I109850) );
nand I_6337 (I109859,I110404,I110130);
DFFARX1 I_6338  ( .D(I110404), .CLK(I2702), .RSTB(I109867), .Q(I109829) );
not I_6339 (I110513,I2709);
not I_6340 (I110530,I592304);
nor I_6341 (I110547,I592289,I592316);
nand I_6342 (I110564,I110547,I592292);
DFFARX1 I_6343  ( .D(I110564), .CLK(I2702), .RSTB(I110513), .Q(I110487) );
nor I_6344 (I110595,I110530,I592289);
nand I_6345 (I110612,I110595,I592307);
not I_6346 (I110502,I110612);
DFFARX1 I_6347  ( .D(I110612), .CLK(I2702), .RSTB(I110513), .Q(I110484) );
not I_6348 (I110657,I592289);
not I_6349 (I110674,I110657);
not I_6350 (I110691,I592319);
nor I_6351 (I110708,I110691,I592301);
and I_6352 (I110725,I110708,I592310);
or I_6353 (I110742,I110725,I592295);
DFFARX1 I_6354  ( .D(I110742), .CLK(I2702), .RSTB(I110513), .Q(I110759) );
nor I_6355 (I110776,I110759,I110612);
nor I_6356 (I110793,I110759,I110674);
nand I_6357 (I110499,I110564,I110793);
nand I_6358 (I110824,I110530,I592319);
nand I_6359 (I110841,I110824,I110759);
and I_6360 (I110858,I110824,I110841);
DFFARX1 I_6361  ( .D(I110858), .CLK(I2702), .RSTB(I110513), .Q(I110481) );
DFFARX1 I_6362  ( .D(I110824), .CLK(I2702), .RSTB(I110513), .Q(I110889) );
and I_6363 (I110478,I110657,I110889);
DFFARX1 I_6364  ( .D(I592298), .CLK(I2702), .RSTB(I110513), .Q(I110920) );
not I_6365 (I110937,I110920);
nor I_6366 (I110954,I110612,I110937);
and I_6367 (I110971,I110920,I110954);
nand I_6368 (I110493,I110920,I110674);
DFFARX1 I_6369  ( .D(I110920), .CLK(I2702), .RSTB(I110513), .Q(I111002) );
not I_6370 (I110490,I111002);
DFFARX1 I_6371  ( .D(I592313), .CLK(I2702), .RSTB(I110513), .Q(I111033) );
not I_6372 (I111050,I111033);
or I_6373 (I111067,I111050,I110971);
DFFARX1 I_6374  ( .D(I111067), .CLK(I2702), .RSTB(I110513), .Q(I110496) );
nand I_6375 (I110505,I111050,I110776);
DFFARX1 I_6376  ( .D(I111050), .CLK(I2702), .RSTB(I110513), .Q(I110475) );
not I_6377 (I111159,I2709);
not I_6378 (I111176,I619965);
nor I_6379 (I111193,I619980,I619995);
nand I_6380 (I111210,I111193,I619983);
DFFARX1 I_6381  ( .D(I111210), .CLK(I2702), .RSTB(I111159), .Q(I111133) );
nor I_6382 (I111241,I111176,I619980);
nand I_6383 (I111258,I111241,I619986);
not I_6384 (I111148,I111258);
DFFARX1 I_6385  ( .D(I111258), .CLK(I2702), .RSTB(I111159), .Q(I111130) );
not I_6386 (I111303,I619980);
not I_6387 (I111320,I111303);
not I_6388 (I111337,I619992);
nor I_6389 (I111354,I111337,I619989);
and I_6390 (I111371,I111354,I619968);
or I_6391 (I111388,I111371,I619977);
DFFARX1 I_6392  ( .D(I111388), .CLK(I2702), .RSTB(I111159), .Q(I111405) );
nor I_6393 (I111422,I111405,I111258);
nor I_6394 (I111439,I111405,I111320);
nand I_6395 (I111145,I111210,I111439);
nand I_6396 (I111470,I111176,I619992);
nand I_6397 (I111487,I111470,I111405);
and I_6398 (I111504,I111470,I111487);
DFFARX1 I_6399  ( .D(I111504), .CLK(I2702), .RSTB(I111159), .Q(I111127) );
DFFARX1 I_6400  ( .D(I111470), .CLK(I2702), .RSTB(I111159), .Q(I111535) );
and I_6401 (I111124,I111303,I111535);
DFFARX1 I_6402  ( .D(I619974), .CLK(I2702), .RSTB(I111159), .Q(I111566) );
not I_6403 (I111583,I111566);
nor I_6404 (I111600,I111258,I111583);
and I_6405 (I111617,I111566,I111600);
nand I_6406 (I111139,I111566,I111320);
DFFARX1 I_6407  ( .D(I111566), .CLK(I2702), .RSTB(I111159), .Q(I111648) );
not I_6408 (I111136,I111648);
DFFARX1 I_6409  ( .D(I619971), .CLK(I2702), .RSTB(I111159), .Q(I111679) );
not I_6410 (I111696,I111679);
or I_6411 (I111713,I111696,I111617);
DFFARX1 I_6412  ( .D(I111713), .CLK(I2702), .RSTB(I111159), .Q(I111142) );
nand I_6413 (I111151,I111696,I111422);
DFFARX1 I_6414  ( .D(I111696), .CLK(I2702), .RSTB(I111159), .Q(I111121) );
not I_6415 (I111805,I2709);
not I_6416 (I111822,I39741);
nor I_6417 (I111839,I39753,I39738);
nand I_6418 (I111856,I111839,I39750);
DFFARX1 I_6419  ( .D(I111856), .CLK(I2702), .RSTB(I111805), .Q(I111779) );
nor I_6420 (I111887,I111822,I39753);
nand I_6421 (I111904,I111887,I39768);
not I_6422 (I111794,I111904);
DFFARX1 I_6423  ( .D(I111904), .CLK(I2702), .RSTB(I111805), .Q(I111776) );
not I_6424 (I111949,I39753);
not I_6425 (I111966,I111949);
not I_6426 (I111983,I39744);
nor I_6427 (I112000,I111983,I39756);
and I_6428 (I112017,I112000,I39747);
or I_6429 (I112034,I112017,I39762);
DFFARX1 I_6430  ( .D(I112034), .CLK(I2702), .RSTB(I111805), .Q(I112051) );
nor I_6431 (I112068,I112051,I111904);
nor I_6432 (I112085,I112051,I111966);
nand I_6433 (I111791,I111856,I112085);
nand I_6434 (I112116,I111822,I39744);
nand I_6435 (I112133,I112116,I112051);
and I_6436 (I112150,I112116,I112133);
DFFARX1 I_6437  ( .D(I112150), .CLK(I2702), .RSTB(I111805), .Q(I111773) );
DFFARX1 I_6438  ( .D(I112116), .CLK(I2702), .RSTB(I111805), .Q(I112181) );
and I_6439 (I111770,I111949,I112181);
DFFARX1 I_6440  ( .D(I39765), .CLK(I2702), .RSTB(I111805), .Q(I112212) );
not I_6441 (I112229,I112212);
nor I_6442 (I112246,I111904,I112229);
and I_6443 (I112263,I112212,I112246);
nand I_6444 (I111785,I112212,I111966);
DFFARX1 I_6445  ( .D(I112212), .CLK(I2702), .RSTB(I111805), .Q(I112294) );
not I_6446 (I111782,I112294);
DFFARX1 I_6447  ( .D(I39759), .CLK(I2702), .RSTB(I111805), .Q(I112325) );
not I_6448 (I112342,I112325);
or I_6449 (I112359,I112342,I112263);
DFFARX1 I_6450  ( .D(I112359), .CLK(I2702), .RSTB(I111805), .Q(I111788) );
nand I_6451 (I111797,I112342,I112068);
DFFARX1 I_6452  ( .D(I112342), .CLK(I2702), .RSTB(I111805), .Q(I111767) );
not I_6453 (I112451,I2709);
not I_6454 (I112468,I261555);
nor I_6455 (I112485,I261552,I261540);
nand I_6456 (I112502,I112485,I261543);
DFFARX1 I_6457  ( .D(I112502), .CLK(I2702), .RSTB(I112451), .Q(I112425) );
nor I_6458 (I112533,I112468,I261552);
nand I_6459 (I112550,I112533,I261549);
not I_6460 (I112440,I112550);
DFFARX1 I_6461  ( .D(I112550), .CLK(I2702), .RSTB(I112451), .Q(I112422) );
not I_6462 (I112595,I261552);
not I_6463 (I112612,I112595);
not I_6464 (I112629,I261561);
nor I_6465 (I112646,I112629,I261537);
and I_6466 (I112663,I112646,I261558);
or I_6467 (I112680,I112663,I261546);
DFFARX1 I_6468  ( .D(I112680), .CLK(I2702), .RSTB(I112451), .Q(I112697) );
nor I_6469 (I112714,I112697,I112550);
nor I_6470 (I112731,I112697,I112612);
nand I_6471 (I112437,I112502,I112731);
nand I_6472 (I112762,I112468,I261561);
nand I_6473 (I112779,I112762,I112697);
and I_6474 (I112796,I112762,I112779);
DFFARX1 I_6475  ( .D(I112796), .CLK(I2702), .RSTB(I112451), .Q(I112419) );
DFFARX1 I_6476  ( .D(I112762), .CLK(I2702), .RSTB(I112451), .Q(I112827) );
and I_6477 (I112416,I112595,I112827);
DFFARX1 I_6478  ( .D(I261567), .CLK(I2702), .RSTB(I112451), .Q(I112858) );
not I_6479 (I112875,I112858);
nor I_6480 (I112892,I112550,I112875);
and I_6481 (I112909,I112858,I112892);
nand I_6482 (I112431,I112858,I112612);
DFFARX1 I_6483  ( .D(I112858), .CLK(I2702), .RSTB(I112451), .Q(I112940) );
not I_6484 (I112428,I112940);
DFFARX1 I_6485  ( .D(I261564), .CLK(I2702), .RSTB(I112451), .Q(I112971) );
not I_6486 (I112988,I112971);
or I_6487 (I113005,I112988,I112909);
DFFARX1 I_6488  ( .D(I113005), .CLK(I2702), .RSTB(I112451), .Q(I112434) );
nand I_6489 (I112443,I112988,I112714);
DFFARX1 I_6490  ( .D(I112988), .CLK(I2702), .RSTB(I112451), .Q(I112413) );
not I_6491 (I113097,I2709);
not I_6492 (I113114,I183984);
nor I_6493 (I113131,I183972,I183978);
nand I_6494 (I113148,I113131,I183987);
DFFARX1 I_6495  ( .D(I113148), .CLK(I2702), .RSTB(I113097), .Q(I113071) );
nor I_6496 (I113179,I113114,I183972);
nand I_6497 (I113196,I113179,I183975);
not I_6498 (I113086,I113196);
DFFARX1 I_6499  ( .D(I113196), .CLK(I2702), .RSTB(I113097), .Q(I113068) );
not I_6500 (I113241,I183972);
not I_6501 (I113258,I113241);
not I_6502 (I113275,I183996);
nor I_6503 (I113292,I113275,I183969);
and I_6504 (I113309,I113292,I183990);
or I_6505 (I113326,I113309,I183981);
DFFARX1 I_6506  ( .D(I113326), .CLK(I2702), .RSTB(I113097), .Q(I113343) );
nor I_6507 (I113360,I113343,I113196);
nor I_6508 (I113377,I113343,I113258);
nand I_6509 (I113083,I113148,I113377);
nand I_6510 (I113408,I113114,I183996);
nand I_6511 (I113425,I113408,I113343);
and I_6512 (I113442,I113408,I113425);
DFFARX1 I_6513  ( .D(I113442), .CLK(I2702), .RSTB(I113097), .Q(I113065) );
DFFARX1 I_6514  ( .D(I113408), .CLK(I2702), .RSTB(I113097), .Q(I113473) );
and I_6515 (I113062,I113241,I113473);
DFFARX1 I_6516  ( .D(I183966), .CLK(I2702), .RSTB(I113097), .Q(I113504) );
not I_6517 (I113521,I113504);
nor I_6518 (I113538,I113196,I113521);
and I_6519 (I113555,I113504,I113538);
nand I_6520 (I113077,I113504,I113258);
DFFARX1 I_6521  ( .D(I113504), .CLK(I2702), .RSTB(I113097), .Q(I113586) );
not I_6522 (I113074,I113586);
DFFARX1 I_6523  ( .D(I183993), .CLK(I2702), .RSTB(I113097), .Q(I113617) );
not I_6524 (I113634,I113617);
or I_6525 (I113651,I113634,I113555);
DFFARX1 I_6526  ( .D(I113651), .CLK(I2702), .RSTB(I113097), .Q(I113080) );
nand I_6527 (I113089,I113634,I113360);
DFFARX1 I_6528  ( .D(I113634), .CLK(I2702), .RSTB(I113097), .Q(I113059) );
not I_6529 (I113743,I2709);
not I_6530 (I113760,I400343);
nor I_6531 (I113777,I400355,I400337);
nand I_6532 (I113794,I113777,I400352);
DFFARX1 I_6533  ( .D(I113794), .CLK(I2702), .RSTB(I113743), .Q(I113717) );
nor I_6534 (I113825,I113760,I400355);
nand I_6535 (I113842,I113825,I400340);
not I_6536 (I113732,I113842);
DFFARX1 I_6537  ( .D(I113842), .CLK(I2702), .RSTB(I113743), .Q(I113714) );
not I_6538 (I113887,I400355);
not I_6539 (I113904,I113887);
not I_6540 (I113921,I400349);
nor I_6541 (I113938,I113921,I400328);
and I_6542 (I113955,I113938,I400331);
or I_6543 (I113972,I113955,I400334);
DFFARX1 I_6544  ( .D(I113972), .CLK(I2702), .RSTB(I113743), .Q(I113989) );
nor I_6545 (I114006,I113989,I113842);
nor I_6546 (I114023,I113989,I113904);
nand I_6547 (I113729,I113794,I114023);
nand I_6548 (I114054,I113760,I400349);
nand I_6549 (I114071,I114054,I113989);
and I_6550 (I114088,I114054,I114071);
DFFARX1 I_6551  ( .D(I114088), .CLK(I2702), .RSTB(I113743), .Q(I113711) );
DFFARX1 I_6552  ( .D(I114054), .CLK(I2702), .RSTB(I113743), .Q(I114119) );
and I_6553 (I113708,I113887,I114119);
DFFARX1 I_6554  ( .D(I400325), .CLK(I2702), .RSTB(I113743), .Q(I114150) );
not I_6555 (I114167,I114150);
nor I_6556 (I114184,I113842,I114167);
and I_6557 (I114201,I114150,I114184);
nand I_6558 (I113723,I114150,I113904);
DFFARX1 I_6559  ( .D(I114150), .CLK(I2702), .RSTB(I113743), .Q(I114232) );
not I_6560 (I113720,I114232);
DFFARX1 I_6561  ( .D(I400346), .CLK(I2702), .RSTB(I113743), .Q(I114263) );
not I_6562 (I114280,I114263);
or I_6563 (I114297,I114280,I114201);
DFFARX1 I_6564  ( .D(I114297), .CLK(I2702), .RSTB(I113743), .Q(I113726) );
nand I_6565 (I113735,I114280,I114006);
DFFARX1 I_6566  ( .D(I114280), .CLK(I2702), .RSTB(I113743), .Q(I113705) );
not I_6567 (I114389,I2709);
not I_6568 (I114406,I242724);
nor I_6569 (I114423,I242745,I242718);
nand I_6570 (I114440,I114423,I242733);
DFFARX1 I_6571  ( .D(I114440), .CLK(I2702), .RSTB(I114389), .Q(I114363) );
nor I_6572 (I114471,I114406,I242745);
nand I_6573 (I114488,I114471,I242748);
not I_6574 (I114378,I114488);
DFFARX1 I_6575  ( .D(I114488), .CLK(I2702), .RSTB(I114389), .Q(I114360) );
not I_6576 (I114533,I242745);
not I_6577 (I114550,I114533);
not I_6578 (I114567,I242721);
nor I_6579 (I114584,I114567,I242739);
and I_6580 (I114601,I114584,I242727);
or I_6581 (I114618,I114601,I242730);
DFFARX1 I_6582  ( .D(I114618), .CLK(I2702), .RSTB(I114389), .Q(I114635) );
nor I_6583 (I114652,I114635,I114488);
nor I_6584 (I114669,I114635,I114550);
nand I_6585 (I114375,I114440,I114669);
nand I_6586 (I114700,I114406,I242721);
nand I_6587 (I114717,I114700,I114635);
and I_6588 (I114734,I114700,I114717);
DFFARX1 I_6589  ( .D(I114734), .CLK(I2702), .RSTB(I114389), .Q(I114357) );
DFFARX1 I_6590  ( .D(I114700), .CLK(I2702), .RSTB(I114389), .Q(I114765) );
and I_6591 (I114354,I114533,I114765);
DFFARX1 I_6592  ( .D(I242742), .CLK(I2702), .RSTB(I114389), .Q(I114796) );
not I_6593 (I114813,I114796);
nor I_6594 (I114830,I114488,I114813);
and I_6595 (I114847,I114796,I114830);
nand I_6596 (I114369,I114796,I114550);
DFFARX1 I_6597  ( .D(I114796), .CLK(I2702), .RSTB(I114389), .Q(I114878) );
not I_6598 (I114366,I114878);
DFFARX1 I_6599  ( .D(I242736), .CLK(I2702), .RSTB(I114389), .Q(I114909) );
not I_6600 (I114926,I114909);
or I_6601 (I114943,I114926,I114847);
DFFARX1 I_6602  ( .D(I114943), .CLK(I2702), .RSTB(I114389), .Q(I114372) );
nand I_6603 (I114381,I114926,I114652);
DFFARX1 I_6604  ( .D(I114926), .CLK(I2702), .RSTB(I114389), .Q(I114351) );
not I_6605 (I115035,I2709);
not I_6606 (I115052,I565541);
nor I_6607 (I115069,I565517,I565523);
nand I_6608 (I115086,I115069,I565526);
DFFARX1 I_6609  ( .D(I115086), .CLK(I2702), .RSTB(I115035), .Q(I115009) );
nor I_6610 (I115117,I115052,I565517);
nand I_6611 (I115134,I115117,I565535);
not I_6612 (I115024,I115134);
DFFARX1 I_6613  ( .D(I115134), .CLK(I2702), .RSTB(I115035), .Q(I115006) );
not I_6614 (I115179,I565517);
not I_6615 (I115196,I115179);
not I_6616 (I115213,I565514);
nor I_6617 (I115230,I115213,I565529);
and I_6618 (I115247,I115230,I565520);
or I_6619 (I115264,I115247,I565532);
DFFARX1 I_6620  ( .D(I115264), .CLK(I2702), .RSTB(I115035), .Q(I115281) );
nor I_6621 (I115298,I115281,I115134);
nor I_6622 (I115315,I115281,I115196);
nand I_6623 (I115021,I115086,I115315);
nand I_6624 (I115346,I115052,I565514);
nand I_6625 (I115363,I115346,I115281);
and I_6626 (I115380,I115346,I115363);
DFFARX1 I_6627  ( .D(I115380), .CLK(I2702), .RSTB(I115035), .Q(I115003) );
DFFARX1 I_6628  ( .D(I115346), .CLK(I2702), .RSTB(I115035), .Q(I115411) );
and I_6629 (I115000,I115179,I115411);
DFFARX1 I_6630  ( .D(I565544), .CLK(I2702), .RSTB(I115035), .Q(I115442) );
not I_6631 (I115459,I115442);
nor I_6632 (I115476,I115134,I115459);
and I_6633 (I115493,I115442,I115476);
nand I_6634 (I115015,I115442,I115196);
DFFARX1 I_6635  ( .D(I115442), .CLK(I2702), .RSTB(I115035), .Q(I115524) );
not I_6636 (I115012,I115524);
DFFARX1 I_6637  ( .D(I565538), .CLK(I2702), .RSTB(I115035), .Q(I115555) );
not I_6638 (I115572,I115555);
or I_6639 (I115589,I115572,I115493);
DFFARX1 I_6640  ( .D(I115589), .CLK(I2702), .RSTB(I115035), .Q(I115018) );
nand I_6641 (I115027,I115572,I115298);
DFFARX1 I_6642  ( .D(I115572), .CLK(I2702), .RSTB(I115035), .Q(I114997) );
not I_6643 (I115681,I2709);
not I_6644 (I115698,I438488);
nor I_6645 (I115715,I438476,I438482);
nand I_6646 (I115732,I115715,I438473);
DFFARX1 I_6647  ( .D(I115732), .CLK(I2702), .RSTB(I115681), .Q(I115655) );
nor I_6648 (I115763,I115698,I438476);
nand I_6649 (I115780,I115763,I438479);
not I_6650 (I115670,I115780);
DFFARX1 I_6651  ( .D(I115780), .CLK(I2702), .RSTB(I115681), .Q(I115652) );
not I_6652 (I115825,I438476);
not I_6653 (I115842,I115825);
not I_6654 (I115859,I438491);
nor I_6655 (I115876,I115859,I438503);
and I_6656 (I115893,I115876,I438485);
or I_6657 (I115910,I115893,I438500);
DFFARX1 I_6658  ( .D(I115910), .CLK(I2702), .RSTB(I115681), .Q(I115927) );
nor I_6659 (I115944,I115927,I115780);
nor I_6660 (I115961,I115927,I115842);
nand I_6661 (I115667,I115732,I115961);
nand I_6662 (I115992,I115698,I438491);
nand I_6663 (I116009,I115992,I115927);
and I_6664 (I116026,I115992,I116009);
DFFARX1 I_6665  ( .D(I116026), .CLK(I2702), .RSTB(I115681), .Q(I115649) );
DFFARX1 I_6666  ( .D(I115992), .CLK(I2702), .RSTB(I115681), .Q(I116057) );
and I_6667 (I115646,I115825,I116057);
DFFARX1 I_6668  ( .D(I438494), .CLK(I2702), .RSTB(I115681), .Q(I116088) );
not I_6669 (I116105,I116088);
nor I_6670 (I116122,I115780,I116105);
and I_6671 (I116139,I116088,I116122);
nand I_6672 (I115661,I116088,I115842);
DFFARX1 I_6673  ( .D(I116088), .CLK(I2702), .RSTB(I115681), .Q(I116170) );
not I_6674 (I115658,I116170);
DFFARX1 I_6675  ( .D(I438497), .CLK(I2702), .RSTB(I115681), .Q(I116201) );
not I_6676 (I116218,I116201);
or I_6677 (I116235,I116218,I116139);
DFFARX1 I_6678  ( .D(I116235), .CLK(I2702), .RSTB(I115681), .Q(I115664) );
nand I_6679 (I115673,I116218,I115944);
DFFARX1 I_6680  ( .D(I116218), .CLK(I2702), .RSTB(I115681), .Q(I115643) );
not I_6681 (I116327,I2709);
not I_6682 (I116344,I360291);
nor I_6683 (I116361,I360303,I360285);
nand I_6684 (I116378,I116361,I360300);
DFFARX1 I_6685  ( .D(I116378), .CLK(I2702), .RSTB(I116327), .Q(I116301) );
nor I_6686 (I116409,I116344,I360303);
nand I_6687 (I116426,I116409,I360288);
not I_6688 (I116316,I116426);
DFFARX1 I_6689  ( .D(I116426), .CLK(I2702), .RSTB(I116327), .Q(I116298) );
not I_6690 (I116471,I360303);
not I_6691 (I116488,I116471);
not I_6692 (I116505,I360297);
nor I_6693 (I116522,I116505,I360276);
and I_6694 (I116539,I116522,I360279);
or I_6695 (I116556,I116539,I360282);
DFFARX1 I_6696  ( .D(I116556), .CLK(I2702), .RSTB(I116327), .Q(I116573) );
nor I_6697 (I116590,I116573,I116426);
nor I_6698 (I116607,I116573,I116488);
nand I_6699 (I116313,I116378,I116607);
nand I_6700 (I116638,I116344,I360297);
nand I_6701 (I116655,I116638,I116573);
and I_6702 (I116672,I116638,I116655);
DFFARX1 I_6703  ( .D(I116672), .CLK(I2702), .RSTB(I116327), .Q(I116295) );
DFFARX1 I_6704  ( .D(I116638), .CLK(I2702), .RSTB(I116327), .Q(I116703) );
and I_6705 (I116292,I116471,I116703);
DFFARX1 I_6706  ( .D(I360273), .CLK(I2702), .RSTB(I116327), .Q(I116734) );
not I_6707 (I116751,I116734);
nor I_6708 (I116768,I116426,I116751);
and I_6709 (I116785,I116734,I116768);
nand I_6710 (I116307,I116734,I116488);
DFFARX1 I_6711  ( .D(I116734), .CLK(I2702), .RSTB(I116327), .Q(I116816) );
not I_6712 (I116304,I116816);
DFFARX1 I_6713  ( .D(I360294), .CLK(I2702), .RSTB(I116327), .Q(I116847) );
not I_6714 (I116864,I116847);
or I_6715 (I116881,I116864,I116785);
DFFARX1 I_6716  ( .D(I116881), .CLK(I2702), .RSTB(I116327), .Q(I116310) );
nand I_6717 (I116319,I116864,I116590);
DFFARX1 I_6718  ( .D(I116864), .CLK(I2702), .RSTB(I116327), .Q(I116289) );
not I_6719 (I116973,I2709);
not I_6720 (I116990,I375149);
nor I_6721 (I117007,I375161,I375143);
nand I_6722 (I117024,I117007,I375158);
DFFARX1 I_6723  ( .D(I117024), .CLK(I2702), .RSTB(I116973), .Q(I116947) );
nor I_6724 (I117055,I116990,I375161);
nand I_6725 (I117072,I117055,I375146);
not I_6726 (I116962,I117072);
DFFARX1 I_6727  ( .D(I117072), .CLK(I2702), .RSTB(I116973), .Q(I116944) );
not I_6728 (I117117,I375161);
not I_6729 (I117134,I117117);
not I_6730 (I117151,I375155);
nor I_6731 (I117168,I117151,I375134);
and I_6732 (I117185,I117168,I375137);
or I_6733 (I117202,I117185,I375140);
DFFARX1 I_6734  ( .D(I117202), .CLK(I2702), .RSTB(I116973), .Q(I117219) );
nor I_6735 (I117236,I117219,I117072);
nor I_6736 (I117253,I117219,I117134);
nand I_6737 (I116959,I117024,I117253);
nand I_6738 (I117284,I116990,I375155);
nand I_6739 (I117301,I117284,I117219);
and I_6740 (I117318,I117284,I117301);
DFFARX1 I_6741  ( .D(I117318), .CLK(I2702), .RSTB(I116973), .Q(I116941) );
DFFARX1 I_6742  ( .D(I117284), .CLK(I2702), .RSTB(I116973), .Q(I117349) );
and I_6743 (I116938,I117117,I117349);
DFFARX1 I_6744  ( .D(I375131), .CLK(I2702), .RSTB(I116973), .Q(I117380) );
not I_6745 (I117397,I117380);
nor I_6746 (I117414,I117072,I117397);
and I_6747 (I117431,I117380,I117414);
nand I_6748 (I116953,I117380,I117134);
DFFARX1 I_6749  ( .D(I117380), .CLK(I2702), .RSTB(I116973), .Q(I117462) );
not I_6750 (I116950,I117462);
DFFARX1 I_6751  ( .D(I375152), .CLK(I2702), .RSTB(I116973), .Q(I117493) );
not I_6752 (I117510,I117493);
or I_6753 (I117527,I117510,I117431);
DFFARX1 I_6754  ( .D(I117527), .CLK(I2702), .RSTB(I116973), .Q(I116956) );
nand I_6755 (I116965,I117510,I117236);
DFFARX1 I_6756  ( .D(I117510), .CLK(I2702), .RSTB(I116973), .Q(I116935) );
not I_6757 (I117619,I2709);
not I_6758 (I117636,I512586);
nor I_6759 (I117653,I512562,I512568);
nand I_6760 (I117670,I117653,I512571);
DFFARX1 I_6761  ( .D(I117670), .CLK(I2702), .RSTB(I117619), .Q(I117593) );
nor I_6762 (I117701,I117636,I512562);
nand I_6763 (I117718,I117701,I512580);
not I_6764 (I117608,I117718);
DFFARX1 I_6765  ( .D(I117718), .CLK(I2702), .RSTB(I117619), .Q(I117590) );
not I_6766 (I117763,I512562);
not I_6767 (I117780,I117763);
not I_6768 (I117797,I512559);
nor I_6769 (I117814,I117797,I512574);
and I_6770 (I117831,I117814,I512565);
or I_6771 (I117848,I117831,I512577);
DFFARX1 I_6772  ( .D(I117848), .CLK(I2702), .RSTB(I117619), .Q(I117865) );
nor I_6773 (I117882,I117865,I117718);
nor I_6774 (I117899,I117865,I117780);
nand I_6775 (I117605,I117670,I117899);
nand I_6776 (I117930,I117636,I512559);
nand I_6777 (I117947,I117930,I117865);
and I_6778 (I117964,I117930,I117947);
DFFARX1 I_6779  ( .D(I117964), .CLK(I2702), .RSTB(I117619), .Q(I117587) );
DFFARX1 I_6780  ( .D(I117930), .CLK(I2702), .RSTB(I117619), .Q(I117995) );
and I_6781 (I117584,I117763,I117995);
DFFARX1 I_6782  ( .D(I512589), .CLK(I2702), .RSTB(I117619), .Q(I118026) );
not I_6783 (I118043,I118026);
nor I_6784 (I118060,I117718,I118043);
and I_6785 (I118077,I118026,I118060);
nand I_6786 (I117599,I118026,I117780);
DFFARX1 I_6787  ( .D(I118026), .CLK(I2702), .RSTB(I117619), .Q(I118108) );
not I_6788 (I117596,I118108);
DFFARX1 I_6789  ( .D(I512583), .CLK(I2702), .RSTB(I117619), .Q(I118139) );
not I_6790 (I118156,I118139);
or I_6791 (I118173,I118156,I118077);
DFFARX1 I_6792  ( .D(I118173), .CLK(I2702), .RSTB(I117619), .Q(I117602) );
nand I_6793 (I117611,I118156,I117882);
DFFARX1 I_6794  ( .D(I118156), .CLK(I2702), .RSTB(I117619), .Q(I117581) );
not I_6795 (I118265,I2709);
not I_6796 (I118282,I49839);
nor I_6797 (I118299,I49851,I49836);
nand I_6798 (I118316,I118299,I49848);
DFFARX1 I_6799  ( .D(I118316), .CLK(I2702), .RSTB(I118265), .Q(I118239) );
nor I_6800 (I118347,I118282,I49851);
nand I_6801 (I118364,I118347,I49866);
not I_6802 (I118254,I118364);
DFFARX1 I_6803  ( .D(I118364), .CLK(I2702), .RSTB(I118265), .Q(I118236) );
not I_6804 (I118409,I49851);
not I_6805 (I118426,I118409);
not I_6806 (I118443,I49842);
nor I_6807 (I118460,I118443,I49854);
and I_6808 (I118477,I118460,I49845);
or I_6809 (I118494,I118477,I49860);
DFFARX1 I_6810  ( .D(I118494), .CLK(I2702), .RSTB(I118265), .Q(I118511) );
nor I_6811 (I118528,I118511,I118364);
nor I_6812 (I118545,I118511,I118426);
nand I_6813 (I118251,I118316,I118545);
nand I_6814 (I118576,I118282,I49842);
nand I_6815 (I118593,I118576,I118511);
and I_6816 (I118610,I118576,I118593);
DFFARX1 I_6817  ( .D(I118610), .CLK(I2702), .RSTB(I118265), .Q(I118233) );
DFFARX1 I_6818  ( .D(I118576), .CLK(I2702), .RSTB(I118265), .Q(I118641) );
and I_6819 (I118230,I118409,I118641);
DFFARX1 I_6820  ( .D(I49863), .CLK(I2702), .RSTB(I118265), .Q(I118672) );
not I_6821 (I118689,I118672);
nor I_6822 (I118706,I118364,I118689);
and I_6823 (I118723,I118672,I118706);
nand I_6824 (I118245,I118672,I118426);
DFFARX1 I_6825  ( .D(I118672), .CLK(I2702), .RSTB(I118265), .Q(I118754) );
not I_6826 (I118242,I118754);
DFFARX1 I_6827  ( .D(I49857), .CLK(I2702), .RSTB(I118265), .Q(I118785) );
not I_6828 (I118802,I118785);
or I_6829 (I118819,I118802,I118723);
DFFARX1 I_6830  ( .D(I118819), .CLK(I2702), .RSTB(I118265), .Q(I118248) );
nand I_6831 (I118257,I118802,I118528);
DFFARX1 I_6832  ( .D(I118802), .CLK(I2702), .RSTB(I118265), .Q(I118227) );
not I_6833 (I118911,I2709);
not I_6834 (I118928,I665882);
nor I_6835 (I118945,I665897,I665912);
nand I_6836 (I118962,I118945,I665900);
DFFARX1 I_6837  ( .D(I118962), .CLK(I2702), .RSTB(I118911), .Q(I118885) );
nor I_6838 (I118993,I118928,I665897);
nand I_6839 (I119010,I118993,I665903);
not I_6840 (I118900,I119010);
DFFARX1 I_6841  ( .D(I119010), .CLK(I2702), .RSTB(I118911), .Q(I118882) );
not I_6842 (I119055,I665897);
not I_6843 (I119072,I119055);
not I_6844 (I119089,I665909);
nor I_6845 (I119106,I119089,I665906);
and I_6846 (I119123,I119106,I665885);
or I_6847 (I119140,I119123,I665894);
DFFARX1 I_6848  ( .D(I119140), .CLK(I2702), .RSTB(I118911), .Q(I119157) );
nor I_6849 (I119174,I119157,I119010);
nor I_6850 (I119191,I119157,I119072);
nand I_6851 (I118897,I118962,I119191);
nand I_6852 (I119222,I118928,I665909);
nand I_6853 (I119239,I119222,I119157);
and I_6854 (I119256,I119222,I119239);
DFFARX1 I_6855  ( .D(I119256), .CLK(I2702), .RSTB(I118911), .Q(I118879) );
DFFARX1 I_6856  ( .D(I119222), .CLK(I2702), .RSTB(I118911), .Q(I119287) );
and I_6857 (I118876,I119055,I119287);
DFFARX1 I_6858  ( .D(I665891), .CLK(I2702), .RSTB(I118911), .Q(I119318) );
not I_6859 (I119335,I119318);
nor I_6860 (I119352,I119010,I119335);
and I_6861 (I119369,I119318,I119352);
nand I_6862 (I118891,I119318,I119072);
DFFARX1 I_6863  ( .D(I119318), .CLK(I2702), .RSTB(I118911), .Q(I119400) );
not I_6864 (I118888,I119400);
DFFARX1 I_6865  ( .D(I665888), .CLK(I2702), .RSTB(I118911), .Q(I119431) );
not I_6866 (I119448,I119431);
or I_6867 (I119465,I119448,I119369);
DFFARX1 I_6868  ( .D(I119465), .CLK(I2702), .RSTB(I118911), .Q(I118894) );
nand I_6869 (I118903,I119448,I119174);
DFFARX1 I_6870  ( .D(I119448), .CLK(I2702), .RSTB(I118911), .Q(I118873) );
not I_6871 (I119557,I2709);
not I_6872 (I119574,I152160);
nor I_6873 (I119591,I152148,I152154);
nand I_6874 (I119608,I119591,I152163);
DFFARX1 I_6875  ( .D(I119608), .CLK(I2702), .RSTB(I119557), .Q(I119531) );
nor I_6876 (I119639,I119574,I152148);
nand I_6877 (I119656,I119639,I152151);
not I_6878 (I119546,I119656);
DFFARX1 I_6879  ( .D(I119656), .CLK(I2702), .RSTB(I119557), .Q(I119528) );
not I_6880 (I119701,I152148);
not I_6881 (I119718,I119701);
not I_6882 (I119735,I152172);
nor I_6883 (I119752,I119735,I152145);
and I_6884 (I119769,I119752,I152166);
or I_6885 (I119786,I119769,I152157);
DFFARX1 I_6886  ( .D(I119786), .CLK(I2702), .RSTB(I119557), .Q(I119803) );
nor I_6887 (I119820,I119803,I119656);
nor I_6888 (I119837,I119803,I119718);
nand I_6889 (I119543,I119608,I119837);
nand I_6890 (I119868,I119574,I152172);
nand I_6891 (I119885,I119868,I119803);
and I_6892 (I119902,I119868,I119885);
DFFARX1 I_6893  ( .D(I119902), .CLK(I2702), .RSTB(I119557), .Q(I119525) );
DFFARX1 I_6894  ( .D(I119868), .CLK(I2702), .RSTB(I119557), .Q(I119933) );
and I_6895 (I119522,I119701,I119933);
DFFARX1 I_6896  ( .D(I152142), .CLK(I2702), .RSTB(I119557), .Q(I119964) );
not I_6897 (I119981,I119964);
nor I_6898 (I119998,I119656,I119981);
and I_6899 (I120015,I119964,I119998);
nand I_6900 (I119537,I119964,I119718);
DFFARX1 I_6901  ( .D(I119964), .CLK(I2702), .RSTB(I119557), .Q(I120046) );
not I_6902 (I119534,I120046);
DFFARX1 I_6903  ( .D(I152169), .CLK(I2702), .RSTB(I119557), .Q(I120077) );
not I_6904 (I120094,I120077);
or I_6905 (I120111,I120094,I120015);
DFFARX1 I_6906  ( .D(I120111), .CLK(I2702), .RSTB(I119557), .Q(I119540) );
nand I_6907 (I119549,I120094,I119820);
DFFARX1 I_6908  ( .D(I120094), .CLK(I2702), .RSTB(I119557), .Q(I119519) );
not I_6909 (I120203,I2709);
not I_6910 (I120220,I358353);
nor I_6911 (I120237,I358365,I358347);
nand I_6912 (I120254,I120237,I358362);
DFFARX1 I_6913  ( .D(I120254), .CLK(I2702), .RSTB(I120203), .Q(I120177) );
nor I_6914 (I120285,I120220,I358365);
nand I_6915 (I120302,I120285,I358350);
not I_6916 (I120192,I120302);
DFFARX1 I_6917  ( .D(I120302), .CLK(I2702), .RSTB(I120203), .Q(I120174) );
not I_6918 (I120347,I358365);
not I_6919 (I120364,I120347);
not I_6920 (I120381,I358359);
nor I_6921 (I120398,I120381,I358338);
and I_6922 (I120415,I120398,I358341);
or I_6923 (I120432,I120415,I358344);
DFFARX1 I_6924  ( .D(I120432), .CLK(I2702), .RSTB(I120203), .Q(I120449) );
nor I_6925 (I120466,I120449,I120302);
nor I_6926 (I120483,I120449,I120364);
nand I_6927 (I120189,I120254,I120483);
nand I_6928 (I120514,I120220,I358359);
nand I_6929 (I120531,I120514,I120449);
and I_6930 (I120548,I120514,I120531);
DFFARX1 I_6931  ( .D(I120548), .CLK(I2702), .RSTB(I120203), .Q(I120171) );
DFFARX1 I_6932  ( .D(I120514), .CLK(I2702), .RSTB(I120203), .Q(I120579) );
and I_6933 (I120168,I120347,I120579);
DFFARX1 I_6934  ( .D(I358335), .CLK(I2702), .RSTB(I120203), .Q(I120610) );
not I_6935 (I120627,I120610);
nor I_6936 (I120644,I120302,I120627);
and I_6937 (I120661,I120610,I120644);
nand I_6938 (I120183,I120610,I120364);
DFFARX1 I_6939  ( .D(I120610), .CLK(I2702), .RSTB(I120203), .Q(I120692) );
not I_6940 (I120180,I120692);
DFFARX1 I_6941  ( .D(I358356), .CLK(I2702), .RSTB(I120203), .Q(I120723) );
not I_6942 (I120740,I120723);
or I_6943 (I120757,I120740,I120661);
DFFARX1 I_6944  ( .D(I120757), .CLK(I2702), .RSTB(I120203), .Q(I120186) );
nand I_6945 (I120195,I120740,I120466);
DFFARX1 I_6946  ( .D(I120740), .CLK(I2702), .RSTB(I120203), .Q(I120165) );
not I_6947 (I120849,I2709);
not I_6948 (I120866,I607774);
nor I_6949 (I120883,I607759,I607786);
nand I_6950 (I120900,I120883,I607762);
DFFARX1 I_6951  ( .D(I120900), .CLK(I2702), .RSTB(I120849), .Q(I120823) );
nor I_6952 (I120931,I120866,I607759);
nand I_6953 (I120948,I120931,I607777);
not I_6954 (I120838,I120948);
DFFARX1 I_6955  ( .D(I120948), .CLK(I2702), .RSTB(I120849), .Q(I120820) );
not I_6956 (I120993,I607759);
not I_6957 (I121010,I120993);
not I_6958 (I121027,I607789);
nor I_6959 (I121044,I121027,I607771);
and I_6960 (I121061,I121044,I607780);
or I_6961 (I121078,I121061,I607765);
DFFARX1 I_6962  ( .D(I121078), .CLK(I2702), .RSTB(I120849), .Q(I121095) );
nor I_6963 (I121112,I121095,I120948);
nor I_6964 (I121129,I121095,I121010);
nand I_6965 (I120835,I120900,I121129);
nand I_6966 (I121160,I120866,I607789);
nand I_6967 (I121177,I121160,I121095);
and I_6968 (I121194,I121160,I121177);
DFFARX1 I_6969  ( .D(I121194), .CLK(I2702), .RSTB(I120849), .Q(I120817) );
DFFARX1 I_6970  ( .D(I121160), .CLK(I2702), .RSTB(I120849), .Q(I121225) );
and I_6971 (I120814,I120993,I121225);
DFFARX1 I_6972  ( .D(I607768), .CLK(I2702), .RSTB(I120849), .Q(I121256) );
not I_6973 (I121273,I121256);
nor I_6974 (I121290,I120948,I121273);
and I_6975 (I121307,I121256,I121290);
nand I_6976 (I120829,I121256,I121010);
DFFARX1 I_6977  ( .D(I121256), .CLK(I2702), .RSTB(I120849), .Q(I121338) );
not I_6978 (I120826,I121338);
DFFARX1 I_6979  ( .D(I607783), .CLK(I2702), .RSTB(I120849), .Q(I121369) );
not I_6980 (I121386,I121369);
or I_6981 (I121403,I121386,I121307);
DFFARX1 I_6982  ( .D(I121403), .CLK(I2702), .RSTB(I120849), .Q(I120832) );
nand I_6983 (I120841,I121386,I121112);
DFFARX1 I_6984  ( .D(I121386), .CLK(I2702), .RSTB(I120849), .Q(I120811) );
not I_6985 (I121495,I2709);
not I_6986 (I121512,I339619);
nor I_6987 (I121529,I339631,I339613);
nand I_6988 (I121546,I121529,I339628);
DFFARX1 I_6989  ( .D(I121546), .CLK(I2702), .RSTB(I121495), .Q(I121469) );
nor I_6990 (I121577,I121512,I339631);
nand I_6991 (I121594,I121577,I339616);
not I_6992 (I121484,I121594);
DFFARX1 I_6993  ( .D(I121594), .CLK(I2702), .RSTB(I121495), .Q(I121466) );
not I_6994 (I121639,I339631);
not I_6995 (I121656,I121639);
not I_6996 (I121673,I339625);
nor I_6997 (I121690,I121673,I339604);
and I_6998 (I121707,I121690,I339607);
or I_6999 (I121724,I121707,I339610);
DFFARX1 I_7000  ( .D(I121724), .CLK(I2702), .RSTB(I121495), .Q(I121741) );
nor I_7001 (I121758,I121741,I121594);
nor I_7002 (I121775,I121741,I121656);
nand I_7003 (I121481,I121546,I121775);
nand I_7004 (I121806,I121512,I339625);
nand I_7005 (I121823,I121806,I121741);
and I_7006 (I121840,I121806,I121823);
DFFARX1 I_7007  ( .D(I121840), .CLK(I2702), .RSTB(I121495), .Q(I121463) );
DFFARX1 I_7008  ( .D(I121806), .CLK(I2702), .RSTB(I121495), .Q(I121871) );
and I_7009 (I121460,I121639,I121871);
DFFARX1 I_7010  ( .D(I339601), .CLK(I2702), .RSTB(I121495), .Q(I121902) );
not I_7011 (I121919,I121902);
nor I_7012 (I121936,I121594,I121919);
and I_7013 (I121953,I121902,I121936);
nand I_7014 (I121475,I121902,I121656);
DFFARX1 I_7015  ( .D(I121902), .CLK(I2702), .RSTB(I121495), .Q(I121984) );
not I_7016 (I121472,I121984);
DFFARX1 I_7017  ( .D(I339622), .CLK(I2702), .RSTB(I121495), .Q(I122015) );
not I_7018 (I122032,I122015);
or I_7019 (I122049,I122032,I121953);
DFFARX1 I_7020  ( .D(I122049), .CLK(I2702), .RSTB(I121495), .Q(I121478) );
nand I_7021 (I121487,I122032,I121758);
DFFARX1 I_7022  ( .D(I122032), .CLK(I2702), .RSTB(I121495), .Q(I121457) );
not I_7023 (I122141,I2709);
not I_7024 (I122158,I2715);
nor I_7025 (I122175,I2727,I2712);
nand I_7026 (I122192,I122175,I2724);
DFFARX1 I_7027  ( .D(I122192), .CLK(I2702), .RSTB(I122141), .Q(I122115) );
nor I_7028 (I122223,I122158,I2727);
nand I_7029 (I122240,I122223,I2742);
not I_7030 (I122130,I122240);
DFFARX1 I_7031  ( .D(I122240), .CLK(I2702), .RSTB(I122141), .Q(I122112) );
not I_7032 (I122285,I2727);
not I_7033 (I122302,I122285);
not I_7034 (I122319,I2718);
nor I_7035 (I122336,I122319,I2730);
and I_7036 (I122353,I122336,I2721);
or I_7037 (I122370,I122353,I2736);
DFFARX1 I_7038  ( .D(I122370), .CLK(I2702), .RSTB(I122141), .Q(I122387) );
nor I_7039 (I122404,I122387,I122240);
nor I_7040 (I122421,I122387,I122302);
nand I_7041 (I122127,I122192,I122421);
nand I_7042 (I122452,I122158,I2718);
nand I_7043 (I122469,I122452,I122387);
and I_7044 (I122486,I122452,I122469);
DFFARX1 I_7045  ( .D(I122486), .CLK(I2702), .RSTB(I122141), .Q(I122109) );
DFFARX1 I_7046  ( .D(I122452), .CLK(I2702), .RSTB(I122141), .Q(I122517) );
and I_7047 (I122106,I122285,I122517);
DFFARX1 I_7048  ( .D(I2739), .CLK(I2702), .RSTB(I122141), .Q(I122548) );
not I_7049 (I122565,I122548);
nor I_7050 (I122582,I122240,I122565);
and I_7051 (I122599,I122548,I122582);
nand I_7052 (I122121,I122548,I122302);
DFFARX1 I_7053  ( .D(I122548), .CLK(I2702), .RSTB(I122141), .Q(I122630) );
not I_7054 (I122118,I122630);
DFFARX1 I_7055  ( .D(I2733), .CLK(I2702), .RSTB(I122141), .Q(I122661) );
not I_7056 (I122678,I122661);
or I_7057 (I122695,I122678,I122599);
DFFARX1 I_7058  ( .D(I122695), .CLK(I2702), .RSTB(I122141), .Q(I122124) );
nand I_7059 (I122133,I122678,I122404);
DFFARX1 I_7060  ( .D(I122678), .CLK(I2702), .RSTB(I122141), .Q(I122103) );
not I_7061 (I122787,I2709);
not I_7062 (I122804,I432130);
nor I_7063 (I122821,I432118,I432124);
nand I_7064 (I122838,I122821,I432115);
DFFARX1 I_7065  ( .D(I122838), .CLK(I2702), .RSTB(I122787), .Q(I122761) );
nor I_7066 (I122869,I122804,I432118);
nand I_7067 (I122886,I122869,I432121);
not I_7068 (I122776,I122886);
DFFARX1 I_7069  ( .D(I122886), .CLK(I2702), .RSTB(I122787), .Q(I122758) );
not I_7070 (I122931,I432118);
not I_7071 (I122948,I122931);
not I_7072 (I122965,I432133);
nor I_7073 (I122982,I122965,I432145);
and I_7074 (I122999,I122982,I432127);
or I_7075 (I123016,I122999,I432142);
DFFARX1 I_7076  ( .D(I123016), .CLK(I2702), .RSTB(I122787), .Q(I123033) );
nor I_7077 (I123050,I123033,I122886);
nor I_7078 (I123067,I123033,I122948);
nand I_7079 (I122773,I122838,I123067);
nand I_7080 (I123098,I122804,I432133);
nand I_7081 (I123115,I123098,I123033);
and I_7082 (I123132,I123098,I123115);
DFFARX1 I_7083  ( .D(I123132), .CLK(I2702), .RSTB(I122787), .Q(I122755) );
DFFARX1 I_7084  ( .D(I123098), .CLK(I2702), .RSTB(I122787), .Q(I123163) );
and I_7085 (I122752,I122931,I123163);
DFFARX1 I_7086  ( .D(I432136), .CLK(I2702), .RSTB(I122787), .Q(I123194) );
not I_7087 (I123211,I123194);
nor I_7088 (I123228,I122886,I123211);
and I_7089 (I123245,I123194,I123228);
nand I_7090 (I122767,I123194,I122948);
DFFARX1 I_7091  ( .D(I123194), .CLK(I2702), .RSTB(I122787), .Q(I123276) );
not I_7092 (I122764,I123276);
DFFARX1 I_7093  ( .D(I432139), .CLK(I2702), .RSTB(I122787), .Q(I123307) );
not I_7094 (I123324,I123307);
or I_7095 (I123341,I123324,I123245);
DFFARX1 I_7096  ( .D(I123341), .CLK(I2702), .RSTB(I122787), .Q(I122770) );
nand I_7097 (I122779,I123324,I123050);
DFFARX1 I_7098  ( .D(I123324), .CLK(I2702), .RSTB(I122787), .Q(I122749) );
not I_7099 (I123433,I2709);
not I_7100 (I123450,I290064);
nor I_7101 (I123467,I290061,I290049);
nand I_7102 (I123484,I123467,I290052);
DFFARX1 I_7103  ( .D(I123484), .CLK(I2702), .RSTB(I123433), .Q(I123407) );
nor I_7104 (I123515,I123450,I290061);
nand I_7105 (I123532,I123515,I290058);
not I_7106 (I123422,I123532);
DFFARX1 I_7107  ( .D(I123532), .CLK(I2702), .RSTB(I123433), .Q(I123404) );
not I_7108 (I123577,I290061);
not I_7109 (I123594,I123577);
not I_7110 (I123611,I290070);
nor I_7111 (I123628,I123611,I290046);
and I_7112 (I123645,I123628,I290067);
or I_7113 (I123662,I123645,I290055);
DFFARX1 I_7114  ( .D(I123662), .CLK(I2702), .RSTB(I123433), .Q(I123679) );
nor I_7115 (I123696,I123679,I123532);
nor I_7116 (I123713,I123679,I123594);
nand I_7117 (I123419,I123484,I123713);
nand I_7118 (I123744,I123450,I290070);
nand I_7119 (I123761,I123744,I123679);
and I_7120 (I123778,I123744,I123761);
DFFARX1 I_7121  ( .D(I123778), .CLK(I2702), .RSTB(I123433), .Q(I123401) );
DFFARX1 I_7122  ( .D(I123744), .CLK(I2702), .RSTB(I123433), .Q(I123809) );
and I_7123 (I123398,I123577,I123809);
DFFARX1 I_7124  ( .D(I290076), .CLK(I2702), .RSTB(I123433), .Q(I123840) );
not I_7125 (I123857,I123840);
nor I_7126 (I123874,I123532,I123857);
and I_7127 (I123891,I123840,I123874);
nand I_7128 (I123413,I123840,I123594);
DFFARX1 I_7129  ( .D(I123840), .CLK(I2702), .RSTB(I123433), .Q(I123922) );
not I_7130 (I123410,I123922);
DFFARX1 I_7131  ( .D(I290073), .CLK(I2702), .RSTB(I123433), .Q(I123953) );
not I_7132 (I123970,I123953);
or I_7133 (I123987,I123970,I123891);
DFFARX1 I_7134  ( .D(I123987), .CLK(I2702), .RSTB(I123433), .Q(I123416) );
nand I_7135 (I123425,I123970,I123696);
DFFARX1 I_7136  ( .D(I123970), .CLK(I2702), .RSTB(I123433), .Q(I123395) );
not I_7137 (I124079,I2709);
not I_7138 (I124096,I162105);
nor I_7139 (I124113,I162093,I162099);
nand I_7140 (I124130,I124113,I162108);
DFFARX1 I_7141  ( .D(I124130), .CLK(I2702), .RSTB(I124079), .Q(I124053) );
nor I_7142 (I124161,I124096,I162093);
nand I_7143 (I124178,I124161,I162096);
not I_7144 (I124068,I124178);
DFFARX1 I_7145  ( .D(I124178), .CLK(I2702), .RSTB(I124079), .Q(I124050) );
not I_7146 (I124223,I162093);
not I_7147 (I124240,I124223);
not I_7148 (I124257,I162117);
nor I_7149 (I124274,I124257,I162090);
and I_7150 (I124291,I124274,I162111);
or I_7151 (I124308,I124291,I162102);
DFFARX1 I_7152  ( .D(I124308), .CLK(I2702), .RSTB(I124079), .Q(I124325) );
nor I_7153 (I124342,I124325,I124178);
nor I_7154 (I124359,I124325,I124240);
nand I_7155 (I124065,I124130,I124359);
nand I_7156 (I124390,I124096,I162117);
nand I_7157 (I124407,I124390,I124325);
and I_7158 (I124424,I124390,I124407);
DFFARX1 I_7159  ( .D(I124424), .CLK(I2702), .RSTB(I124079), .Q(I124047) );
DFFARX1 I_7160  ( .D(I124390), .CLK(I2702), .RSTB(I124079), .Q(I124455) );
and I_7161 (I124044,I124223,I124455);
DFFARX1 I_7162  ( .D(I162087), .CLK(I2702), .RSTB(I124079), .Q(I124486) );
not I_7163 (I124503,I124486);
nor I_7164 (I124520,I124178,I124503);
and I_7165 (I124537,I124486,I124520);
nand I_7166 (I124059,I124486,I124240);
DFFARX1 I_7167  ( .D(I124486), .CLK(I2702), .RSTB(I124079), .Q(I124568) );
not I_7168 (I124056,I124568);
DFFARX1 I_7169  ( .D(I162114), .CLK(I2702), .RSTB(I124079), .Q(I124599) );
not I_7170 (I124616,I124599);
or I_7171 (I124633,I124616,I124537);
DFFARX1 I_7172  ( .D(I124633), .CLK(I2702), .RSTB(I124079), .Q(I124062) );
nand I_7173 (I124071,I124616,I124342);
DFFARX1 I_7174  ( .D(I124616), .CLK(I2702), .RSTB(I124079), .Q(I124041) );
not I_7175 (I124725,I2709);
not I_7176 (I124742,I313932);
nor I_7177 (I124759,I313929,I313917);
nand I_7178 (I124776,I124759,I313920);
DFFARX1 I_7179  ( .D(I124776), .CLK(I2702), .RSTB(I124725), .Q(I124699) );
nor I_7180 (I124807,I124742,I313929);
nand I_7181 (I124824,I124807,I313926);
not I_7182 (I124714,I124824);
DFFARX1 I_7183  ( .D(I124824), .CLK(I2702), .RSTB(I124725), .Q(I124696) );
not I_7184 (I124869,I313929);
not I_7185 (I124886,I124869);
not I_7186 (I124903,I313938);
nor I_7187 (I124920,I124903,I313914);
and I_7188 (I124937,I124920,I313935);
or I_7189 (I124954,I124937,I313923);
DFFARX1 I_7190  ( .D(I124954), .CLK(I2702), .RSTB(I124725), .Q(I124971) );
nor I_7191 (I124988,I124971,I124824);
nor I_7192 (I125005,I124971,I124886);
nand I_7193 (I124711,I124776,I125005);
nand I_7194 (I125036,I124742,I313938);
nand I_7195 (I125053,I125036,I124971);
and I_7196 (I125070,I125036,I125053);
DFFARX1 I_7197  ( .D(I125070), .CLK(I2702), .RSTB(I124725), .Q(I124693) );
DFFARX1 I_7198  ( .D(I125036), .CLK(I2702), .RSTB(I124725), .Q(I125101) );
and I_7199 (I124690,I124869,I125101);
DFFARX1 I_7200  ( .D(I313944), .CLK(I2702), .RSTB(I124725), .Q(I125132) );
not I_7201 (I125149,I125132);
nor I_7202 (I125166,I124824,I125149);
and I_7203 (I125183,I125132,I125166);
nand I_7204 (I124705,I125132,I124886);
DFFARX1 I_7205  ( .D(I125132), .CLK(I2702), .RSTB(I124725), .Q(I125214) );
not I_7206 (I124702,I125214);
DFFARX1 I_7207  ( .D(I313941), .CLK(I2702), .RSTB(I124725), .Q(I125245) );
not I_7208 (I125262,I125245);
or I_7209 (I125279,I125262,I125183);
DFFARX1 I_7210  ( .D(I125279), .CLK(I2702), .RSTB(I124725), .Q(I124708) );
nand I_7211 (I124717,I125262,I124988);
DFFARX1 I_7212  ( .D(I125262), .CLK(I2702), .RSTB(I124725), .Q(I124687) );
not I_7213 (I125371,I2709);
not I_7214 (I125388,I493169);
nor I_7215 (I125405,I493151,I493160);
nand I_7216 (I125422,I125405,I493172);
DFFARX1 I_7217  ( .D(I125422), .CLK(I2702), .RSTB(I125371), .Q(I125345) );
nor I_7218 (I125453,I125388,I493151);
nand I_7219 (I125470,I125453,I493157);
not I_7220 (I125360,I125470);
DFFARX1 I_7221  ( .D(I125470), .CLK(I2702), .RSTB(I125371), .Q(I125342) );
not I_7222 (I125515,I493151);
not I_7223 (I125532,I125515);
not I_7224 (I125549,I493148);
nor I_7225 (I125566,I125549,I493166);
and I_7226 (I125583,I125566,I493154);
or I_7227 (I125600,I125583,I493175);
DFFARX1 I_7228  ( .D(I125600), .CLK(I2702), .RSTB(I125371), .Q(I125617) );
nor I_7229 (I125634,I125617,I125470);
nor I_7230 (I125651,I125617,I125532);
nand I_7231 (I125357,I125422,I125651);
nand I_7232 (I125682,I125388,I493148);
nand I_7233 (I125699,I125682,I125617);
and I_7234 (I125716,I125682,I125699);
DFFARX1 I_7235  ( .D(I125716), .CLK(I2702), .RSTB(I125371), .Q(I125339) );
DFFARX1 I_7236  ( .D(I125682), .CLK(I2702), .RSTB(I125371), .Q(I125747) );
and I_7237 (I125336,I125515,I125747);
DFFARX1 I_7238  ( .D(I493163), .CLK(I2702), .RSTB(I125371), .Q(I125778) );
not I_7239 (I125795,I125778);
nor I_7240 (I125812,I125470,I125795);
and I_7241 (I125829,I125778,I125812);
nand I_7242 (I125351,I125778,I125532);
DFFARX1 I_7243  ( .D(I125778), .CLK(I2702), .RSTB(I125371), .Q(I125860) );
not I_7244 (I125348,I125860);
DFFARX1 I_7245  ( .D(I493145), .CLK(I2702), .RSTB(I125371), .Q(I125891) );
not I_7246 (I125908,I125891);
or I_7247 (I125925,I125908,I125829);
DFFARX1 I_7248  ( .D(I125925), .CLK(I2702), .RSTB(I125371), .Q(I125354) );
nand I_7249 (I125363,I125908,I125634);
DFFARX1 I_7250  ( .D(I125908), .CLK(I2702), .RSTB(I125371), .Q(I125333) );
not I_7251 (I126017,I2709);
not I_7252 (I126034,I417479);
nor I_7253 (I126051,I417461,I417476);
nand I_7254 (I126068,I126051,I417485);
DFFARX1 I_7255  ( .D(I126068), .CLK(I2702), .RSTB(I126017), .Q(I125991) );
nor I_7256 (I126099,I126034,I417461);
nand I_7257 (I126116,I126099,I417488);
not I_7258 (I126006,I126116);
DFFARX1 I_7259  ( .D(I126116), .CLK(I2702), .RSTB(I126017), .Q(I125988) );
not I_7260 (I126161,I417461);
not I_7261 (I126178,I126161);
not I_7262 (I126195,I417491);
nor I_7263 (I126212,I126195,I417467);
and I_7264 (I126229,I126212,I417470);
or I_7265 (I126246,I126229,I417464);
DFFARX1 I_7266  ( .D(I126246), .CLK(I2702), .RSTB(I126017), .Q(I126263) );
nor I_7267 (I126280,I126263,I126116);
nor I_7268 (I126297,I126263,I126178);
nand I_7269 (I126003,I126068,I126297);
nand I_7270 (I126328,I126034,I417491);
nand I_7271 (I126345,I126328,I126263);
and I_7272 (I126362,I126328,I126345);
DFFARX1 I_7273  ( .D(I126362), .CLK(I2702), .RSTB(I126017), .Q(I125985) );
DFFARX1 I_7274  ( .D(I126328), .CLK(I2702), .RSTB(I126017), .Q(I126393) );
and I_7275 (I125982,I126161,I126393);
DFFARX1 I_7276  ( .D(I417473), .CLK(I2702), .RSTB(I126017), .Q(I126424) );
not I_7277 (I126441,I126424);
nor I_7278 (I126458,I126116,I126441);
and I_7279 (I126475,I126424,I126458);
nand I_7280 (I125997,I126424,I126178);
DFFARX1 I_7281  ( .D(I126424), .CLK(I2702), .RSTB(I126017), .Q(I126506) );
not I_7282 (I125994,I126506);
DFFARX1 I_7283  ( .D(I417482), .CLK(I2702), .RSTB(I126017), .Q(I126537) );
not I_7284 (I126554,I126537);
or I_7285 (I126571,I126554,I126475);
DFFARX1 I_7286  ( .D(I126571), .CLK(I2702), .RSTB(I126017), .Q(I126000) );
nand I_7287 (I126009,I126554,I126280);
DFFARX1 I_7288  ( .D(I126554), .CLK(I2702), .RSTB(I126017), .Q(I125979) );
not I_7289 (I126663,I2709);
not I_7290 (I126680,I334451);
nor I_7291 (I126697,I334463,I334445);
nand I_7292 (I126714,I126697,I334460);
DFFARX1 I_7293  ( .D(I126714), .CLK(I2702), .RSTB(I126663), .Q(I126637) );
nor I_7294 (I126745,I126680,I334463);
nand I_7295 (I126762,I126745,I334448);
not I_7296 (I126652,I126762);
DFFARX1 I_7297  ( .D(I126762), .CLK(I2702), .RSTB(I126663), .Q(I126634) );
not I_7298 (I126807,I334463);
not I_7299 (I126824,I126807);
not I_7300 (I126841,I334457);
nor I_7301 (I126858,I126841,I334436);
and I_7302 (I126875,I126858,I334439);
or I_7303 (I126892,I126875,I334442);
DFFARX1 I_7304  ( .D(I126892), .CLK(I2702), .RSTB(I126663), .Q(I126909) );
nor I_7305 (I126926,I126909,I126762);
nor I_7306 (I126943,I126909,I126824);
nand I_7307 (I126649,I126714,I126943);
nand I_7308 (I126974,I126680,I334457);
nand I_7309 (I126991,I126974,I126909);
and I_7310 (I127008,I126974,I126991);
DFFARX1 I_7311  ( .D(I127008), .CLK(I2702), .RSTB(I126663), .Q(I126631) );
DFFARX1 I_7312  ( .D(I126974), .CLK(I2702), .RSTB(I126663), .Q(I127039) );
and I_7313 (I126628,I126807,I127039);
DFFARX1 I_7314  ( .D(I334433), .CLK(I2702), .RSTB(I126663), .Q(I127070) );
not I_7315 (I127087,I127070);
nor I_7316 (I127104,I126762,I127087);
and I_7317 (I127121,I127070,I127104);
nand I_7318 (I126643,I127070,I126824);
DFFARX1 I_7319  ( .D(I127070), .CLK(I2702), .RSTB(I126663), .Q(I127152) );
not I_7320 (I126640,I127152);
DFFARX1 I_7321  ( .D(I334454), .CLK(I2702), .RSTB(I126663), .Q(I127183) );
not I_7322 (I127200,I127183);
or I_7323 (I127217,I127200,I127121);
DFFARX1 I_7324  ( .D(I127217), .CLK(I2702), .RSTB(I126663), .Q(I126646) );
nand I_7325 (I126655,I127200,I126926);
DFFARX1 I_7326  ( .D(I127200), .CLK(I2702), .RSTB(I126663), .Q(I126625) );
not I_7327 (I127309,I2709);
not I_7328 (I127326,I17862);
nor I_7329 (I127343,I17874,I17859);
nand I_7330 (I127360,I127343,I17871);
DFFARX1 I_7331  ( .D(I127360), .CLK(I2702), .RSTB(I127309), .Q(I127283) );
nor I_7332 (I127391,I127326,I17874);
nand I_7333 (I127408,I127391,I17889);
not I_7334 (I127298,I127408);
DFFARX1 I_7335  ( .D(I127408), .CLK(I2702), .RSTB(I127309), .Q(I127280) );
not I_7336 (I127453,I17874);
not I_7337 (I127470,I127453);
not I_7338 (I127487,I17865);
nor I_7339 (I127504,I127487,I17877);
and I_7340 (I127521,I127504,I17868);
or I_7341 (I127538,I127521,I17883);
DFFARX1 I_7342  ( .D(I127538), .CLK(I2702), .RSTB(I127309), .Q(I127555) );
nor I_7343 (I127572,I127555,I127408);
nor I_7344 (I127589,I127555,I127470);
nand I_7345 (I127295,I127360,I127589);
nand I_7346 (I127620,I127326,I17865);
nand I_7347 (I127637,I127620,I127555);
and I_7348 (I127654,I127620,I127637);
DFFARX1 I_7349  ( .D(I127654), .CLK(I2702), .RSTB(I127309), .Q(I127277) );
DFFARX1 I_7350  ( .D(I127620), .CLK(I2702), .RSTB(I127309), .Q(I127685) );
and I_7351 (I127274,I127453,I127685);
DFFARX1 I_7352  ( .D(I17886), .CLK(I2702), .RSTB(I127309), .Q(I127716) );
not I_7353 (I127733,I127716);
nor I_7354 (I127750,I127408,I127733);
and I_7355 (I127767,I127716,I127750);
nand I_7356 (I127289,I127716,I127470);
DFFARX1 I_7357  ( .D(I127716), .CLK(I2702), .RSTB(I127309), .Q(I127798) );
not I_7358 (I127286,I127798);
DFFARX1 I_7359  ( .D(I17880), .CLK(I2702), .RSTB(I127309), .Q(I127829) );
not I_7360 (I127846,I127829);
or I_7361 (I127863,I127846,I127767);
DFFARX1 I_7362  ( .D(I127863), .CLK(I2702), .RSTB(I127309), .Q(I127292) );
nand I_7363 (I127301,I127846,I127572);
DFFARX1 I_7364  ( .D(I127846), .CLK(I2702), .RSTB(I127309), .Q(I127271) );
not I_7365 (I127955,I2709);
not I_7366 (I127972,I662108);
nor I_7367 (I127989,I662123,I662138);
nand I_7368 (I128006,I127989,I662126);
DFFARX1 I_7369  ( .D(I128006), .CLK(I2702), .RSTB(I127955), .Q(I127929) );
nor I_7370 (I128037,I127972,I662123);
nand I_7371 (I128054,I128037,I662129);
not I_7372 (I127944,I128054);
DFFARX1 I_7373  ( .D(I128054), .CLK(I2702), .RSTB(I127955), .Q(I127926) );
not I_7374 (I128099,I662123);
not I_7375 (I128116,I128099);
not I_7376 (I128133,I662135);
nor I_7377 (I128150,I128133,I662132);
and I_7378 (I128167,I128150,I662111);
or I_7379 (I128184,I128167,I662120);
DFFARX1 I_7380  ( .D(I128184), .CLK(I2702), .RSTB(I127955), .Q(I128201) );
nor I_7381 (I128218,I128201,I128054);
nor I_7382 (I128235,I128201,I128116);
nand I_7383 (I127941,I128006,I128235);
nand I_7384 (I128266,I127972,I662135);
nand I_7385 (I128283,I128266,I128201);
and I_7386 (I128300,I128266,I128283);
DFFARX1 I_7387  ( .D(I128300), .CLK(I2702), .RSTB(I127955), .Q(I127923) );
DFFARX1 I_7388  ( .D(I128266), .CLK(I2702), .RSTB(I127955), .Q(I128331) );
and I_7389 (I127920,I128099,I128331);
DFFARX1 I_7390  ( .D(I662117), .CLK(I2702), .RSTB(I127955), .Q(I128362) );
not I_7391 (I128379,I128362);
nor I_7392 (I128396,I128054,I128379);
and I_7393 (I128413,I128362,I128396);
nand I_7394 (I127935,I128362,I128116);
DFFARX1 I_7395  ( .D(I128362), .CLK(I2702), .RSTB(I127955), .Q(I128444) );
not I_7396 (I127932,I128444);
DFFARX1 I_7397  ( .D(I662114), .CLK(I2702), .RSTB(I127955), .Q(I128475) );
not I_7398 (I128492,I128475);
or I_7399 (I128509,I128492,I128413);
DFFARX1 I_7400  ( .D(I128509), .CLK(I2702), .RSTB(I127955), .Q(I127938) );
nand I_7401 (I127947,I128492,I128218);
DFFARX1 I_7402  ( .D(I128492), .CLK(I2702), .RSTB(I127955), .Q(I127917) );
not I_7403 (I128601,I2709);
not I_7404 (I128618,I191277);
nor I_7405 (I128635,I191265,I191271);
nand I_7406 (I128652,I128635,I191280);
DFFARX1 I_7407  ( .D(I128652), .CLK(I2702), .RSTB(I128601), .Q(I128575) );
nor I_7408 (I128683,I128618,I191265);
nand I_7409 (I128700,I128683,I191268);
not I_7410 (I128590,I128700);
DFFARX1 I_7411  ( .D(I128700), .CLK(I2702), .RSTB(I128601), .Q(I128572) );
not I_7412 (I128745,I191265);
not I_7413 (I128762,I128745);
not I_7414 (I128779,I191289);
nor I_7415 (I128796,I128779,I191262);
and I_7416 (I128813,I128796,I191283);
or I_7417 (I128830,I128813,I191274);
DFFARX1 I_7418  ( .D(I128830), .CLK(I2702), .RSTB(I128601), .Q(I128847) );
nor I_7419 (I128864,I128847,I128700);
nor I_7420 (I128881,I128847,I128762);
nand I_7421 (I128587,I128652,I128881);
nand I_7422 (I128912,I128618,I191289);
nand I_7423 (I128929,I128912,I128847);
and I_7424 (I128946,I128912,I128929);
DFFARX1 I_7425  ( .D(I128946), .CLK(I2702), .RSTB(I128601), .Q(I128569) );
DFFARX1 I_7426  ( .D(I128912), .CLK(I2702), .RSTB(I128601), .Q(I128977) );
and I_7427 (I128566,I128745,I128977);
DFFARX1 I_7428  ( .D(I191259), .CLK(I2702), .RSTB(I128601), .Q(I129008) );
not I_7429 (I129025,I129008);
nor I_7430 (I129042,I128700,I129025);
and I_7431 (I129059,I129008,I129042);
nand I_7432 (I128581,I129008,I128762);
DFFARX1 I_7433  ( .D(I129008), .CLK(I2702), .RSTB(I128601), .Q(I129090) );
not I_7434 (I128578,I129090);
DFFARX1 I_7435  ( .D(I191286), .CLK(I2702), .RSTB(I128601), .Q(I129121) );
not I_7436 (I129138,I129121);
or I_7437 (I129155,I129138,I129059);
DFFARX1 I_7438  ( .D(I129155), .CLK(I2702), .RSTB(I128601), .Q(I128584) );
nand I_7439 (I128593,I129138,I128864);
DFFARX1 I_7440  ( .D(I129138), .CLK(I2702), .RSTB(I128601), .Q(I128563) );
not I_7441 (I129247,I2709);
not I_7442 (I129264,I641980);
nor I_7443 (I129281,I641995,I642010);
nand I_7444 (I129298,I129281,I641998);
DFFARX1 I_7445  ( .D(I129298), .CLK(I2702), .RSTB(I129247), .Q(I129221) );
nor I_7446 (I129329,I129264,I641995);
nand I_7447 (I129346,I129329,I642001);
not I_7448 (I129236,I129346);
DFFARX1 I_7449  ( .D(I129346), .CLK(I2702), .RSTB(I129247), .Q(I129218) );
not I_7450 (I129391,I641995);
not I_7451 (I129408,I129391);
not I_7452 (I129425,I642007);
nor I_7453 (I129442,I129425,I642004);
and I_7454 (I129459,I129442,I641983);
or I_7455 (I129476,I129459,I641992);
DFFARX1 I_7456  ( .D(I129476), .CLK(I2702), .RSTB(I129247), .Q(I129493) );
nor I_7457 (I129510,I129493,I129346);
nor I_7458 (I129527,I129493,I129408);
nand I_7459 (I129233,I129298,I129527);
nand I_7460 (I129558,I129264,I642007);
nand I_7461 (I129575,I129558,I129493);
and I_7462 (I129592,I129558,I129575);
DFFARX1 I_7463  ( .D(I129592), .CLK(I2702), .RSTB(I129247), .Q(I129215) );
DFFARX1 I_7464  ( .D(I129558), .CLK(I2702), .RSTB(I129247), .Q(I129623) );
and I_7465 (I129212,I129391,I129623);
DFFARX1 I_7466  ( .D(I641989), .CLK(I2702), .RSTB(I129247), .Q(I129654) );
not I_7467 (I129671,I129654);
nor I_7468 (I129688,I129346,I129671);
and I_7469 (I129705,I129654,I129688);
nand I_7470 (I129227,I129654,I129408);
DFFARX1 I_7471  ( .D(I129654), .CLK(I2702), .RSTB(I129247), .Q(I129736) );
not I_7472 (I129224,I129736);
DFFARX1 I_7473  ( .D(I641986), .CLK(I2702), .RSTB(I129247), .Q(I129767) );
not I_7474 (I129784,I129767);
or I_7475 (I129801,I129784,I129705);
DFFARX1 I_7476  ( .D(I129801), .CLK(I2702), .RSTB(I129247), .Q(I129230) );
nand I_7477 (I129239,I129784,I129510);
DFFARX1 I_7478  ( .D(I129784), .CLK(I2702), .RSTB(I129247), .Q(I129209) );
not I_7479 (I129893,I2709);
not I_7480 (I129910,I170724);
nor I_7481 (I129927,I170712,I170718);
nand I_7482 (I129944,I129927,I170727);
DFFARX1 I_7483  ( .D(I129944), .CLK(I2702), .RSTB(I129893), .Q(I129867) );
nor I_7484 (I129975,I129910,I170712);
nand I_7485 (I129992,I129975,I170715);
not I_7486 (I129882,I129992);
DFFARX1 I_7487  ( .D(I129992), .CLK(I2702), .RSTB(I129893), .Q(I129864) );
not I_7488 (I130037,I170712);
not I_7489 (I130054,I130037);
not I_7490 (I130071,I170736);
nor I_7491 (I130088,I130071,I170709);
and I_7492 (I130105,I130088,I170730);
or I_7493 (I130122,I130105,I170721);
DFFARX1 I_7494  ( .D(I130122), .CLK(I2702), .RSTB(I129893), .Q(I130139) );
nor I_7495 (I130156,I130139,I129992);
nor I_7496 (I130173,I130139,I130054);
nand I_7497 (I129879,I129944,I130173);
nand I_7498 (I130204,I129910,I170736);
nand I_7499 (I130221,I130204,I130139);
and I_7500 (I130238,I130204,I130221);
DFFARX1 I_7501  ( .D(I130238), .CLK(I2702), .RSTB(I129893), .Q(I129861) );
DFFARX1 I_7502  ( .D(I130204), .CLK(I2702), .RSTB(I129893), .Q(I130269) );
and I_7503 (I129858,I130037,I130269);
DFFARX1 I_7504  ( .D(I170706), .CLK(I2702), .RSTB(I129893), .Q(I130300) );
not I_7505 (I130317,I130300);
nor I_7506 (I130334,I129992,I130317);
and I_7507 (I130351,I130300,I130334);
nand I_7508 (I129873,I130300,I130054);
DFFARX1 I_7509  ( .D(I130300), .CLK(I2702), .RSTB(I129893), .Q(I130382) );
not I_7510 (I129870,I130382);
DFFARX1 I_7511  ( .D(I170733), .CLK(I2702), .RSTB(I129893), .Q(I130413) );
not I_7512 (I130430,I130413);
or I_7513 (I130447,I130430,I130351);
DFFARX1 I_7514  ( .D(I130447), .CLK(I2702), .RSTB(I129893), .Q(I129876) );
nand I_7515 (I129885,I130430,I130156);
DFFARX1 I_7516  ( .D(I130430), .CLK(I2702), .RSTB(I129893), .Q(I129855) );
not I_7517 (I130539,I2709);
not I_7518 (I130556,I427883);
nor I_7519 (I130573,I427865,I427880);
nand I_7520 (I130590,I130573,I427889);
DFFARX1 I_7521  ( .D(I130590), .CLK(I2702), .RSTB(I130539), .Q(I130513) );
nor I_7522 (I130621,I130556,I427865);
nand I_7523 (I130638,I130621,I427892);
not I_7524 (I130528,I130638);
DFFARX1 I_7525  ( .D(I130638), .CLK(I2702), .RSTB(I130539), .Q(I130510) );
not I_7526 (I130683,I427865);
not I_7527 (I130700,I130683);
not I_7528 (I130717,I427895);
nor I_7529 (I130734,I130717,I427871);
and I_7530 (I130751,I130734,I427874);
or I_7531 (I130768,I130751,I427868);
DFFARX1 I_7532  ( .D(I130768), .CLK(I2702), .RSTB(I130539), .Q(I130785) );
nor I_7533 (I130802,I130785,I130638);
nor I_7534 (I130819,I130785,I130700);
nand I_7535 (I130525,I130590,I130819);
nand I_7536 (I130850,I130556,I427895);
nand I_7537 (I130867,I130850,I130785);
and I_7538 (I130884,I130850,I130867);
DFFARX1 I_7539  ( .D(I130884), .CLK(I2702), .RSTB(I130539), .Q(I130507) );
DFFARX1 I_7540  ( .D(I130850), .CLK(I2702), .RSTB(I130539), .Q(I130915) );
and I_7541 (I130504,I130683,I130915);
DFFARX1 I_7542  ( .D(I427877), .CLK(I2702), .RSTB(I130539), .Q(I130946) );
not I_7543 (I130963,I130946);
nor I_7544 (I130980,I130638,I130963);
and I_7545 (I130997,I130946,I130980);
nand I_7546 (I130519,I130946,I130700);
DFFARX1 I_7547  ( .D(I130946), .CLK(I2702), .RSTB(I130539), .Q(I131028) );
not I_7548 (I130516,I131028);
DFFARX1 I_7549  ( .D(I427886), .CLK(I2702), .RSTB(I130539), .Q(I131059) );
not I_7550 (I131076,I131059);
or I_7551 (I131093,I131076,I130997);
DFFARX1 I_7552  ( .D(I131093), .CLK(I2702), .RSTB(I130539), .Q(I130522) );
nand I_7553 (I130531,I131076,I130802);
DFFARX1 I_7554  ( .D(I131076), .CLK(I2702), .RSTB(I130539), .Q(I130501) );
not I_7555 (I131185,I2709);
not I_7556 (I131202,I633174);
nor I_7557 (I131219,I633189,I633204);
nand I_7558 (I131236,I131219,I633192);
DFFARX1 I_7559  ( .D(I131236), .CLK(I2702), .RSTB(I131185), .Q(I131159) );
nor I_7560 (I131267,I131202,I633189);
nand I_7561 (I131284,I131267,I633195);
not I_7562 (I131174,I131284);
DFFARX1 I_7563  ( .D(I131284), .CLK(I2702), .RSTB(I131185), .Q(I131156) );
not I_7564 (I131329,I633189);
not I_7565 (I131346,I131329);
not I_7566 (I131363,I633201);
nor I_7567 (I131380,I131363,I633198);
and I_7568 (I131397,I131380,I633177);
or I_7569 (I131414,I131397,I633186);
DFFARX1 I_7570  ( .D(I131414), .CLK(I2702), .RSTB(I131185), .Q(I131431) );
nor I_7571 (I131448,I131431,I131284);
nor I_7572 (I131465,I131431,I131346);
nand I_7573 (I131171,I131236,I131465);
nand I_7574 (I131496,I131202,I633201);
nand I_7575 (I131513,I131496,I131431);
and I_7576 (I131530,I131496,I131513);
DFFARX1 I_7577  ( .D(I131530), .CLK(I2702), .RSTB(I131185), .Q(I131153) );
DFFARX1 I_7578  ( .D(I131496), .CLK(I2702), .RSTB(I131185), .Q(I131561) );
and I_7579 (I131150,I131329,I131561);
DFFARX1 I_7580  ( .D(I633183), .CLK(I2702), .RSTB(I131185), .Q(I131592) );
not I_7581 (I131609,I131592);
nor I_7582 (I131626,I131284,I131609);
and I_7583 (I131643,I131592,I131626);
nand I_7584 (I131165,I131592,I131346);
DFFARX1 I_7585  ( .D(I131592), .CLK(I2702), .RSTB(I131185), .Q(I131674) );
not I_7586 (I131162,I131674);
DFFARX1 I_7587  ( .D(I633180), .CLK(I2702), .RSTB(I131185), .Q(I131705) );
not I_7588 (I131722,I131705);
or I_7589 (I131739,I131722,I131643);
DFFARX1 I_7590  ( .D(I131739), .CLK(I2702), .RSTB(I131185), .Q(I131168) );
nand I_7591 (I131177,I131722,I131448);
DFFARX1 I_7592  ( .D(I131722), .CLK(I2702), .RSTB(I131185), .Q(I131147) );
not I_7593 (I131831,I2709);
not I_7594 (I131848,I616191);
nor I_7595 (I131865,I616206,I616221);
nand I_7596 (I131882,I131865,I616209);
DFFARX1 I_7597  ( .D(I131882), .CLK(I2702), .RSTB(I131831), .Q(I131805) );
nor I_7598 (I131913,I131848,I616206);
nand I_7599 (I131930,I131913,I616212);
not I_7600 (I131820,I131930);
DFFARX1 I_7601  ( .D(I131930), .CLK(I2702), .RSTB(I131831), .Q(I131802) );
not I_7602 (I131975,I616206);
not I_7603 (I131992,I131975);
not I_7604 (I132009,I616218);
nor I_7605 (I132026,I132009,I616215);
and I_7606 (I132043,I132026,I616194);
or I_7607 (I132060,I132043,I616203);
DFFARX1 I_7608  ( .D(I132060), .CLK(I2702), .RSTB(I131831), .Q(I132077) );
nor I_7609 (I132094,I132077,I131930);
nor I_7610 (I132111,I132077,I131992);
nand I_7611 (I131817,I131882,I132111);
nand I_7612 (I132142,I131848,I616218);
nand I_7613 (I132159,I132142,I132077);
and I_7614 (I132176,I132142,I132159);
DFFARX1 I_7615  ( .D(I132176), .CLK(I2702), .RSTB(I131831), .Q(I131799) );
DFFARX1 I_7616  ( .D(I132142), .CLK(I2702), .RSTB(I131831), .Q(I132207) );
and I_7617 (I131796,I131975,I132207);
DFFARX1 I_7618  ( .D(I616200), .CLK(I2702), .RSTB(I131831), .Q(I132238) );
not I_7619 (I132255,I132238);
nor I_7620 (I132272,I131930,I132255);
and I_7621 (I132289,I132238,I132272);
nand I_7622 (I131811,I132238,I131992);
DFFARX1 I_7623  ( .D(I132238), .CLK(I2702), .RSTB(I131831), .Q(I132320) );
not I_7624 (I131808,I132320);
DFFARX1 I_7625  ( .D(I616197), .CLK(I2702), .RSTB(I131831), .Q(I132351) );
not I_7626 (I132368,I132351);
or I_7627 (I132385,I132368,I132289);
DFFARX1 I_7628  ( .D(I132385), .CLK(I2702), .RSTB(I131831), .Q(I131814) );
nand I_7629 (I131823,I132368,I132094);
DFFARX1 I_7630  ( .D(I132368), .CLK(I2702), .RSTB(I131831), .Q(I131793) );
not I_7631 (I132477,I2709);
not I_7632 (I132494,I651415);
nor I_7633 (I132511,I651430,I651445);
nand I_7634 (I132528,I132511,I651433);
DFFARX1 I_7635  ( .D(I132528), .CLK(I2702), .RSTB(I132477), .Q(I132451) );
nor I_7636 (I132559,I132494,I651430);
nand I_7637 (I132576,I132559,I651436);
not I_7638 (I132466,I132576);
DFFARX1 I_7639  ( .D(I132576), .CLK(I2702), .RSTB(I132477), .Q(I132448) );
not I_7640 (I132621,I651430);
not I_7641 (I132638,I132621);
not I_7642 (I132655,I651442);
nor I_7643 (I132672,I132655,I651439);
and I_7644 (I132689,I132672,I651418);
or I_7645 (I132706,I132689,I651427);
DFFARX1 I_7646  ( .D(I132706), .CLK(I2702), .RSTB(I132477), .Q(I132723) );
nor I_7647 (I132740,I132723,I132576);
nor I_7648 (I132757,I132723,I132638);
nand I_7649 (I132463,I132528,I132757);
nand I_7650 (I132788,I132494,I651442);
nand I_7651 (I132805,I132788,I132723);
and I_7652 (I132822,I132788,I132805);
DFFARX1 I_7653  ( .D(I132822), .CLK(I2702), .RSTB(I132477), .Q(I132445) );
DFFARX1 I_7654  ( .D(I132788), .CLK(I2702), .RSTB(I132477), .Q(I132853) );
and I_7655 (I132442,I132621,I132853);
DFFARX1 I_7656  ( .D(I651424), .CLK(I2702), .RSTB(I132477), .Q(I132884) );
not I_7657 (I132901,I132884);
nor I_7658 (I132918,I132576,I132901);
and I_7659 (I132935,I132884,I132918);
nand I_7660 (I132457,I132884,I132638);
DFFARX1 I_7661  ( .D(I132884), .CLK(I2702), .RSTB(I132477), .Q(I132966) );
not I_7662 (I132454,I132966);
DFFARX1 I_7663  ( .D(I651421), .CLK(I2702), .RSTB(I132477), .Q(I132997) );
not I_7664 (I133014,I132997);
or I_7665 (I133031,I133014,I132935);
DFFARX1 I_7666  ( .D(I133031), .CLK(I2702), .RSTB(I132477), .Q(I132460) );
nand I_7667 (I132469,I133014,I132740);
DFFARX1 I_7668  ( .D(I133014), .CLK(I2702), .RSTB(I132477), .Q(I132439) );
not I_7669 (I133123,I2709);
not I_7670 (I133140,I364167);
nor I_7671 (I133157,I364179,I364161);
nand I_7672 (I133174,I133157,I364176);
DFFARX1 I_7673  ( .D(I133174), .CLK(I2702), .RSTB(I133123), .Q(I133097) );
nor I_7674 (I133205,I133140,I364179);
nand I_7675 (I133222,I133205,I364164);
not I_7676 (I133112,I133222);
DFFARX1 I_7677  ( .D(I133222), .CLK(I2702), .RSTB(I133123), .Q(I133094) );
not I_7678 (I133267,I364179);
not I_7679 (I133284,I133267);
not I_7680 (I133301,I364173);
nor I_7681 (I133318,I133301,I364152);
and I_7682 (I133335,I133318,I364155);
or I_7683 (I133352,I133335,I364158);
DFFARX1 I_7684  ( .D(I133352), .CLK(I2702), .RSTB(I133123), .Q(I133369) );
nor I_7685 (I133386,I133369,I133222);
nor I_7686 (I133403,I133369,I133284);
nand I_7687 (I133109,I133174,I133403);
nand I_7688 (I133434,I133140,I364173);
nand I_7689 (I133451,I133434,I133369);
and I_7690 (I133468,I133434,I133451);
DFFARX1 I_7691  ( .D(I133468), .CLK(I2702), .RSTB(I133123), .Q(I133091) );
DFFARX1 I_7692  ( .D(I133434), .CLK(I2702), .RSTB(I133123), .Q(I133499) );
and I_7693 (I133088,I133267,I133499);
DFFARX1 I_7694  ( .D(I364149), .CLK(I2702), .RSTB(I133123), .Q(I133530) );
not I_7695 (I133547,I133530);
nor I_7696 (I133564,I133222,I133547);
and I_7697 (I133581,I133530,I133564);
nand I_7698 (I133103,I133530,I133284);
DFFARX1 I_7699  ( .D(I133530), .CLK(I2702), .RSTB(I133123), .Q(I133612) );
not I_7700 (I133100,I133612);
DFFARX1 I_7701  ( .D(I364170), .CLK(I2702), .RSTB(I133123), .Q(I133643) );
not I_7702 (I133660,I133643);
or I_7703 (I133677,I133660,I133581);
DFFARX1 I_7704  ( .D(I133677), .CLK(I2702), .RSTB(I133123), .Q(I133106) );
nand I_7705 (I133115,I133660,I133386);
DFFARX1 I_7706  ( .D(I133660), .CLK(I2702), .RSTB(I133123), .Q(I133085) );
not I_7707 (I133769,I2709);
not I_7708 (I133786,I5520);
nor I_7709 (I133803,I5532,I5517);
nand I_7710 (I133820,I133803,I5529);
DFFARX1 I_7711  ( .D(I133820), .CLK(I2702), .RSTB(I133769), .Q(I133743) );
nor I_7712 (I133851,I133786,I5532);
nand I_7713 (I133868,I133851,I5547);
not I_7714 (I133758,I133868);
DFFARX1 I_7715  ( .D(I133868), .CLK(I2702), .RSTB(I133769), .Q(I133740) );
not I_7716 (I133913,I5532);
not I_7717 (I133930,I133913);
not I_7718 (I133947,I5523);
nor I_7719 (I133964,I133947,I5535);
and I_7720 (I133981,I133964,I5526);
or I_7721 (I133998,I133981,I5541);
DFFARX1 I_7722  ( .D(I133998), .CLK(I2702), .RSTB(I133769), .Q(I134015) );
nor I_7723 (I134032,I134015,I133868);
nor I_7724 (I134049,I134015,I133930);
nand I_7725 (I133755,I133820,I134049);
nand I_7726 (I134080,I133786,I5523);
nand I_7727 (I134097,I134080,I134015);
and I_7728 (I134114,I134080,I134097);
DFFARX1 I_7729  ( .D(I134114), .CLK(I2702), .RSTB(I133769), .Q(I133737) );
DFFARX1 I_7730  ( .D(I134080), .CLK(I2702), .RSTB(I133769), .Q(I134145) );
and I_7731 (I133734,I133913,I134145);
DFFARX1 I_7732  ( .D(I5544), .CLK(I2702), .RSTB(I133769), .Q(I134176) );
not I_7733 (I134193,I134176);
nor I_7734 (I134210,I133868,I134193);
and I_7735 (I134227,I134176,I134210);
nand I_7736 (I133749,I134176,I133930);
DFFARX1 I_7737  ( .D(I134176), .CLK(I2702), .RSTB(I133769), .Q(I134258) );
not I_7738 (I133746,I134258);
DFFARX1 I_7739  ( .D(I5538), .CLK(I2702), .RSTB(I133769), .Q(I134289) );
not I_7740 (I134306,I134289);
or I_7741 (I134323,I134306,I134227);
DFFARX1 I_7742  ( .D(I134323), .CLK(I2702), .RSTB(I133769), .Q(I133752) );
nand I_7743 (I133761,I134306,I134032);
DFFARX1 I_7744  ( .D(I134306), .CLK(I2702), .RSTB(I133769), .Q(I133731) );
not I_7745 (I134415,I2709);
not I_7746 (I134432,I469700);
nor I_7747 (I134449,I469688,I469694);
nand I_7748 (I134466,I134449,I469685);
DFFARX1 I_7749  ( .D(I134466), .CLK(I2702), .RSTB(I134415), .Q(I134389) );
nor I_7750 (I134497,I134432,I469688);
nand I_7751 (I134514,I134497,I469691);
not I_7752 (I134404,I134514);
DFFARX1 I_7753  ( .D(I134514), .CLK(I2702), .RSTB(I134415), .Q(I134386) );
not I_7754 (I134559,I469688);
not I_7755 (I134576,I134559);
not I_7756 (I134593,I469703);
nor I_7757 (I134610,I134593,I469715);
and I_7758 (I134627,I134610,I469697);
or I_7759 (I134644,I134627,I469712);
DFFARX1 I_7760  ( .D(I134644), .CLK(I2702), .RSTB(I134415), .Q(I134661) );
nor I_7761 (I134678,I134661,I134514);
nor I_7762 (I134695,I134661,I134576);
nand I_7763 (I134401,I134466,I134695);
nand I_7764 (I134726,I134432,I469703);
nand I_7765 (I134743,I134726,I134661);
and I_7766 (I134760,I134726,I134743);
DFFARX1 I_7767  ( .D(I134760), .CLK(I2702), .RSTB(I134415), .Q(I134383) );
DFFARX1 I_7768  ( .D(I134726), .CLK(I2702), .RSTB(I134415), .Q(I134791) );
and I_7769 (I134380,I134559,I134791);
DFFARX1 I_7770  ( .D(I469706), .CLK(I2702), .RSTB(I134415), .Q(I134822) );
not I_7771 (I134839,I134822);
nor I_7772 (I134856,I134514,I134839);
and I_7773 (I134873,I134822,I134856);
nand I_7774 (I134395,I134822,I134576);
DFFARX1 I_7775  ( .D(I134822), .CLK(I2702), .RSTB(I134415), .Q(I134904) );
not I_7776 (I134392,I134904);
DFFARX1 I_7777  ( .D(I469709), .CLK(I2702), .RSTB(I134415), .Q(I134935) );
not I_7778 (I134952,I134935);
or I_7779 (I134969,I134952,I134873);
DFFARX1 I_7780  ( .D(I134969), .CLK(I2702), .RSTB(I134415), .Q(I134398) );
nand I_7781 (I134407,I134952,I134678);
DFFARX1 I_7782  ( .D(I134952), .CLK(I2702), .RSTB(I134415), .Q(I134377) );
not I_7783 (I135061,I2709);
not I_7784 (I135078,I347371);
nor I_7785 (I135095,I347383,I347365);
nand I_7786 (I135112,I135095,I347380);
DFFARX1 I_7787  ( .D(I135112), .CLK(I2702), .RSTB(I135061), .Q(I135035) );
nor I_7788 (I135143,I135078,I347383);
nand I_7789 (I135160,I135143,I347368);
not I_7790 (I135050,I135160);
DFFARX1 I_7791  ( .D(I135160), .CLK(I2702), .RSTB(I135061), .Q(I135032) );
not I_7792 (I135205,I347383);
not I_7793 (I135222,I135205);
not I_7794 (I135239,I347377);
nor I_7795 (I135256,I135239,I347356);
and I_7796 (I135273,I135256,I347359);
or I_7797 (I135290,I135273,I347362);
DFFARX1 I_7798  ( .D(I135290), .CLK(I2702), .RSTB(I135061), .Q(I135307) );
nor I_7799 (I135324,I135307,I135160);
nor I_7800 (I135341,I135307,I135222);
nand I_7801 (I135047,I135112,I135341);
nand I_7802 (I135372,I135078,I347377);
nand I_7803 (I135389,I135372,I135307);
and I_7804 (I135406,I135372,I135389);
DFFARX1 I_7805  ( .D(I135406), .CLK(I2702), .RSTB(I135061), .Q(I135029) );
DFFARX1 I_7806  ( .D(I135372), .CLK(I2702), .RSTB(I135061), .Q(I135437) );
and I_7807 (I135026,I135205,I135437);
DFFARX1 I_7808  ( .D(I347353), .CLK(I2702), .RSTB(I135061), .Q(I135468) );
not I_7809 (I135485,I135468);
nor I_7810 (I135502,I135160,I135485);
and I_7811 (I135519,I135468,I135502);
nand I_7812 (I135041,I135468,I135222);
DFFARX1 I_7813  ( .D(I135468), .CLK(I2702), .RSTB(I135061), .Q(I135550) );
not I_7814 (I135038,I135550);
DFFARX1 I_7815  ( .D(I347374), .CLK(I2702), .RSTB(I135061), .Q(I135581) );
not I_7816 (I135598,I135581);
or I_7817 (I135615,I135598,I135519);
DFFARX1 I_7818  ( .D(I135615), .CLK(I2702), .RSTB(I135061), .Q(I135044) );
nand I_7819 (I135053,I135598,I135324);
DFFARX1 I_7820  ( .D(I135598), .CLK(I2702), .RSTB(I135061), .Q(I135023) );
not I_7821 (I135707,I2709);
not I_7822 (I135724,I199878);
nor I_7823 (I135741,I199908,I199887);
nand I_7824 (I135758,I135741,I199899);
DFFARX1 I_7825  ( .D(I135758), .CLK(I2702), .RSTB(I135707), .Q(I135681) );
nor I_7826 (I135789,I135724,I199908);
nand I_7827 (I135806,I135789,I199881);
not I_7828 (I135696,I135806);
DFFARX1 I_7829  ( .D(I135806), .CLK(I2702), .RSTB(I135707), .Q(I135678) );
not I_7830 (I135851,I199908);
not I_7831 (I135868,I135851);
not I_7832 (I135885,I199884);
nor I_7833 (I135902,I135885,I199902);
and I_7834 (I135919,I135902,I199893);
or I_7835 (I135936,I135919,I199890);
DFFARX1 I_7836  ( .D(I135936), .CLK(I2702), .RSTB(I135707), .Q(I135953) );
nor I_7837 (I135970,I135953,I135806);
nor I_7838 (I135987,I135953,I135868);
nand I_7839 (I135693,I135758,I135987);
nand I_7840 (I136018,I135724,I199884);
nand I_7841 (I136035,I136018,I135953);
and I_7842 (I136052,I136018,I136035);
DFFARX1 I_7843  ( .D(I136052), .CLK(I2702), .RSTB(I135707), .Q(I135675) );
DFFARX1 I_7844  ( .D(I136018), .CLK(I2702), .RSTB(I135707), .Q(I136083) );
and I_7845 (I135672,I135851,I136083);
DFFARX1 I_7846  ( .D(I199896), .CLK(I2702), .RSTB(I135707), .Q(I136114) );
not I_7847 (I136131,I136114);
nor I_7848 (I136148,I135806,I136131);
and I_7849 (I136165,I136114,I136148);
nand I_7850 (I135687,I136114,I135868);
DFFARX1 I_7851  ( .D(I136114), .CLK(I2702), .RSTB(I135707), .Q(I136196) );
not I_7852 (I135684,I136196);
DFFARX1 I_7853  ( .D(I199905), .CLK(I2702), .RSTB(I135707), .Q(I136227) );
not I_7854 (I136244,I136227);
or I_7855 (I136261,I136244,I136165);
DFFARX1 I_7856  ( .D(I136261), .CLK(I2702), .RSTB(I135707), .Q(I135690) );
nand I_7857 (I135699,I136244,I135970);
DFFARX1 I_7858  ( .D(I136244), .CLK(I2702), .RSTB(I135707), .Q(I135669) );
not I_7859 (I136353,I2709);
not I_7860 (I136370,I566136);
nor I_7861 (I136387,I566112,I566118);
nand I_7862 (I136404,I136387,I566121);
DFFARX1 I_7863  ( .D(I136404), .CLK(I2702), .RSTB(I136353), .Q(I136327) );
nor I_7864 (I136435,I136370,I566112);
nand I_7865 (I136452,I136435,I566130);
not I_7866 (I136342,I136452);
DFFARX1 I_7867  ( .D(I136452), .CLK(I2702), .RSTB(I136353), .Q(I136324) );
not I_7868 (I136497,I566112);
not I_7869 (I136514,I136497);
not I_7870 (I136531,I566109);
nor I_7871 (I136548,I136531,I566124);
and I_7872 (I136565,I136548,I566115);
or I_7873 (I136582,I136565,I566127);
DFFARX1 I_7874  ( .D(I136582), .CLK(I2702), .RSTB(I136353), .Q(I136599) );
nor I_7875 (I136616,I136599,I136452);
nor I_7876 (I136633,I136599,I136514);
nand I_7877 (I136339,I136404,I136633);
nand I_7878 (I136664,I136370,I566109);
nand I_7879 (I136681,I136664,I136599);
and I_7880 (I136698,I136664,I136681);
DFFARX1 I_7881  ( .D(I136698), .CLK(I2702), .RSTB(I136353), .Q(I136321) );
DFFARX1 I_7882  ( .D(I136664), .CLK(I2702), .RSTB(I136353), .Q(I136729) );
and I_7883 (I136318,I136497,I136729);
DFFARX1 I_7884  ( .D(I566139), .CLK(I2702), .RSTB(I136353), .Q(I136760) );
not I_7885 (I136777,I136760);
nor I_7886 (I136794,I136452,I136777);
and I_7887 (I136811,I136760,I136794);
nand I_7888 (I136333,I136760,I136514);
DFFARX1 I_7889  ( .D(I136760), .CLK(I2702), .RSTB(I136353), .Q(I136842) );
not I_7890 (I136330,I136842);
DFFARX1 I_7891  ( .D(I566133), .CLK(I2702), .RSTB(I136353), .Q(I136873) );
not I_7892 (I136890,I136873);
or I_7893 (I136907,I136890,I136811);
DFFARX1 I_7894  ( .D(I136907), .CLK(I2702), .RSTB(I136353), .Q(I136336) );
nand I_7895 (I136345,I136890,I136616);
DFFARX1 I_7896  ( .D(I136890), .CLK(I2702), .RSTB(I136353), .Q(I136315) );
not I_7897 (I136999,I2709);
not I_7898 (I137016,I516751);
nor I_7899 (I137033,I516727,I516733);
nand I_7900 (I137050,I137033,I516736);
DFFARX1 I_7901  ( .D(I137050), .CLK(I2702), .RSTB(I136999), .Q(I136973) );
nor I_7902 (I137081,I137016,I516727);
nand I_7903 (I137098,I137081,I516745);
not I_7904 (I136988,I137098);
DFFARX1 I_7905  ( .D(I137098), .CLK(I2702), .RSTB(I136999), .Q(I136970) );
not I_7906 (I137143,I516727);
not I_7907 (I137160,I137143);
not I_7908 (I137177,I516724);
nor I_7909 (I137194,I137177,I516739);
and I_7910 (I137211,I137194,I516730);
or I_7911 (I137228,I137211,I516742);
DFFARX1 I_7912  ( .D(I137228), .CLK(I2702), .RSTB(I136999), .Q(I137245) );
nor I_7913 (I137262,I137245,I137098);
nor I_7914 (I137279,I137245,I137160);
nand I_7915 (I136985,I137050,I137279);
nand I_7916 (I137310,I137016,I516724);
nand I_7917 (I137327,I137310,I137245);
and I_7918 (I137344,I137310,I137327);
DFFARX1 I_7919  ( .D(I137344), .CLK(I2702), .RSTB(I136999), .Q(I136967) );
DFFARX1 I_7920  ( .D(I137310), .CLK(I2702), .RSTB(I136999), .Q(I137375) );
and I_7921 (I136964,I137143,I137375);
DFFARX1 I_7922  ( .D(I516754), .CLK(I2702), .RSTB(I136999), .Q(I137406) );
not I_7923 (I137423,I137406);
nor I_7924 (I137440,I137098,I137423);
and I_7925 (I137457,I137406,I137440);
nand I_7926 (I136979,I137406,I137160);
DFFARX1 I_7927  ( .D(I137406), .CLK(I2702), .RSTB(I136999), .Q(I137488) );
not I_7928 (I136976,I137488);
DFFARX1 I_7929  ( .D(I516748), .CLK(I2702), .RSTB(I136999), .Q(I137519) );
not I_7930 (I137536,I137519);
or I_7931 (I137553,I137536,I137457);
DFFARX1 I_7932  ( .D(I137553), .CLK(I2702), .RSTB(I136999), .Q(I136982) );
nand I_7933 (I136991,I137536,I137262);
DFFARX1 I_7934  ( .D(I137536), .CLK(I2702), .RSTB(I136999), .Q(I136961) );
not I_7935 (I137645,I2709);
not I_7936 (I137662,I671543);
nor I_7937 (I137679,I671558,I671573);
nand I_7938 (I137696,I137679,I671561);
DFFARX1 I_7939  ( .D(I137696), .CLK(I2702), .RSTB(I137645), .Q(I137619) );
nor I_7940 (I137727,I137662,I671558);
nand I_7941 (I137744,I137727,I671564);
not I_7942 (I137634,I137744);
DFFARX1 I_7943  ( .D(I137744), .CLK(I2702), .RSTB(I137645), .Q(I137616) );
not I_7944 (I137789,I671558);
not I_7945 (I137806,I137789);
not I_7946 (I137823,I671570);
nor I_7947 (I137840,I137823,I671567);
and I_7948 (I137857,I137840,I671546);
or I_7949 (I137874,I137857,I671555);
DFFARX1 I_7950  ( .D(I137874), .CLK(I2702), .RSTB(I137645), .Q(I137891) );
nor I_7951 (I137908,I137891,I137744);
nor I_7952 (I137925,I137891,I137806);
nand I_7953 (I137631,I137696,I137925);
nand I_7954 (I137956,I137662,I671570);
nand I_7955 (I137973,I137956,I137891);
and I_7956 (I137990,I137956,I137973);
DFFARX1 I_7957  ( .D(I137990), .CLK(I2702), .RSTB(I137645), .Q(I137613) );
DFFARX1 I_7958  ( .D(I137956), .CLK(I2702), .RSTB(I137645), .Q(I138021) );
and I_7959 (I137610,I137789,I138021);
DFFARX1 I_7960  ( .D(I671552), .CLK(I2702), .RSTB(I137645), .Q(I138052) );
not I_7961 (I138069,I138052);
nor I_7962 (I138086,I137744,I138069);
and I_7963 (I138103,I138052,I138086);
nand I_7964 (I137625,I138052,I137806);
DFFARX1 I_7965  ( .D(I138052), .CLK(I2702), .RSTB(I137645), .Q(I138134) );
not I_7966 (I137622,I138134);
DFFARX1 I_7967  ( .D(I671549), .CLK(I2702), .RSTB(I137645), .Q(I138165) );
not I_7968 (I138182,I138165);
or I_7969 (I138199,I138182,I138103);
DFFARX1 I_7970  ( .D(I138199), .CLK(I2702), .RSTB(I137645), .Q(I137628) );
nand I_7971 (I137637,I138182,I137908);
DFFARX1 I_7972  ( .D(I138182), .CLK(I2702), .RSTB(I137645), .Q(I137607) );
not I_7973 (I138291,I2709);
not I_7974 (I138308,I300672);
nor I_7975 (I138325,I300669,I300657);
nand I_7976 (I138342,I138325,I300660);
DFFARX1 I_7977  ( .D(I138342), .CLK(I2702), .RSTB(I138291), .Q(I138265) );
nor I_7978 (I138373,I138308,I300669);
nand I_7979 (I138390,I138373,I300666);
not I_7980 (I138280,I138390);
DFFARX1 I_7981  ( .D(I138390), .CLK(I2702), .RSTB(I138291), .Q(I138262) );
not I_7982 (I138435,I300669);
not I_7983 (I138452,I138435);
not I_7984 (I138469,I300678);
nor I_7985 (I138486,I138469,I300654);
and I_7986 (I138503,I138486,I300675);
or I_7987 (I138520,I138503,I300663);
DFFARX1 I_7988  ( .D(I138520), .CLK(I2702), .RSTB(I138291), .Q(I138537) );
nor I_7989 (I138554,I138537,I138390);
nor I_7990 (I138571,I138537,I138452);
nand I_7991 (I138277,I138342,I138571);
nand I_7992 (I138602,I138308,I300678);
nand I_7993 (I138619,I138602,I138537);
and I_7994 (I138636,I138602,I138619);
DFFARX1 I_7995  ( .D(I138636), .CLK(I2702), .RSTB(I138291), .Q(I138259) );
DFFARX1 I_7996  ( .D(I138602), .CLK(I2702), .RSTB(I138291), .Q(I138667) );
and I_7997 (I138256,I138435,I138667);
DFFARX1 I_7998  ( .D(I300684), .CLK(I2702), .RSTB(I138291), .Q(I138698) );
not I_7999 (I138715,I138698);
nor I_8000 (I138732,I138390,I138715);
and I_8001 (I138749,I138698,I138732);
nand I_8002 (I138271,I138698,I138452);
DFFARX1 I_8003  ( .D(I138698), .CLK(I2702), .RSTB(I138291), .Q(I138780) );
not I_8004 (I138268,I138780);
DFFARX1 I_8005  ( .D(I300681), .CLK(I2702), .RSTB(I138291), .Q(I138811) );
not I_8006 (I138828,I138811);
or I_8007 (I138845,I138828,I138749);
DFFARX1 I_8008  ( .D(I138845), .CLK(I2702), .RSTB(I138291), .Q(I138274) );
nand I_8009 (I138283,I138828,I138554);
DFFARX1 I_8010  ( .D(I138828), .CLK(I2702), .RSTB(I138291), .Q(I138253) );
not I_8011 (I138937,I2709);
not I_8012 (I138954,I49278);
nor I_8013 (I138971,I49290,I49275);
nand I_8014 (I138988,I138971,I49287);
DFFARX1 I_8015  ( .D(I138988), .CLK(I2702), .RSTB(I138937), .Q(I138911) );
nor I_8016 (I139019,I138954,I49290);
nand I_8017 (I139036,I139019,I49305);
not I_8018 (I138926,I139036);
DFFARX1 I_8019  ( .D(I139036), .CLK(I2702), .RSTB(I138937), .Q(I138908) );
not I_8020 (I139081,I49290);
not I_8021 (I139098,I139081);
not I_8022 (I139115,I49281);
nor I_8023 (I139132,I139115,I49293);
and I_8024 (I139149,I139132,I49284);
or I_8025 (I139166,I139149,I49299);
DFFARX1 I_8026  ( .D(I139166), .CLK(I2702), .RSTB(I138937), .Q(I139183) );
nor I_8027 (I139200,I139183,I139036);
nor I_8028 (I139217,I139183,I139098);
nand I_8029 (I138923,I138988,I139217);
nand I_8030 (I139248,I138954,I49281);
nand I_8031 (I139265,I139248,I139183);
and I_8032 (I139282,I139248,I139265);
DFFARX1 I_8033  ( .D(I139282), .CLK(I2702), .RSTB(I138937), .Q(I138905) );
DFFARX1 I_8034  ( .D(I139248), .CLK(I2702), .RSTB(I138937), .Q(I139313) );
and I_8035 (I138902,I139081,I139313);
DFFARX1 I_8036  ( .D(I49302), .CLK(I2702), .RSTB(I138937), .Q(I139344) );
not I_8037 (I139361,I139344);
nor I_8038 (I139378,I139036,I139361);
and I_8039 (I139395,I139344,I139378);
nand I_8040 (I138917,I139344,I139098);
DFFARX1 I_8041  ( .D(I139344), .CLK(I2702), .RSTB(I138937), .Q(I139426) );
not I_8042 (I138914,I139426);
DFFARX1 I_8043  ( .D(I49296), .CLK(I2702), .RSTB(I138937), .Q(I139457) );
not I_8044 (I139474,I139457);
or I_8045 (I139491,I139474,I139395);
DFFARX1 I_8046  ( .D(I139491), .CLK(I2702), .RSTB(I138937), .Q(I138920) );
nand I_8047 (I138929,I139474,I139200);
DFFARX1 I_8048  ( .D(I139474), .CLK(I2702), .RSTB(I138937), .Q(I138899) );
not I_8049 (I139583,I2709);
not I_8050 (I139600,I528044);
nor I_8051 (I139617,I528056,I528059);
nand I_8052 (I139634,I139617,I528047);
DFFARX1 I_8053  ( .D(I139634), .CLK(I2702), .RSTB(I139583), .Q(I139554) );
nor I_8054 (I139665,I139600,I528056);
nand I_8055 (I139682,I139665,I528032);
nand I_8056 (I139699,I139682,I139634);
not I_8057 (I139716,I528056);
not I_8058 (I139733,I528035);
nor I_8059 (I139750,I139733,I528038);
and I_8060 (I139767,I139750,I528041);
or I_8061 (I139784,I139767,I528050);
DFFARX1 I_8062  ( .D(I139784), .CLK(I2702), .RSTB(I139583), .Q(I139801) );
nor I_8063 (I139818,I139801,I139682);
nand I_8064 (I139569,I139716,I139818);
not I_8065 (I139566,I139801);
and I_8066 (I139863,I139801,I139699);
DFFARX1 I_8067  ( .D(I139863), .CLK(I2702), .RSTB(I139583), .Q(I139551) );
DFFARX1 I_8068  ( .D(I139801), .CLK(I2702), .RSTB(I139583), .Q(I139894) );
and I_8069 (I139548,I139716,I139894);
nand I_8070 (I139925,I139600,I528035);
not I_8071 (I139942,I139925);
nor I_8072 (I139959,I139801,I139942);
DFFARX1 I_8073  ( .D(I528053), .CLK(I2702), .RSTB(I139583), .Q(I139976) );
nand I_8074 (I139993,I139976,I139925);
and I_8075 (I140010,I139716,I139993);
DFFARX1 I_8076  ( .D(I140010), .CLK(I2702), .RSTB(I139583), .Q(I139575) );
not I_8077 (I140041,I139976);
nand I_8078 (I139563,I139976,I139959);
nand I_8079 (I139557,I139976,I139942);
DFFARX1 I_8080  ( .D(I528029), .CLK(I2702), .RSTB(I139583), .Q(I140086) );
not I_8081 (I140103,I140086);
nor I_8082 (I139572,I139976,I140103);
nor I_8083 (I140134,I140103,I140041);
and I_8084 (I140151,I139682,I140134);
or I_8085 (I140168,I139925,I140151);
DFFARX1 I_8086  ( .D(I140168), .CLK(I2702), .RSTB(I139583), .Q(I139560) );
DFFARX1 I_8087  ( .D(I140103), .CLK(I2702), .RSTB(I139583), .Q(I139545) );
not I_8088 (I140246,I2709);
not I_8089 (I140263,I415025);
nor I_8090 (I140280,I415043,I415031);
nand I_8091 (I140297,I140280,I415037);
DFFARX1 I_8092  ( .D(I140297), .CLK(I2702), .RSTB(I140246), .Q(I140217) );
nor I_8093 (I140328,I140263,I415043);
nand I_8094 (I140345,I140328,I415040);
nand I_8095 (I140362,I140345,I140297);
not I_8096 (I140379,I415043);
not I_8097 (I140396,I415019);
nor I_8098 (I140413,I140396,I415013);
and I_8099 (I140430,I140413,I415022);
or I_8100 (I140447,I140430,I415034);
DFFARX1 I_8101  ( .D(I140447), .CLK(I2702), .RSTB(I140246), .Q(I140464) );
nor I_8102 (I140481,I140464,I140345);
nand I_8103 (I140232,I140379,I140481);
not I_8104 (I140229,I140464);
and I_8105 (I140526,I140464,I140362);
DFFARX1 I_8106  ( .D(I140526), .CLK(I2702), .RSTB(I140246), .Q(I140214) );
DFFARX1 I_8107  ( .D(I140464), .CLK(I2702), .RSTB(I140246), .Q(I140557) );
and I_8108 (I140211,I140379,I140557);
nand I_8109 (I140588,I140263,I415019);
not I_8110 (I140605,I140588);
nor I_8111 (I140622,I140464,I140605);
DFFARX1 I_8112  ( .D(I415028), .CLK(I2702), .RSTB(I140246), .Q(I140639) );
nand I_8113 (I140656,I140639,I140588);
and I_8114 (I140673,I140379,I140656);
DFFARX1 I_8115  ( .D(I140673), .CLK(I2702), .RSTB(I140246), .Q(I140238) );
not I_8116 (I140704,I140639);
nand I_8117 (I140226,I140639,I140622);
nand I_8118 (I140220,I140639,I140605);
DFFARX1 I_8119  ( .D(I415016), .CLK(I2702), .RSTB(I140246), .Q(I140749) );
not I_8120 (I140766,I140749);
nor I_8121 (I140235,I140639,I140766);
nor I_8122 (I140797,I140766,I140704);
and I_8123 (I140814,I140345,I140797);
or I_8124 (I140831,I140588,I140814);
DFFARX1 I_8125  ( .D(I140831), .CLK(I2702), .RSTB(I140246), .Q(I140223) );
DFFARX1 I_8126  ( .D(I140766), .CLK(I2702), .RSTB(I140246), .Q(I140208) );
not I_8127 (I140909,I2709);
not I_8128 (I140926,I494987);
nor I_8129 (I140943,I494993,I494984);
nand I_8130 (I140960,I140943,I495002);
DFFARX1 I_8131  ( .D(I140960), .CLK(I2702), .RSTB(I140909), .Q(I140880) );
nor I_8132 (I140991,I140926,I494993);
nand I_8133 (I141008,I140991,I494981);
nand I_8134 (I141025,I141008,I140960);
not I_8135 (I141042,I494993);
not I_8136 (I141059,I495011);
nor I_8137 (I141076,I141059,I494990);
and I_8138 (I141093,I141076,I494999);
or I_8139 (I141110,I141093,I495005);
DFFARX1 I_8140  ( .D(I141110), .CLK(I2702), .RSTB(I140909), .Q(I141127) );
nor I_8141 (I141144,I141127,I141008);
nand I_8142 (I140895,I141042,I141144);
not I_8143 (I140892,I141127);
and I_8144 (I141189,I141127,I141025);
DFFARX1 I_8145  ( .D(I141189), .CLK(I2702), .RSTB(I140909), .Q(I140877) );
DFFARX1 I_8146  ( .D(I141127), .CLK(I2702), .RSTB(I140909), .Q(I141220) );
and I_8147 (I140874,I141042,I141220);
nand I_8148 (I141251,I140926,I495011);
not I_8149 (I141268,I141251);
nor I_8150 (I141285,I141127,I141268);
DFFARX1 I_8151  ( .D(I494996), .CLK(I2702), .RSTB(I140909), .Q(I141302) );
nand I_8152 (I141319,I141302,I141251);
and I_8153 (I141336,I141042,I141319);
DFFARX1 I_8154  ( .D(I141336), .CLK(I2702), .RSTB(I140909), .Q(I140901) );
not I_8155 (I141367,I141302);
nand I_8156 (I140889,I141302,I141285);
nand I_8157 (I140883,I141302,I141268);
DFFARX1 I_8158  ( .D(I495008), .CLK(I2702), .RSTB(I140909), .Q(I141412) );
not I_8159 (I141429,I141412);
nor I_8160 (I140898,I141302,I141429);
nor I_8161 (I141460,I141429,I141367);
and I_8162 (I141477,I141008,I141460);
or I_8163 (I141494,I141251,I141477);
DFFARX1 I_8164  ( .D(I141494), .CLK(I2702), .RSTB(I140909), .Q(I140886) );
DFFARX1 I_8165  ( .D(I141429), .CLK(I2702), .RSTB(I140909), .Q(I140871) );
not I_8166 (I141572,I2709);
not I_8167 (I141589,I604790);
nor I_8168 (I141606,I604805,I604787);
nand I_8169 (I141623,I141606,I604799);
DFFARX1 I_8170  ( .D(I141623), .CLK(I2702), .RSTB(I141572), .Q(I141543) );
nor I_8171 (I141654,I141589,I604805);
nand I_8172 (I141671,I141654,I604796);
nand I_8173 (I141688,I141671,I141623);
not I_8174 (I141705,I604805);
not I_8175 (I141722,I604814);
nor I_8176 (I141739,I141722,I604784);
and I_8177 (I141756,I141739,I604793);
or I_8178 (I141773,I141756,I604811);
DFFARX1 I_8179  ( .D(I141773), .CLK(I2702), .RSTB(I141572), .Q(I141790) );
nor I_8180 (I141807,I141790,I141671);
nand I_8181 (I141558,I141705,I141807);
not I_8182 (I141555,I141790);
and I_8183 (I141852,I141790,I141688);
DFFARX1 I_8184  ( .D(I141852), .CLK(I2702), .RSTB(I141572), .Q(I141540) );
DFFARX1 I_8185  ( .D(I141790), .CLK(I2702), .RSTB(I141572), .Q(I141883) );
and I_8186 (I141537,I141705,I141883);
nand I_8187 (I141914,I141589,I604814);
not I_8188 (I141931,I141914);
nor I_8189 (I141948,I141790,I141931);
DFFARX1 I_8190  ( .D(I604802), .CLK(I2702), .RSTB(I141572), .Q(I141965) );
nand I_8191 (I141982,I141965,I141914);
and I_8192 (I141999,I141705,I141982);
DFFARX1 I_8193  ( .D(I141999), .CLK(I2702), .RSTB(I141572), .Q(I141564) );
not I_8194 (I142030,I141965);
nand I_8195 (I141552,I141965,I141948);
nand I_8196 (I141546,I141965,I141931);
DFFARX1 I_8197  ( .D(I604808), .CLK(I2702), .RSTB(I141572), .Q(I142075) );
not I_8198 (I142092,I142075);
nor I_8199 (I141561,I141965,I142092);
nor I_8200 (I142123,I142092,I142030);
and I_8201 (I142140,I141671,I142123);
or I_8202 (I142157,I141914,I142140);
DFFARX1 I_8203  ( .D(I142157), .CLK(I2702), .RSTB(I141572), .Q(I141549) );
DFFARX1 I_8204  ( .D(I142092), .CLK(I2702), .RSTB(I141572), .Q(I141534) );
not I_8205 (I142235,I2709);
not I_8206 (I142252,I503107);
nor I_8207 (I142269,I503119,I503122);
nand I_8208 (I142286,I142269,I503128);
DFFARX1 I_8209  ( .D(I142286), .CLK(I2702), .RSTB(I142235), .Q(I142206) );
nor I_8210 (I142317,I142252,I503119);
nand I_8211 (I142334,I142317,I503131);
nand I_8212 (I142351,I142334,I142286);
not I_8213 (I142368,I503119);
not I_8214 (I142385,I503110);
nor I_8215 (I142402,I142385,I503125);
and I_8216 (I142419,I142402,I503134);
or I_8217 (I142436,I142419,I503137);
DFFARX1 I_8218  ( .D(I142436), .CLK(I2702), .RSTB(I142235), .Q(I142453) );
nor I_8219 (I142470,I142453,I142334);
nand I_8220 (I142221,I142368,I142470);
not I_8221 (I142218,I142453);
and I_8222 (I142515,I142453,I142351);
DFFARX1 I_8223  ( .D(I142515), .CLK(I2702), .RSTB(I142235), .Q(I142203) );
DFFARX1 I_8224  ( .D(I142453), .CLK(I2702), .RSTB(I142235), .Q(I142546) );
and I_8225 (I142200,I142368,I142546);
nand I_8226 (I142577,I142252,I503110);
not I_8227 (I142594,I142577);
nor I_8228 (I142611,I142453,I142594);
DFFARX1 I_8229  ( .D(I503113), .CLK(I2702), .RSTB(I142235), .Q(I142628) );
nand I_8230 (I142645,I142628,I142577);
and I_8231 (I142662,I142368,I142645);
DFFARX1 I_8232  ( .D(I142662), .CLK(I2702), .RSTB(I142235), .Q(I142227) );
not I_8233 (I142693,I142628);
nand I_8234 (I142215,I142628,I142611);
nand I_8235 (I142209,I142628,I142594);
DFFARX1 I_8236  ( .D(I503116), .CLK(I2702), .RSTB(I142235), .Q(I142738) );
not I_8237 (I142755,I142738);
nor I_8238 (I142224,I142628,I142755);
nor I_8239 (I142786,I142755,I142693);
and I_8240 (I142803,I142334,I142786);
or I_8241 (I142820,I142577,I142803);
DFFARX1 I_8242  ( .D(I142820), .CLK(I2702), .RSTB(I142235), .Q(I142212) );
DFFARX1 I_8243  ( .D(I142755), .CLK(I2702), .RSTB(I142235), .Q(I142197) );
not I_8244 (I142898,I2709);
not I_8245 (I142915,I506624);
nor I_8246 (I142932,I506636,I506639);
nand I_8247 (I142949,I142932,I506627);
DFFARX1 I_8248  ( .D(I142949), .CLK(I2702), .RSTB(I142898), .Q(I142869) );
nor I_8249 (I142980,I142915,I506636);
nand I_8250 (I142997,I142980,I506612);
nand I_8251 (I143014,I142997,I142949);
not I_8252 (I143031,I506636);
not I_8253 (I143048,I506615);
nor I_8254 (I143065,I143048,I506618);
and I_8255 (I143082,I143065,I506621);
or I_8256 (I143099,I143082,I506630);
DFFARX1 I_8257  ( .D(I143099), .CLK(I2702), .RSTB(I142898), .Q(I143116) );
nor I_8258 (I143133,I143116,I142997);
nand I_8259 (I142884,I143031,I143133);
not I_8260 (I142881,I143116);
and I_8261 (I143178,I143116,I143014);
DFFARX1 I_8262  ( .D(I143178), .CLK(I2702), .RSTB(I142898), .Q(I142866) );
DFFARX1 I_8263  ( .D(I143116), .CLK(I2702), .RSTB(I142898), .Q(I143209) );
and I_8264 (I142863,I143031,I143209);
nand I_8265 (I143240,I142915,I506615);
not I_8266 (I143257,I143240);
nor I_8267 (I143274,I143116,I143257);
DFFARX1 I_8268  ( .D(I506633), .CLK(I2702), .RSTB(I142898), .Q(I143291) );
nand I_8269 (I143308,I143291,I143240);
and I_8270 (I143325,I143031,I143308);
DFFARX1 I_8271  ( .D(I143325), .CLK(I2702), .RSTB(I142898), .Q(I142890) );
not I_8272 (I143356,I143291);
nand I_8273 (I142878,I143291,I143274);
nand I_8274 (I142872,I143291,I143257);
DFFARX1 I_8275  ( .D(I506609), .CLK(I2702), .RSTB(I142898), .Q(I143401) );
not I_8276 (I143418,I143401);
nor I_8277 (I142887,I143291,I143418);
nor I_8278 (I143449,I143418,I143356);
and I_8279 (I143466,I142997,I143449);
or I_8280 (I143483,I143240,I143466);
DFFARX1 I_8281  ( .D(I143483), .CLK(I2702), .RSTB(I142898), .Q(I142875) );
DFFARX1 I_8282  ( .D(I143418), .CLK(I2702), .RSTB(I142898), .Q(I142860) );
not I_8283 (I143561,I2709);
not I_8284 (I143578,I84650);
nor I_8285 (I143595,I84638,I84662);
nand I_8286 (I143612,I143595,I84647);
DFFARX1 I_8287  ( .D(I143612), .CLK(I2702), .RSTB(I143561), .Q(I143532) );
nor I_8288 (I143643,I143578,I84638);
nand I_8289 (I143660,I143643,I84665);
nand I_8290 (I143677,I143660,I143612);
not I_8291 (I143694,I84638);
not I_8292 (I143711,I84635);
nor I_8293 (I143728,I143711,I84644);
and I_8294 (I143745,I143728,I84659);
or I_8295 (I143762,I143745,I84641);
DFFARX1 I_8296  ( .D(I143762), .CLK(I2702), .RSTB(I143561), .Q(I143779) );
nor I_8297 (I143796,I143779,I143660);
nand I_8298 (I143547,I143694,I143796);
not I_8299 (I143544,I143779);
and I_8300 (I143841,I143779,I143677);
DFFARX1 I_8301  ( .D(I143841), .CLK(I2702), .RSTB(I143561), .Q(I143529) );
DFFARX1 I_8302  ( .D(I143779), .CLK(I2702), .RSTB(I143561), .Q(I143872) );
and I_8303 (I143526,I143694,I143872);
nand I_8304 (I143903,I143578,I84635);
not I_8305 (I143920,I143903);
nor I_8306 (I143937,I143779,I143920);
DFFARX1 I_8307  ( .D(I84656), .CLK(I2702), .RSTB(I143561), .Q(I143954) );
nand I_8308 (I143971,I143954,I143903);
and I_8309 (I143988,I143694,I143971);
DFFARX1 I_8310  ( .D(I143988), .CLK(I2702), .RSTB(I143561), .Q(I143553) );
not I_8311 (I144019,I143954);
nand I_8312 (I143541,I143954,I143937);
nand I_8313 (I143535,I143954,I143920);
DFFARX1 I_8314  ( .D(I84653), .CLK(I2702), .RSTB(I143561), .Q(I144064) );
not I_8315 (I144081,I144064);
nor I_8316 (I143550,I143954,I144081);
nor I_8317 (I144112,I144081,I144019);
and I_8318 (I144129,I143660,I144112);
or I_8319 (I144146,I143903,I144129);
DFFARX1 I_8320  ( .D(I144146), .CLK(I2702), .RSTB(I143561), .Q(I143538) );
DFFARX1 I_8321  ( .D(I144081), .CLK(I2702), .RSTB(I143561), .Q(I143523) );
not I_8322 (I144224,I2709);
not I_8323 (I144241,I221917);
nor I_8324 (I144258,I221899,I221893);
nand I_8325 (I144275,I144258,I221896);
DFFARX1 I_8326  ( .D(I144275), .CLK(I2702), .RSTB(I144224), .Q(I144195) );
nor I_8327 (I144306,I144241,I221899);
nand I_8328 (I144323,I144306,I221905);
nand I_8329 (I144340,I144323,I144275);
not I_8330 (I144357,I221899);
not I_8331 (I144374,I221914);
nor I_8332 (I144391,I144374,I221902);
and I_8333 (I144408,I144391,I221908);
or I_8334 (I144425,I144408,I221923);
DFFARX1 I_8335  ( .D(I144425), .CLK(I2702), .RSTB(I144224), .Q(I144442) );
nor I_8336 (I144459,I144442,I144323);
nand I_8337 (I144210,I144357,I144459);
not I_8338 (I144207,I144442);
and I_8339 (I144504,I144442,I144340);
DFFARX1 I_8340  ( .D(I144504), .CLK(I2702), .RSTB(I144224), .Q(I144192) );
DFFARX1 I_8341  ( .D(I144442), .CLK(I2702), .RSTB(I144224), .Q(I144535) );
and I_8342 (I144189,I144357,I144535);
nand I_8343 (I144566,I144241,I221914);
not I_8344 (I144583,I144566);
nor I_8345 (I144600,I144442,I144583);
DFFARX1 I_8346  ( .D(I221911), .CLK(I2702), .RSTB(I144224), .Q(I144617) );
nand I_8347 (I144634,I144617,I144566);
and I_8348 (I144651,I144357,I144634);
DFFARX1 I_8349  ( .D(I144651), .CLK(I2702), .RSTB(I144224), .Q(I144216) );
not I_8350 (I144682,I144617);
nand I_8351 (I144204,I144617,I144600);
nand I_8352 (I144198,I144617,I144583);
DFFARX1 I_8353  ( .D(I221920), .CLK(I2702), .RSTB(I144224), .Q(I144727) );
not I_8354 (I144744,I144727);
nor I_8355 (I144213,I144617,I144744);
nor I_8356 (I144775,I144744,I144682);
and I_8357 (I144792,I144323,I144775);
or I_8358 (I144809,I144566,I144792);
DFFARX1 I_8359  ( .D(I144809), .CLK(I2702), .RSTB(I144224), .Q(I144201) );
DFFARX1 I_8360  ( .D(I144744), .CLK(I2702), .RSTB(I144224), .Q(I144186) );
not I_8361 (I144887,I2709);
not I_8362 (I144904,I338973);
nor I_8363 (I144921,I338982,I338955);
nand I_8364 (I144938,I144921,I338967);
DFFARX1 I_8365  ( .D(I144938), .CLK(I2702), .RSTB(I144887), .Q(I144858) );
nor I_8366 (I144969,I144904,I338982);
nand I_8367 (I144986,I144969,I338979);
nand I_8368 (I145003,I144986,I144938);
not I_8369 (I145020,I338982);
not I_8370 (I145037,I338958);
nor I_8371 (I145054,I145037,I338964);
and I_8372 (I145071,I145054,I338976);
or I_8373 (I145088,I145071,I338961);
DFFARX1 I_8374  ( .D(I145088), .CLK(I2702), .RSTB(I144887), .Q(I145105) );
nor I_8375 (I145122,I145105,I144986);
nand I_8376 (I144873,I145020,I145122);
not I_8377 (I144870,I145105);
and I_8378 (I145167,I145105,I145003);
DFFARX1 I_8379  ( .D(I145167), .CLK(I2702), .RSTB(I144887), .Q(I144855) );
DFFARX1 I_8380  ( .D(I145105), .CLK(I2702), .RSTB(I144887), .Q(I145198) );
and I_8381 (I144852,I145020,I145198);
nand I_8382 (I145229,I144904,I338958);
not I_8383 (I145246,I145229);
nor I_8384 (I145263,I145105,I145246);
DFFARX1 I_8385  ( .D(I338985), .CLK(I2702), .RSTB(I144887), .Q(I145280) );
nand I_8386 (I145297,I145280,I145229);
and I_8387 (I145314,I145020,I145297);
DFFARX1 I_8388  ( .D(I145314), .CLK(I2702), .RSTB(I144887), .Q(I144879) );
not I_8389 (I145345,I145280);
nand I_8390 (I144867,I145280,I145263);
nand I_8391 (I144861,I145280,I145246);
DFFARX1 I_8392  ( .D(I338970), .CLK(I2702), .RSTB(I144887), .Q(I145390) );
not I_8393 (I145407,I145390);
nor I_8394 (I144876,I145280,I145407);
nor I_8395 (I145438,I145407,I145345);
and I_8396 (I145455,I144986,I145438);
or I_8397 (I145472,I145229,I145455);
DFFARX1 I_8398  ( .D(I145472), .CLK(I2702), .RSTB(I144887), .Q(I144864) );
DFFARX1 I_8399  ( .D(I145407), .CLK(I2702), .RSTB(I144887), .Q(I144849) );
not I_8400 (I145550,I2709);
not I_8401 (I145567,I73668);
nor I_8402 (I145584,I73656,I73680);
nand I_8403 (I145601,I145584,I73665);
DFFARX1 I_8404  ( .D(I145601), .CLK(I2702), .RSTB(I145550), .Q(I145521) );
nor I_8405 (I145632,I145567,I73656);
nand I_8406 (I145649,I145632,I73683);
nand I_8407 (I145666,I145649,I145601);
not I_8408 (I145683,I73656);
not I_8409 (I145700,I73653);
nor I_8410 (I145717,I145700,I73662);
and I_8411 (I145734,I145717,I73677);
or I_8412 (I145751,I145734,I73659);
DFFARX1 I_8413  ( .D(I145751), .CLK(I2702), .RSTB(I145550), .Q(I145768) );
nor I_8414 (I145785,I145768,I145649);
nand I_8415 (I145536,I145683,I145785);
not I_8416 (I145533,I145768);
and I_8417 (I145830,I145768,I145666);
DFFARX1 I_8418  ( .D(I145830), .CLK(I2702), .RSTB(I145550), .Q(I145518) );
DFFARX1 I_8419  ( .D(I145768), .CLK(I2702), .RSTB(I145550), .Q(I145861) );
and I_8420 (I145515,I145683,I145861);
nand I_8421 (I145892,I145567,I73653);
not I_8422 (I145909,I145892);
nor I_8423 (I145926,I145768,I145909);
DFFARX1 I_8424  ( .D(I73674), .CLK(I2702), .RSTB(I145550), .Q(I145943) );
nand I_8425 (I145960,I145943,I145892);
and I_8426 (I145977,I145683,I145960);
DFFARX1 I_8427  ( .D(I145977), .CLK(I2702), .RSTB(I145550), .Q(I145542) );
not I_8428 (I146008,I145943);
nand I_8429 (I145530,I145943,I145926);
nand I_8430 (I145524,I145943,I145909);
DFFARX1 I_8431  ( .D(I73671), .CLK(I2702), .RSTB(I145550), .Q(I146053) );
not I_8432 (I146070,I146053);
nor I_8433 (I145539,I145943,I146070);
nor I_8434 (I146101,I146070,I146008);
and I_8435 (I146118,I145649,I146101);
or I_8436 (I146135,I145892,I146118);
DFFARX1 I_8437  ( .D(I146135), .CLK(I2702), .RSTB(I145550), .Q(I145527) );
DFFARX1 I_8438  ( .D(I146070), .CLK(I2702), .RSTB(I145550), .Q(I145512) );
not I_8439 (I146213,I2709);
not I_8440 (I146230,I62040);
nor I_8441 (I146247,I62028,I62052);
nand I_8442 (I146264,I146247,I62037);
DFFARX1 I_8443  ( .D(I146264), .CLK(I2702), .RSTB(I146213), .Q(I146184) );
nor I_8444 (I146295,I146230,I62028);
nand I_8445 (I146312,I146295,I62055);
nand I_8446 (I146329,I146312,I146264);
not I_8447 (I146346,I62028);
not I_8448 (I146363,I62025);
nor I_8449 (I146380,I146363,I62034);
and I_8450 (I146397,I146380,I62049);
or I_8451 (I146414,I146397,I62031);
DFFARX1 I_8452  ( .D(I146414), .CLK(I2702), .RSTB(I146213), .Q(I146431) );
nor I_8453 (I146448,I146431,I146312);
nand I_8454 (I146199,I146346,I146448);
not I_8455 (I146196,I146431);
and I_8456 (I146493,I146431,I146329);
DFFARX1 I_8457  ( .D(I146493), .CLK(I2702), .RSTB(I146213), .Q(I146181) );
DFFARX1 I_8458  ( .D(I146431), .CLK(I2702), .RSTB(I146213), .Q(I146524) );
and I_8459 (I146178,I146346,I146524);
nand I_8460 (I146555,I146230,I62025);
not I_8461 (I146572,I146555);
nor I_8462 (I146589,I146431,I146572);
DFFARX1 I_8463  ( .D(I62046), .CLK(I2702), .RSTB(I146213), .Q(I146606) );
nand I_8464 (I146623,I146606,I146555);
and I_8465 (I146640,I146346,I146623);
DFFARX1 I_8466  ( .D(I146640), .CLK(I2702), .RSTB(I146213), .Q(I146205) );
not I_8467 (I146671,I146606);
nand I_8468 (I146193,I146606,I146589);
nand I_8469 (I146187,I146606,I146572);
DFFARX1 I_8470  ( .D(I62043), .CLK(I2702), .RSTB(I146213), .Q(I146716) );
not I_8471 (I146733,I146716);
nor I_8472 (I146202,I146606,I146733);
nor I_8473 (I146764,I146733,I146671);
and I_8474 (I146781,I146312,I146764);
or I_8475 (I146798,I146555,I146781);
DFFARX1 I_8476  ( .D(I146798), .CLK(I2702), .RSTB(I146213), .Q(I146190) );
DFFARX1 I_8477  ( .D(I146733), .CLK(I2702), .RSTB(I146213), .Q(I146175) );
not I_8478 (I146876,I2709);
not I_8479 (I146893,I366105);
nor I_8480 (I146910,I366114,I366087);
nand I_8481 (I146927,I146910,I366099);
DFFARX1 I_8482  ( .D(I146927), .CLK(I2702), .RSTB(I146876), .Q(I146847) );
nor I_8483 (I146958,I146893,I366114);
nand I_8484 (I146975,I146958,I366111);
nand I_8485 (I146992,I146975,I146927);
not I_8486 (I147009,I366114);
not I_8487 (I147026,I366090);
nor I_8488 (I147043,I147026,I366096);
and I_8489 (I147060,I147043,I366108);
or I_8490 (I147077,I147060,I366093);
DFFARX1 I_8491  ( .D(I147077), .CLK(I2702), .RSTB(I146876), .Q(I147094) );
nor I_8492 (I147111,I147094,I146975);
nand I_8493 (I146862,I147009,I147111);
not I_8494 (I146859,I147094);
and I_8495 (I147156,I147094,I146992);
DFFARX1 I_8496  ( .D(I147156), .CLK(I2702), .RSTB(I146876), .Q(I146844) );
DFFARX1 I_8497  ( .D(I147094), .CLK(I2702), .RSTB(I146876), .Q(I147187) );
and I_8498 (I146841,I147009,I147187);
nand I_8499 (I147218,I146893,I366090);
not I_8500 (I147235,I147218);
nor I_8501 (I147252,I147094,I147235);
DFFARX1 I_8502  ( .D(I366117), .CLK(I2702), .RSTB(I146876), .Q(I147269) );
nand I_8503 (I147286,I147269,I147218);
and I_8504 (I147303,I147009,I147286);
DFFARX1 I_8505  ( .D(I147303), .CLK(I2702), .RSTB(I146876), .Q(I146868) );
not I_8506 (I147334,I147269);
nand I_8507 (I146856,I147269,I147252);
nand I_8508 (I146850,I147269,I147235);
DFFARX1 I_8509  ( .D(I366102), .CLK(I2702), .RSTB(I146876), .Q(I147379) );
not I_8510 (I147396,I147379);
nor I_8511 (I146865,I147269,I147396);
nor I_8512 (I147427,I147396,I147334);
and I_8513 (I147444,I146975,I147427);
or I_8514 (I147461,I147218,I147444);
DFFARX1 I_8515  ( .D(I147461), .CLK(I2702), .RSTB(I146876), .Q(I146853) );
DFFARX1 I_8516  ( .D(I147396), .CLK(I2702), .RSTB(I146876), .Q(I146838) );
not I_8517 (I147539,I2709);
not I_8518 (I147556,I520904);
nor I_8519 (I147573,I520916,I520919);
nand I_8520 (I147590,I147573,I520907);
DFFARX1 I_8521  ( .D(I147590), .CLK(I2702), .RSTB(I147539), .Q(I147510) );
nor I_8522 (I147621,I147556,I520916);
nand I_8523 (I147638,I147621,I520892);
nand I_8524 (I147655,I147638,I147590);
not I_8525 (I147672,I520916);
not I_8526 (I147689,I520895);
nor I_8527 (I147706,I147689,I520898);
and I_8528 (I147723,I147706,I520901);
or I_8529 (I147740,I147723,I520910);
DFFARX1 I_8530  ( .D(I147740), .CLK(I2702), .RSTB(I147539), .Q(I147757) );
nor I_8531 (I147774,I147757,I147638);
nand I_8532 (I147525,I147672,I147774);
not I_8533 (I147522,I147757);
and I_8534 (I147819,I147757,I147655);
DFFARX1 I_8535  ( .D(I147819), .CLK(I2702), .RSTB(I147539), .Q(I147507) );
DFFARX1 I_8536  ( .D(I147757), .CLK(I2702), .RSTB(I147539), .Q(I147850) );
and I_8537 (I147504,I147672,I147850);
nand I_8538 (I147881,I147556,I520895);
not I_8539 (I147898,I147881);
nor I_8540 (I147915,I147757,I147898);
DFFARX1 I_8541  ( .D(I520913), .CLK(I2702), .RSTB(I147539), .Q(I147932) );
nand I_8542 (I147949,I147932,I147881);
and I_8543 (I147966,I147672,I147949);
DFFARX1 I_8544  ( .D(I147966), .CLK(I2702), .RSTB(I147539), .Q(I147531) );
not I_8545 (I147997,I147932);
nand I_8546 (I147519,I147932,I147915);
nand I_8547 (I147513,I147932,I147898);
DFFARX1 I_8548  ( .D(I520889), .CLK(I2702), .RSTB(I147539), .Q(I148042) );
not I_8549 (I148059,I148042);
nor I_8550 (I147528,I147932,I148059);
nor I_8551 (I148090,I148059,I147997);
and I_8552 (I148107,I147638,I148090);
or I_8553 (I148124,I147881,I148107);
DFFARX1 I_8554  ( .D(I148124), .CLK(I2702), .RSTB(I147539), .Q(I147516) );
DFFARX1 I_8555  ( .D(I148059), .CLK(I2702), .RSTB(I147539), .Q(I147501) );
not I_8556 (I148202,I2709);
not I_8557 (I148219,I513764);
nor I_8558 (I148236,I513776,I513779);
nand I_8559 (I148253,I148236,I513767);
DFFARX1 I_8560  ( .D(I148253), .CLK(I2702), .RSTB(I148202), .Q(I148173) );
nor I_8561 (I148284,I148219,I513776);
nand I_8562 (I148301,I148284,I513752);
nand I_8563 (I148318,I148301,I148253);
not I_8564 (I148335,I513776);
not I_8565 (I148352,I513755);
nor I_8566 (I148369,I148352,I513758);
and I_8567 (I148386,I148369,I513761);
or I_8568 (I148403,I148386,I513770);
DFFARX1 I_8569  ( .D(I148403), .CLK(I2702), .RSTB(I148202), .Q(I148420) );
nor I_8570 (I148437,I148420,I148301);
nand I_8571 (I148188,I148335,I148437);
not I_8572 (I148185,I148420);
and I_8573 (I148482,I148420,I148318);
DFFARX1 I_8574  ( .D(I148482), .CLK(I2702), .RSTB(I148202), .Q(I148170) );
DFFARX1 I_8575  ( .D(I148420), .CLK(I2702), .RSTB(I148202), .Q(I148513) );
and I_8576 (I148167,I148335,I148513);
nand I_8577 (I148544,I148219,I513755);
not I_8578 (I148561,I148544);
nor I_8579 (I148578,I148420,I148561);
DFFARX1 I_8580  ( .D(I513773), .CLK(I2702), .RSTB(I148202), .Q(I148595) );
nand I_8581 (I148612,I148595,I148544);
and I_8582 (I148629,I148335,I148612);
DFFARX1 I_8583  ( .D(I148629), .CLK(I2702), .RSTB(I148202), .Q(I148194) );
not I_8584 (I148660,I148595);
nand I_8585 (I148182,I148595,I148578);
nand I_8586 (I148176,I148595,I148561);
DFFARX1 I_8587  ( .D(I513749), .CLK(I2702), .RSTB(I148202), .Q(I148705) );
not I_8588 (I148722,I148705);
nor I_8589 (I148191,I148595,I148722);
nor I_8590 (I148753,I148722,I148660);
and I_8591 (I148770,I148301,I148753);
or I_8592 (I148787,I148544,I148770);
DFFARX1 I_8593  ( .D(I148787), .CLK(I2702), .RSTB(I148202), .Q(I148179) );
DFFARX1 I_8594  ( .D(I148722), .CLK(I2702), .RSTB(I148202), .Q(I148164) );
not I_8595 (I148865,I2709);
not I_8596 (I148882,I386777);
nor I_8597 (I148899,I386786,I386759);
nand I_8598 (I148916,I148899,I386771);
DFFARX1 I_8599  ( .D(I148916), .CLK(I2702), .RSTB(I148865), .Q(I148836) );
nor I_8600 (I148947,I148882,I386786);
nand I_8601 (I148964,I148947,I386783);
nand I_8602 (I148981,I148964,I148916);
not I_8603 (I148998,I386786);
not I_8604 (I149015,I386762);
nor I_8605 (I149032,I149015,I386768);
and I_8606 (I149049,I149032,I386780);
or I_8607 (I149066,I149049,I386765);
DFFARX1 I_8608  ( .D(I149066), .CLK(I2702), .RSTB(I148865), .Q(I149083) );
nor I_8609 (I149100,I149083,I148964);
nand I_8610 (I148851,I148998,I149100);
not I_8611 (I148848,I149083);
and I_8612 (I149145,I149083,I148981);
DFFARX1 I_8613  ( .D(I149145), .CLK(I2702), .RSTB(I148865), .Q(I148833) );
DFFARX1 I_8614  ( .D(I149083), .CLK(I2702), .RSTB(I148865), .Q(I149176) );
and I_8615 (I148830,I148998,I149176);
nand I_8616 (I149207,I148882,I386762);
not I_8617 (I149224,I149207);
nor I_8618 (I149241,I149083,I149224);
DFFARX1 I_8619  ( .D(I386789), .CLK(I2702), .RSTB(I148865), .Q(I149258) );
nand I_8620 (I149275,I149258,I149207);
and I_8621 (I149292,I148998,I149275);
DFFARX1 I_8622  ( .D(I149292), .CLK(I2702), .RSTB(I148865), .Q(I148857) );
not I_8623 (I149323,I149258);
nand I_8624 (I148845,I149258,I149241);
nand I_8625 (I148839,I149258,I149224);
DFFARX1 I_8626  ( .D(I386774), .CLK(I2702), .RSTB(I148865), .Q(I149368) );
not I_8627 (I149385,I149368);
nor I_8628 (I148854,I149258,I149385);
nor I_8629 (I149416,I149385,I149323);
and I_8630 (I149433,I148964,I149416);
or I_8631 (I149450,I149207,I149433);
DFFARX1 I_8632  ( .D(I149450), .CLK(I2702), .RSTB(I148865), .Q(I148842) );
DFFARX1 I_8633  ( .D(I149385), .CLK(I2702), .RSTB(I148865), .Q(I148827) );
not I_8634 (I149528,I2709);
not I_8635 (I149545,I327174);
nor I_8636 (I149562,I327183,I327195);
nand I_8637 (I149579,I149562,I327186);
DFFARX1 I_8638  ( .D(I149579), .CLK(I2702), .RSTB(I149528), .Q(I149499) );
nor I_8639 (I149610,I149545,I327183);
nand I_8640 (I149627,I149610,I327198);
nand I_8641 (I149644,I149627,I149579);
not I_8642 (I149661,I327183);
not I_8643 (I149678,I327204);
nor I_8644 (I149695,I149678,I327180);
and I_8645 (I149712,I149695,I327189);
or I_8646 (I149729,I149712,I327177);
DFFARX1 I_8647  ( .D(I149729), .CLK(I2702), .RSTB(I149528), .Q(I149746) );
nor I_8648 (I149763,I149746,I149627);
nand I_8649 (I149514,I149661,I149763);
not I_8650 (I149511,I149746);
and I_8651 (I149808,I149746,I149644);
DFFARX1 I_8652  ( .D(I149808), .CLK(I2702), .RSTB(I149528), .Q(I149496) );
DFFARX1 I_8653  ( .D(I149746), .CLK(I2702), .RSTB(I149528), .Q(I149839) );
and I_8654 (I149493,I149661,I149839);
nand I_8655 (I149870,I149545,I327204);
not I_8656 (I149887,I149870);
nor I_8657 (I149904,I149746,I149887);
DFFARX1 I_8658  ( .D(I327201), .CLK(I2702), .RSTB(I149528), .Q(I149921) );
nand I_8659 (I149938,I149921,I149870);
and I_8660 (I149955,I149661,I149938);
DFFARX1 I_8661  ( .D(I149955), .CLK(I2702), .RSTB(I149528), .Q(I149520) );
not I_8662 (I149986,I149921);
nand I_8663 (I149508,I149921,I149904);
nand I_8664 (I149502,I149921,I149887);
DFFARX1 I_8665  ( .D(I327192), .CLK(I2702), .RSTB(I149528), .Q(I150031) );
not I_8666 (I150048,I150031);
nor I_8667 (I149517,I149921,I150048);
nor I_8668 (I150079,I150048,I149986);
and I_8669 (I150096,I149627,I150079);
or I_8670 (I150113,I149870,I150096);
DFFARX1 I_8671  ( .D(I150113), .CLK(I2702), .RSTB(I149528), .Q(I149505) );
DFFARX1 I_8672  ( .D(I150048), .CLK(I2702), .RSTB(I149528), .Q(I149490) );
not I_8673 (I150191,I2709);
not I_8674 (I150208,I475465);
nor I_8675 (I150225,I475471,I475468);
nand I_8676 (I150242,I150225,I475486);
DFFARX1 I_8677  ( .D(I150242), .CLK(I2702), .RSTB(I150191), .Q(I150162) );
nor I_8678 (I150273,I150208,I475471);
nand I_8679 (I150290,I150273,I475495);
nand I_8680 (I150307,I150290,I150242);
not I_8681 (I150324,I475471);
not I_8682 (I150341,I475489);
nor I_8683 (I150358,I150341,I475480);
and I_8684 (I150375,I150358,I475483);
or I_8685 (I150392,I150375,I475474);
DFFARX1 I_8686  ( .D(I150392), .CLK(I2702), .RSTB(I150191), .Q(I150409) );
nor I_8687 (I150426,I150409,I150290);
nand I_8688 (I150177,I150324,I150426);
not I_8689 (I150174,I150409);
and I_8690 (I150471,I150409,I150307);
DFFARX1 I_8691  ( .D(I150471), .CLK(I2702), .RSTB(I150191), .Q(I150159) );
DFFARX1 I_8692  ( .D(I150409), .CLK(I2702), .RSTB(I150191), .Q(I150502) );
and I_8693 (I150156,I150324,I150502);
nand I_8694 (I150533,I150208,I475489);
not I_8695 (I150550,I150533);
nor I_8696 (I150567,I150409,I150550);
DFFARX1 I_8697  ( .D(I475492), .CLK(I2702), .RSTB(I150191), .Q(I150584) );
nand I_8698 (I150601,I150584,I150533);
and I_8699 (I150618,I150324,I150601);
DFFARX1 I_8700  ( .D(I150618), .CLK(I2702), .RSTB(I150191), .Q(I150183) );
not I_8701 (I150649,I150584);
nand I_8702 (I150171,I150584,I150567);
nand I_8703 (I150165,I150584,I150550);
DFFARX1 I_8704  ( .D(I475477), .CLK(I2702), .RSTB(I150191), .Q(I150694) );
not I_8705 (I150711,I150694);
nor I_8706 (I150180,I150584,I150711);
nor I_8707 (I150742,I150711,I150649);
and I_8708 (I150759,I150290,I150742);
or I_8709 (I150776,I150533,I150759);
DFFARX1 I_8710  ( .D(I150776), .CLK(I2702), .RSTB(I150191), .Q(I150168) );
DFFARX1 I_8711  ( .D(I150711), .CLK(I2702), .RSTB(I150191), .Q(I150153) );
not I_8712 (I150854,I2709);
not I_8713 (I150871,I716974);
nor I_8714 (I150888,I716953,I716965);
nand I_8715 (I150905,I150888,I716959);
DFFARX1 I_8716  ( .D(I150905), .CLK(I2702), .RSTB(I150854), .Q(I150825) );
nor I_8717 (I150936,I150871,I716953);
nand I_8718 (I150953,I150936,I716980);
nand I_8719 (I150970,I150953,I150905);
not I_8720 (I150987,I716953);
not I_8721 (I151004,I716956);
nor I_8722 (I151021,I151004,I716968);
and I_8723 (I151038,I151021,I716971);
or I_8724 (I151055,I151038,I716977);
DFFARX1 I_8725  ( .D(I151055), .CLK(I2702), .RSTB(I150854), .Q(I151072) );
nor I_8726 (I151089,I151072,I150953);
nand I_8727 (I150840,I150987,I151089);
not I_8728 (I150837,I151072);
and I_8729 (I151134,I151072,I150970);
DFFARX1 I_8730  ( .D(I151134), .CLK(I2702), .RSTB(I150854), .Q(I150822) );
DFFARX1 I_8731  ( .D(I151072), .CLK(I2702), .RSTB(I150854), .Q(I151165) );
and I_8732 (I150819,I150987,I151165);
nand I_8733 (I151196,I150871,I716956);
not I_8734 (I151213,I151196);
nor I_8735 (I151230,I151072,I151213);
DFFARX1 I_8736  ( .D(I716950), .CLK(I2702), .RSTB(I150854), .Q(I151247) );
nand I_8737 (I151264,I151247,I151196);
and I_8738 (I151281,I150987,I151264);
DFFARX1 I_8739  ( .D(I151281), .CLK(I2702), .RSTB(I150854), .Q(I150846) );
not I_8740 (I151312,I151247);
nand I_8741 (I150834,I151247,I151230);
nand I_8742 (I150828,I151247,I151213);
DFFARX1 I_8743  ( .D(I716962), .CLK(I2702), .RSTB(I150854), .Q(I151357) );
not I_8744 (I151374,I151357);
nor I_8745 (I150843,I151247,I151374);
nor I_8746 (I151405,I151374,I151312);
and I_8747 (I151422,I150953,I151405);
or I_8748 (I151439,I151196,I151422);
DFFARX1 I_8749  ( .D(I151439), .CLK(I2702), .RSTB(I150854), .Q(I150831) );
DFFARX1 I_8750  ( .D(I151374), .CLK(I2702), .RSTB(I150854), .Q(I150816) );
not I_8751 (I151517,I2709);
not I_8752 (I151534,I529234);
nor I_8753 (I151551,I529246,I529249);
nand I_8754 (I151568,I151551,I529237);
DFFARX1 I_8755  ( .D(I151568), .CLK(I2702), .RSTB(I151517), .Q(I151488) );
nor I_8756 (I151599,I151534,I529246);
nand I_8757 (I151616,I151599,I529222);
nand I_8758 (I151633,I151616,I151568);
not I_8759 (I151650,I529246);
not I_8760 (I151667,I529225);
nor I_8761 (I151684,I151667,I529228);
and I_8762 (I151701,I151684,I529231);
or I_8763 (I151718,I151701,I529240);
DFFARX1 I_8764  ( .D(I151718), .CLK(I2702), .RSTB(I151517), .Q(I151735) );
nor I_8765 (I151752,I151735,I151616);
nand I_8766 (I151503,I151650,I151752);
not I_8767 (I151500,I151735);
and I_8768 (I151797,I151735,I151633);
DFFARX1 I_8769  ( .D(I151797), .CLK(I2702), .RSTB(I151517), .Q(I151485) );
DFFARX1 I_8770  ( .D(I151735), .CLK(I2702), .RSTB(I151517), .Q(I151828) );
and I_8771 (I151482,I151650,I151828);
nand I_8772 (I151859,I151534,I529225);
not I_8773 (I151876,I151859);
nor I_8774 (I151893,I151735,I151876);
DFFARX1 I_8775  ( .D(I529243), .CLK(I2702), .RSTB(I151517), .Q(I151910) );
nand I_8776 (I151927,I151910,I151859);
and I_8777 (I151944,I151650,I151927);
DFFARX1 I_8778  ( .D(I151944), .CLK(I2702), .RSTB(I151517), .Q(I151509) );
not I_8779 (I151975,I151910);
nand I_8780 (I151497,I151910,I151893);
nand I_8781 (I151491,I151910,I151876);
DFFARX1 I_8782  ( .D(I529219), .CLK(I2702), .RSTB(I151517), .Q(I152020) );
not I_8783 (I152037,I152020);
nor I_8784 (I151506,I151910,I152037);
nor I_8785 (I152068,I152037,I151975);
and I_8786 (I152085,I151616,I152068);
or I_8787 (I152102,I151859,I152085);
DFFARX1 I_8788  ( .D(I152102), .CLK(I2702), .RSTB(I151517), .Q(I151494) );
DFFARX1 I_8789  ( .D(I152037), .CLK(I2702), .RSTB(I151517), .Q(I151479) );
not I_8790 (I152180,I2709);
not I_8791 (I152197,I252918);
nor I_8792 (I152214,I252927,I252939);
nand I_8793 (I152231,I152214,I252930);
DFFARX1 I_8794  ( .D(I152231), .CLK(I2702), .RSTB(I152180), .Q(I152151) );
nor I_8795 (I152262,I152197,I252927);
nand I_8796 (I152279,I152262,I252942);
nand I_8797 (I152296,I152279,I152231);
not I_8798 (I152313,I252927);
not I_8799 (I152330,I252948);
nor I_8800 (I152347,I152330,I252924);
and I_8801 (I152364,I152347,I252933);
or I_8802 (I152381,I152364,I252921);
DFFARX1 I_8803  ( .D(I152381), .CLK(I2702), .RSTB(I152180), .Q(I152398) );
nor I_8804 (I152415,I152398,I152279);
nand I_8805 (I152166,I152313,I152415);
not I_8806 (I152163,I152398);
and I_8807 (I152460,I152398,I152296);
DFFARX1 I_8808  ( .D(I152460), .CLK(I2702), .RSTB(I152180), .Q(I152148) );
DFFARX1 I_8809  ( .D(I152398), .CLK(I2702), .RSTB(I152180), .Q(I152491) );
and I_8810 (I152145,I152313,I152491);
nand I_8811 (I152522,I152197,I252948);
not I_8812 (I152539,I152522);
nor I_8813 (I152556,I152398,I152539);
DFFARX1 I_8814  ( .D(I252945), .CLK(I2702), .RSTB(I152180), .Q(I152573) );
nand I_8815 (I152590,I152573,I152522);
and I_8816 (I152607,I152313,I152590);
DFFARX1 I_8817  ( .D(I152607), .CLK(I2702), .RSTB(I152180), .Q(I152172) );
not I_8818 (I152638,I152573);
nand I_8819 (I152160,I152573,I152556);
nand I_8820 (I152154,I152573,I152539);
DFFARX1 I_8821  ( .D(I252936), .CLK(I2702), .RSTB(I152180), .Q(I152683) );
not I_8822 (I152700,I152683);
nor I_8823 (I152169,I152573,I152700);
nor I_8824 (I152731,I152700,I152638);
and I_8825 (I152748,I152279,I152731);
or I_8826 (I152765,I152522,I152748);
DFFARX1 I_8827  ( .D(I152765), .CLK(I2702), .RSTB(I152180), .Q(I152157) );
DFFARX1 I_8828  ( .D(I152700), .CLK(I2702), .RSTB(I152180), .Q(I152142) );
not I_8829 (I152843,I2709);
not I_8830 (I152860,I251592);
nor I_8831 (I152877,I251601,I251613);
nand I_8832 (I152894,I152877,I251604);
DFFARX1 I_8833  ( .D(I152894), .CLK(I2702), .RSTB(I152843), .Q(I152814) );
nor I_8834 (I152925,I152860,I251601);
nand I_8835 (I152942,I152925,I251616);
nand I_8836 (I152959,I152942,I152894);
not I_8837 (I152976,I251601);
not I_8838 (I152993,I251622);
nor I_8839 (I153010,I152993,I251598);
and I_8840 (I153027,I153010,I251607);
or I_8841 (I153044,I153027,I251595);
DFFARX1 I_8842  ( .D(I153044), .CLK(I2702), .RSTB(I152843), .Q(I153061) );
nor I_8843 (I153078,I153061,I152942);
nand I_8844 (I152829,I152976,I153078);
not I_8845 (I152826,I153061);
and I_8846 (I153123,I153061,I152959);
DFFARX1 I_8847  ( .D(I153123), .CLK(I2702), .RSTB(I152843), .Q(I152811) );
DFFARX1 I_8848  ( .D(I153061), .CLK(I2702), .RSTB(I152843), .Q(I153154) );
and I_8849 (I152808,I152976,I153154);
nand I_8850 (I153185,I152860,I251622);
not I_8851 (I153202,I153185);
nor I_8852 (I153219,I153061,I153202);
DFFARX1 I_8853  ( .D(I251619), .CLK(I2702), .RSTB(I152843), .Q(I153236) );
nand I_8854 (I153253,I153236,I153185);
and I_8855 (I153270,I152976,I153253);
DFFARX1 I_8856  ( .D(I153270), .CLK(I2702), .RSTB(I152843), .Q(I152835) );
not I_8857 (I153301,I153236);
nand I_8858 (I152823,I153236,I153219);
nand I_8859 (I152817,I153236,I153202);
DFFARX1 I_8860  ( .D(I251610), .CLK(I2702), .RSTB(I152843), .Q(I153346) );
not I_8861 (I153363,I153346);
nor I_8862 (I152832,I153236,I153363);
nor I_8863 (I153394,I153363,I153301);
and I_8864 (I153411,I152942,I153394);
or I_8865 (I153428,I153185,I153411);
DFFARX1 I_8866  ( .D(I153428), .CLK(I2702), .RSTB(I152843), .Q(I152820) );
DFFARX1 I_8867  ( .D(I153363), .CLK(I2702), .RSTB(I152843), .Q(I152805) );
not I_8868 (I153506,I2709);
not I_8869 (I153523,I680990);
nor I_8870 (I153540,I680996,I681008);
nand I_8871 (I153557,I153540,I680999);
DFFARX1 I_8872  ( .D(I153557), .CLK(I2702), .RSTB(I153506), .Q(I153477) );
nor I_8873 (I153588,I153523,I680996);
nand I_8874 (I153605,I153588,I680978);
nand I_8875 (I153622,I153605,I153557);
not I_8876 (I153639,I680996);
not I_8877 (I153656,I680993);
nor I_8878 (I153673,I153656,I680981);
and I_8879 (I153690,I153673,I681002);
or I_8880 (I153707,I153690,I680984);
DFFARX1 I_8881  ( .D(I153707), .CLK(I2702), .RSTB(I153506), .Q(I153724) );
nor I_8882 (I153741,I153724,I153605);
nand I_8883 (I153492,I153639,I153741);
not I_8884 (I153489,I153724);
and I_8885 (I153786,I153724,I153622);
DFFARX1 I_8886  ( .D(I153786), .CLK(I2702), .RSTB(I153506), .Q(I153474) );
DFFARX1 I_8887  ( .D(I153724), .CLK(I2702), .RSTB(I153506), .Q(I153817) );
and I_8888 (I153471,I153639,I153817);
nand I_8889 (I153848,I153523,I680993);
not I_8890 (I153865,I153848);
nor I_8891 (I153882,I153724,I153865);
DFFARX1 I_8892  ( .D(I681005), .CLK(I2702), .RSTB(I153506), .Q(I153899) );
nand I_8893 (I153916,I153899,I153848);
and I_8894 (I153933,I153639,I153916);
DFFARX1 I_8895  ( .D(I153933), .CLK(I2702), .RSTB(I153506), .Q(I153498) );
not I_8896 (I153964,I153899);
nand I_8897 (I153486,I153899,I153882);
nand I_8898 (I153480,I153899,I153865);
DFFARX1 I_8899  ( .D(I680987), .CLK(I2702), .RSTB(I153506), .Q(I154009) );
not I_8900 (I154026,I154009);
nor I_8901 (I153495,I153899,I154026);
nor I_8902 (I154057,I154026,I153964);
and I_8903 (I154074,I153605,I154057);
or I_8904 (I154091,I153848,I154074);
DFFARX1 I_8905  ( .D(I154091), .CLK(I2702), .RSTB(I153506), .Q(I153483) );
DFFARX1 I_8906  ( .D(I154026), .CLK(I2702), .RSTB(I153506), .Q(I153468) );
not I_8907 (I154169,I2709);
not I_8908 (I154186,I713506);
nor I_8909 (I154203,I713485,I713497);
nand I_8910 (I154220,I154203,I713491);
DFFARX1 I_8911  ( .D(I154220), .CLK(I2702), .RSTB(I154169), .Q(I154140) );
nor I_8912 (I154251,I154186,I713485);
nand I_8913 (I154268,I154251,I713512);
nand I_8914 (I154285,I154268,I154220);
not I_8915 (I154302,I713485);
not I_8916 (I154319,I713488);
nor I_8917 (I154336,I154319,I713500);
and I_8918 (I154353,I154336,I713503);
or I_8919 (I154370,I154353,I713509);
DFFARX1 I_8920  ( .D(I154370), .CLK(I2702), .RSTB(I154169), .Q(I154387) );
nor I_8921 (I154404,I154387,I154268);
nand I_8922 (I154155,I154302,I154404);
not I_8923 (I154152,I154387);
and I_8924 (I154449,I154387,I154285);
DFFARX1 I_8925  ( .D(I154449), .CLK(I2702), .RSTB(I154169), .Q(I154137) );
DFFARX1 I_8926  ( .D(I154387), .CLK(I2702), .RSTB(I154169), .Q(I154480) );
and I_8927 (I154134,I154302,I154480);
nand I_8928 (I154511,I154186,I713488);
not I_8929 (I154528,I154511);
nor I_8930 (I154545,I154387,I154528);
DFFARX1 I_8931  ( .D(I713482), .CLK(I2702), .RSTB(I154169), .Q(I154562) );
nand I_8932 (I154579,I154562,I154511);
and I_8933 (I154596,I154302,I154579);
DFFARX1 I_8934  ( .D(I154596), .CLK(I2702), .RSTB(I154169), .Q(I154161) );
not I_8935 (I154627,I154562);
nand I_8936 (I154149,I154562,I154545);
nand I_8937 (I154143,I154562,I154528);
DFFARX1 I_8938  ( .D(I713494), .CLK(I2702), .RSTB(I154169), .Q(I154672) );
not I_8939 (I154689,I154672);
nor I_8940 (I154158,I154562,I154689);
nor I_8941 (I154720,I154689,I154627);
and I_8942 (I154737,I154268,I154720);
or I_8943 (I154754,I154511,I154737);
DFFARX1 I_8944  ( .D(I154754), .CLK(I2702), .RSTB(I154169), .Q(I154146) );
DFFARX1 I_8945  ( .D(I154689), .CLK(I2702), .RSTB(I154169), .Q(I154131) );
not I_8946 (I154832,I2709);
not I_8947 (I154849,I588725);
nor I_8948 (I154866,I588740,I588722);
nand I_8949 (I154883,I154866,I588734);
DFFARX1 I_8950  ( .D(I154883), .CLK(I2702), .RSTB(I154832), .Q(I154803) );
nor I_8951 (I154914,I154849,I588740);
nand I_8952 (I154931,I154914,I588731);
nand I_8953 (I154948,I154931,I154883);
not I_8954 (I154965,I588740);
not I_8955 (I154982,I588749);
nor I_8956 (I154999,I154982,I588719);
and I_8957 (I155016,I154999,I588728);
or I_8958 (I155033,I155016,I588746);
DFFARX1 I_8959  ( .D(I155033), .CLK(I2702), .RSTB(I154832), .Q(I155050) );
nor I_8960 (I155067,I155050,I154931);
nand I_8961 (I154818,I154965,I155067);
not I_8962 (I154815,I155050);
and I_8963 (I155112,I155050,I154948);
DFFARX1 I_8964  ( .D(I155112), .CLK(I2702), .RSTB(I154832), .Q(I154800) );
DFFARX1 I_8965  ( .D(I155050), .CLK(I2702), .RSTB(I154832), .Q(I155143) );
and I_8966 (I154797,I154965,I155143);
nand I_8967 (I155174,I154849,I588749);
not I_8968 (I155191,I155174);
nor I_8969 (I155208,I155050,I155191);
DFFARX1 I_8970  ( .D(I588737), .CLK(I2702), .RSTB(I154832), .Q(I155225) );
nand I_8971 (I155242,I155225,I155174);
and I_8972 (I155259,I154965,I155242);
DFFARX1 I_8973  ( .D(I155259), .CLK(I2702), .RSTB(I154832), .Q(I154824) );
not I_8974 (I155290,I155225);
nand I_8975 (I154812,I155225,I155208);
nand I_8976 (I154806,I155225,I155191);
DFFARX1 I_8977  ( .D(I588743), .CLK(I2702), .RSTB(I154832), .Q(I155335) );
not I_8978 (I155352,I155335);
nor I_8979 (I154821,I155225,I155352);
nor I_8980 (I155383,I155352,I155290);
and I_8981 (I155400,I154931,I155383);
or I_8982 (I155417,I155174,I155400);
DFFARX1 I_8983  ( .D(I155417), .CLK(I2702), .RSTB(I154832), .Q(I154809) );
DFFARX1 I_8984  ( .D(I155352), .CLK(I2702), .RSTB(I154832), .Q(I154794) );
not I_8985 (I155495,I2709);
not I_8986 (I155512,I100154);
nor I_8987 (I155529,I100142,I100166);
nand I_8988 (I155546,I155529,I100151);
DFFARX1 I_8989  ( .D(I155546), .CLK(I2702), .RSTB(I155495), .Q(I155466) );
nor I_8990 (I155577,I155512,I100142);
nand I_8991 (I155594,I155577,I100169);
nand I_8992 (I155611,I155594,I155546);
not I_8993 (I155628,I100142);
not I_8994 (I155645,I100139);
nor I_8995 (I155662,I155645,I100148);
and I_8996 (I155679,I155662,I100163);
or I_8997 (I155696,I155679,I100145);
DFFARX1 I_8998  ( .D(I155696), .CLK(I2702), .RSTB(I155495), .Q(I155713) );
nor I_8999 (I155730,I155713,I155594);
nand I_9000 (I155481,I155628,I155730);
not I_9001 (I155478,I155713);
and I_9002 (I155775,I155713,I155611);
DFFARX1 I_9003  ( .D(I155775), .CLK(I2702), .RSTB(I155495), .Q(I155463) );
DFFARX1 I_9004  ( .D(I155713), .CLK(I2702), .RSTB(I155495), .Q(I155806) );
and I_9005 (I155460,I155628,I155806);
nand I_9006 (I155837,I155512,I100139);
not I_9007 (I155854,I155837);
nor I_9008 (I155871,I155713,I155854);
DFFARX1 I_9009  ( .D(I100160), .CLK(I2702), .RSTB(I155495), .Q(I155888) );
nand I_9010 (I155905,I155888,I155837);
and I_9011 (I155922,I155628,I155905);
DFFARX1 I_9012  ( .D(I155922), .CLK(I2702), .RSTB(I155495), .Q(I155487) );
not I_9013 (I155953,I155888);
nand I_9014 (I155475,I155888,I155871);
nand I_9015 (I155469,I155888,I155854);
DFFARX1 I_9016  ( .D(I100157), .CLK(I2702), .RSTB(I155495), .Q(I155998) );
not I_9017 (I156015,I155998);
nor I_9018 (I155484,I155888,I156015);
nor I_9019 (I156046,I156015,I155953);
and I_9020 (I156063,I155594,I156046);
or I_9021 (I156080,I155837,I156063);
DFFARX1 I_9022  ( .D(I156080), .CLK(I2702), .RSTB(I155495), .Q(I155472) );
DFFARX1 I_9023  ( .D(I156015), .CLK(I2702), .RSTB(I155495), .Q(I155457) );
not I_9024 (I156158,I2709);
not I_9025 (I156175,I236780);
nor I_9026 (I156192,I236774,I236792);
nand I_9027 (I156209,I156192,I236768);
DFFARX1 I_9028  ( .D(I156209), .CLK(I2702), .RSTB(I156158), .Q(I156129) );
nor I_9029 (I156240,I156175,I236774);
nand I_9030 (I156257,I156240,I236783);
nand I_9031 (I156274,I156257,I156209);
not I_9032 (I156291,I236774);
not I_9033 (I156308,I236798);
nor I_9034 (I156325,I156308,I236789);
and I_9035 (I156342,I156325,I236777);
or I_9036 (I156359,I156342,I236795);
DFFARX1 I_9037  ( .D(I156359), .CLK(I2702), .RSTB(I156158), .Q(I156376) );
nor I_9038 (I156393,I156376,I156257);
nand I_9039 (I156144,I156291,I156393);
not I_9040 (I156141,I156376);
and I_9041 (I156438,I156376,I156274);
DFFARX1 I_9042  ( .D(I156438), .CLK(I2702), .RSTB(I156158), .Q(I156126) );
DFFARX1 I_9043  ( .D(I156376), .CLK(I2702), .RSTB(I156158), .Q(I156469) );
and I_9044 (I156123,I156291,I156469);
nand I_9045 (I156500,I156175,I236798);
not I_9046 (I156517,I156500);
nor I_9047 (I156534,I156376,I156517);
DFFARX1 I_9048  ( .D(I236786), .CLK(I2702), .RSTB(I156158), .Q(I156551) );
nand I_9049 (I156568,I156551,I156500);
and I_9050 (I156585,I156291,I156568);
DFFARX1 I_9051  ( .D(I156585), .CLK(I2702), .RSTB(I156158), .Q(I156150) );
not I_9052 (I156616,I156551);
nand I_9053 (I156138,I156551,I156534);
nand I_9054 (I156132,I156551,I156517);
DFFARX1 I_9055  ( .D(I236771), .CLK(I2702), .RSTB(I156158), .Q(I156661) );
not I_9056 (I156678,I156661);
nor I_9057 (I156147,I156551,I156678);
nor I_9058 (I156709,I156678,I156616);
and I_9059 (I156726,I156257,I156709);
or I_9060 (I156743,I156500,I156726);
DFFARX1 I_9061  ( .D(I156743), .CLK(I2702), .RSTB(I156158), .Q(I156135) );
DFFARX1 I_9062  ( .D(I156678), .CLK(I2702), .RSTB(I156158), .Q(I156120) );
not I_9063 (I156821,I2709);
not I_9064 (I156838,I683506);
nor I_9065 (I156855,I683512,I683524);
nand I_9066 (I156872,I156855,I683515);
DFFARX1 I_9067  ( .D(I156872), .CLK(I2702), .RSTB(I156821), .Q(I156792) );
nor I_9068 (I156903,I156838,I683512);
nand I_9069 (I156920,I156903,I683494);
nand I_9070 (I156937,I156920,I156872);
not I_9071 (I156954,I683512);
not I_9072 (I156971,I683509);
nor I_9073 (I156988,I156971,I683497);
and I_9074 (I157005,I156988,I683518);
or I_9075 (I157022,I157005,I683500);
DFFARX1 I_9076  ( .D(I157022), .CLK(I2702), .RSTB(I156821), .Q(I157039) );
nor I_9077 (I157056,I157039,I156920);
nand I_9078 (I156807,I156954,I157056);
not I_9079 (I156804,I157039);
and I_9080 (I157101,I157039,I156937);
DFFARX1 I_9081  ( .D(I157101), .CLK(I2702), .RSTB(I156821), .Q(I156789) );
DFFARX1 I_9082  ( .D(I157039), .CLK(I2702), .RSTB(I156821), .Q(I157132) );
and I_9083 (I156786,I156954,I157132);
nand I_9084 (I157163,I156838,I683509);
not I_9085 (I157180,I157163);
nor I_9086 (I157197,I157039,I157180);
DFFARX1 I_9087  ( .D(I683521), .CLK(I2702), .RSTB(I156821), .Q(I157214) );
nand I_9088 (I157231,I157214,I157163);
and I_9089 (I157248,I156954,I157231);
DFFARX1 I_9090  ( .D(I157248), .CLK(I2702), .RSTB(I156821), .Q(I156813) );
not I_9091 (I157279,I157214);
nand I_9092 (I156801,I157214,I157197);
nand I_9093 (I156795,I157214,I157180);
DFFARX1 I_9094  ( .D(I683503), .CLK(I2702), .RSTB(I156821), .Q(I157324) );
not I_9095 (I157341,I157324);
nor I_9096 (I156810,I157214,I157341);
nor I_9097 (I157372,I157341,I157279);
and I_9098 (I157389,I156920,I157372);
or I_9099 (I157406,I157163,I157389);
DFFARX1 I_9100  ( .D(I157406), .CLK(I2702), .RSTB(I156821), .Q(I156798) );
DFFARX1 I_9101  ( .D(I157341), .CLK(I2702), .RSTB(I156821), .Q(I156783) );
not I_9102 (I157484,I2709);
not I_9103 (I157501,I657088);
nor I_9104 (I157518,I657094,I657106);
nand I_9105 (I157535,I157518,I657097);
DFFARX1 I_9106  ( .D(I157535), .CLK(I2702), .RSTB(I157484), .Q(I157455) );
nor I_9107 (I157566,I157501,I657094);
nand I_9108 (I157583,I157566,I657076);
nand I_9109 (I157600,I157583,I157535);
not I_9110 (I157617,I657094);
not I_9111 (I157634,I657091);
nor I_9112 (I157651,I157634,I657079);
and I_9113 (I157668,I157651,I657100);
or I_9114 (I157685,I157668,I657082);
DFFARX1 I_9115  ( .D(I157685), .CLK(I2702), .RSTB(I157484), .Q(I157702) );
nor I_9116 (I157719,I157702,I157583);
nand I_9117 (I157470,I157617,I157719);
not I_9118 (I157467,I157702);
and I_9119 (I157764,I157702,I157600);
DFFARX1 I_9120  ( .D(I157764), .CLK(I2702), .RSTB(I157484), .Q(I157452) );
DFFARX1 I_9121  ( .D(I157702), .CLK(I2702), .RSTB(I157484), .Q(I157795) );
and I_9122 (I157449,I157617,I157795);
nand I_9123 (I157826,I157501,I657091);
not I_9124 (I157843,I157826);
nor I_9125 (I157860,I157702,I157843);
DFFARX1 I_9126  ( .D(I657103), .CLK(I2702), .RSTB(I157484), .Q(I157877) );
nand I_9127 (I157894,I157877,I157826);
and I_9128 (I157911,I157617,I157894);
DFFARX1 I_9129  ( .D(I157911), .CLK(I2702), .RSTB(I157484), .Q(I157476) );
not I_9130 (I157942,I157877);
nand I_9131 (I157464,I157877,I157860);
nand I_9132 (I157458,I157877,I157843);
DFFARX1 I_9133  ( .D(I657085), .CLK(I2702), .RSTB(I157484), .Q(I157987) );
not I_9134 (I158004,I157987);
nor I_9135 (I157473,I157877,I158004);
nor I_9136 (I158035,I158004,I157942);
and I_9137 (I158052,I157583,I158035);
or I_9138 (I158069,I157826,I158052);
DFFARX1 I_9139  ( .D(I158069), .CLK(I2702), .RSTB(I157484), .Q(I157461) );
DFFARX1 I_9140  ( .D(I158004), .CLK(I2702), .RSTB(I157484), .Q(I157446) );
not I_9141 (I158147,I2709);
not I_9142 (I158164,I211802);
nor I_9143 (I158181,I211784,I211778);
nand I_9144 (I158198,I158181,I211781);
DFFARX1 I_9145  ( .D(I158198), .CLK(I2702), .RSTB(I158147), .Q(I158118) );
nor I_9146 (I158229,I158164,I211784);
nand I_9147 (I158246,I158229,I211790);
nand I_9148 (I158263,I158246,I158198);
not I_9149 (I158280,I211784);
not I_9150 (I158297,I211799);
nor I_9151 (I158314,I158297,I211787);
and I_9152 (I158331,I158314,I211793);
or I_9153 (I158348,I158331,I211808);
DFFARX1 I_9154  ( .D(I158348), .CLK(I2702), .RSTB(I158147), .Q(I158365) );
nor I_9155 (I158382,I158365,I158246);
nand I_9156 (I158133,I158280,I158382);
not I_9157 (I158130,I158365);
and I_9158 (I158427,I158365,I158263);
DFFARX1 I_9159  ( .D(I158427), .CLK(I2702), .RSTB(I158147), .Q(I158115) );
DFFARX1 I_9160  ( .D(I158365), .CLK(I2702), .RSTB(I158147), .Q(I158458) );
and I_9161 (I158112,I158280,I158458);
nand I_9162 (I158489,I158164,I211799);
not I_9163 (I158506,I158489);
nor I_9164 (I158523,I158365,I158506);
DFFARX1 I_9165  ( .D(I211796), .CLK(I2702), .RSTB(I158147), .Q(I158540) );
nand I_9166 (I158557,I158540,I158489);
and I_9167 (I158574,I158280,I158557);
DFFARX1 I_9168  ( .D(I158574), .CLK(I2702), .RSTB(I158147), .Q(I158139) );
not I_9169 (I158605,I158540);
nand I_9170 (I158127,I158540,I158523);
nand I_9171 (I158121,I158540,I158506);
DFFARX1 I_9172  ( .D(I211805), .CLK(I2702), .RSTB(I158147), .Q(I158650) );
not I_9173 (I158667,I158650);
nor I_9174 (I158136,I158540,I158667);
nor I_9175 (I158698,I158667,I158605);
and I_9176 (I158715,I158246,I158698);
or I_9177 (I158732,I158489,I158715);
DFFARX1 I_9178  ( .D(I158732), .CLK(I2702), .RSTB(I158147), .Q(I158124) );
DFFARX1 I_9179  ( .D(I158667), .CLK(I2702), .RSTB(I158147), .Q(I158109) );
not I_9180 (I158810,I2709);
not I_9181 (I158827,I459859);
nor I_9182 (I158844,I459865,I459862);
nand I_9183 (I158861,I158844,I459880);
DFFARX1 I_9184  ( .D(I158861), .CLK(I2702), .RSTB(I158810), .Q(I158781) );
nor I_9185 (I158892,I158827,I459865);
nand I_9186 (I158909,I158892,I459889);
nand I_9187 (I158926,I158909,I158861);
not I_9188 (I158943,I459865);
not I_9189 (I158960,I459883);
nor I_9190 (I158977,I158960,I459874);
and I_9191 (I158994,I158977,I459877);
or I_9192 (I159011,I158994,I459868);
DFFARX1 I_9193  ( .D(I159011), .CLK(I2702), .RSTB(I158810), .Q(I159028) );
nor I_9194 (I159045,I159028,I158909);
nand I_9195 (I158796,I158943,I159045);
not I_9196 (I158793,I159028);
and I_9197 (I159090,I159028,I158926);
DFFARX1 I_9198  ( .D(I159090), .CLK(I2702), .RSTB(I158810), .Q(I158778) );
DFFARX1 I_9199  ( .D(I159028), .CLK(I2702), .RSTB(I158810), .Q(I159121) );
and I_9200 (I158775,I158943,I159121);
nand I_9201 (I159152,I158827,I459883);
not I_9202 (I159169,I159152);
nor I_9203 (I159186,I159028,I159169);
DFFARX1 I_9204  ( .D(I459886), .CLK(I2702), .RSTB(I158810), .Q(I159203) );
nand I_9205 (I159220,I159203,I159152);
and I_9206 (I159237,I158943,I159220);
DFFARX1 I_9207  ( .D(I159237), .CLK(I2702), .RSTB(I158810), .Q(I158802) );
not I_9208 (I159268,I159203);
nand I_9209 (I158790,I159203,I159186);
nand I_9210 (I158784,I159203,I159169);
DFFARX1 I_9211  ( .D(I459871), .CLK(I2702), .RSTB(I158810), .Q(I159313) );
not I_9212 (I159330,I159313);
nor I_9213 (I158799,I159203,I159330);
nor I_9214 (I159361,I159330,I159268);
and I_9215 (I159378,I158909,I159361);
or I_9216 (I159395,I159152,I159378);
DFFARX1 I_9217  ( .D(I159395), .CLK(I2702), .RSTB(I158810), .Q(I158787) );
DFFARX1 I_9218  ( .D(I159330), .CLK(I2702), .RSTB(I158810), .Q(I158772) );
not I_9219 (I159473,I2709);
not I_9220 (I159490,I516144);
nor I_9221 (I159507,I516156,I516159);
nand I_9222 (I159524,I159507,I516147);
DFFARX1 I_9223  ( .D(I159524), .CLK(I2702), .RSTB(I159473), .Q(I159444) );
nor I_9224 (I159555,I159490,I516156);
nand I_9225 (I159572,I159555,I516132);
nand I_9226 (I159589,I159572,I159524);
not I_9227 (I159606,I516156);
not I_9228 (I159623,I516135);
nor I_9229 (I159640,I159623,I516138);
and I_9230 (I159657,I159640,I516141);
or I_9231 (I159674,I159657,I516150);
DFFARX1 I_9232  ( .D(I159674), .CLK(I2702), .RSTB(I159473), .Q(I159691) );
nor I_9233 (I159708,I159691,I159572);
nand I_9234 (I159459,I159606,I159708);
not I_9235 (I159456,I159691);
and I_9236 (I159753,I159691,I159589);
DFFARX1 I_9237  ( .D(I159753), .CLK(I2702), .RSTB(I159473), .Q(I159441) );
DFFARX1 I_9238  ( .D(I159691), .CLK(I2702), .RSTB(I159473), .Q(I159784) );
and I_9239 (I159438,I159606,I159784);
nand I_9240 (I159815,I159490,I516135);
not I_9241 (I159832,I159815);
nor I_9242 (I159849,I159691,I159832);
DFFARX1 I_9243  ( .D(I516153), .CLK(I2702), .RSTB(I159473), .Q(I159866) );
nand I_9244 (I159883,I159866,I159815);
and I_9245 (I159900,I159606,I159883);
DFFARX1 I_9246  ( .D(I159900), .CLK(I2702), .RSTB(I159473), .Q(I159465) );
not I_9247 (I159931,I159866);
nand I_9248 (I159453,I159866,I159849);
nand I_9249 (I159447,I159866,I159832);
DFFARX1 I_9250  ( .D(I516129), .CLK(I2702), .RSTB(I159473), .Q(I159976) );
not I_9251 (I159993,I159976);
nor I_9252 (I159462,I159866,I159993);
nor I_9253 (I160024,I159993,I159931);
and I_9254 (I160041,I159572,I160024);
or I_9255 (I160058,I159815,I160041);
DFFARX1 I_9256  ( .D(I160058), .CLK(I2702), .RSTB(I159473), .Q(I159450) );
DFFARX1 I_9257  ( .D(I159993), .CLK(I2702), .RSTB(I159473), .Q(I159435) );
not I_9258 (I160136,I2709);
not I_9259 (I160153,I660862);
nor I_9260 (I160170,I660868,I660880);
nand I_9261 (I160187,I160170,I660871);
DFFARX1 I_9262  ( .D(I160187), .CLK(I2702), .RSTB(I160136), .Q(I160107) );
nor I_9263 (I160218,I160153,I660868);
nand I_9264 (I160235,I160218,I660850);
nand I_9265 (I160252,I160235,I160187);
not I_9266 (I160269,I660868);
not I_9267 (I160286,I660865);
nor I_9268 (I160303,I160286,I660853);
and I_9269 (I160320,I160303,I660874);
or I_9270 (I160337,I160320,I660856);
DFFARX1 I_9271  ( .D(I160337), .CLK(I2702), .RSTB(I160136), .Q(I160354) );
nor I_9272 (I160371,I160354,I160235);
nand I_9273 (I160122,I160269,I160371);
not I_9274 (I160119,I160354);
and I_9275 (I160416,I160354,I160252);
DFFARX1 I_9276  ( .D(I160416), .CLK(I2702), .RSTB(I160136), .Q(I160104) );
DFFARX1 I_9277  ( .D(I160354), .CLK(I2702), .RSTB(I160136), .Q(I160447) );
and I_9278 (I160101,I160269,I160447);
nand I_9279 (I160478,I160153,I660865);
not I_9280 (I160495,I160478);
nor I_9281 (I160512,I160354,I160495);
DFFARX1 I_9282  ( .D(I660877), .CLK(I2702), .RSTB(I160136), .Q(I160529) );
nand I_9283 (I160546,I160529,I160478);
and I_9284 (I160563,I160269,I160546);
DFFARX1 I_9285  ( .D(I160563), .CLK(I2702), .RSTB(I160136), .Q(I160128) );
not I_9286 (I160594,I160529);
nand I_9287 (I160116,I160529,I160512);
nand I_9288 (I160110,I160529,I160495);
DFFARX1 I_9289  ( .D(I660859), .CLK(I2702), .RSTB(I160136), .Q(I160639) );
not I_9290 (I160656,I160639);
nor I_9291 (I160125,I160529,I160656);
nor I_9292 (I160687,I160656,I160594);
and I_9293 (I160704,I160235,I160687);
or I_9294 (I160721,I160478,I160704);
DFFARX1 I_9295  ( .D(I160721), .CLK(I2702), .RSTB(I160136), .Q(I160113) );
DFFARX1 I_9296  ( .D(I160656), .CLK(I2702), .RSTB(I160136), .Q(I160098) );
not I_9297 (I160799,I2709);
not I_9298 (I160816,I93048);
nor I_9299 (I160833,I93036,I93060);
nand I_9300 (I160850,I160833,I93045);
DFFARX1 I_9301  ( .D(I160850), .CLK(I2702), .RSTB(I160799), .Q(I160770) );
nor I_9302 (I160881,I160816,I93036);
nand I_9303 (I160898,I160881,I93063);
nand I_9304 (I160915,I160898,I160850);
not I_9305 (I160932,I93036);
not I_9306 (I160949,I93033);
nor I_9307 (I160966,I160949,I93042);
and I_9308 (I160983,I160966,I93057);
or I_9309 (I161000,I160983,I93039);
DFFARX1 I_9310  ( .D(I161000), .CLK(I2702), .RSTB(I160799), .Q(I161017) );
nor I_9311 (I161034,I161017,I160898);
nand I_9312 (I160785,I160932,I161034);
not I_9313 (I160782,I161017);
and I_9314 (I161079,I161017,I160915);
DFFARX1 I_9315  ( .D(I161079), .CLK(I2702), .RSTB(I160799), .Q(I160767) );
DFFARX1 I_9316  ( .D(I161017), .CLK(I2702), .RSTB(I160799), .Q(I161110) );
and I_9317 (I160764,I160932,I161110);
nand I_9318 (I161141,I160816,I93033);
not I_9319 (I161158,I161141);
nor I_9320 (I161175,I161017,I161158);
DFFARX1 I_9321  ( .D(I93054), .CLK(I2702), .RSTB(I160799), .Q(I161192) );
nand I_9322 (I161209,I161192,I161141);
and I_9323 (I161226,I160932,I161209);
DFFARX1 I_9324  ( .D(I161226), .CLK(I2702), .RSTB(I160799), .Q(I160791) );
not I_9325 (I161257,I161192);
nand I_9326 (I160779,I161192,I161175);
nand I_9327 (I160773,I161192,I161158);
DFFARX1 I_9328  ( .D(I93051), .CLK(I2702), .RSTB(I160799), .Q(I161302) );
not I_9329 (I161319,I161302);
nor I_9330 (I160788,I161192,I161319);
nor I_9331 (I161350,I161319,I161257);
and I_9332 (I161367,I160898,I161350);
or I_9333 (I161384,I161141,I161367);
DFFARX1 I_9334  ( .D(I161384), .CLK(I2702), .RSTB(I160799), .Q(I160776) );
DFFARX1 I_9335  ( .D(I161319), .CLK(I2702), .RSTB(I160799), .Q(I160761) );
not I_9336 (I161462,I2709);
not I_9337 (I161479,I566719);
nor I_9338 (I161496,I566731,I566734);
nand I_9339 (I161513,I161496,I566722);
DFFARX1 I_9340  ( .D(I161513), .CLK(I2702), .RSTB(I161462), .Q(I161433) );
nor I_9341 (I161544,I161479,I566731);
nand I_9342 (I161561,I161544,I566707);
nand I_9343 (I161578,I161561,I161513);
not I_9344 (I161595,I566731);
not I_9345 (I161612,I566710);
nor I_9346 (I161629,I161612,I566713);
and I_9347 (I161646,I161629,I566716);
or I_9348 (I161663,I161646,I566725);
DFFARX1 I_9349  ( .D(I161663), .CLK(I2702), .RSTB(I161462), .Q(I161680) );
nor I_9350 (I161697,I161680,I161561);
nand I_9351 (I161448,I161595,I161697);
not I_9352 (I161445,I161680);
and I_9353 (I161742,I161680,I161578);
DFFARX1 I_9354  ( .D(I161742), .CLK(I2702), .RSTB(I161462), .Q(I161430) );
DFFARX1 I_9355  ( .D(I161680), .CLK(I2702), .RSTB(I161462), .Q(I161773) );
and I_9356 (I161427,I161595,I161773);
nand I_9357 (I161804,I161479,I566710);
not I_9358 (I161821,I161804);
nor I_9359 (I161838,I161680,I161821);
DFFARX1 I_9360  ( .D(I566728), .CLK(I2702), .RSTB(I161462), .Q(I161855) );
nand I_9361 (I161872,I161855,I161804);
and I_9362 (I161889,I161595,I161872);
DFFARX1 I_9363  ( .D(I161889), .CLK(I2702), .RSTB(I161462), .Q(I161454) );
not I_9364 (I161920,I161855);
nand I_9365 (I161442,I161855,I161838);
nand I_9366 (I161436,I161855,I161821);
DFFARX1 I_9367  ( .D(I566704), .CLK(I2702), .RSTB(I161462), .Q(I161965) );
not I_9368 (I161982,I161965);
nor I_9369 (I161451,I161855,I161982);
nor I_9370 (I162013,I161982,I161920);
and I_9371 (I162030,I161561,I162013);
or I_9372 (I162047,I161804,I162030);
DFFARX1 I_9373  ( .D(I162047), .CLK(I2702), .RSTB(I161462), .Q(I161439) );
DFFARX1 I_9374  ( .D(I161982), .CLK(I2702), .RSTB(I161462), .Q(I161424) );
not I_9375 (I162125,I2709);
not I_9376 (I162142,I11142);
nor I_9377 (I162159,I11130,I11133);
nand I_9378 (I162176,I162159,I11148);
DFFARX1 I_9379  ( .D(I162176), .CLK(I2702), .RSTB(I162125), .Q(I162096) );
nor I_9380 (I162207,I162142,I11130);
nand I_9381 (I162224,I162207,I11139);
nand I_9382 (I162241,I162224,I162176);
not I_9383 (I162258,I11130);
not I_9384 (I162275,I11151);
nor I_9385 (I162292,I162275,I11127);
and I_9386 (I162309,I162292,I11136);
or I_9387 (I162326,I162309,I11145);
DFFARX1 I_9388  ( .D(I162326), .CLK(I2702), .RSTB(I162125), .Q(I162343) );
nor I_9389 (I162360,I162343,I162224);
nand I_9390 (I162111,I162258,I162360);
not I_9391 (I162108,I162343);
and I_9392 (I162405,I162343,I162241);
DFFARX1 I_9393  ( .D(I162405), .CLK(I2702), .RSTB(I162125), .Q(I162093) );
DFFARX1 I_9394  ( .D(I162343), .CLK(I2702), .RSTB(I162125), .Q(I162436) );
and I_9395 (I162090,I162258,I162436);
nand I_9396 (I162467,I162142,I11151);
not I_9397 (I162484,I162467);
nor I_9398 (I162501,I162343,I162484);
DFFARX1 I_9399  ( .D(I11157), .CLK(I2702), .RSTB(I162125), .Q(I162518) );
nand I_9400 (I162535,I162518,I162467);
and I_9401 (I162552,I162258,I162535);
DFFARX1 I_9402  ( .D(I162552), .CLK(I2702), .RSTB(I162125), .Q(I162117) );
not I_9403 (I162583,I162518);
nand I_9404 (I162105,I162518,I162501);
nand I_9405 (I162099,I162518,I162484);
DFFARX1 I_9406  ( .D(I11154), .CLK(I2702), .RSTB(I162125), .Q(I162628) );
not I_9407 (I162645,I162628);
nor I_9408 (I162114,I162518,I162645);
nor I_9409 (I162676,I162645,I162583);
and I_9410 (I162693,I162224,I162676);
or I_9411 (I162710,I162467,I162693);
DFFARX1 I_9412  ( .D(I162710), .CLK(I2702), .RSTB(I162125), .Q(I162102) );
DFFARX1 I_9413  ( .D(I162645), .CLK(I2702), .RSTB(I162125), .Q(I162087) );
not I_9414 (I162788,I2709);
not I_9415 (I162805,I640105);
nor I_9416 (I162822,I640111,I640123);
nand I_9417 (I162839,I162822,I640114);
DFFARX1 I_9418  ( .D(I162839), .CLK(I2702), .RSTB(I162788), .Q(I162759) );
nor I_9419 (I162870,I162805,I640111);
nand I_9420 (I162887,I162870,I640093);
nand I_9421 (I162904,I162887,I162839);
not I_9422 (I162921,I640111);
not I_9423 (I162938,I640108);
nor I_9424 (I162955,I162938,I640096);
and I_9425 (I162972,I162955,I640117);
or I_9426 (I162989,I162972,I640099);
DFFARX1 I_9427  ( .D(I162989), .CLK(I2702), .RSTB(I162788), .Q(I163006) );
nor I_9428 (I163023,I163006,I162887);
nand I_9429 (I162774,I162921,I163023);
not I_9430 (I162771,I163006);
and I_9431 (I163068,I163006,I162904);
DFFARX1 I_9432  ( .D(I163068), .CLK(I2702), .RSTB(I162788), .Q(I162756) );
DFFARX1 I_9433  ( .D(I163006), .CLK(I2702), .RSTB(I162788), .Q(I163099) );
and I_9434 (I162753,I162921,I163099);
nand I_9435 (I163130,I162805,I640108);
not I_9436 (I163147,I163130);
nor I_9437 (I163164,I163006,I163147);
DFFARX1 I_9438  ( .D(I640120), .CLK(I2702), .RSTB(I162788), .Q(I163181) );
nand I_9439 (I163198,I163181,I163130);
and I_9440 (I163215,I162921,I163198);
DFFARX1 I_9441  ( .D(I163215), .CLK(I2702), .RSTB(I162788), .Q(I162780) );
not I_9442 (I163246,I163181);
nand I_9443 (I162768,I163181,I163164);
nand I_9444 (I162762,I163181,I163147);
DFFARX1 I_9445  ( .D(I640102), .CLK(I2702), .RSTB(I162788), .Q(I163291) );
not I_9446 (I163308,I163291);
nor I_9447 (I162777,I163181,I163308);
nor I_9448 (I163339,I163308,I163246);
and I_9449 (I163356,I162887,I163339);
or I_9450 (I163373,I163130,I163356);
DFFARX1 I_9451  ( .D(I163373), .CLK(I2702), .RSTB(I162788), .Q(I162765) );
DFFARX1 I_9452  ( .D(I163308), .CLK(I2702), .RSTB(I162788), .Q(I162750) );
not I_9453 (I163451,I2709);
not I_9454 (I163468,I367397);
nor I_9455 (I163485,I367406,I367379);
nand I_9456 (I163502,I163485,I367391);
DFFARX1 I_9457  ( .D(I163502), .CLK(I2702), .RSTB(I163451), .Q(I163422) );
nor I_9458 (I163533,I163468,I367406);
nand I_9459 (I163550,I163533,I367403);
nand I_9460 (I163567,I163550,I163502);
not I_9461 (I163584,I367406);
not I_9462 (I163601,I367382);
nor I_9463 (I163618,I163601,I367388);
and I_9464 (I163635,I163618,I367400);
or I_9465 (I163652,I163635,I367385);
DFFARX1 I_9466  ( .D(I163652), .CLK(I2702), .RSTB(I163451), .Q(I163669) );
nor I_9467 (I163686,I163669,I163550);
nand I_9468 (I163437,I163584,I163686);
not I_9469 (I163434,I163669);
and I_9470 (I163731,I163669,I163567);
DFFARX1 I_9471  ( .D(I163731), .CLK(I2702), .RSTB(I163451), .Q(I163419) );
DFFARX1 I_9472  ( .D(I163669), .CLK(I2702), .RSTB(I163451), .Q(I163762) );
and I_9473 (I163416,I163584,I163762);
nand I_9474 (I163793,I163468,I367382);
not I_9475 (I163810,I163793);
nor I_9476 (I163827,I163669,I163810);
DFFARX1 I_9477  ( .D(I367409), .CLK(I2702), .RSTB(I163451), .Q(I163844) );
nand I_9478 (I163861,I163844,I163793);
and I_9479 (I163878,I163584,I163861);
DFFARX1 I_9480  ( .D(I163878), .CLK(I2702), .RSTB(I163451), .Q(I163443) );
not I_9481 (I163909,I163844);
nand I_9482 (I163431,I163844,I163827);
nand I_9483 (I163425,I163844,I163810);
DFFARX1 I_9484  ( .D(I367394), .CLK(I2702), .RSTB(I163451), .Q(I163954) );
not I_9485 (I163971,I163954);
nor I_9486 (I163440,I163844,I163971);
nor I_9487 (I164002,I163971,I163909);
and I_9488 (I164019,I163550,I164002);
or I_9489 (I164036,I163793,I164019);
DFFARX1 I_9490  ( .D(I164036), .CLK(I2702), .RSTB(I163451), .Q(I163428) );
DFFARX1 I_9491  ( .D(I163971), .CLK(I2702), .RSTB(I163451), .Q(I163413) );
not I_9492 (I164114,I2709);
not I_9493 (I164131,I276123);
nor I_9494 (I164148,I276132,I276144);
nand I_9495 (I164165,I164148,I276135);
DFFARX1 I_9496  ( .D(I164165), .CLK(I2702), .RSTB(I164114), .Q(I164085) );
nor I_9497 (I164196,I164131,I276132);
nand I_9498 (I164213,I164196,I276147);
nand I_9499 (I164230,I164213,I164165);
not I_9500 (I164247,I276132);
not I_9501 (I164264,I276153);
nor I_9502 (I164281,I164264,I276129);
and I_9503 (I164298,I164281,I276138);
or I_9504 (I164315,I164298,I276126);
DFFARX1 I_9505  ( .D(I164315), .CLK(I2702), .RSTB(I164114), .Q(I164332) );
nor I_9506 (I164349,I164332,I164213);
nand I_9507 (I164100,I164247,I164349);
not I_9508 (I164097,I164332);
and I_9509 (I164394,I164332,I164230);
DFFARX1 I_9510  ( .D(I164394), .CLK(I2702), .RSTB(I164114), .Q(I164082) );
DFFARX1 I_9511  ( .D(I164332), .CLK(I2702), .RSTB(I164114), .Q(I164425) );
and I_9512 (I164079,I164247,I164425);
nand I_9513 (I164456,I164131,I276153);
not I_9514 (I164473,I164456);
nor I_9515 (I164490,I164332,I164473);
DFFARX1 I_9516  ( .D(I276150), .CLK(I2702), .RSTB(I164114), .Q(I164507) );
nand I_9517 (I164524,I164507,I164456);
and I_9518 (I164541,I164247,I164524);
DFFARX1 I_9519  ( .D(I164541), .CLK(I2702), .RSTB(I164114), .Q(I164106) );
not I_9520 (I164572,I164507);
nand I_9521 (I164094,I164507,I164490);
nand I_9522 (I164088,I164507,I164473);
DFFARX1 I_9523  ( .D(I276141), .CLK(I2702), .RSTB(I164114), .Q(I164617) );
not I_9524 (I164634,I164617);
nor I_9525 (I164103,I164507,I164634);
nor I_9526 (I164665,I164634,I164572);
and I_9527 (I164682,I164213,I164665);
or I_9528 (I164699,I164456,I164682);
DFFARX1 I_9529  ( .D(I164699), .CLK(I2702), .RSTB(I164114), .Q(I164091) );
DFFARX1 I_9530  ( .D(I164634), .CLK(I2702), .RSTB(I164114), .Q(I164076) );
not I_9531 (I164777,I2709);
not I_9532 (I164794,I42558);
nor I_9533 (I164811,I42546,I42549);
nand I_9534 (I164828,I164811,I42564);
DFFARX1 I_9535  ( .D(I164828), .CLK(I2702), .RSTB(I164777), .Q(I164748) );
nor I_9536 (I164859,I164794,I42546);
nand I_9537 (I164876,I164859,I42555);
nand I_9538 (I164893,I164876,I164828);
not I_9539 (I164910,I42546);
not I_9540 (I164927,I42567);
nor I_9541 (I164944,I164927,I42543);
and I_9542 (I164961,I164944,I42552);
or I_9543 (I164978,I164961,I42561);
DFFARX1 I_9544  ( .D(I164978), .CLK(I2702), .RSTB(I164777), .Q(I164995) );
nor I_9545 (I165012,I164995,I164876);
nand I_9546 (I164763,I164910,I165012);
not I_9547 (I164760,I164995);
and I_9548 (I165057,I164995,I164893);
DFFARX1 I_9549  ( .D(I165057), .CLK(I2702), .RSTB(I164777), .Q(I164745) );
DFFARX1 I_9550  ( .D(I164995), .CLK(I2702), .RSTB(I164777), .Q(I165088) );
and I_9551 (I164742,I164910,I165088);
nand I_9552 (I165119,I164794,I42567);
not I_9553 (I165136,I165119);
nor I_9554 (I165153,I164995,I165136);
DFFARX1 I_9555  ( .D(I42573), .CLK(I2702), .RSTB(I164777), .Q(I165170) );
nand I_9556 (I165187,I165170,I165119);
and I_9557 (I165204,I164910,I165187);
DFFARX1 I_9558  ( .D(I165204), .CLK(I2702), .RSTB(I164777), .Q(I164769) );
not I_9559 (I165235,I165170);
nand I_9560 (I164757,I165170,I165153);
nand I_9561 (I164751,I165170,I165136);
DFFARX1 I_9562  ( .D(I42570), .CLK(I2702), .RSTB(I164777), .Q(I165280) );
not I_9563 (I165297,I165280);
nor I_9564 (I164766,I165170,I165297);
nor I_9565 (I165328,I165297,I165235);
and I_9566 (I165345,I164876,I165328);
or I_9567 (I165362,I165119,I165345);
DFFARX1 I_9568  ( .D(I165362), .CLK(I2702), .RSTB(I164777), .Q(I164754) );
DFFARX1 I_9569  ( .D(I165297), .CLK(I2702), .RSTB(I164777), .Q(I164739) );
not I_9570 (I165440,I2709);
not I_9571 (I165457,I657717);
nor I_9572 (I165474,I657723,I657735);
nand I_9573 (I165491,I165474,I657726);
DFFARX1 I_9574  ( .D(I165491), .CLK(I2702), .RSTB(I165440), .Q(I165411) );
nor I_9575 (I165522,I165457,I657723);
nand I_9576 (I165539,I165522,I657705);
nand I_9577 (I165556,I165539,I165491);
not I_9578 (I165573,I657723);
not I_9579 (I165590,I657720);
nor I_9580 (I165607,I165590,I657708);
and I_9581 (I165624,I165607,I657729);
or I_9582 (I165641,I165624,I657711);
DFFARX1 I_9583  ( .D(I165641), .CLK(I2702), .RSTB(I165440), .Q(I165658) );
nor I_9584 (I165675,I165658,I165539);
nand I_9585 (I165426,I165573,I165675);
not I_9586 (I165423,I165658);
and I_9587 (I165720,I165658,I165556);
DFFARX1 I_9588  ( .D(I165720), .CLK(I2702), .RSTB(I165440), .Q(I165408) );
DFFARX1 I_9589  ( .D(I165658), .CLK(I2702), .RSTB(I165440), .Q(I165751) );
and I_9590 (I165405,I165573,I165751);
nand I_9591 (I165782,I165457,I657720);
not I_9592 (I165799,I165782);
nor I_9593 (I165816,I165658,I165799);
DFFARX1 I_9594  ( .D(I657732), .CLK(I2702), .RSTB(I165440), .Q(I165833) );
nand I_9595 (I165850,I165833,I165782);
and I_9596 (I165867,I165573,I165850);
DFFARX1 I_9597  ( .D(I165867), .CLK(I2702), .RSTB(I165440), .Q(I165432) );
not I_9598 (I165898,I165833);
nand I_9599 (I165420,I165833,I165816);
nand I_9600 (I165414,I165833,I165799);
DFFARX1 I_9601  ( .D(I657714), .CLK(I2702), .RSTB(I165440), .Q(I165943) );
not I_9602 (I165960,I165943);
nor I_9603 (I165429,I165833,I165960);
nor I_9604 (I165991,I165960,I165898);
and I_9605 (I166008,I165539,I165991);
or I_9606 (I166025,I165782,I166008);
DFFARX1 I_9607  ( .D(I166025), .CLK(I2702), .RSTB(I165440), .Q(I165417) );
DFFARX1 I_9608  ( .D(I165960), .CLK(I2702), .RSTB(I165440), .Q(I165402) );
not I_9609 (I166103,I2709);
not I_9610 (I166120,I384839);
nor I_9611 (I166137,I384848,I384821);
nand I_9612 (I166154,I166137,I384833);
DFFARX1 I_9613  ( .D(I166154), .CLK(I2702), .RSTB(I166103), .Q(I166074) );
nor I_9614 (I166185,I166120,I384848);
nand I_9615 (I166202,I166185,I384845);
nand I_9616 (I166219,I166202,I166154);
not I_9617 (I166236,I384848);
not I_9618 (I166253,I384824);
nor I_9619 (I166270,I166253,I384830);
and I_9620 (I166287,I166270,I384842);
or I_9621 (I166304,I166287,I384827);
DFFARX1 I_9622  ( .D(I166304), .CLK(I2702), .RSTB(I166103), .Q(I166321) );
nor I_9623 (I166338,I166321,I166202);
nand I_9624 (I166089,I166236,I166338);
not I_9625 (I166086,I166321);
and I_9626 (I166383,I166321,I166219);
DFFARX1 I_9627  ( .D(I166383), .CLK(I2702), .RSTB(I166103), .Q(I166071) );
DFFARX1 I_9628  ( .D(I166321), .CLK(I2702), .RSTB(I166103), .Q(I166414) );
and I_9629 (I166068,I166236,I166414);
nand I_9630 (I166445,I166120,I384824);
not I_9631 (I166462,I166445);
nor I_9632 (I166479,I166321,I166462);
DFFARX1 I_9633  ( .D(I384851), .CLK(I2702), .RSTB(I166103), .Q(I166496) );
nand I_9634 (I166513,I166496,I166445);
and I_9635 (I166530,I166236,I166513);
DFFARX1 I_9636  ( .D(I166530), .CLK(I2702), .RSTB(I166103), .Q(I166095) );
not I_9637 (I166561,I166496);
nand I_9638 (I166083,I166496,I166479);
nand I_9639 (I166077,I166496,I166462);
DFFARX1 I_9640  ( .D(I384836), .CLK(I2702), .RSTB(I166103), .Q(I166606) );
not I_9641 (I166623,I166606);
nor I_9642 (I166092,I166496,I166623);
nor I_9643 (I166654,I166623,I166561);
and I_9644 (I166671,I166202,I166654);
or I_9645 (I166688,I166445,I166671);
DFFARX1 I_9646  ( .D(I166688), .CLK(I2702), .RSTB(I166103), .Q(I166080) );
DFFARX1 I_9647  ( .D(I166623), .CLK(I2702), .RSTB(I166103), .Q(I166065) );
not I_9648 (I166766,I2709);
not I_9649 (I166783,I647653);
nor I_9650 (I166800,I647659,I647671);
nand I_9651 (I166817,I166800,I647662);
DFFARX1 I_9652  ( .D(I166817), .CLK(I2702), .RSTB(I166766), .Q(I166737) );
nor I_9653 (I166848,I166783,I647659);
nand I_9654 (I166865,I166848,I647641);
nand I_9655 (I166882,I166865,I166817);
not I_9656 (I166899,I647659);
not I_9657 (I166916,I647656);
nor I_9658 (I166933,I166916,I647644);
and I_9659 (I166950,I166933,I647665);
or I_9660 (I166967,I166950,I647647);
DFFARX1 I_9661  ( .D(I166967), .CLK(I2702), .RSTB(I166766), .Q(I166984) );
nor I_9662 (I167001,I166984,I166865);
nand I_9663 (I166752,I166899,I167001);
not I_9664 (I166749,I166984);
and I_9665 (I167046,I166984,I166882);
DFFARX1 I_9666  ( .D(I167046), .CLK(I2702), .RSTB(I166766), .Q(I166734) );
DFFARX1 I_9667  ( .D(I166984), .CLK(I2702), .RSTB(I166766), .Q(I167077) );
and I_9668 (I166731,I166899,I167077);
nand I_9669 (I167108,I166783,I647656);
not I_9670 (I167125,I167108);
nor I_9671 (I167142,I166984,I167125);
DFFARX1 I_9672  ( .D(I647668), .CLK(I2702), .RSTB(I166766), .Q(I167159) );
nand I_9673 (I167176,I167159,I167108);
and I_9674 (I167193,I166899,I167176);
DFFARX1 I_9675  ( .D(I167193), .CLK(I2702), .RSTB(I166766), .Q(I166758) );
not I_9676 (I167224,I167159);
nand I_9677 (I166746,I167159,I167142);
nand I_9678 (I166740,I167159,I167125);
DFFARX1 I_9679  ( .D(I647650), .CLK(I2702), .RSTB(I166766), .Q(I167269) );
not I_9680 (I167286,I167269);
nor I_9681 (I166755,I167159,I167286);
nor I_9682 (I167317,I167286,I167224);
and I_9683 (I167334,I166865,I167317);
or I_9684 (I167351,I167108,I167334);
DFFARX1 I_9685  ( .D(I167351), .CLK(I2702), .RSTB(I166766), .Q(I166743) );
DFFARX1 I_9686  ( .D(I167286), .CLK(I2702), .RSTB(I166766), .Q(I166728) );
not I_9687 (I167429,I2709);
not I_9688 (I167446,I585750);
nor I_9689 (I167463,I585765,I585747);
nand I_9690 (I167480,I167463,I585759);
DFFARX1 I_9691  ( .D(I167480), .CLK(I2702), .RSTB(I167429), .Q(I167400) );
nor I_9692 (I167511,I167446,I585765);
nand I_9693 (I167528,I167511,I585756);
nand I_9694 (I167545,I167528,I167480);
not I_9695 (I167562,I585765);
not I_9696 (I167579,I585774);
nor I_9697 (I167596,I167579,I585744);
and I_9698 (I167613,I167596,I585753);
or I_9699 (I167630,I167613,I585771);
DFFARX1 I_9700  ( .D(I167630), .CLK(I2702), .RSTB(I167429), .Q(I167647) );
nor I_9701 (I167664,I167647,I167528);
nand I_9702 (I167415,I167562,I167664);
not I_9703 (I167412,I167647);
and I_9704 (I167709,I167647,I167545);
DFFARX1 I_9705  ( .D(I167709), .CLK(I2702), .RSTB(I167429), .Q(I167397) );
DFFARX1 I_9706  ( .D(I167647), .CLK(I2702), .RSTB(I167429), .Q(I167740) );
and I_9707 (I167394,I167562,I167740);
nand I_9708 (I167771,I167446,I585774);
not I_9709 (I167788,I167771);
nor I_9710 (I167805,I167647,I167788);
DFFARX1 I_9711  ( .D(I585762), .CLK(I2702), .RSTB(I167429), .Q(I167822) );
nand I_9712 (I167839,I167822,I167771);
and I_9713 (I167856,I167562,I167839);
DFFARX1 I_9714  ( .D(I167856), .CLK(I2702), .RSTB(I167429), .Q(I167421) );
not I_9715 (I167887,I167822);
nand I_9716 (I167409,I167822,I167805);
nand I_9717 (I167403,I167822,I167788);
DFFARX1 I_9718  ( .D(I585768), .CLK(I2702), .RSTB(I167429), .Q(I167932) );
not I_9719 (I167949,I167932);
nor I_9720 (I167418,I167822,I167949);
nor I_9721 (I167980,I167949,I167887);
and I_9722 (I167997,I167528,I167980);
or I_9723 (I168014,I167771,I167997);
DFFARX1 I_9724  ( .D(I168014), .CLK(I2702), .RSTB(I167429), .Q(I167406) );
DFFARX1 I_9725  ( .D(I167949), .CLK(I2702), .RSTB(I167429), .Q(I167391) );
not I_9726 (I168092,I2709);
not I_9727 (I168109,I85296);
nor I_9728 (I168126,I85284,I85308);
nand I_9729 (I168143,I168126,I85293);
DFFARX1 I_9730  ( .D(I168143), .CLK(I2702), .RSTB(I168092), .Q(I168063) );
nor I_9731 (I168174,I168109,I85284);
nand I_9732 (I168191,I168174,I85311);
nand I_9733 (I168208,I168191,I168143);
not I_9734 (I168225,I85284);
not I_9735 (I168242,I85281);
nor I_9736 (I168259,I168242,I85290);
and I_9737 (I168276,I168259,I85305);
or I_9738 (I168293,I168276,I85287);
DFFARX1 I_9739  ( .D(I168293), .CLK(I2702), .RSTB(I168092), .Q(I168310) );
nor I_9740 (I168327,I168310,I168191);
nand I_9741 (I168078,I168225,I168327);
not I_9742 (I168075,I168310);
and I_9743 (I168372,I168310,I168208);
DFFARX1 I_9744  ( .D(I168372), .CLK(I2702), .RSTB(I168092), .Q(I168060) );
DFFARX1 I_9745  ( .D(I168310), .CLK(I2702), .RSTB(I168092), .Q(I168403) );
and I_9746 (I168057,I168225,I168403);
nand I_9747 (I168434,I168109,I85281);
not I_9748 (I168451,I168434);
nor I_9749 (I168468,I168310,I168451);
DFFARX1 I_9750  ( .D(I85302), .CLK(I2702), .RSTB(I168092), .Q(I168485) );
nand I_9751 (I168502,I168485,I168434);
and I_9752 (I168519,I168225,I168502);
DFFARX1 I_9753  ( .D(I168519), .CLK(I2702), .RSTB(I168092), .Q(I168084) );
not I_9754 (I168550,I168485);
nand I_9755 (I168072,I168485,I168468);
nand I_9756 (I168066,I168485,I168451);
DFFARX1 I_9757  ( .D(I85299), .CLK(I2702), .RSTB(I168092), .Q(I168595) );
not I_9758 (I168612,I168595);
nor I_9759 (I168081,I168485,I168612);
nor I_9760 (I168643,I168612,I168550);
and I_9761 (I168660,I168191,I168643);
or I_9762 (I168677,I168434,I168660);
DFFARX1 I_9763  ( .D(I168677), .CLK(I2702), .RSTB(I168092), .Q(I168069) );
DFFARX1 I_9764  ( .D(I168612), .CLK(I2702), .RSTB(I168092), .Q(I168054) );
not I_9765 (I168755,I2709);
not I_9766 (I168772,I353831);
nor I_9767 (I168789,I353840,I353813);
nand I_9768 (I168806,I168789,I353825);
DFFARX1 I_9769  ( .D(I168806), .CLK(I2702), .RSTB(I168755), .Q(I168726) );
nor I_9770 (I168837,I168772,I353840);
nand I_9771 (I168854,I168837,I353837);
nand I_9772 (I168871,I168854,I168806);
not I_9773 (I168888,I353840);
not I_9774 (I168905,I353816);
nor I_9775 (I168922,I168905,I353822);
and I_9776 (I168939,I168922,I353834);
or I_9777 (I168956,I168939,I353819);
DFFARX1 I_9778  ( .D(I168956), .CLK(I2702), .RSTB(I168755), .Q(I168973) );
nor I_9779 (I168990,I168973,I168854);
nand I_9780 (I168741,I168888,I168990);
not I_9781 (I168738,I168973);
and I_9782 (I169035,I168973,I168871);
DFFARX1 I_9783  ( .D(I169035), .CLK(I2702), .RSTB(I168755), .Q(I168723) );
DFFARX1 I_9784  ( .D(I168973), .CLK(I2702), .RSTB(I168755), .Q(I169066) );
and I_9785 (I168720,I168888,I169066);
nand I_9786 (I169097,I168772,I353816);
not I_9787 (I169114,I169097);
nor I_9788 (I169131,I168973,I169114);
DFFARX1 I_9789  ( .D(I353843), .CLK(I2702), .RSTB(I168755), .Q(I169148) );
nand I_9790 (I169165,I169148,I169097);
and I_9791 (I169182,I168888,I169165);
DFFARX1 I_9792  ( .D(I169182), .CLK(I2702), .RSTB(I168755), .Q(I168747) );
not I_9793 (I169213,I169148);
nand I_9794 (I168735,I169148,I169131);
nand I_9795 (I168729,I169148,I169114);
DFFARX1 I_9796  ( .D(I353828), .CLK(I2702), .RSTB(I168755), .Q(I169258) );
not I_9797 (I169275,I169258);
nor I_9798 (I168744,I169148,I169275);
nor I_9799 (I169306,I169275,I169213);
and I_9800 (I169323,I168854,I169306);
or I_9801 (I169340,I169097,I169323);
DFFARX1 I_9802  ( .D(I169340), .CLK(I2702), .RSTB(I168755), .Q(I168732) );
DFFARX1 I_9803  ( .D(I169275), .CLK(I2702), .RSTB(I168755), .Q(I168717) );
not I_9804 (I169418,I2709);
not I_9805 (I169435,I82712);
nor I_9806 (I169452,I82700,I82724);
nand I_9807 (I169469,I169452,I82709);
DFFARX1 I_9808  ( .D(I169469), .CLK(I2702), .RSTB(I169418), .Q(I169389) );
nor I_9809 (I169500,I169435,I82700);
nand I_9810 (I169517,I169500,I82727);
nand I_9811 (I169534,I169517,I169469);
not I_9812 (I169551,I82700);
not I_9813 (I169568,I82697);
nor I_9814 (I169585,I169568,I82706);
and I_9815 (I169602,I169585,I82721);
or I_9816 (I169619,I169602,I82703);
DFFARX1 I_9817  ( .D(I169619), .CLK(I2702), .RSTB(I169418), .Q(I169636) );
nor I_9818 (I169653,I169636,I169517);
nand I_9819 (I169404,I169551,I169653);
not I_9820 (I169401,I169636);
and I_9821 (I169698,I169636,I169534);
DFFARX1 I_9822  ( .D(I169698), .CLK(I2702), .RSTB(I169418), .Q(I169386) );
DFFARX1 I_9823  ( .D(I169636), .CLK(I2702), .RSTB(I169418), .Q(I169729) );
and I_9824 (I169383,I169551,I169729);
nand I_9825 (I169760,I169435,I82697);
not I_9826 (I169777,I169760);
nor I_9827 (I169794,I169636,I169777);
DFFARX1 I_9828  ( .D(I82718), .CLK(I2702), .RSTB(I169418), .Q(I169811) );
nand I_9829 (I169828,I169811,I169760);
and I_9830 (I169845,I169551,I169828);
DFFARX1 I_9831  ( .D(I169845), .CLK(I2702), .RSTB(I169418), .Q(I169410) );
not I_9832 (I169876,I169811);
nand I_9833 (I169398,I169811,I169794);
nand I_9834 (I169392,I169811,I169777);
DFFARX1 I_9835  ( .D(I82715), .CLK(I2702), .RSTB(I169418), .Q(I169921) );
not I_9836 (I169938,I169921);
nor I_9837 (I169407,I169811,I169938);
nor I_9838 (I169969,I169938,I169876);
and I_9839 (I169986,I169517,I169969);
or I_9840 (I170003,I169760,I169986);
DFFARX1 I_9841  ( .D(I170003), .CLK(I2702), .RSTB(I169418), .Q(I169395) );
DFFARX1 I_9842  ( .D(I169938), .CLK(I2702), .RSTB(I169418), .Q(I169380) );
not I_9843 (I170081,I2709);
not I_9844 (I170098,I659604);
nor I_9845 (I170115,I659610,I659622);
nand I_9846 (I170132,I170115,I659613);
DFFARX1 I_9847  ( .D(I170132), .CLK(I2702), .RSTB(I170081), .Q(I170052) );
nor I_9848 (I170163,I170098,I659610);
nand I_9849 (I170180,I170163,I659592);
nand I_9850 (I170197,I170180,I170132);
not I_9851 (I170214,I659610);
not I_9852 (I170231,I659607);
nor I_9853 (I170248,I170231,I659595);
and I_9854 (I170265,I170248,I659616);
or I_9855 (I170282,I170265,I659598);
DFFARX1 I_9856  ( .D(I170282), .CLK(I2702), .RSTB(I170081), .Q(I170299) );
nor I_9857 (I170316,I170299,I170180);
nand I_9858 (I170067,I170214,I170316);
not I_9859 (I170064,I170299);
and I_9860 (I170361,I170299,I170197);
DFFARX1 I_9861  ( .D(I170361), .CLK(I2702), .RSTB(I170081), .Q(I170049) );
DFFARX1 I_9862  ( .D(I170299), .CLK(I2702), .RSTB(I170081), .Q(I170392) );
and I_9863 (I170046,I170214,I170392);
nand I_9864 (I170423,I170098,I659607);
not I_9865 (I170440,I170423);
nor I_9866 (I170457,I170299,I170440);
DFFARX1 I_9867  ( .D(I659619), .CLK(I2702), .RSTB(I170081), .Q(I170474) );
nand I_9868 (I170491,I170474,I170423);
and I_9869 (I170508,I170214,I170491);
DFFARX1 I_9870  ( .D(I170508), .CLK(I2702), .RSTB(I170081), .Q(I170073) );
not I_9871 (I170539,I170474);
nand I_9872 (I170061,I170474,I170457);
nand I_9873 (I170055,I170474,I170440);
DFFARX1 I_9874  ( .D(I659601), .CLK(I2702), .RSTB(I170081), .Q(I170584) );
not I_9875 (I170601,I170584);
nor I_9876 (I170070,I170474,I170601);
nor I_9877 (I170632,I170601,I170539);
and I_9878 (I170649,I170180,I170632);
or I_9879 (I170666,I170423,I170649);
DFFARX1 I_9880  ( .D(I170666), .CLK(I2702), .RSTB(I170081), .Q(I170058) );
DFFARX1 I_9881  ( .D(I170601), .CLK(I2702), .RSTB(I170081), .Q(I170043) );
not I_9882 (I170744,I2709);
not I_9883 (I170761,I223702);
nor I_9884 (I170778,I223684,I223678);
nand I_9885 (I170795,I170778,I223681);
DFFARX1 I_9886  ( .D(I170795), .CLK(I2702), .RSTB(I170744), .Q(I170715) );
nor I_9887 (I170826,I170761,I223684);
nand I_9888 (I170843,I170826,I223690);
nand I_9889 (I170860,I170843,I170795);
not I_9890 (I170877,I223684);
not I_9891 (I170894,I223699);
nor I_9892 (I170911,I170894,I223687);
and I_9893 (I170928,I170911,I223693);
or I_9894 (I170945,I170928,I223708);
DFFARX1 I_9895  ( .D(I170945), .CLK(I2702), .RSTB(I170744), .Q(I170962) );
nor I_9896 (I170979,I170962,I170843);
nand I_9897 (I170730,I170877,I170979);
not I_9898 (I170727,I170962);
and I_9899 (I171024,I170962,I170860);
DFFARX1 I_9900  ( .D(I171024), .CLK(I2702), .RSTB(I170744), .Q(I170712) );
DFFARX1 I_9901  ( .D(I170962), .CLK(I2702), .RSTB(I170744), .Q(I171055) );
and I_9902 (I170709,I170877,I171055);
nand I_9903 (I171086,I170761,I223699);
not I_9904 (I171103,I171086);
nor I_9905 (I171120,I170962,I171103);
DFFARX1 I_9906  ( .D(I223696), .CLK(I2702), .RSTB(I170744), .Q(I171137) );
nand I_9907 (I171154,I171137,I171086);
and I_9908 (I171171,I170877,I171154);
DFFARX1 I_9909  ( .D(I171171), .CLK(I2702), .RSTB(I170744), .Q(I170736) );
not I_9910 (I171202,I171137);
nand I_9911 (I170724,I171137,I171120);
nand I_9912 (I170718,I171137,I171103);
DFFARX1 I_9913  ( .D(I223705), .CLK(I2702), .RSTB(I170744), .Q(I171247) );
not I_9914 (I171264,I171247);
nor I_9915 (I170733,I171137,I171264);
nor I_9916 (I171295,I171264,I171202);
and I_9917 (I171312,I170843,I171295);
or I_9918 (I171329,I171086,I171312);
DFFARX1 I_9919  ( .D(I171329), .CLK(I2702), .RSTB(I170744), .Q(I170721) );
DFFARX1 I_9920  ( .D(I171264), .CLK(I2702), .RSTB(I170744), .Q(I170706) );
not I_9921 (I171407,I2709);
not I_9922 (I171424,I136976);
nor I_9923 (I171441,I136964,I136988);
nand I_9924 (I171458,I171441,I136973);
DFFARX1 I_9925  ( .D(I171458), .CLK(I2702), .RSTB(I171407), .Q(I171378) );
nor I_9926 (I171489,I171424,I136964);
nand I_9927 (I171506,I171489,I136991);
nand I_9928 (I171523,I171506,I171458);
not I_9929 (I171540,I136964);
not I_9930 (I171557,I136961);
nor I_9931 (I171574,I171557,I136970);
and I_9932 (I171591,I171574,I136985);
or I_9933 (I171608,I171591,I136967);
DFFARX1 I_9934  ( .D(I171608), .CLK(I2702), .RSTB(I171407), .Q(I171625) );
nor I_9935 (I171642,I171625,I171506);
nand I_9936 (I171393,I171540,I171642);
not I_9937 (I171390,I171625);
and I_9938 (I171687,I171625,I171523);
DFFARX1 I_9939  ( .D(I171687), .CLK(I2702), .RSTB(I171407), .Q(I171375) );
DFFARX1 I_9940  ( .D(I171625), .CLK(I2702), .RSTB(I171407), .Q(I171718) );
and I_9941 (I171372,I171540,I171718);
nand I_9942 (I171749,I171424,I136961);
not I_9943 (I171766,I171749);
nor I_9944 (I171783,I171625,I171766);
DFFARX1 I_9945  ( .D(I136982), .CLK(I2702), .RSTB(I171407), .Q(I171800) );
nand I_9946 (I171817,I171800,I171749);
and I_9947 (I171834,I171540,I171817);
DFFARX1 I_9948  ( .D(I171834), .CLK(I2702), .RSTB(I171407), .Q(I171399) );
not I_9949 (I171865,I171800);
nand I_9950 (I171387,I171800,I171783);
nand I_9951 (I171381,I171800,I171766);
DFFARX1 I_9952  ( .D(I136979), .CLK(I2702), .RSTB(I171407), .Q(I171910) );
not I_9953 (I171927,I171910);
nor I_9954 (I171396,I171800,I171927);
nor I_9955 (I171958,I171927,I171865);
and I_9956 (I171975,I171506,I171958);
or I_9957 (I171992,I171749,I171975);
DFFARX1 I_9958  ( .D(I171992), .CLK(I2702), .RSTB(I171407), .Q(I171384) );
DFFARX1 I_9959  ( .D(I171927), .CLK(I2702), .RSTB(I171407), .Q(I171369) );
not I_9960 (I172070,I2709);
not I_9961 (I172087,I519119);
nor I_9962 (I172104,I519131,I519134);
nand I_9963 (I172121,I172104,I519122);
DFFARX1 I_9964  ( .D(I172121), .CLK(I2702), .RSTB(I172070), .Q(I172041) );
nor I_9965 (I172152,I172087,I519131);
nand I_9966 (I172169,I172152,I519107);
nand I_9967 (I172186,I172169,I172121);
not I_9968 (I172203,I519131);
not I_9969 (I172220,I519110);
nor I_9970 (I172237,I172220,I519113);
and I_9971 (I172254,I172237,I519116);
or I_9972 (I172271,I172254,I519125);
DFFARX1 I_9973  ( .D(I172271), .CLK(I2702), .RSTB(I172070), .Q(I172288) );
nor I_9974 (I172305,I172288,I172169);
nand I_9975 (I172056,I172203,I172305);
not I_9976 (I172053,I172288);
and I_9977 (I172350,I172288,I172186);
DFFARX1 I_9978  ( .D(I172350), .CLK(I2702), .RSTB(I172070), .Q(I172038) );
DFFARX1 I_9979  ( .D(I172288), .CLK(I2702), .RSTB(I172070), .Q(I172381) );
and I_9980 (I172035,I172203,I172381);
nand I_9981 (I172412,I172087,I519110);
not I_9982 (I172429,I172412);
nor I_9983 (I172446,I172288,I172429);
DFFARX1 I_9984  ( .D(I519128), .CLK(I2702), .RSTB(I172070), .Q(I172463) );
nand I_9985 (I172480,I172463,I172412);
and I_9986 (I172497,I172203,I172480);
DFFARX1 I_9987  ( .D(I172497), .CLK(I2702), .RSTB(I172070), .Q(I172062) );
not I_9988 (I172528,I172463);
nand I_9989 (I172050,I172463,I172446);
nand I_9990 (I172044,I172463,I172429);
DFFARX1 I_9991  ( .D(I519104), .CLK(I2702), .RSTB(I172070), .Q(I172573) );
not I_9992 (I172590,I172573);
nor I_9993 (I172059,I172463,I172590);
nor I_9994 (I172621,I172590,I172528);
and I_9995 (I172638,I172169,I172621);
or I_9996 (I172655,I172412,I172638);
DFFARX1 I_9997  ( .D(I172655), .CLK(I2702), .RSTB(I172070), .Q(I172047) );
DFFARX1 I_9998  ( .D(I172590), .CLK(I2702), .RSTB(I172070), .Q(I172032) );
not I_9999 (I172733,I2709);
not I_10000 (I172750,I297339);
nor I_10001 (I172767,I297348,I297360);
nand I_10002 (I172784,I172767,I297351);
DFFARX1 I_10003  ( .D(I172784), .CLK(I2702), .RSTB(I172733), .Q(I172704) );
nor I_10004 (I172815,I172750,I297348);
nand I_10005 (I172832,I172815,I297363);
nand I_10006 (I172849,I172832,I172784);
not I_10007 (I172866,I297348);
not I_10008 (I172883,I297369);
nor I_10009 (I172900,I172883,I297345);
and I_10010 (I172917,I172900,I297354);
or I_10011 (I172934,I172917,I297342);
DFFARX1 I_10012  ( .D(I172934), .CLK(I2702), .RSTB(I172733), .Q(I172951) );
nor I_10013 (I172968,I172951,I172832);
nand I_10014 (I172719,I172866,I172968);
not I_10015 (I172716,I172951);
and I_10016 (I173013,I172951,I172849);
DFFARX1 I_10017  ( .D(I173013), .CLK(I2702), .RSTB(I172733), .Q(I172701) );
DFFARX1 I_10018  ( .D(I172951), .CLK(I2702), .RSTB(I172733), .Q(I173044) );
and I_10019 (I172698,I172866,I173044);
nand I_10020 (I173075,I172750,I297369);
not I_10021 (I173092,I173075);
nor I_10022 (I173109,I172951,I173092);
DFFARX1 I_10023  ( .D(I297366), .CLK(I2702), .RSTB(I172733), .Q(I173126) );
nand I_10024 (I173143,I173126,I173075);
and I_10025 (I173160,I172866,I173143);
DFFARX1 I_10026  ( .D(I173160), .CLK(I2702), .RSTB(I172733), .Q(I172725) );
not I_10027 (I173191,I173126);
nand I_10028 (I172713,I173126,I173109);
nand I_10029 (I172707,I173126,I173092);
DFFARX1 I_10030  ( .D(I297357), .CLK(I2702), .RSTB(I172733), .Q(I173236) );
not I_10031 (I173253,I173236);
nor I_10032 (I172722,I173126,I173253);
nor I_10033 (I173284,I173253,I173191);
and I_10034 (I173301,I172832,I173284);
or I_10035 (I173318,I173075,I173301);
DFFARX1 I_10036  ( .D(I173318), .CLK(I2702), .RSTB(I172733), .Q(I172710) );
DFFARX1 I_10037  ( .D(I173253), .CLK(I2702), .RSTB(I172733), .Q(I172695) );
not I_10038 (I173396,I2709);
not I_10039 (I173413,I560174);
nor I_10040 (I173430,I560186,I560189);
nand I_10041 (I173447,I173430,I560177);
DFFARX1 I_10042  ( .D(I173447), .CLK(I2702), .RSTB(I173396), .Q(I173367) );
nor I_10043 (I173478,I173413,I560186);
nand I_10044 (I173495,I173478,I560162);
nand I_10045 (I173512,I173495,I173447);
not I_10046 (I173529,I560186);
not I_10047 (I173546,I560165);
nor I_10048 (I173563,I173546,I560168);
and I_10049 (I173580,I173563,I560171);
or I_10050 (I173597,I173580,I560180);
DFFARX1 I_10051  ( .D(I173597), .CLK(I2702), .RSTB(I173396), .Q(I173614) );
nor I_10052 (I173631,I173614,I173495);
nand I_10053 (I173382,I173529,I173631);
not I_10054 (I173379,I173614);
and I_10055 (I173676,I173614,I173512);
DFFARX1 I_10056  ( .D(I173676), .CLK(I2702), .RSTB(I173396), .Q(I173364) );
DFFARX1 I_10057  ( .D(I173614), .CLK(I2702), .RSTB(I173396), .Q(I173707) );
and I_10058 (I173361,I173529,I173707);
nand I_10059 (I173738,I173413,I560165);
not I_10060 (I173755,I173738);
nor I_10061 (I173772,I173614,I173755);
DFFARX1 I_10062  ( .D(I560183), .CLK(I2702), .RSTB(I173396), .Q(I173789) );
nand I_10063 (I173806,I173789,I173738);
and I_10064 (I173823,I173529,I173806);
DFFARX1 I_10065  ( .D(I173823), .CLK(I2702), .RSTB(I173396), .Q(I173388) );
not I_10066 (I173854,I173789);
nand I_10067 (I173376,I173789,I173772);
nand I_10068 (I173370,I173789,I173755);
DFFARX1 I_10069  ( .D(I560159), .CLK(I2702), .RSTB(I173396), .Q(I173899) );
not I_10070 (I173916,I173899);
nor I_10071 (I173385,I173789,I173916);
nor I_10072 (I173947,I173916,I173854);
and I_10073 (I173964,I173495,I173947);
or I_10074 (I173981,I173738,I173964);
DFFARX1 I_10075  ( .D(I173981), .CLK(I2702), .RSTB(I173396), .Q(I173373) );
DFFARX1 I_10076  ( .D(I173916), .CLK(I2702), .RSTB(I173396), .Q(I173358) );
not I_10077 (I174059,I2709);
not I_10078 (I174076,I537564);
nor I_10079 (I174093,I537576,I537579);
nand I_10080 (I174110,I174093,I537567);
DFFARX1 I_10081  ( .D(I174110), .CLK(I2702), .RSTB(I174059), .Q(I174030) );
nor I_10082 (I174141,I174076,I537576);
nand I_10083 (I174158,I174141,I537552);
nand I_10084 (I174175,I174158,I174110);
not I_10085 (I174192,I537576);
not I_10086 (I174209,I537555);
nor I_10087 (I174226,I174209,I537558);
and I_10088 (I174243,I174226,I537561);
or I_10089 (I174260,I174243,I537570);
DFFARX1 I_10090  ( .D(I174260), .CLK(I2702), .RSTB(I174059), .Q(I174277) );
nor I_10091 (I174294,I174277,I174158);
nand I_10092 (I174045,I174192,I174294);
not I_10093 (I174042,I174277);
and I_10094 (I174339,I174277,I174175);
DFFARX1 I_10095  ( .D(I174339), .CLK(I2702), .RSTB(I174059), .Q(I174027) );
DFFARX1 I_10096  ( .D(I174277), .CLK(I2702), .RSTB(I174059), .Q(I174370) );
and I_10097 (I174024,I174192,I174370);
nand I_10098 (I174401,I174076,I537555);
not I_10099 (I174418,I174401);
nor I_10100 (I174435,I174277,I174418);
DFFARX1 I_10101  ( .D(I537573), .CLK(I2702), .RSTB(I174059), .Q(I174452) );
nand I_10102 (I174469,I174452,I174401);
and I_10103 (I174486,I174192,I174469);
DFFARX1 I_10104  ( .D(I174486), .CLK(I2702), .RSTB(I174059), .Q(I174051) );
not I_10105 (I174517,I174452);
nand I_10106 (I174039,I174452,I174435);
nand I_10107 (I174033,I174452,I174418);
DFFARX1 I_10108  ( .D(I537549), .CLK(I2702), .RSTB(I174059), .Q(I174562) );
not I_10109 (I174579,I174562);
nor I_10110 (I174048,I174452,I174579);
nor I_10111 (I174610,I174579,I174517);
and I_10112 (I174627,I174158,I174610);
or I_10113 (I174644,I174401,I174627);
DFFARX1 I_10114  ( .D(I174644), .CLK(I2702), .RSTB(I174059), .Q(I174036) );
DFFARX1 I_10115  ( .D(I174579), .CLK(I2702), .RSTB(I174059), .Q(I174021) );
not I_10116 (I174722,I2709);
not I_10117 (I174739,I482401);
nor I_10118 (I174756,I482407,I482404);
nand I_10119 (I174773,I174756,I482422);
DFFARX1 I_10120  ( .D(I174773), .CLK(I2702), .RSTB(I174722), .Q(I174693) );
nor I_10121 (I174804,I174739,I482407);
nand I_10122 (I174821,I174804,I482431);
nand I_10123 (I174838,I174821,I174773);
not I_10124 (I174855,I482407);
not I_10125 (I174872,I482425);
nor I_10126 (I174889,I174872,I482416);
and I_10127 (I174906,I174889,I482419);
or I_10128 (I174923,I174906,I482410);
DFFARX1 I_10129  ( .D(I174923), .CLK(I2702), .RSTB(I174722), .Q(I174940) );
nor I_10130 (I174957,I174940,I174821);
nand I_10131 (I174708,I174855,I174957);
not I_10132 (I174705,I174940);
and I_10133 (I175002,I174940,I174838);
DFFARX1 I_10134  ( .D(I175002), .CLK(I2702), .RSTB(I174722), .Q(I174690) );
DFFARX1 I_10135  ( .D(I174940), .CLK(I2702), .RSTB(I174722), .Q(I175033) );
and I_10136 (I174687,I174855,I175033);
nand I_10137 (I175064,I174739,I482425);
not I_10138 (I175081,I175064);
nor I_10139 (I175098,I174940,I175081);
DFFARX1 I_10140  ( .D(I482428), .CLK(I2702), .RSTB(I174722), .Q(I175115) );
nand I_10141 (I175132,I175115,I175064);
and I_10142 (I175149,I174855,I175132);
DFFARX1 I_10143  ( .D(I175149), .CLK(I2702), .RSTB(I174722), .Q(I174714) );
not I_10144 (I175180,I175115);
nand I_10145 (I174702,I175115,I175098);
nand I_10146 (I174696,I175115,I175081);
DFFARX1 I_10147  ( .D(I482413), .CLK(I2702), .RSTB(I174722), .Q(I175225) );
not I_10148 (I175242,I175225);
nor I_10149 (I174711,I175115,I175242);
nor I_10150 (I175273,I175242,I175180);
and I_10151 (I175290,I174821,I175273);
or I_10152 (I175307,I175064,I175290);
DFFARX1 I_10153  ( .D(I175307), .CLK(I2702), .RSTB(I174722), .Q(I174699) );
DFFARX1 I_10154  ( .D(I175242), .CLK(I2702), .RSTB(I174722), .Q(I174684) );
not I_10155 (I175385,I2709);
not I_10156 (I175402,I419921);
nor I_10157 (I175419,I419939,I419927);
nand I_10158 (I175436,I175419,I419933);
DFFARX1 I_10159  ( .D(I175436), .CLK(I2702), .RSTB(I175385), .Q(I175356) );
nor I_10160 (I175467,I175402,I419939);
nand I_10161 (I175484,I175467,I419936);
nand I_10162 (I175501,I175484,I175436);
not I_10163 (I175518,I419939);
not I_10164 (I175535,I419915);
nor I_10165 (I175552,I175535,I419909);
and I_10166 (I175569,I175552,I419918);
or I_10167 (I175586,I175569,I419930);
DFFARX1 I_10168  ( .D(I175586), .CLK(I2702), .RSTB(I175385), .Q(I175603) );
nor I_10169 (I175620,I175603,I175484);
nand I_10170 (I175371,I175518,I175620);
not I_10171 (I175368,I175603);
and I_10172 (I175665,I175603,I175501);
DFFARX1 I_10173  ( .D(I175665), .CLK(I2702), .RSTB(I175385), .Q(I175353) );
DFFARX1 I_10174  ( .D(I175603), .CLK(I2702), .RSTB(I175385), .Q(I175696) );
and I_10175 (I175350,I175518,I175696);
nand I_10176 (I175727,I175402,I419915);
not I_10177 (I175744,I175727);
nor I_10178 (I175761,I175603,I175744);
DFFARX1 I_10179  ( .D(I419924), .CLK(I2702), .RSTB(I175385), .Q(I175778) );
nand I_10180 (I175795,I175778,I175727);
and I_10181 (I175812,I175518,I175795);
DFFARX1 I_10182  ( .D(I175812), .CLK(I2702), .RSTB(I175385), .Q(I175377) );
not I_10183 (I175843,I175778);
nand I_10184 (I175365,I175778,I175761);
nand I_10185 (I175359,I175778,I175744);
DFFARX1 I_10186  ( .D(I419912), .CLK(I2702), .RSTB(I175385), .Q(I175888) );
not I_10187 (I175905,I175888);
nor I_10188 (I175374,I175778,I175905);
nor I_10189 (I175936,I175905,I175843);
and I_10190 (I175953,I175484,I175936);
or I_10191 (I175970,I175727,I175953);
DFFARX1 I_10192  ( .D(I175970), .CLK(I2702), .RSTB(I175385), .Q(I175362) );
DFFARX1 I_10193  ( .D(I175905), .CLK(I2702), .RSTB(I175385), .Q(I175347) );
not I_10194 (I176048,I2709);
not I_10195 (I176065,I623751);
nor I_10196 (I176082,I623757,I623769);
nand I_10197 (I176099,I176082,I623760);
DFFARX1 I_10198  ( .D(I176099), .CLK(I2702), .RSTB(I176048), .Q(I176019) );
nor I_10199 (I176130,I176065,I623757);
nand I_10200 (I176147,I176130,I623739);
nand I_10201 (I176164,I176147,I176099);
not I_10202 (I176181,I623757);
not I_10203 (I176198,I623754);
nor I_10204 (I176215,I176198,I623742);
and I_10205 (I176232,I176215,I623763);
or I_10206 (I176249,I176232,I623745);
DFFARX1 I_10207  ( .D(I176249), .CLK(I2702), .RSTB(I176048), .Q(I176266) );
nor I_10208 (I176283,I176266,I176147);
nand I_10209 (I176034,I176181,I176283);
not I_10210 (I176031,I176266);
and I_10211 (I176328,I176266,I176164);
DFFARX1 I_10212  ( .D(I176328), .CLK(I2702), .RSTB(I176048), .Q(I176016) );
DFFARX1 I_10213  ( .D(I176266), .CLK(I2702), .RSTB(I176048), .Q(I176359) );
and I_10214 (I176013,I176181,I176359);
nand I_10215 (I176390,I176065,I623754);
not I_10216 (I176407,I176390);
nor I_10217 (I176424,I176266,I176407);
DFFARX1 I_10218  ( .D(I623766), .CLK(I2702), .RSTB(I176048), .Q(I176441) );
nand I_10219 (I176458,I176441,I176390);
and I_10220 (I176475,I176181,I176458);
DFFARX1 I_10221  ( .D(I176475), .CLK(I2702), .RSTB(I176048), .Q(I176040) );
not I_10222 (I176506,I176441);
nand I_10223 (I176028,I176441,I176424);
nand I_10224 (I176022,I176441,I176407);
DFFARX1 I_10225  ( .D(I623748), .CLK(I2702), .RSTB(I176048), .Q(I176551) );
not I_10226 (I176568,I176551);
nor I_10227 (I176037,I176441,I176568);
nor I_10228 (I176599,I176568,I176506);
and I_10229 (I176616,I176147,I176599);
or I_10230 (I176633,I176390,I176616);
DFFARX1 I_10231  ( .D(I176633), .CLK(I2702), .RSTB(I176048), .Q(I176025) );
DFFARX1 I_10232  ( .D(I176568), .CLK(I2702), .RSTB(I176048), .Q(I176010) );
not I_10233 (I176711,I2709);
not I_10234 (I176728,I621235);
nor I_10235 (I176745,I621241,I621253);
nand I_10236 (I176762,I176745,I621244);
DFFARX1 I_10237  ( .D(I176762), .CLK(I2702), .RSTB(I176711), .Q(I176682) );
nor I_10238 (I176793,I176728,I621241);
nand I_10239 (I176810,I176793,I621223);
nand I_10240 (I176827,I176810,I176762);
not I_10241 (I176844,I621241);
not I_10242 (I176861,I621238);
nor I_10243 (I176878,I176861,I621226);
and I_10244 (I176895,I176878,I621247);
or I_10245 (I176912,I176895,I621229);
DFFARX1 I_10246  ( .D(I176912), .CLK(I2702), .RSTB(I176711), .Q(I176929) );
nor I_10247 (I176946,I176929,I176810);
nand I_10248 (I176697,I176844,I176946);
not I_10249 (I176694,I176929);
and I_10250 (I176991,I176929,I176827);
DFFARX1 I_10251  ( .D(I176991), .CLK(I2702), .RSTB(I176711), .Q(I176679) );
DFFARX1 I_10252  ( .D(I176929), .CLK(I2702), .RSTB(I176711), .Q(I177022) );
and I_10253 (I176676,I176844,I177022);
nand I_10254 (I177053,I176728,I621238);
not I_10255 (I177070,I177053);
nor I_10256 (I177087,I176929,I177070);
DFFARX1 I_10257  ( .D(I621250), .CLK(I2702), .RSTB(I176711), .Q(I177104) );
nand I_10258 (I177121,I177104,I177053);
and I_10259 (I177138,I176844,I177121);
DFFARX1 I_10260  ( .D(I177138), .CLK(I2702), .RSTB(I176711), .Q(I176703) );
not I_10261 (I177169,I177104);
nand I_10262 (I176691,I177104,I177087);
nand I_10263 (I176685,I177104,I177070);
DFFARX1 I_10264  ( .D(I621232), .CLK(I2702), .RSTB(I176711), .Q(I177214) );
not I_10265 (I177231,I177214);
nor I_10266 (I176700,I177104,I177231);
nor I_10267 (I177262,I177231,I177169);
and I_10268 (I177279,I176810,I177262);
or I_10269 (I177296,I177053,I177279);
DFFARX1 I_10270  ( .D(I177296), .CLK(I2702), .RSTB(I176711), .Q(I176688) );
DFFARX1 I_10271  ( .D(I177231), .CLK(I2702), .RSTB(I176711), .Q(I176673) );
not I_10272 (I177374,I2709);
not I_10273 (I177391,I635073);
nor I_10274 (I177408,I635079,I635091);
nand I_10275 (I177425,I177408,I635082);
DFFARX1 I_10276  ( .D(I177425), .CLK(I2702), .RSTB(I177374), .Q(I177345) );
nor I_10277 (I177456,I177391,I635079);
nand I_10278 (I177473,I177456,I635061);
nand I_10279 (I177490,I177473,I177425);
not I_10280 (I177507,I635079);
not I_10281 (I177524,I635076);
nor I_10282 (I177541,I177524,I635064);
and I_10283 (I177558,I177541,I635085);
or I_10284 (I177575,I177558,I635067);
DFFARX1 I_10285  ( .D(I177575), .CLK(I2702), .RSTB(I177374), .Q(I177592) );
nor I_10286 (I177609,I177592,I177473);
nand I_10287 (I177360,I177507,I177609);
not I_10288 (I177357,I177592);
and I_10289 (I177654,I177592,I177490);
DFFARX1 I_10290  ( .D(I177654), .CLK(I2702), .RSTB(I177374), .Q(I177342) );
DFFARX1 I_10291  ( .D(I177592), .CLK(I2702), .RSTB(I177374), .Q(I177685) );
and I_10292 (I177339,I177507,I177685);
nand I_10293 (I177716,I177391,I635076);
not I_10294 (I177733,I177716);
nor I_10295 (I177750,I177592,I177733);
DFFARX1 I_10296  ( .D(I635088), .CLK(I2702), .RSTB(I177374), .Q(I177767) );
nand I_10297 (I177784,I177767,I177716);
and I_10298 (I177801,I177507,I177784);
DFFARX1 I_10299  ( .D(I177801), .CLK(I2702), .RSTB(I177374), .Q(I177366) );
not I_10300 (I177832,I177767);
nand I_10301 (I177354,I177767,I177750);
nand I_10302 (I177348,I177767,I177733);
DFFARX1 I_10303  ( .D(I635070), .CLK(I2702), .RSTB(I177374), .Q(I177877) );
not I_10304 (I177894,I177877);
nor I_10305 (I177363,I177767,I177894);
nor I_10306 (I177925,I177894,I177832);
and I_10307 (I177942,I177473,I177925);
or I_10308 (I177959,I177716,I177942);
DFFARX1 I_10309  ( .D(I177959), .CLK(I2702), .RSTB(I177374), .Q(I177351) );
DFFARX1 I_10310  ( .D(I177894), .CLK(I2702), .RSTB(I177374), .Q(I177336) );
not I_10311 (I178037,I2709);
not I_10312 (I178054,I460437);
nor I_10313 (I178071,I460443,I460440);
nand I_10314 (I178088,I178071,I460458);
DFFARX1 I_10315  ( .D(I178088), .CLK(I2702), .RSTB(I178037), .Q(I178008) );
nor I_10316 (I178119,I178054,I460443);
nand I_10317 (I178136,I178119,I460467);
nand I_10318 (I178153,I178136,I178088);
not I_10319 (I178170,I460443);
not I_10320 (I178187,I460461);
nor I_10321 (I178204,I178187,I460452);
and I_10322 (I178221,I178204,I460455);
or I_10323 (I178238,I178221,I460446);
DFFARX1 I_10324  ( .D(I178238), .CLK(I2702), .RSTB(I178037), .Q(I178255) );
nor I_10325 (I178272,I178255,I178136);
nand I_10326 (I178023,I178170,I178272);
not I_10327 (I178020,I178255);
and I_10328 (I178317,I178255,I178153);
DFFARX1 I_10329  ( .D(I178317), .CLK(I2702), .RSTB(I178037), .Q(I178005) );
DFFARX1 I_10330  ( .D(I178255), .CLK(I2702), .RSTB(I178037), .Q(I178348) );
and I_10331 (I178002,I178170,I178348);
nand I_10332 (I178379,I178054,I460461);
not I_10333 (I178396,I178379);
nor I_10334 (I178413,I178255,I178396);
DFFARX1 I_10335  ( .D(I460464), .CLK(I2702), .RSTB(I178037), .Q(I178430) );
nand I_10336 (I178447,I178430,I178379);
and I_10337 (I178464,I178170,I178447);
DFFARX1 I_10338  ( .D(I178464), .CLK(I2702), .RSTB(I178037), .Q(I178029) );
not I_10339 (I178495,I178430);
nand I_10340 (I178017,I178430,I178413);
nand I_10341 (I178011,I178430,I178396);
DFFARX1 I_10342  ( .D(I460449), .CLK(I2702), .RSTB(I178037), .Q(I178540) );
not I_10343 (I178557,I178540);
nor I_10344 (I178026,I178430,I178557);
nor I_10345 (I178588,I178557,I178495);
and I_10346 (I178605,I178136,I178588);
or I_10347 (I178622,I178379,I178605);
DFFARX1 I_10348  ( .D(I178622), .CLK(I2702), .RSTB(I178037), .Q(I178014) );
DFFARX1 I_10349  ( .D(I178557), .CLK(I2702), .RSTB(I178037), .Q(I177999) );
not I_10350 (I178700,I2709);
not I_10351 (I178717,I290709);
nor I_10352 (I178734,I290718,I290730);
nand I_10353 (I178751,I178734,I290721);
DFFARX1 I_10354  ( .D(I178751), .CLK(I2702), .RSTB(I178700), .Q(I178671) );
nor I_10355 (I178782,I178717,I290718);
nand I_10356 (I178799,I178782,I290733);
nand I_10357 (I178816,I178799,I178751);
not I_10358 (I178833,I290718);
not I_10359 (I178850,I290739);
nor I_10360 (I178867,I178850,I290715);
and I_10361 (I178884,I178867,I290724);
or I_10362 (I178901,I178884,I290712);
DFFARX1 I_10363  ( .D(I178901), .CLK(I2702), .RSTB(I178700), .Q(I178918) );
nor I_10364 (I178935,I178918,I178799);
nand I_10365 (I178686,I178833,I178935);
not I_10366 (I178683,I178918);
and I_10367 (I178980,I178918,I178816);
DFFARX1 I_10368  ( .D(I178980), .CLK(I2702), .RSTB(I178700), .Q(I178668) );
DFFARX1 I_10369  ( .D(I178918), .CLK(I2702), .RSTB(I178700), .Q(I179011) );
and I_10370 (I178665,I178833,I179011);
nand I_10371 (I179042,I178717,I290739);
not I_10372 (I179059,I179042);
nor I_10373 (I179076,I178918,I179059);
DFFARX1 I_10374  ( .D(I290736), .CLK(I2702), .RSTB(I178700), .Q(I179093) );
nand I_10375 (I179110,I179093,I179042);
and I_10376 (I179127,I178833,I179110);
DFFARX1 I_10377  ( .D(I179127), .CLK(I2702), .RSTB(I178700), .Q(I178692) );
not I_10378 (I179158,I179093);
nand I_10379 (I178680,I179093,I179076);
nand I_10380 (I178674,I179093,I179059);
DFFARX1 I_10381  ( .D(I290727), .CLK(I2702), .RSTB(I178700), .Q(I179203) );
not I_10382 (I179220,I179203);
nor I_10383 (I178689,I179093,I179220);
nor I_10384 (I179251,I179220,I179158);
and I_10385 (I179268,I178799,I179251);
or I_10386 (I179285,I179042,I179268);
DFFARX1 I_10387  ( .D(I179285), .CLK(I2702), .RSTB(I178700), .Q(I178677) );
DFFARX1 I_10388  ( .D(I179220), .CLK(I2702), .RSTB(I178700), .Q(I178662) );
not I_10389 (I179363,I2709);
not I_10390 (I179380,I257559);
nor I_10391 (I179397,I257568,I257580);
nand I_10392 (I179414,I179397,I257571);
DFFARX1 I_10393  ( .D(I179414), .CLK(I2702), .RSTB(I179363), .Q(I179334) );
nor I_10394 (I179445,I179380,I257568);
nand I_10395 (I179462,I179445,I257583);
nand I_10396 (I179479,I179462,I179414);
not I_10397 (I179496,I257568);
not I_10398 (I179513,I257589);
nor I_10399 (I179530,I179513,I257565);
and I_10400 (I179547,I179530,I257574);
or I_10401 (I179564,I179547,I257562);
DFFARX1 I_10402  ( .D(I179564), .CLK(I2702), .RSTB(I179363), .Q(I179581) );
nor I_10403 (I179598,I179581,I179462);
nand I_10404 (I179349,I179496,I179598);
not I_10405 (I179346,I179581);
and I_10406 (I179643,I179581,I179479);
DFFARX1 I_10407  ( .D(I179643), .CLK(I2702), .RSTB(I179363), .Q(I179331) );
DFFARX1 I_10408  ( .D(I179581), .CLK(I2702), .RSTB(I179363), .Q(I179674) );
and I_10409 (I179328,I179496,I179674);
nand I_10410 (I179705,I179380,I257589);
not I_10411 (I179722,I179705);
nor I_10412 (I179739,I179581,I179722);
DFFARX1 I_10413  ( .D(I257586), .CLK(I2702), .RSTB(I179363), .Q(I179756) );
nand I_10414 (I179773,I179756,I179705);
and I_10415 (I179790,I179496,I179773);
DFFARX1 I_10416  ( .D(I179790), .CLK(I2702), .RSTB(I179363), .Q(I179355) );
not I_10417 (I179821,I179756);
nand I_10418 (I179343,I179756,I179739);
nand I_10419 (I179337,I179756,I179722);
DFFARX1 I_10420  ( .D(I257577), .CLK(I2702), .RSTB(I179363), .Q(I179866) );
not I_10421 (I179883,I179866);
nor I_10422 (I179352,I179756,I179883);
nor I_10423 (I179914,I179883,I179821);
and I_10424 (I179931,I179462,I179914);
or I_10425 (I179948,I179705,I179931);
DFFARX1 I_10426  ( .D(I179948), .CLK(I2702), .RSTB(I179363), .Q(I179340) );
DFFARX1 I_10427  ( .D(I179883), .CLK(I2702), .RSTB(I179363), .Q(I179325) );
not I_10428 (I180026,I2709);
not I_10429 (I180043,I557199);
nor I_10430 (I180060,I557211,I557214);
nand I_10431 (I180077,I180060,I557202);
DFFARX1 I_10432  ( .D(I180077), .CLK(I2702), .RSTB(I180026), .Q(I179997) );
nor I_10433 (I180108,I180043,I557211);
nand I_10434 (I180125,I180108,I557187);
nand I_10435 (I180142,I180125,I180077);
not I_10436 (I180159,I557211);
not I_10437 (I180176,I557190);
nor I_10438 (I180193,I180176,I557193);
and I_10439 (I180210,I180193,I557196);
or I_10440 (I180227,I180210,I557205);
DFFARX1 I_10441  ( .D(I180227), .CLK(I2702), .RSTB(I180026), .Q(I180244) );
nor I_10442 (I180261,I180244,I180125);
nand I_10443 (I180012,I180159,I180261);
not I_10444 (I180009,I180244);
and I_10445 (I180306,I180244,I180142);
DFFARX1 I_10446  ( .D(I180306), .CLK(I2702), .RSTB(I180026), .Q(I179994) );
DFFARX1 I_10447  ( .D(I180244), .CLK(I2702), .RSTB(I180026), .Q(I180337) );
and I_10448 (I179991,I180159,I180337);
nand I_10449 (I180368,I180043,I557190);
not I_10450 (I180385,I180368);
nor I_10451 (I180402,I180244,I180385);
DFFARX1 I_10452  ( .D(I557208), .CLK(I2702), .RSTB(I180026), .Q(I180419) );
nand I_10453 (I180436,I180419,I180368);
and I_10454 (I180453,I180159,I180436);
DFFARX1 I_10455  ( .D(I180453), .CLK(I2702), .RSTB(I180026), .Q(I180018) );
not I_10456 (I180484,I180419);
nand I_10457 (I180006,I180419,I180402);
nand I_10458 (I180000,I180419,I180385);
DFFARX1 I_10459  ( .D(I557184), .CLK(I2702), .RSTB(I180026), .Q(I180529) );
not I_10460 (I180546,I180529);
nor I_10461 (I180015,I180419,I180546);
nor I_10462 (I180577,I180546,I180484);
and I_10463 (I180594,I180125,I180577);
or I_10464 (I180611,I180368,I180594);
DFFARX1 I_10465  ( .D(I180611), .CLK(I2702), .RSTB(I180026), .Q(I180003) );
DFFARX1 I_10466  ( .D(I180546), .CLK(I2702), .RSTB(I180026), .Q(I179988) );
not I_10467 (I180689,I2709);
not I_10468 (I180706,I337035);
nor I_10469 (I180723,I337044,I337017);
nand I_10470 (I180740,I180723,I337029);
DFFARX1 I_10471  ( .D(I180740), .CLK(I2702), .RSTB(I180689), .Q(I180660) );
nor I_10472 (I180771,I180706,I337044);
nand I_10473 (I180788,I180771,I337041);
nand I_10474 (I180805,I180788,I180740);
not I_10475 (I180822,I337044);
not I_10476 (I180839,I337020);
nor I_10477 (I180856,I180839,I337026);
and I_10478 (I180873,I180856,I337038);
or I_10479 (I180890,I180873,I337023);
DFFARX1 I_10480  ( .D(I180890), .CLK(I2702), .RSTB(I180689), .Q(I180907) );
nor I_10481 (I180924,I180907,I180788);
nand I_10482 (I180675,I180822,I180924);
not I_10483 (I180672,I180907);
and I_10484 (I180969,I180907,I180805);
DFFARX1 I_10485  ( .D(I180969), .CLK(I2702), .RSTB(I180689), .Q(I180657) );
DFFARX1 I_10486  ( .D(I180907), .CLK(I2702), .RSTB(I180689), .Q(I181000) );
and I_10487 (I180654,I180822,I181000);
nand I_10488 (I181031,I180706,I337020);
not I_10489 (I181048,I181031);
nor I_10490 (I181065,I180907,I181048);
DFFARX1 I_10491  ( .D(I337047), .CLK(I2702), .RSTB(I180689), .Q(I181082) );
nand I_10492 (I181099,I181082,I181031);
and I_10493 (I181116,I180822,I181099);
DFFARX1 I_10494  ( .D(I181116), .CLK(I2702), .RSTB(I180689), .Q(I180681) );
not I_10495 (I181147,I181082);
nand I_10496 (I180669,I181082,I181065);
nand I_10497 (I180663,I181082,I181048);
DFFARX1 I_10498  ( .D(I337032), .CLK(I2702), .RSTB(I180689), .Q(I181192) );
not I_10499 (I181209,I181192);
nor I_10500 (I180678,I181082,I181209);
nor I_10501 (I181240,I181209,I181147);
and I_10502 (I181257,I180788,I181240);
or I_10503 (I181274,I181031,I181257);
DFFARX1 I_10504  ( .D(I181274), .CLK(I2702), .RSTB(I180689), .Q(I180666) );
DFFARX1 I_10505  ( .D(I181209), .CLK(I2702), .RSTB(I180689), .Q(I180651) );
not I_10506 (I181352,I2709);
not I_10507 (I181369,I91756);
nor I_10508 (I181386,I91744,I91768);
nand I_10509 (I181403,I181386,I91753);
DFFARX1 I_10510  ( .D(I181403), .CLK(I2702), .RSTB(I181352), .Q(I181323) );
nor I_10511 (I181434,I181369,I91744);
nand I_10512 (I181451,I181434,I91771);
nand I_10513 (I181468,I181451,I181403);
not I_10514 (I181485,I91744);
not I_10515 (I181502,I91741);
nor I_10516 (I181519,I181502,I91750);
and I_10517 (I181536,I181519,I91765);
or I_10518 (I181553,I181536,I91747);
DFFARX1 I_10519  ( .D(I181553), .CLK(I2702), .RSTB(I181352), .Q(I181570) );
nor I_10520 (I181587,I181570,I181451);
nand I_10521 (I181338,I181485,I181587);
not I_10522 (I181335,I181570);
and I_10523 (I181632,I181570,I181468);
DFFARX1 I_10524  ( .D(I181632), .CLK(I2702), .RSTB(I181352), .Q(I181320) );
DFFARX1 I_10525  ( .D(I181570), .CLK(I2702), .RSTB(I181352), .Q(I181663) );
and I_10526 (I181317,I181485,I181663);
nand I_10527 (I181694,I181369,I91741);
not I_10528 (I181711,I181694);
nor I_10529 (I181728,I181570,I181711);
DFFARX1 I_10530  ( .D(I91762), .CLK(I2702), .RSTB(I181352), .Q(I181745) );
nand I_10531 (I181762,I181745,I181694);
and I_10532 (I181779,I181485,I181762);
DFFARX1 I_10533  ( .D(I181779), .CLK(I2702), .RSTB(I181352), .Q(I181344) );
not I_10534 (I181810,I181745);
nand I_10535 (I181332,I181745,I181728);
nand I_10536 (I181326,I181745,I181711);
DFFARX1 I_10537  ( .D(I91759), .CLK(I2702), .RSTB(I181352), .Q(I181855) );
not I_10538 (I181872,I181855);
nor I_10539 (I181341,I181745,I181872);
nor I_10540 (I181903,I181872,I181810);
and I_10541 (I181920,I181451,I181903);
or I_10542 (I181937,I181694,I181920);
DFFARX1 I_10543  ( .D(I181937), .CLK(I2702), .RSTB(I181352), .Q(I181329) );
DFFARX1 I_10544  ( .D(I181872), .CLK(I2702), .RSTB(I181352), .Q(I181314) );
not I_10545 (I182015,I2709);
not I_10546 (I182032,I246951);
nor I_10547 (I182049,I246960,I246972);
nand I_10548 (I182066,I182049,I246963);
DFFARX1 I_10549  ( .D(I182066), .CLK(I2702), .RSTB(I182015), .Q(I181986) );
nor I_10550 (I182097,I182032,I246960);
nand I_10551 (I182114,I182097,I246975);
nand I_10552 (I182131,I182114,I182066);
not I_10553 (I182148,I246960);
not I_10554 (I182165,I246981);
nor I_10555 (I182182,I182165,I246957);
and I_10556 (I182199,I182182,I246966);
or I_10557 (I182216,I182199,I246954);
DFFARX1 I_10558  ( .D(I182216), .CLK(I2702), .RSTB(I182015), .Q(I182233) );
nor I_10559 (I182250,I182233,I182114);
nand I_10560 (I182001,I182148,I182250);
not I_10561 (I181998,I182233);
and I_10562 (I182295,I182233,I182131);
DFFARX1 I_10563  ( .D(I182295), .CLK(I2702), .RSTB(I182015), .Q(I181983) );
DFFARX1 I_10564  ( .D(I182233), .CLK(I2702), .RSTB(I182015), .Q(I182326) );
and I_10565 (I181980,I182148,I182326);
nand I_10566 (I182357,I182032,I246981);
not I_10567 (I182374,I182357);
nor I_10568 (I182391,I182233,I182374);
DFFARX1 I_10569  ( .D(I246978), .CLK(I2702), .RSTB(I182015), .Q(I182408) );
nand I_10570 (I182425,I182408,I182357);
and I_10571 (I182442,I182148,I182425);
DFFARX1 I_10572  ( .D(I182442), .CLK(I2702), .RSTB(I182015), .Q(I182007) );
not I_10573 (I182473,I182408);
nand I_10574 (I181995,I182408,I182391);
nand I_10575 (I181989,I182408,I182374);
DFFARX1 I_10576  ( .D(I246969), .CLK(I2702), .RSTB(I182015), .Q(I182518) );
not I_10577 (I182535,I182518);
nor I_10578 (I182004,I182408,I182535);
nor I_10579 (I182566,I182535,I182473);
and I_10580 (I182583,I182114,I182566);
or I_10581 (I182600,I182357,I182583);
DFFARX1 I_10582  ( .D(I182600), .CLK(I2702), .RSTB(I182015), .Q(I181992) );
DFFARX1 I_10583  ( .D(I182535), .CLK(I2702), .RSTB(I182015), .Q(I181977) );
not I_10584 (I182678,I2709);
not I_10585 (I182695,I115012);
nor I_10586 (I182712,I115000,I115024);
nand I_10587 (I182729,I182712,I115009);
DFFARX1 I_10588  ( .D(I182729), .CLK(I2702), .RSTB(I182678), .Q(I182649) );
nor I_10589 (I182760,I182695,I115000);
nand I_10590 (I182777,I182760,I115027);
nand I_10591 (I182794,I182777,I182729);
not I_10592 (I182811,I115000);
not I_10593 (I182828,I114997);
nor I_10594 (I182845,I182828,I115006);
and I_10595 (I182862,I182845,I115021);
or I_10596 (I182879,I182862,I115003);
DFFARX1 I_10597  ( .D(I182879), .CLK(I2702), .RSTB(I182678), .Q(I182896) );
nor I_10598 (I182913,I182896,I182777);
nand I_10599 (I182664,I182811,I182913);
not I_10600 (I182661,I182896);
and I_10601 (I182958,I182896,I182794);
DFFARX1 I_10602  ( .D(I182958), .CLK(I2702), .RSTB(I182678), .Q(I182646) );
DFFARX1 I_10603  ( .D(I182896), .CLK(I2702), .RSTB(I182678), .Q(I182989) );
and I_10604 (I182643,I182811,I182989);
nand I_10605 (I183020,I182695,I114997);
not I_10606 (I183037,I183020);
nor I_10607 (I183054,I182896,I183037);
DFFARX1 I_10608  ( .D(I115018), .CLK(I2702), .RSTB(I182678), .Q(I183071) );
nand I_10609 (I183088,I183071,I183020);
and I_10610 (I183105,I182811,I183088);
DFFARX1 I_10611  ( .D(I183105), .CLK(I2702), .RSTB(I182678), .Q(I182670) );
not I_10612 (I183136,I183071);
nand I_10613 (I182658,I183071,I183054);
nand I_10614 (I182652,I183071,I183037);
DFFARX1 I_10615  ( .D(I115015), .CLK(I2702), .RSTB(I182678), .Q(I183181) );
not I_10616 (I183198,I183181);
nor I_10617 (I182667,I183071,I183198);
nor I_10618 (I183229,I183198,I183136);
and I_10619 (I183246,I182777,I183229);
or I_10620 (I183263,I183020,I183246);
DFFARX1 I_10621  ( .D(I183263), .CLK(I2702), .RSTB(I182678), .Q(I182655) );
DFFARX1 I_10622  ( .D(I183198), .CLK(I2702), .RSTB(I182678), .Q(I182640) );
not I_10623 (I183341,I2709);
not I_10624 (I183358,I34143);
nor I_10625 (I183375,I34131,I34134);
nand I_10626 (I183392,I183375,I34149);
DFFARX1 I_10627  ( .D(I183392), .CLK(I2702), .RSTB(I183341), .Q(I183312) );
nor I_10628 (I183423,I183358,I34131);
nand I_10629 (I183440,I183423,I34140);
nand I_10630 (I183457,I183440,I183392);
not I_10631 (I183474,I34131);
not I_10632 (I183491,I34152);
nor I_10633 (I183508,I183491,I34128);
and I_10634 (I183525,I183508,I34137);
or I_10635 (I183542,I183525,I34146);
DFFARX1 I_10636  ( .D(I183542), .CLK(I2702), .RSTB(I183341), .Q(I183559) );
nor I_10637 (I183576,I183559,I183440);
nand I_10638 (I183327,I183474,I183576);
not I_10639 (I183324,I183559);
and I_10640 (I183621,I183559,I183457);
DFFARX1 I_10641  ( .D(I183621), .CLK(I2702), .RSTB(I183341), .Q(I183309) );
DFFARX1 I_10642  ( .D(I183559), .CLK(I2702), .RSTB(I183341), .Q(I183652) );
and I_10643 (I183306,I183474,I183652);
nand I_10644 (I183683,I183358,I34152);
not I_10645 (I183700,I183683);
nor I_10646 (I183717,I183559,I183700);
DFFARX1 I_10647  ( .D(I34158), .CLK(I2702), .RSTB(I183341), .Q(I183734) );
nand I_10648 (I183751,I183734,I183683);
and I_10649 (I183768,I183474,I183751);
DFFARX1 I_10650  ( .D(I183768), .CLK(I2702), .RSTB(I183341), .Q(I183333) );
not I_10651 (I183799,I183734);
nand I_10652 (I183321,I183734,I183717);
nand I_10653 (I183315,I183734,I183700);
DFFARX1 I_10654  ( .D(I34155), .CLK(I2702), .RSTB(I183341), .Q(I183844) );
not I_10655 (I183861,I183844);
nor I_10656 (I183330,I183734,I183861);
nor I_10657 (I183892,I183861,I183799);
and I_10658 (I183909,I183440,I183892);
or I_10659 (I183926,I183683,I183909);
DFFARX1 I_10660  ( .D(I183926), .CLK(I2702), .RSTB(I183341), .Q(I183318) );
DFFARX1 I_10661  ( .D(I183861), .CLK(I2702), .RSTB(I183341), .Q(I183303) );
not I_10662 (I184004,I2709);
not I_10663 (I184021,I605385);
nor I_10664 (I184038,I605400,I605382);
nand I_10665 (I184055,I184038,I605394);
DFFARX1 I_10666  ( .D(I184055), .CLK(I2702), .RSTB(I184004), .Q(I183975) );
nor I_10667 (I184086,I184021,I605400);
nand I_10668 (I184103,I184086,I605391);
nand I_10669 (I184120,I184103,I184055);
not I_10670 (I184137,I605400);
not I_10671 (I184154,I605409);
nor I_10672 (I184171,I184154,I605379);
and I_10673 (I184188,I184171,I605388);
or I_10674 (I184205,I184188,I605406);
DFFARX1 I_10675  ( .D(I184205), .CLK(I2702), .RSTB(I184004), .Q(I184222) );
nor I_10676 (I184239,I184222,I184103);
nand I_10677 (I183990,I184137,I184239);
not I_10678 (I183987,I184222);
and I_10679 (I184284,I184222,I184120);
DFFARX1 I_10680  ( .D(I184284), .CLK(I2702), .RSTB(I184004), .Q(I183972) );
DFFARX1 I_10681  ( .D(I184222), .CLK(I2702), .RSTB(I184004), .Q(I184315) );
and I_10682 (I183969,I184137,I184315);
nand I_10683 (I184346,I184021,I605409);
not I_10684 (I184363,I184346);
nor I_10685 (I184380,I184222,I184363);
DFFARX1 I_10686  ( .D(I605397), .CLK(I2702), .RSTB(I184004), .Q(I184397) );
nand I_10687 (I184414,I184397,I184346);
and I_10688 (I184431,I184137,I184414);
DFFARX1 I_10689  ( .D(I184431), .CLK(I2702), .RSTB(I184004), .Q(I183996) );
not I_10690 (I184462,I184397);
nand I_10691 (I183984,I184397,I184380);
nand I_10692 (I183978,I184397,I184363);
DFFARX1 I_10693  ( .D(I605403), .CLK(I2702), .RSTB(I184004), .Q(I184507) );
not I_10694 (I184524,I184507);
nor I_10695 (I183993,I184397,I184524);
nor I_10696 (I184555,I184524,I184462);
and I_10697 (I184572,I184103,I184555);
or I_10698 (I184589,I184346,I184572);
DFFARX1 I_10699  ( .D(I184589), .CLK(I2702), .RSTB(I184004), .Q(I183981) );
DFFARX1 I_10700  ( .D(I184524), .CLK(I2702), .RSTB(I184004), .Q(I183966) );
not I_10701 (I184667,I2709);
not I_10702 (I184684,I217752);
nor I_10703 (I184701,I217734,I217728);
nand I_10704 (I184718,I184701,I217731);
DFFARX1 I_10705  ( .D(I184718), .CLK(I2702), .RSTB(I184667), .Q(I184638) );
nor I_10706 (I184749,I184684,I217734);
nand I_10707 (I184766,I184749,I217740);
nand I_10708 (I184783,I184766,I184718);
not I_10709 (I184800,I217734);
not I_10710 (I184817,I217749);
nor I_10711 (I184834,I184817,I217737);
and I_10712 (I184851,I184834,I217743);
or I_10713 (I184868,I184851,I217758);
DFFARX1 I_10714  ( .D(I184868), .CLK(I2702), .RSTB(I184667), .Q(I184885) );
nor I_10715 (I184902,I184885,I184766);
nand I_10716 (I184653,I184800,I184902);
not I_10717 (I184650,I184885);
and I_10718 (I184947,I184885,I184783);
DFFARX1 I_10719  ( .D(I184947), .CLK(I2702), .RSTB(I184667), .Q(I184635) );
DFFARX1 I_10720  ( .D(I184885), .CLK(I2702), .RSTB(I184667), .Q(I184978) );
and I_10721 (I184632,I184800,I184978);
nand I_10722 (I185009,I184684,I217749);
not I_10723 (I185026,I185009);
nor I_10724 (I185043,I184885,I185026);
DFFARX1 I_10725  ( .D(I217746), .CLK(I2702), .RSTB(I184667), .Q(I185060) );
nand I_10726 (I185077,I185060,I185009);
and I_10727 (I185094,I184800,I185077);
DFFARX1 I_10728  ( .D(I185094), .CLK(I2702), .RSTB(I184667), .Q(I184659) );
not I_10729 (I185125,I185060);
nand I_10730 (I184647,I185060,I185043);
nand I_10731 (I184641,I185060,I185026);
DFFARX1 I_10732  ( .D(I217755), .CLK(I2702), .RSTB(I184667), .Q(I185170) );
not I_10733 (I185187,I185170);
nor I_10734 (I184656,I185060,I185187);
nor I_10735 (I185218,I185187,I185125);
and I_10736 (I185235,I184766,I185218);
or I_10737 (I185252,I185009,I185235);
DFFARX1 I_10738  ( .D(I185252), .CLK(I2702), .RSTB(I184667), .Q(I184644) );
DFFARX1 I_10739  ( .D(I185187), .CLK(I2702), .RSTB(I184667), .Q(I184629) );
not I_10740 (I185330,I2709);
not I_10741 (I185347,I539349);
nor I_10742 (I185364,I539361,I539364);
nand I_10743 (I185381,I185364,I539352);
DFFARX1 I_10744  ( .D(I185381), .CLK(I2702), .RSTB(I185330), .Q(I185301) );
nor I_10745 (I185412,I185347,I539361);
nand I_10746 (I185429,I185412,I539337);
nand I_10747 (I185446,I185429,I185381);
not I_10748 (I185463,I539361);
not I_10749 (I185480,I539340);
nor I_10750 (I185497,I185480,I539343);
and I_10751 (I185514,I185497,I539346);
or I_10752 (I185531,I185514,I539355);
DFFARX1 I_10753  ( .D(I185531), .CLK(I2702), .RSTB(I185330), .Q(I185548) );
nor I_10754 (I185565,I185548,I185429);
nand I_10755 (I185316,I185463,I185565);
not I_10756 (I185313,I185548);
and I_10757 (I185610,I185548,I185446);
DFFARX1 I_10758  ( .D(I185610), .CLK(I2702), .RSTB(I185330), .Q(I185298) );
DFFARX1 I_10759  ( .D(I185548), .CLK(I2702), .RSTB(I185330), .Q(I185641) );
and I_10760 (I185295,I185463,I185641);
nand I_10761 (I185672,I185347,I539340);
not I_10762 (I185689,I185672);
nor I_10763 (I185706,I185548,I185689);
DFFARX1 I_10764  ( .D(I539358), .CLK(I2702), .RSTB(I185330), .Q(I185723) );
nand I_10765 (I185740,I185723,I185672);
and I_10766 (I185757,I185463,I185740);
DFFARX1 I_10767  ( .D(I185757), .CLK(I2702), .RSTB(I185330), .Q(I185322) );
not I_10768 (I185788,I185723);
nand I_10769 (I185310,I185723,I185706);
nand I_10770 (I185304,I185723,I185689);
DFFARX1 I_10771  ( .D(I539334), .CLK(I2702), .RSTB(I185330), .Q(I185833) );
not I_10772 (I185850,I185833);
nor I_10773 (I185319,I185723,I185850);
nor I_10774 (I185881,I185850,I185788);
and I_10775 (I185898,I185429,I185881);
or I_10776 (I185915,I185672,I185898);
DFFARX1 I_10777  ( .D(I185915), .CLK(I2702), .RSTB(I185330), .Q(I185307) );
DFFARX1 I_10778  ( .D(I185850), .CLK(I2702), .RSTB(I185330), .Q(I185292) );
not I_10779 (I185993,I2709);
not I_10780 (I186010,I662749);
nor I_10781 (I186027,I662755,I662767);
nand I_10782 (I186044,I186027,I662758);
DFFARX1 I_10783  ( .D(I186044), .CLK(I2702), .RSTB(I185993), .Q(I185964) );
nor I_10784 (I186075,I186010,I662755);
nand I_10785 (I186092,I186075,I662737);
nand I_10786 (I186109,I186092,I186044);
not I_10787 (I186126,I662755);
not I_10788 (I186143,I662752);
nor I_10789 (I186160,I186143,I662740);
and I_10790 (I186177,I186160,I662761);
or I_10791 (I186194,I186177,I662743);
DFFARX1 I_10792  ( .D(I186194), .CLK(I2702), .RSTB(I185993), .Q(I186211) );
nor I_10793 (I186228,I186211,I186092);
nand I_10794 (I185979,I186126,I186228);
not I_10795 (I185976,I186211);
and I_10796 (I186273,I186211,I186109);
DFFARX1 I_10797  ( .D(I186273), .CLK(I2702), .RSTB(I185993), .Q(I185961) );
DFFARX1 I_10798  ( .D(I186211), .CLK(I2702), .RSTB(I185993), .Q(I186304) );
and I_10799 (I185958,I186126,I186304);
nand I_10800 (I186335,I186010,I662752);
not I_10801 (I186352,I186335);
nor I_10802 (I186369,I186211,I186352);
DFFARX1 I_10803  ( .D(I662764), .CLK(I2702), .RSTB(I185993), .Q(I186386) );
nand I_10804 (I186403,I186386,I186335);
and I_10805 (I186420,I186126,I186403);
DFFARX1 I_10806  ( .D(I186420), .CLK(I2702), .RSTB(I185993), .Q(I185985) );
not I_10807 (I186451,I186386);
nand I_10808 (I185973,I186386,I186369);
nand I_10809 (I185967,I186386,I186352);
DFFARX1 I_10810  ( .D(I662746), .CLK(I2702), .RSTB(I185993), .Q(I186496) );
not I_10811 (I186513,I186496);
nor I_10812 (I185982,I186386,I186513);
nor I_10813 (I186544,I186513,I186451);
and I_10814 (I186561,I186092,I186544);
or I_10815 (I186578,I186335,I186561);
DFFARX1 I_10816  ( .D(I186578), .CLK(I2702), .RSTB(I185993), .Q(I185970) );
DFFARX1 I_10817  ( .D(I186513), .CLK(I2702), .RSTB(I185993), .Q(I185955) );
not I_10818 (I186656,I2709);
not I_10819 (I186673,I68500);
nor I_10820 (I186690,I68488,I68512);
nand I_10821 (I186707,I186690,I68497);
DFFARX1 I_10822  ( .D(I186707), .CLK(I2702), .RSTB(I186656), .Q(I186627) );
nor I_10823 (I186738,I186673,I68488);
nand I_10824 (I186755,I186738,I68515);
nand I_10825 (I186772,I186755,I186707);
not I_10826 (I186789,I68488);
not I_10827 (I186806,I68485);
nor I_10828 (I186823,I186806,I68494);
and I_10829 (I186840,I186823,I68509);
or I_10830 (I186857,I186840,I68491);
DFFARX1 I_10831  ( .D(I186857), .CLK(I2702), .RSTB(I186656), .Q(I186874) );
nor I_10832 (I186891,I186874,I186755);
nand I_10833 (I186642,I186789,I186891);
not I_10834 (I186639,I186874);
and I_10835 (I186936,I186874,I186772);
DFFARX1 I_10836  ( .D(I186936), .CLK(I2702), .RSTB(I186656), .Q(I186624) );
DFFARX1 I_10837  ( .D(I186874), .CLK(I2702), .RSTB(I186656), .Q(I186967) );
and I_10838 (I186621,I186789,I186967);
nand I_10839 (I186998,I186673,I68485);
not I_10840 (I187015,I186998);
nor I_10841 (I187032,I186874,I187015);
DFFARX1 I_10842  ( .D(I68506), .CLK(I2702), .RSTB(I186656), .Q(I187049) );
nand I_10843 (I187066,I187049,I186998);
and I_10844 (I187083,I186789,I187066);
DFFARX1 I_10845  ( .D(I187083), .CLK(I2702), .RSTB(I186656), .Q(I186648) );
not I_10846 (I187114,I187049);
nand I_10847 (I186636,I187049,I187032);
nand I_10848 (I186630,I187049,I187015);
DFFARX1 I_10849  ( .D(I68503), .CLK(I2702), .RSTB(I186656), .Q(I187159) );
not I_10850 (I187176,I187159);
nor I_10851 (I186645,I187049,I187176);
nor I_10852 (I187207,I187176,I187114);
and I_10853 (I187224,I186755,I187207);
or I_10854 (I187241,I186998,I187224);
DFFARX1 I_10855  ( .D(I187241), .CLK(I2702), .RSTB(I186656), .Q(I186633) );
DFFARX1 I_10856  ( .D(I187176), .CLK(I2702), .RSTB(I186656), .Q(I186618) );
not I_10857 (I187319,I2709);
not I_10858 (I187336,I487643);
nor I_10859 (I187353,I487649,I487640);
nand I_10860 (I187370,I187353,I487658);
DFFARX1 I_10861  ( .D(I187370), .CLK(I2702), .RSTB(I187319), .Q(I187290) );
nor I_10862 (I187401,I187336,I487649);
nand I_10863 (I187418,I187401,I487637);
nand I_10864 (I187435,I187418,I187370);
not I_10865 (I187452,I487649);
not I_10866 (I187469,I487667);
nor I_10867 (I187486,I187469,I487646);
and I_10868 (I187503,I187486,I487655);
or I_10869 (I187520,I187503,I487661);
DFFARX1 I_10870  ( .D(I187520), .CLK(I2702), .RSTB(I187319), .Q(I187537) );
nor I_10871 (I187554,I187537,I187418);
nand I_10872 (I187305,I187452,I187554);
not I_10873 (I187302,I187537);
and I_10874 (I187599,I187537,I187435);
DFFARX1 I_10875  ( .D(I187599), .CLK(I2702), .RSTB(I187319), .Q(I187287) );
DFFARX1 I_10876  ( .D(I187537), .CLK(I2702), .RSTB(I187319), .Q(I187630) );
and I_10877 (I187284,I187452,I187630);
nand I_10878 (I187661,I187336,I487667);
not I_10879 (I187678,I187661);
nor I_10880 (I187695,I187537,I187678);
DFFARX1 I_10881  ( .D(I487652), .CLK(I2702), .RSTB(I187319), .Q(I187712) );
nand I_10882 (I187729,I187712,I187661);
and I_10883 (I187746,I187452,I187729);
DFFARX1 I_10884  ( .D(I187746), .CLK(I2702), .RSTB(I187319), .Q(I187311) );
not I_10885 (I187777,I187712);
nand I_10886 (I187299,I187712,I187695);
nand I_10887 (I187293,I187712,I187678);
DFFARX1 I_10888  ( .D(I487664), .CLK(I2702), .RSTB(I187319), .Q(I187822) );
not I_10889 (I187839,I187822);
nor I_10890 (I187308,I187712,I187839);
nor I_10891 (I187870,I187839,I187777);
and I_10892 (I187887,I187418,I187870);
or I_10893 (I187904,I187661,I187887);
DFFARX1 I_10894  ( .D(I187904), .CLK(I2702), .RSTB(I187319), .Q(I187296) );
DFFARX1 I_10895  ( .D(I187839), .CLK(I2702), .RSTB(I187319), .Q(I187281) );
not I_10896 (I187982,I2709);
not I_10897 (I187999,I452923);
nor I_10898 (I188016,I452929,I452926);
nand I_10899 (I188033,I188016,I452944);
DFFARX1 I_10900  ( .D(I188033), .CLK(I2702), .RSTB(I187982), .Q(I187953) );
nor I_10901 (I188064,I187999,I452929);
nand I_10902 (I188081,I188064,I452953);
nand I_10903 (I188098,I188081,I188033);
not I_10904 (I188115,I452929);
not I_10905 (I188132,I452947);
nor I_10906 (I188149,I188132,I452938);
and I_10907 (I188166,I188149,I452941);
or I_10908 (I188183,I188166,I452932);
DFFARX1 I_10909  ( .D(I188183), .CLK(I2702), .RSTB(I187982), .Q(I188200) );
nor I_10910 (I188217,I188200,I188081);
nand I_10911 (I187968,I188115,I188217);
not I_10912 (I187965,I188200);
and I_10913 (I188262,I188200,I188098);
DFFARX1 I_10914  ( .D(I188262), .CLK(I2702), .RSTB(I187982), .Q(I187950) );
DFFARX1 I_10915  ( .D(I188200), .CLK(I2702), .RSTB(I187982), .Q(I188293) );
and I_10916 (I187947,I188115,I188293);
nand I_10917 (I188324,I187999,I452947);
not I_10918 (I188341,I188324);
nor I_10919 (I188358,I188200,I188341);
DFFARX1 I_10920  ( .D(I452950), .CLK(I2702), .RSTB(I187982), .Q(I188375) );
nand I_10921 (I188392,I188375,I188324);
and I_10922 (I188409,I188115,I188392);
DFFARX1 I_10923  ( .D(I188409), .CLK(I2702), .RSTB(I187982), .Q(I187974) );
not I_10924 (I188440,I188375);
nand I_10925 (I187962,I188375,I188358);
nand I_10926 (I187956,I188375,I188341);
DFFARX1 I_10927  ( .D(I452935), .CLK(I2702), .RSTB(I187982), .Q(I188485) );
not I_10928 (I188502,I188485);
nor I_10929 (I187971,I188375,I188502);
nor I_10930 (I188533,I188502,I188440);
and I_10931 (I188550,I188081,I188533);
or I_10932 (I188567,I188324,I188550);
DFFARX1 I_10933  ( .D(I188567), .CLK(I2702), .RSTB(I187982), .Q(I187959) );
DFFARX1 I_10934  ( .D(I188502), .CLK(I2702), .RSTB(I187982), .Q(I187944) );
not I_10935 (I188645,I2709);
not I_10936 (I188662,I322533);
nor I_10937 (I188679,I322542,I322554);
nand I_10938 (I188696,I188679,I322545);
DFFARX1 I_10939  ( .D(I188696), .CLK(I2702), .RSTB(I188645), .Q(I188616) );
nor I_10940 (I188727,I188662,I322542);
nand I_10941 (I188744,I188727,I322557);
nand I_10942 (I188761,I188744,I188696);
not I_10943 (I188778,I322542);
not I_10944 (I188795,I322563);
nor I_10945 (I188812,I188795,I322539);
and I_10946 (I188829,I188812,I322548);
or I_10947 (I188846,I188829,I322536);
DFFARX1 I_10948  ( .D(I188846), .CLK(I2702), .RSTB(I188645), .Q(I188863) );
nor I_10949 (I188880,I188863,I188744);
nand I_10950 (I188631,I188778,I188880);
not I_10951 (I188628,I188863);
and I_10952 (I188925,I188863,I188761);
DFFARX1 I_10953  ( .D(I188925), .CLK(I2702), .RSTB(I188645), .Q(I188613) );
DFFARX1 I_10954  ( .D(I188863), .CLK(I2702), .RSTB(I188645), .Q(I188956) );
and I_10955 (I188610,I188778,I188956);
nand I_10956 (I188987,I188662,I322563);
not I_10957 (I189004,I188987);
nor I_10958 (I189021,I188863,I189004);
DFFARX1 I_10959  ( .D(I322560), .CLK(I2702), .RSTB(I188645), .Q(I189038) );
nand I_10960 (I189055,I189038,I188987);
and I_10961 (I189072,I188778,I189055);
DFFARX1 I_10962  ( .D(I189072), .CLK(I2702), .RSTB(I188645), .Q(I188637) );
not I_10963 (I189103,I189038);
nand I_10964 (I188625,I189038,I189021);
nand I_10965 (I188619,I189038,I189004);
DFFARX1 I_10966  ( .D(I322551), .CLK(I2702), .RSTB(I188645), .Q(I189148) );
not I_10967 (I189165,I189148);
nor I_10968 (I188634,I189038,I189165);
nor I_10969 (I189196,I189165,I189103);
and I_10970 (I189213,I188744,I189196);
or I_10971 (I189230,I188987,I189213);
DFFARX1 I_10972  ( .D(I189230), .CLK(I2702), .RSTB(I188645), .Q(I188622) );
DFFARX1 I_10973  ( .D(I189165), .CLK(I2702), .RSTB(I188645), .Q(I188607) );
not I_10974 (I189308,I2709);
not I_10975 (I189325,I362229);
nor I_10976 (I189342,I362238,I362211);
nand I_10977 (I189359,I189342,I362223);
DFFARX1 I_10978  ( .D(I189359), .CLK(I2702), .RSTB(I189308), .Q(I189279) );
nor I_10979 (I189390,I189325,I362238);
nand I_10980 (I189407,I189390,I362235);
nand I_10981 (I189424,I189407,I189359);
not I_10982 (I189441,I362238);
not I_10983 (I189458,I362214);
nor I_10984 (I189475,I189458,I362220);
and I_10985 (I189492,I189475,I362232);
or I_10986 (I189509,I189492,I362217);
DFFARX1 I_10987  ( .D(I189509), .CLK(I2702), .RSTB(I189308), .Q(I189526) );
nor I_10988 (I189543,I189526,I189407);
nand I_10989 (I189294,I189441,I189543);
not I_10990 (I189291,I189526);
and I_10991 (I189588,I189526,I189424);
DFFARX1 I_10992  ( .D(I189588), .CLK(I2702), .RSTB(I189308), .Q(I189276) );
DFFARX1 I_10993  ( .D(I189526), .CLK(I2702), .RSTB(I189308), .Q(I189619) );
and I_10994 (I189273,I189441,I189619);
nand I_10995 (I189650,I189325,I362214);
not I_10996 (I189667,I189650);
nor I_10997 (I189684,I189526,I189667);
DFFARX1 I_10998  ( .D(I362241), .CLK(I2702), .RSTB(I189308), .Q(I189701) );
nand I_10999 (I189718,I189701,I189650);
and I_11000 (I189735,I189441,I189718);
DFFARX1 I_11001  ( .D(I189735), .CLK(I2702), .RSTB(I189308), .Q(I189300) );
not I_11002 (I189766,I189701);
nand I_11003 (I189288,I189701,I189684);
nand I_11004 (I189282,I189701,I189667);
DFFARX1 I_11005  ( .D(I362226), .CLK(I2702), .RSTB(I189308), .Q(I189811) );
not I_11006 (I189828,I189811);
nor I_11007 (I189297,I189701,I189828);
nor I_11008 (I189859,I189828,I189766);
and I_11009 (I189876,I189407,I189859);
or I_11010 (I189893,I189650,I189876);
DFFARX1 I_11011  ( .D(I189893), .CLK(I2702), .RSTB(I189308), .Q(I189285) );
DFFARX1 I_11012  ( .D(I189828), .CLK(I2702), .RSTB(I189308), .Q(I189270) );
not I_11013 (I189971,I2709);
not I_11014 (I189988,I476621);
nor I_11015 (I190005,I476627,I476624);
nand I_11016 (I190022,I190005,I476642);
DFFARX1 I_11017  ( .D(I190022), .CLK(I2702), .RSTB(I189971), .Q(I189942) );
nor I_11018 (I190053,I189988,I476627);
nand I_11019 (I190070,I190053,I476651);
nand I_11020 (I190087,I190070,I190022);
not I_11021 (I190104,I476627);
not I_11022 (I190121,I476645);
nor I_11023 (I190138,I190121,I476636);
and I_11024 (I190155,I190138,I476639);
or I_11025 (I190172,I190155,I476630);
DFFARX1 I_11026  ( .D(I190172), .CLK(I2702), .RSTB(I189971), .Q(I190189) );
nor I_11027 (I190206,I190189,I190070);
nand I_11028 (I189957,I190104,I190206);
not I_11029 (I189954,I190189);
and I_11030 (I190251,I190189,I190087);
DFFARX1 I_11031  ( .D(I190251), .CLK(I2702), .RSTB(I189971), .Q(I189939) );
DFFARX1 I_11032  ( .D(I190189), .CLK(I2702), .RSTB(I189971), .Q(I190282) );
and I_11033 (I189936,I190104,I190282);
nand I_11034 (I190313,I189988,I476645);
not I_11035 (I190330,I190313);
nor I_11036 (I190347,I190189,I190330);
DFFARX1 I_11037  ( .D(I476648), .CLK(I2702), .RSTB(I189971), .Q(I190364) );
nand I_11038 (I190381,I190364,I190313);
and I_11039 (I190398,I190104,I190381);
DFFARX1 I_11040  ( .D(I190398), .CLK(I2702), .RSTB(I189971), .Q(I189963) );
not I_11041 (I190429,I190364);
nand I_11042 (I189951,I190364,I190347);
nand I_11043 (I189945,I190364,I190330);
DFFARX1 I_11044  ( .D(I476633), .CLK(I2702), .RSTB(I189971), .Q(I190474) );
not I_11045 (I190491,I190474);
nor I_11046 (I189960,I190364,I190491);
nor I_11047 (I190522,I190491,I190429);
and I_11048 (I190539,I190070,I190522);
or I_11049 (I190556,I190313,I190539);
DFFARX1 I_11050  ( .D(I190556), .CLK(I2702), .RSTB(I189971), .Q(I189948) );
DFFARX1 I_11051  ( .D(I190491), .CLK(I2702), .RSTB(I189971), .Q(I189933) );
not I_11052 (I190634,I2709);
not I_11053 (I190651,I304632);
nor I_11054 (I190668,I304641,I304653);
nand I_11055 (I190685,I190668,I304644);
DFFARX1 I_11056  ( .D(I190685), .CLK(I2702), .RSTB(I190634), .Q(I190605) );
nor I_11057 (I190716,I190651,I304641);
nand I_11058 (I190733,I190716,I304656);
nand I_11059 (I190750,I190733,I190685);
not I_11060 (I190767,I304641);
not I_11061 (I190784,I304662);
nor I_11062 (I190801,I190784,I304638);
and I_11063 (I190818,I190801,I304647);
or I_11064 (I190835,I190818,I304635);
DFFARX1 I_11065  ( .D(I190835), .CLK(I2702), .RSTB(I190634), .Q(I190852) );
nor I_11066 (I190869,I190852,I190733);
nand I_11067 (I190620,I190767,I190869);
not I_11068 (I190617,I190852);
and I_11069 (I190914,I190852,I190750);
DFFARX1 I_11070  ( .D(I190914), .CLK(I2702), .RSTB(I190634), .Q(I190602) );
DFFARX1 I_11071  ( .D(I190852), .CLK(I2702), .RSTB(I190634), .Q(I190945) );
and I_11072 (I190599,I190767,I190945);
nand I_11073 (I190976,I190651,I304662);
not I_11074 (I190993,I190976);
nor I_11075 (I191010,I190852,I190993);
DFFARX1 I_11076  ( .D(I304659), .CLK(I2702), .RSTB(I190634), .Q(I191027) );
nand I_11077 (I191044,I191027,I190976);
and I_11078 (I191061,I190767,I191044);
DFFARX1 I_11079  ( .D(I191061), .CLK(I2702), .RSTB(I190634), .Q(I190626) );
not I_11080 (I191092,I191027);
nand I_11081 (I190614,I191027,I191010);
nand I_11082 (I190608,I191027,I190993);
DFFARX1 I_11083  ( .D(I304650), .CLK(I2702), .RSTB(I190634), .Q(I191137) );
not I_11084 (I191154,I191137);
nor I_11085 (I190623,I191027,I191154);
nor I_11086 (I191185,I191154,I191092);
and I_11087 (I191202,I190733,I191185);
or I_11088 (I191219,I190976,I191202);
DFFARX1 I_11089  ( .D(I191219), .CLK(I2702), .RSTB(I190634), .Q(I190611) );
DFFARX1 I_11090  ( .D(I191154), .CLK(I2702), .RSTB(I190634), .Q(I190596) );
not I_11091 (I191297,I2709);
not I_11092 (I191314,I462171);
nor I_11093 (I191331,I462177,I462174);
nand I_11094 (I191348,I191331,I462192);
DFFARX1 I_11095  ( .D(I191348), .CLK(I2702), .RSTB(I191297), .Q(I191268) );
nor I_11096 (I191379,I191314,I462177);
nand I_11097 (I191396,I191379,I462201);
nand I_11098 (I191413,I191396,I191348);
not I_11099 (I191430,I462177);
not I_11100 (I191447,I462195);
nor I_11101 (I191464,I191447,I462186);
and I_11102 (I191481,I191464,I462189);
or I_11103 (I191498,I191481,I462180);
DFFARX1 I_11104  ( .D(I191498), .CLK(I2702), .RSTB(I191297), .Q(I191515) );
nor I_11105 (I191532,I191515,I191396);
nand I_11106 (I191283,I191430,I191532);
not I_11107 (I191280,I191515);
and I_11108 (I191577,I191515,I191413);
DFFARX1 I_11109  ( .D(I191577), .CLK(I2702), .RSTB(I191297), .Q(I191265) );
DFFARX1 I_11110  ( .D(I191515), .CLK(I2702), .RSTB(I191297), .Q(I191608) );
and I_11111 (I191262,I191430,I191608);
nand I_11112 (I191639,I191314,I462195);
not I_11113 (I191656,I191639);
nor I_11114 (I191673,I191515,I191656);
DFFARX1 I_11115  ( .D(I462198), .CLK(I2702), .RSTB(I191297), .Q(I191690) );
nand I_11116 (I191707,I191690,I191639);
and I_11117 (I191724,I191430,I191707);
DFFARX1 I_11118  ( .D(I191724), .CLK(I2702), .RSTB(I191297), .Q(I191289) );
not I_11119 (I191755,I191690);
nand I_11120 (I191277,I191690,I191673);
nand I_11121 (I191271,I191690,I191656);
DFFARX1 I_11122  ( .D(I462183), .CLK(I2702), .RSTB(I191297), .Q(I191800) );
not I_11123 (I191817,I191800);
nor I_11124 (I191286,I191690,I191817);
nor I_11125 (I191848,I191817,I191755);
and I_11126 (I191865,I191396,I191848);
or I_11127 (I191882,I191639,I191865);
DFFARX1 I_11128  ( .D(I191882), .CLK(I2702), .RSTB(I191297), .Q(I191274) );
DFFARX1 I_11129  ( .D(I191817), .CLK(I2702), .RSTB(I191297), .Q(I191259) );
not I_11130 (I191960,I2709);
not I_11131 (I191977,I377087);
nor I_11132 (I191994,I377096,I377069);
nand I_11133 (I192011,I191994,I377081);
DFFARX1 I_11134  ( .D(I192011), .CLK(I2702), .RSTB(I191960), .Q(I191931) );
nor I_11135 (I192042,I191977,I377096);
nand I_11136 (I192059,I192042,I377093);
nand I_11137 (I192076,I192059,I192011);
not I_11138 (I192093,I377096);
not I_11139 (I192110,I377072);
nor I_11140 (I192127,I192110,I377078);
and I_11141 (I192144,I192127,I377090);
or I_11142 (I192161,I192144,I377075);
DFFARX1 I_11143  ( .D(I192161), .CLK(I2702), .RSTB(I191960), .Q(I192178) );
nor I_11144 (I192195,I192178,I192059);
nand I_11145 (I191946,I192093,I192195);
not I_11146 (I191943,I192178);
and I_11147 (I192240,I192178,I192076);
DFFARX1 I_11148  ( .D(I192240), .CLK(I2702), .RSTB(I191960), .Q(I191928) );
DFFARX1 I_11149  ( .D(I192178), .CLK(I2702), .RSTB(I191960), .Q(I192271) );
and I_11150 (I191925,I192093,I192271);
nand I_11151 (I192302,I191977,I377072);
not I_11152 (I192319,I192302);
nor I_11153 (I192336,I192178,I192319);
DFFARX1 I_11154  ( .D(I377099), .CLK(I2702), .RSTB(I191960), .Q(I192353) );
nand I_11155 (I192370,I192353,I192302);
and I_11156 (I192387,I192093,I192370);
DFFARX1 I_11157  ( .D(I192387), .CLK(I2702), .RSTB(I191960), .Q(I191952) );
not I_11158 (I192418,I192353);
nand I_11159 (I191940,I192353,I192336);
nand I_11160 (I191934,I192353,I192319);
DFFARX1 I_11161  ( .D(I377084), .CLK(I2702), .RSTB(I191960), .Q(I192463) );
not I_11162 (I192480,I192463);
nor I_11163 (I191949,I192353,I192480);
nor I_11164 (I192511,I192480,I192418);
and I_11165 (I192528,I192059,I192511);
or I_11166 (I192545,I192302,I192528);
DFFARX1 I_11167  ( .D(I192545), .CLK(I2702), .RSTB(I191960), .Q(I191937) );
DFFARX1 I_11168  ( .D(I192480), .CLK(I2702), .RSTB(I191960), .Q(I191922) );
not I_11169 (I192623,I2709);
not I_11170 (I192640,I256896);
nor I_11171 (I192657,I256905,I256917);
nand I_11172 (I192674,I192657,I256908);
DFFARX1 I_11173  ( .D(I192674), .CLK(I2702), .RSTB(I192623), .Q(I192594) );
nor I_11174 (I192705,I192640,I256905);
nand I_11175 (I192722,I192705,I256920);
nand I_11176 (I192739,I192722,I192674);
not I_11177 (I192756,I256905);
not I_11178 (I192773,I256926);
nor I_11179 (I192790,I192773,I256902);
and I_11180 (I192807,I192790,I256911);
or I_11181 (I192824,I192807,I256899);
DFFARX1 I_11182  ( .D(I192824), .CLK(I2702), .RSTB(I192623), .Q(I192841) );
nor I_11183 (I192858,I192841,I192722);
nand I_11184 (I192609,I192756,I192858);
not I_11185 (I192606,I192841);
and I_11186 (I192903,I192841,I192739);
DFFARX1 I_11187  ( .D(I192903), .CLK(I2702), .RSTB(I192623), .Q(I192591) );
DFFARX1 I_11188  ( .D(I192841), .CLK(I2702), .RSTB(I192623), .Q(I192934) );
and I_11189 (I192588,I192756,I192934);
nand I_11190 (I192965,I192640,I256926);
not I_11191 (I192982,I192965);
nor I_11192 (I192999,I192841,I192982);
DFFARX1 I_11193  ( .D(I256923), .CLK(I2702), .RSTB(I192623), .Q(I193016) );
nand I_11194 (I193033,I193016,I192965);
and I_11195 (I193050,I192756,I193033);
DFFARX1 I_11196  ( .D(I193050), .CLK(I2702), .RSTB(I192623), .Q(I192615) );
not I_11197 (I193081,I193016);
nand I_11198 (I192603,I193016,I192999);
nand I_11199 (I192597,I193016,I192982);
DFFARX1 I_11200  ( .D(I256914), .CLK(I2702), .RSTB(I192623), .Q(I193126) );
not I_11201 (I193143,I193126);
nor I_11202 (I192612,I193016,I193143);
nor I_11203 (I193174,I193143,I193081);
and I_11204 (I193191,I192722,I193174);
or I_11205 (I193208,I192965,I193191);
DFFARX1 I_11206  ( .D(I193208), .CLK(I2702), .RSTB(I192623), .Q(I192600) );
DFFARX1 I_11207  ( .D(I193143), .CLK(I2702), .RSTB(I192623), .Q(I192585) );
not I_11208 (I193286,I2709);
not I_11209 (I193303,I572074);
nor I_11210 (I193320,I572086,I572089);
nand I_11211 (I193337,I193320,I572077);
DFFARX1 I_11212  ( .D(I193337), .CLK(I2702), .RSTB(I193286), .Q(I193257) );
nor I_11213 (I193368,I193303,I572086);
nand I_11214 (I193385,I193368,I572062);
nand I_11215 (I193402,I193385,I193337);
not I_11216 (I193419,I572086);
not I_11217 (I193436,I572065);
nor I_11218 (I193453,I193436,I572068);
and I_11219 (I193470,I193453,I572071);
or I_11220 (I193487,I193470,I572080);
DFFARX1 I_11221  ( .D(I193487), .CLK(I2702), .RSTB(I193286), .Q(I193504) );
nor I_11222 (I193521,I193504,I193385);
nand I_11223 (I193272,I193419,I193521);
not I_11224 (I193269,I193504);
and I_11225 (I193566,I193504,I193402);
DFFARX1 I_11226  ( .D(I193566), .CLK(I2702), .RSTB(I193286), .Q(I193254) );
DFFARX1 I_11227  ( .D(I193504), .CLK(I2702), .RSTB(I193286), .Q(I193597) );
and I_11228 (I193251,I193419,I193597);
nand I_11229 (I193628,I193303,I572065);
not I_11230 (I193645,I193628);
nor I_11231 (I193662,I193504,I193645);
DFFARX1 I_11232  ( .D(I572083), .CLK(I2702), .RSTB(I193286), .Q(I193679) );
nand I_11233 (I193696,I193679,I193628);
and I_11234 (I193713,I193419,I193696);
DFFARX1 I_11235  ( .D(I193713), .CLK(I2702), .RSTB(I193286), .Q(I193278) );
not I_11236 (I193744,I193679);
nand I_11237 (I193266,I193679,I193662);
nand I_11238 (I193260,I193679,I193645);
DFFARX1 I_11239  ( .D(I572059), .CLK(I2702), .RSTB(I193286), .Q(I193789) );
not I_11240 (I193806,I193789);
nor I_11241 (I193275,I193679,I193806);
nor I_11242 (I193837,I193806,I193744);
and I_11243 (I193854,I193385,I193837);
or I_11244 (I193871,I193628,I193854);
DFFARX1 I_11245  ( .D(I193871), .CLK(I2702), .RSTB(I193286), .Q(I193263) );
DFFARX1 I_11246  ( .D(I193806), .CLK(I2702), .RSTB(I193286), .Q(I193248) );
not I_11247 (I193949,I2709);
not I_11248 (I193966,I385485);
nor I_11249 (I193983,I385494,I385467);
nand I_11250 (I194000,I193983,I385479);
DFFARX1 I_11251  ( .D(I194000), .CLK(I2702), .RSTB(I193949), .Q(I193920) );
nor I_11252 (I194031,I193966,I385494);
nand I_11253 (I194048,I194031,I385491);
nand I_11254 (I194065,I194048,I194000);
not I_11255 (I194082,I385494);
not I_11256 (I194099,I385470);
nor I_11257 (I194116,I194099,I385476);
and I_11258 (I194133,I194116,I385488);
or I_11259 (I194150,I194133,I385473);
DFFARX1 I_11260  ( .D(I194150), .CLK(I2702), .RSTB(I193949), .Q(I194167) );
nor I_11261 (I194184,I194167,I194048);
nand I_11262 (I193935,I194082,I194184);
not I_11263 (I193932,I194167);
and I_11264 (I194229,I194167,I194065);
DFFARX1 I_11265  ( .D(I194229), .CLK(I2702), .RSTB(I193949), .Q(I193917) );
DFFARX1 I_11266  ( .D(I194167), .CLK(I2702), .RSTB(I193949), .Q(I194260) );
and I_11267 (I193914,I194082,I194260);
nand I_11268 (I194291,I193966,I385470);
not I_11269 (I194308,I194291);
nor I_11270 (I194325,I194167,I194308);
DFFARX1 I_11271  ( .D(I385497), .CLK(I2702), .RSTB(I193949), .Q(I194342) );
nand I_11272 (I194359,I194342,I194291);
and I_11273 (I194376,I194082,I194359);
DFFARX1 I_11274  ( .D(I194376), .CLK(I2702), .RSTB(I193949), .Q(I193941) );
not I_11275 (I194407,I194342);
nand I_11276 (I193929,I194342,I194325);
nand I_11277 (I193923,I194342,I194308);
DFFARX1 I_11278  ( .D(I385482), .CLK(I2702), .RSTB(I193949), .Q(I194452) );
not I_11279 (I194469,I194452);
nor I_11280 (I193938,I194342,I194469);
nor I_11281 (I194500,I194469,I194407);
and I_11282 (I194517,I194048,I194500);
or I_11283 (I194534,I194291,I194517);
DFFARX1 I_11284  ( .D(I194534), .CLK(I2702), .RSTB(I193949), .Q(I193926) );
DFFARX1 I_11285  ( .D(I194469), .CLK(I2702), .RSTB(I193949), .Q(I193911) );
not I_11286 (I194612,I2709);
not I_11287 (I194629,I248940);
nor I_11288 (I194646,I248949,I248961);
nand I_11289 (I194663,I194646,I248952);
DFFARX1 I_11290  ( .D(I194663), .CLK(I2702), .RSTB(I194612), .Q(I194583) );
nor I_11291 (I194694,I194629,I248949);
nand I_11292 (I194711,I194694,I248964);
nand I_11293 (I194728,I194711,I194663);
not I_11294 (I194745,I248949);
not I_11295 (I194762,I248970);
nor I_11296 (I194779,I194762,I248946);
and I_11297 (I194796,I194779,I248955);
or I_11298 (I194813,I194796,I248943);
DFFARX1 I_11299  ( .D(I194813), .CLK(I2702), .RSTB(I194612), .Q(I194830) );
nor I_11300 (I194847,I194830,I194711);
nand I_11301 (I194598,I194745,I194847);
not I_11302 (I194595,I194830);
and I_11303 (I194892,I194830,I194728);
DFFARX1 I_11304  ( .D(I194892), .CLK(I2702), .RSTB(I194612), .Q(I194580) );
DFFARX1 I_11305  ( .D(I194830), .CLK(I2702), .RSTB(I194612), .Q(I194923) );
and I_11306 (I194577,I194745,I194923);
nand I_11307 (I194954,I194629,I248970);
not I_11308 (I194971,I194954);
nor I_11309 (I194988,I194830,I194971);
DFFARX1 I_11310  ( .D(I248967), .CLK(I2702), .RSTB(I194612), .Q(I195005) );
nand I_11311 (I195022,I195005,I194954);
and I_11312 (I195039,I194745,I195022);
DFFARX1 I_11313  ( .D(I195039), .CLK(I2702), .RSTB(I194612), .Q(I194604) );
not I_11314 (I195070,I195005);
nand I_11315 (I194592,I195005,I194988);
nand I_11316 (I194586,I195005,I194971);
DFFARX1 I_11317  ( .D(I248958), .CLK(I2702), .RSTB(I194612), .Q(I195115) );
not I_11318 (I195132,I195115);
nor I_11319 (I194601,I195005,I195132);
nor I_11320 (I195163,I195132,I195070);
and I_11321 (I195180,I194711,I195163);
or I_11322 (I195197,I194954,I195180);
DFFARX1 I_11323  ( .D(I195197), .CLK(I2702), .RSTB(I194612), .Q(I194589) );
DFFARX1 I_11324  ( .D(I195132), .CLK(I2702), .RSTB(I194612), .Q(I194574) );
not I_11325 (I195275,I2709);
not I_11326 (I195292,I448877);
nor I_11327 (I195309,I448883,I448880);
nand I_11328 (I195326,I195309,I448898);
DFFARX1 I_11329  ( .D(I195326), .CLK(I2702), .RSTB(I195275), .Q(I195246) );
nor I_11330 (I195357,I195292,I448883);
nand I_11331 (I195374,I195357,I448907);
nand I_11332 (I195391,I195374,I195326);
not I_11333 (I195408,I448883);
not I_11334 (I195425,I448901);
nor I_11335 (I195442,I195425,I448892);
and I_11336 (I195459,I195442,I448895);
or I_11337 (I195476,I195459,I448886);
DFFARX1 I_11338  ( .D(I195476), .CLK(I2702), .RSTB(I195275), .Q(I195493) );
nor I_11339 (I195510,I195493,I195374);
nand I_11340 (I195261,I195408,I195510);
not I_11341 (I195258,I195493);
and I_11342 (I195555,I195493,I195391);
DFFARX1 I_11343  ( .D(I195555), .CLK(I2702), .RSTB(I195275), .Q(I195243) );
DFFARX1 I_11344  ( .D(I195493), .CLK(I2702), .RSTB(I195275), .Q(I195586) );
and I_11345 (I195240,I195408,I195586);
nand I_11346 (I195617,I195292,I448901);
not I_11347 (I195634,I195617);
nor I_11348 (I195651,I195493,I195634);
DFFARX1 I_11349  ( .D(I448904), .CLK(I2702), .RSTB(I195275), .Q(I195668) );
nand I_11350 (I195685,I195668,I195617);
and I_11351 (I195702,I195408,I195685);
DFFARX1 I_11352  ( .D(I195702), .CLK(I2702), .RSTB(I195275), .Q(I195267) );
not I_11353 (I195733,I195668);
nand I_11354 (I195255,I195668,I195651);
nand I_11355 (I195249,I195668,I195634);
DFFARX1 I_11356  ( .D(I448889), .CLK(I2702), .RSTB(I195275), .Q(I195778) );
not I_11357 (I195795,I195778);
nor I_11358 (I195264,I195668,I195795);
nor I_11359 (I195826,I195795,I195733);
and I_11360 (I195843,I195374,I195826);
or I_11361 (I195860,I195617,I195843);
DFFARX1 I_11362  ( .D(I195860), .CLK(I2702), .RSTB(I195275), .Q(I195252) );
DFFARX1 I_11363  ( .D(I195795), .CLK(I2702), .RSTB(I195275), .Q(I195237) );
not I_11364 (I195938,I2709);
not I_11365 (I195955,I532804);
nor I_11366 (I195972,I532816,I532819);
nand I_11367 (I195989,I195972,I532807);
DFFARX1 I_11368  ( .D(I195989), .CLK(I2702), .RSTB(I195938), .Q(I195909) );
nor I_11369 (I196020,I195955,I532816);
nand I_11370 (I196037,I196020,I532792);
nand I_11371 (I196054,I196037,I195989);
not I_11372 (I196071,I532816);
not I_11373 (I196088,I532795);
nor I_11374 (I196105,I196088,I532798);
and I_11375 (I196122,I196105,I532801);
or I_11376 (I196139,I196122,I532810);
DFFARX1 I_11377  ( .D(I196139), .CLK(I2702), .RSTB(I195938), .Q(I196156) );
nor I_11378 (I196173,I196156,I196037);
nand I_11379 (I195924,I196071,I196173);
not I_11380 (I195921,I196156);
and I_11381 (I196218,I196156,I196054);
DFFARX1 I_11382  ( .D(I196218), .CLK(I2702), .RSTB(I195938), .Q(I195906) );
DFFARX1 I_11383  ( .D(I196156), .CLK(I2702), .RSTB(I195938), .Q(I196249) );
and I_11384 (I195903,I196071,I196249);
nand I_11385 (I196280,I195955,I532795);
not I_11386 (I196297,I196280);
nor I_11387 (I196314,I196156,I196297);
DFFARX1 I_11388  ( .D(I532813), .CLK(I2702), .RSTB(I195938), .Q(I196331) );
nand I_11389 (I196348,I196331,I196280);
and I_11390 (I196365,I196071,I196348);
DFFARX1 I_11391  ( .D(I196365), .CLK(I2702), .RSTB(I195938), .Q(I195930) );
not I_11392 (I196396,I196331);
nand I_11393 (I195918,I196331,I196314);
nand I_11394 (I195912,I196331,I196297);
DFFARX1 I_11395  ( .D(I532789), .CLK(I2702), .RSTB(I195938), .Q(I196441) );
not I_11396 (I196458,I196441);
nor I_11397 (I195927,I196331,I196458);
nor I_11398 (I196489,I196458,I196396);
and I_11399 (I196506,I196037,I196489);
or I_11400 (I196523,I196280,I196506);
DFFARX1 I_11401  ( .D(I196523), .CLK(I2702), .RSTB(I195938), .Q(I195915) );
DFFARX1 I_11402  ( .D(I196458), .CLK(I2702), .RSTB(I195938), .Q(I195900) );
not I_11403 (I196601,I2709);
not I_11404 (I196618,I320544);
nor I_11405 (I196635,I320553,I320565);
nand I_11406 (I196652,I196635,I320556);
DFFARX1 I_11407  ( .D(I196652), .CLK(I2702), .RSTB(I196601), .Q(I196572) );
nor I_11408 (I196683,I196618,I320553);
nand I_11409 (I196700,I196683,I320568);
nand I_11410 (I196717,I196700,I196652);
not I_11411 (I196734,I320553);
not I_11412 (I196751,I320574);
nor I_11413 (I196768,I196751,I320550);
and I_11414 (I196785,I196768,I320559);
or I_11415 (I196802,I196785,I320547);
DFFARX1 I_11416  ( .D(I196802), .CLK(I2702), .RSTB(I196601), .Q(I196819) );
nor I_11417 (I196836,I196819,I196700);
nand I_11418 (I196587,I196734,I196836);
not I_11419 (I196584,I196819);
and I_11420 (I196881,I196819,I196717);
DFFARX1 I_11421  ( .D(I196881), .CLK(I2702), .RSTB(I196601), .Q(I196569) );
DFFARX1 I_11422  ( .D(I196819), .CLK(I2702), .RSTB(I196601), .Q(I196912) );
and I_11423 (I196566,I196734,I196912);
nand I_11424 (I196943,I196618,I320574);
not I_11425 (I196960,I196943);
nor I_11426 (I196977,I196819,I196960);
DFFARX1 I_11427  ( .D(I320571), .CLK(I2702), .RSTB(I196601), .Q(I196994) );
nand I_11428 (I197011,I196994,I196943);
and I_11429 (I197028,I196734,I197011);
DFFARX1 I_11430  ( .D(I197028), .CLK(I2702), .RSTB(I196601), .Q(I196593) );
not I_11431 (I197059,I196994);
nand I_11432 (I196581,I196994,I196977);
nand I_11433 (I196575,I196994,I196960);
DFFARX1 I_11434  ( .D(I320562), .CLK(I2702), .RSTB(I196601), .Q(I197104) );
not I_11435 (I197121,I197104);
nor I_11436 (I196590,I196994,I197121);
nor I_11437 (I197152,I197121,I197059);
and I_11438 (I197169,I196700,I197152);
or I_11439 (I197186,I196943,I197169);
DFFARX1 I_11440  ( .D(I197186), .CLK(I2702), .RSTB(I196601), .Q(I196578) );
DFFARX1 I_11441  ( .D(I197121), .CLK(I2702), .RSTB(I196601), .Q(I196563) );
not I_11442 (I197264,I2709);
not I_11443 (I197281,I576825);
nor I_11444 (I197298,I576840,I576822);
nand I_11445 (I197315,I197298,I576834);
DFFARX1 I_11446  ( .D(I197315), .CLK(I2702), .RSTB(I197264), .Q(I197235) );
nor I_11447 (I197346,I197281,I576840);
nand I_11448 (I197363,I197346,I576831);
nand I_11449 (I197380,I197363,I197315);
not I_11450 (I197397,I576840);
not I_11451 (I197414,I576849);
nor I_11452 (I197431,I197414,I576819);
and I_11453 (I197448,I197431,I576828);
or I_11454 (I197465,I197448,I576846);
DFFARX1 I_11455  ( .D(I197465), .CLK(I2702), .RSTB(I197264), .Q(I197482) );
nor I_11456 (I197499,I197482,I197363);
nand I_11457 (I197250,I197397,I197499);
not I_11458 (I197247,I197482);
and I_11459 (I197544,I197482,I197380);
DFFARX1 I_11460  ( .D(I197544), .CLK(I2702), .RSTB(I197264), .Q(I197232) );
DFFARX1 I_11461  ( .D(I197482), .CLK(I2702), .RSTB(I197264), .Q(I197575) );
and I_11462 (I197229,I197397,I197575);
nand I_11463 (I197606,I197281,I576849);
not I_11464 (I197623,I197606);
nor I_11465 (I197640,I197482,I197623);
DFFARX1 I_11466  ( .D(I576837), .CLK(I2702), .RSTB(I197264), .Q(I197657) );
nand I_11467 (I197674,I197657,I197606);
and I_11468 (I197691,I197397,I197674);
DFFARX1 I_11469  ( .D(I197691), .CLK(I2702), .RSTB(I197264), .Q(I197256) );
not I_11470 (I197722,I197657);
nand I_11471 (I197244,I197657,I197640);
nand I_11472 (I197238,I197657,I197623);
DFFARX1 I_11473  ( .D(I576843), .CLK(I2702), .RSTB(I197264), .Q(I197767) );
not I_11474 (I197784,I197767);
nor I_11475 (I197253,I197657,I197784);
nor I_11476 (I197815,I197784,I197722);
and I_11477 (I197832,I197363,I197815);
or I_11478 (I197849,I197606,I197832);
DFFARX1 I_11479  ( .D(I197849), .CLK(I2702), .RSTB(I197264), .Q(I197241) );
DFFARX1 I_11480  ( .D(I197784), .CLK(I2702), .RSTB(I197264), .Q(I197226) );
not I_11481 (I197927,I2709);
not I_11482 (I197944,I53642);
nor I_11483 (I197961,I53630,I53654);
nand I_11484 (I197978,I197961,I53639);
DFFARX1 I_11485  ( .D(I197978), .CLK(I2702), .RSTB(I197927), .Q(I197898) );
nor I_11486 (I198009,I197944,I53630);
nand I_11487 (I198026,I198009,I53657);
nand I_11488 (I198043,I198026,I197978);
not I_11489 (I198060,I53630);
not I_11490 (I198077,I53627);
nor I_11491 (I198094,I198077,I53636);
and I_11492 (I198111,I198094,I53651);
or I_11493 (I198128,I198111,I53633);
DFFARX1 I_11494  ( .D(I198128), .CLK(I2702), .RSTB(I197927), .Q(I198145) );
nor I_11495 (I198162,I198145,I198026);
nand I_11496 (I197913,I198060,I198162);
not I_11497 (I197910,I198145);
and I_11498 (I198207,I198145,I198043);
DFFARX1 I_11499  ( .D(I198207), .CLK(I2702), .RSTB(I197927), .Q(I197895) );
DFFARX1 I_11500  ( .D(I198145), .CLK(I2702), .RSTB(I197927), .Q(I198238) );
and I_11501 (I197892,I198060,I198238);
nand I_11502 (I198269,I197944,I53627);
not I_11503 (I198286,I198269);
nor I_11504 (I198303,I198145,I198286);
DFFARX1 I_11505  ( .D(I53648), .CLK(I2702), .RSTB(I197927), .Q(I198320) );
nand I_11506 (I198337,I198320,I198269);
and I_11507 (I198354,I198060,I198337);
DFFARX1 I_11508  ( .D(I198354), .CLK(I2702), .RSTB(I197927), .Q(I197919) );
not I_11509 (I198385,I198320);
nand I_11510 (I197907,I198320,I198303);
nand I_11511 (I197901,I198320,I198286);
DFFARX1 I_11512  ( .D(I53645), .CLK(I2702), .RSTB(I197927), .Q(I198430) );
not I_11513 (I198447,I198430);
nor I_11514 (I197916,I198320,I198447);
nor I_11515 (I198478,I198447,I198385);
and I_11516 (I198495,I198026,I198478);
or I_11517 (I198512,I198269,I198495);
DFFARX1 I_11518  ( .D(I198512), .CLK(I2702), .RSTB(I197927), .Q(I197904) );
DFFARX1 I_11519  ( .D(I198447), .CLK(I2702), .RSTB(I197927), .Q(I197889) );
not I_11520 (I198590,I2709);
not I_11521 (I198607,I716396);
nor I_11522 (I198624,I716375,I716387);
nand I_11523 (I198641,I198624,I716381);
DFFARX1 I_11524  ( .D(I198641), .CLK(I2702), .RSTB(I198590), .Q(I198561) );
nor I_11525 (I198672,I198607,I716375);
nand I_11526 (I198689,I198672,I716402);
nand I_11527 (I198706,I198689,I198641);
not I_11528 (I198723,I716375);
not I_11529 (I198740,I716378);
nor I_11530 (I198757,I198740,I716390);
and I_11531 (I198774,I198757,I716393);
or I_11532 (I198791,I198774,I716399);
DFFARX1 I_11533  ( .D(I198791), .CLK(I2702), .RSTB(I198590), .Q(I198808) );
nor I_11534 (I198825,I198808,I198689);
nand I_11535 (I198576,I198723,I198825);
not I_11536 (I198573,I198808);
and I_11537 (I198870,I198808,I198706);
DFFARX1 I_11538  ( .D(I198870), .CLK(I2702), .RSTB(I198590), .Q(I198558) );
DFFARX1 I_11539  ( .D(I198808), .CLK(I2702), .RSTB(I198590), .Q(I198901) );
and I_11540 (I198555,I198723,I198901);
nand I_11541 (I198932,I198607,I716378);
not I_11542 (I198949,I198932);
nor I_11543 (I198966,I198808,I198949);
DFFARX1 I_11544  ( .D(I716372), .CLK(I2702), .RSTB(I198590), .Q(I198983) );
nand I_11545 (I199000,I198983,I198932);
and I_11546 (I199017,I198723,I199000);
DFFARX1 I_11547  ( .D(I199017), .CLK(I2702), .RSTB(I198590), .Q(I198582) );
not I_11548 (I199048,I198983);
nand I_11549 (I198570,I198983,I198966);
nand I_11550 (I198564,I198983,I198949);
DFFARX1 I_11551  ( .D(I716384), .CLK(I2702), .RSTB(I198590), .Q(I199093) );
not I_11552 (I199110,I199093);
nor I_11553 (I198579,I198983,I199110);
nor I_11554 (I199141,I199110,I199048);
and I_11555 (I199158,I198689,I199141);
or I_11556 (I199175,I198932,I199158);
DFFARX1 I_11557  ( .D(I199175), .CLK(I2702), .RSTB(I198590), .Q(I198567) );
DFFARX1 I_11558  ( .D(I199110), .CLK(I2702), .RSTB(I198590), .Q(I198552) );
not I_11559 (I199253,I2709);
not I_11560 (I199270,I439051);
nor I_11561 (I199287,I439057,I439054);
nand I_11562 (I199304,I199287,I439072);
DFFARX1 I_11563  ( .D(I199304), .CLK(I2702), .RSTB(I199253), .Q(I199224) );
nor I_11564 (I199335,I199270,I439057);
nand I_11565 (I199352,I199335,I439081);
nand I_11566 (I199369,I199352,I199304);
not I_11567 (I199386,I439057);
not I_11568 (I199403,I439075);
nor I_11569 (I199420,I199403,I439066);
and I_11570 (I199437,I199420,I439069);
or I_11571 (I199454,I199437,I439060);
DFFARX1 I_11572  ( .D(I199454), .CLK(I2702), .RSTB(I199253), .Q(I199471) );
nor I_11573 (I199488,I199471,I199352);
nand I_11574 (I199239,I199386,I199488);
not I_11575 (I199236,I199471);
and I_11576 (I199533,I199471,I199369);
DFFARX1 I_11577  ( .D(I199533), .CLK(I2702), .RSTB(I199253), .Q(I199221) );
DFFARX1 I_11578  ( .D(I199471), .CLK(I2702), .RSTB(I199253), .Q(I199564) );
and I_11579 (I199218,I199386,I199564);
nand I_11580 (I199595,I199270,I439075);
not I_11581 (I199612,I199595);
nor I_11582 (I199629,I199471,I199612);
DFFARX1 I_11583  ( .D(I439078), .CLK(I2702), .RSTB(I199253), .Q(I199646) );
nand I_11584 (I199663,I199646,I199595);
and I_11585 (I199680,I199386,I199663);
DFFARX1 I_11586  ( .D(I199680), .CLK(I2702), .RSTB(I199253), .Q(I199245) );
not I_11587 (I199711,I199646);
nand I_11588 (I199233,I199646,I199629);
nand I_11589 (I199227,I199646,I199612);
DFFARX1 I_11590  ( .D(I439063), .CLK(I2702), .RSTB(I199253), .Q(I199756) );
not I_11591 (I199773,I199756);
nor I_11592 (I199242,I199646,I199773);
nor I_11593 (I199804,I199773,I199711);
and I_11594 (I199821,I199352,I199804);
or I_11595 (I199838,I199595,I199821);
DFFARX1 I_11596  ( .D(I199838), .CLK(I2702), .RSTB(I199253), .Q(I199230) );
DFFARX1 I_11597  ( .D(I199773), .CLK(I2702), .RSTB(I199253), .Q(I199215) );
not I_11598 (I199916,I2709);
or I_11599 (I199933,I63984,I63978);
or I_11600 (I199950,I63972,I63984);
DFFARX1 I_11601  ( .D(I199950), .CLK(I2702), .RSTB(I199916), .Q(I199890) );
nor I_11602 (I199981,I63990,I63981);
not I_11603 (I199998,I199981);
not I_11604 (I200015,I63990);
and I_11605 (I200032,I200015,I63987);
nor I_11606 (I200049,I200032,I63978);
nor I_11607 (I200066,I63963,I63969);
DFFARX1 I_11608  ( .D(I200066), .CLK(I2702), .RSTB(I199916), .Q(I200083) );
nand I_11609 (I200100,I200083,I199933);
and I_11610 (I200117,I200049,I200100);
DFFARX1 I_11611  ( .D(I200117), .CLK(I2702), .RSTB(I199916), .Q(I199884) );
nor I_11612 (I200148,I63963,I63972);
DFFARX1 I_11613  ( .D(I200148), .CLK(I2702), .RSTB(I199916), .Q(I200165) );
and I_11614 (I199881,I199981,I200165);
DFFARX1 I_11615  ( .D(I63975), .CLK(I2702), .RSTB(I199916), .Q(I200196) );
and I_11616 (I200213,I200196,I63993);
DFFARX1 I_11617  ( .D(I200213), .CLK(I2702), .RSTB(I199916), .Q(I200230) );
not I_11618 (I199893,I200230);
DFFARX1 I_11619  ( .D(I200213), .CLK(I2702), .RSTB(I199916), .Q(I199878) );
DFFARX1 I_11620  ( .D(I63966), .CLK(I2702), .RSTB(I199916), .Q(I200275) );
not I_11621 (I200292,I200275);
nor I_11622 (I200309,I199950,I200292);
and I_11623 (I200326,I200213,I200309);
or I_11624 (I200343,I199933,I200326);
DFFARX1 I_11625  ( .D(I200343), .CLK(I2702), .RSTB(I199916), .Q(I199899) );
nor I_11626 (I200374,I200275,I200083);
nand I_11627 (I199908,I200049,I200374);
nor I_11628 (I200405,I200275,I199998);
nand I_11629 (I199902,I200148,I200405);
not I_11630 (I199905,I200275);
nand I_11631 (I199896,I200275,I199998);
DFFARX1 I_11632  ( .D(I200275), .CLK(I2702), .RSTB(I199916), .Q(I199887) );
not I_11633 (I200511,I2709);
or I_11634 (I200528,I478963,I478948);
or I_11635 (I200545,I478960,I478963);
DFFARX1 I_11636  ( .D(I200545), .CLK(I2702), .RSTB(I200511), .Q(I200485) );
nor I_11637 (I200576,I478942,I478933);
not I_11638 (I200593,I200576);
not I_11639 (I200610,I478942);
and I_11640 (I200627,I200610,I478957);
nor I_11641 (I200644,I200627,I478948);
nor I_11642 (I200661,I478936,I478954);
DFFARX1 I_11643  ( .D(I200661), .CLK(I2702), .RSTB(I200511), .Q(I200678) );
nand I_11644 (I200695,I200678,I200528);
and I_11645 (I200712,I200644,I200695);
DFFARX1 I_11646  ( .D(I200712), .CLK(I2702), .RSTB(I200511), .Q(I200479) );
nor I_11647 (I200743,I478936,I478960);
DFFARX1 I_11648  ( .D(I200743), .CLK(I2702), .RSTB(I200511), .Q(I200760) );
and I_11649 (I200476,I200576,I200760);
DFFARX1 I_11650  ( .D(I478945), .CLK(I2702), .RSTB(I200511), .Q(I200791) );
and I_11651 (I200808,I200791,I478939);
DFFARX1 I_11652  ( .D(I200808), .CLK(I2702), .RSTB(I200511), .Q(I200825) );
not I_11653 (I200488,I200825);
DFFARX1 I_11654  ( .D(I200808), .CLK(I2702), .RSTB(I200511), .Q(I200473) );
DFFARX1 I_11655  ( .D(I478951), .CLK(I2702), .RSTB(I200511), .Q(I200870) );
not I_11656 (I200887,I200870);
nor I_11657 (I200904,I200545,I200887);
and I_11658 (I200921,I200808,I200904);
or I_11659 (I200938,I200528,I200921);
DFFARX1 I_11660  ( .D(I200938), .CLK(I2702), .RSTB(I200511), .Q(I200494) );
nor I_11661 (I200969,I200870,I200678);
nand I_11662 (I200503,I200644,I200969);
nor I_11663 (I201000,I200870,I200593);
nand I_11664 (I200497,I200743,I201000);
not I_11665 (I200500,I200870);
nand I_11666 (I200491,I200870,I200593);
DFFARX1 I_11667  ( .D(I200870), .CLK(I2702), .RSTB(I200511), .Q(I200482) );
not I_11668 (I201106,I2709);
or I_11669 (I201123,I344787,I344784);
or I_11670 (I201140,I344769,I344787);
DFFARX1 I_11671  ( .D(I201140), .CLK(I2702), .RSTB(I201106), .Q(I201080) );
nor I_11672 (I201171,I344778,I344781);
not I_11673 (I201188,I201171);
not I_11674 (I201205,I344778);
and I_11675 (I201222,I201205,I344793);
nor I_11676 (I201239,I201222,I344784);
nor I_11677 (I201256,I344799,I344775);
DFFARX1 I_11678  ( .D(I201256), .CLK(I2702), .RSTB(I201106), .Q(I201273) );
nand I_11679 (I201290,I201273,I201123);
and I_11680 (I201307,I201239,I201290);
DFFARX1 I_11681  ( .D(I201307), .CLK(I2702), .RSTB(I201106), .Q(I201074) );
nor I_11682 (I201338,I344799,I344769);
DFFARX1 I_11683  ( .D(I201338), .CLK(I2702), .RSTB(I201106), .Q(I201355) );
and I_11684 (I201071,I201171,I201355);
DFFARX1 I_11685  ( .D(I344790), .CLK(I2702), .RSTB(I201106), .Q(I201386) );
and I_11686 (I201403,I201386,I344796);
DFFARX1 I_11687  ( .D(I201403), .CLK(I2702), .RSTB(I201106), .Q(I201420) );
not I_11688 (I201083,I201420);
DFFARX1 I_11689  ( .D(I201403), .CLK(I2702), .RSTB(I201106), .Q(I201068) );
DFFARX1 I_11690  ( .D(I344772), .CLK(I2702), .RSTB(I201106), .Q(I201465) );
not I_11691 (I201482,I201465);
nor I_11692 (I201499,I201140,I201482);
and I_11693 (I201516,I201403,I201499);
or I_11694 (I201533,I201123,I201516);
DFFARX1 I_11695  ( .D(I201533), .CLK(I2702), .RSTB(I201106), .Q(I201089) );
nor I_11696 (I201564,I201465,I201273);
nand I_11697 (I201098,I201239,I201564);
nor I_11698 (I201595,I201465,I201188);
nand I_11699 (I201092,I201338,I201595);
not I_11700 (I201095,I201465);
nand I_11701 (I201086,I201465,I201188);
DFFARX1 I_11702  ( .D(I201465), .CLK(I2702), .RSTB(I201106), .Q(I201077) );
not I_11703 (I201701,I2709);
or I_11704 (I201718,I594086,I594080);
or I_11705 (I201735,I594074,I594086);
DFFARX1 I_11706  ( .D(I201735), .CLK(I2702), .RSTB(I201701), .Q(I201675) );
nor I_11707 (I201766,I594077,I594083);
not I_11708 (I201783,I201766);
not I_11709 (I201800,I594077);
and I_11710 (I201817,I201800,I594101);
nor I_11711 (I201834,I201817,I594080);
nor I_11712 (I201851,I594104,I594095);
DFFARX1 I_11713  ( .D(I201851), .CLK(I2702), .RSTB(I201701), .Q(I201868) );
nand I_11714 (I201885,I201868,I201718);
and I_11715 (I201902,I201834,I201885);
DFFARX1 I_11716  ( .D(I201902), .CLK(I2702), .RSTB(I201701), .Q(I201669) );
nor I_11717 (I201933,I594104,I594074);
DFFARX1 I_11718  ( .D(I201933), .CLK(I2702), .RSTB(I201701), .Q(I201950) );
and I_11719 (I201666,I201766,I201950);
DFFARX1 I_11720  ( .D(I594092), .CLK(I2702), .RSTB(I201701), .Q(I201981) );
and I_11721 (I201998,I201981,I594089);
DFFARX1 I_11722  ( .D(I201998), .CLK(I2702), .RSTB(I201701), .Q(I202015) );
not I_11723 (I201678,I202015);
DFFARX1 I_11724  ( .D(I201998), .CLK(I2702), .RSTB(I201701), .Q(I201663) );
DFFARX1 I_11725  ( .D(I594098), .CLK(I2702), .RSTB(I201701), .Q(I202060) );
not I_11726 (I202077,I202060);
nor I_11727 (I202094,I201735,I202077);
and I_11728 (I202111,I201998,I202094);
or I_11729 (I202128,I201718,I202111);
DFFARX1 I_11730  ( .D(I202128), .CLK(I2702), .RSTB(I201701), .Q(I201684) );
nor I_11731 (I202159,I202060,I201868);
nand I_11732 (I201693,I201834,I202159);
nor I_11733 (I202190,I202060,I201783);
nand I_11734 (I201687,I201933,I202190);
not I_11735 (I201690,I202060);
nand I_11736 (I201681,I202060,I201783);
DFFARX1 I_11737  ( .D(I202060), .CLK(I2702), .RSTB(I201701), .Q(I201672) );
not I_11738 (I202296,I2709);
or I_11739 (I202313,I427268,I427253);
or I_11740 (I202330,I427262,I427268);
DFFARX1 I_11741  ( .D(I202330), .CLK(I2702), .RSTB(I202296), .Q(I202270) );
nor I_11742 (I202361,I427274,I427283);
not I_11743 (I202378,I202361);
not I_11744 (I202395,I427274);
and I_11745 (I202412,I202395,I427271);
nor I_11746 (I202429,I202412,I427253);
nor I_11747 (I202446,I427280,I427256);
DFFARX1 I_11748  ( .D(I202446), .CLK(I2702), .RSTB(I202296), .Q(I202463) );
nand I_11749 (I202480,I202463,I202313);
and I_11750 (I202497,I202429,I202480);
DFFARX1 I_11751  ( .D(I202497), .CLK(I2702), .RSTB(I202296), .Q(I202264) );
nor I_11752 (I202528,I427280,I427262);
DFFARX1 I_11753  ( .D(I202528), .CLK(I2702), .RSTB(I202296), .Q(I202545) );
and I_11754 (I202261,I202361,I202545);
DFFARX1 I_11755  ( .D(I427265), .CLK(I2702), .RSTB(I202296), .Q(I202576) );
and I_11756 (I202593,I202576,I427259);
DFFARX1 I_11757  ( .D(I202593), .CLK(I2702), .RSTB(I202296), .Q(I202610) );
not I_11758 (I202273,I202610);
DFFARX1 I_11759  ( .D(I202593), .CLK(I2702), .RSTB(I202296), .Q(I202258) );
DFFARX1 I_11760  ( .D(I427277), .CLK(I2702), .RSTB(I202296), .Q(I202655) );
not I_11761 (I202672,I202655);
nor I_11762 (I202689,I202330,I202672);
and I_11763 (I202706,I202593,I202689);
or I_11764 (I202723,I202313,I202706);
DFFARX1 I_11765  ( .D(I202723), .CLK(I2702), .RSTB(I202296), .Q(I202279) );
nor I_11766 (I202754,I202655,I202463);
nand I_11767 (I202288,I202429,I202754);
nor I_11768 (I202785,I202655,I202378);
nand I_11769 (I202282,I202528,I202785);
not I_11770 (I202285,I202655);
nand I_11771 (I202276,I202655,I202378);
DFFARX1 I_11772  ( .D(I202655), .CLK(I2702), .RSTB(I202296), .Q(I202267) );
not I_11773 (I202891,I2709);
or I_11774 (I202908,I1271,I2495);
or I_11775 (I202925,I1319,I1271);
DFFARX1 I_11776  ( .D(I202925), .CLK(I2702), .RSTB(I202891), .Q(I202865) );
nor I_11777 (I202956,I1695,I1455);
not I_11778 (I202973,I202956);
not I_11779 (I202990,I1695);
and I_11780 (I203007,I202990,I2679);
nor I_11781 (I203024,I203007,I2495);
nor I_11782 (I203041,I2391,I1247);
DFFARX1 I_11783  ( .D(I203041), .CLK(I2702), .RSTB(I202891), .Q(I203058) );
nand I_11784 (I203075,I203058,I202908);
and I_11785 (I203092,I203024,I203075);
DFFARX1 I_11786  ( .D(I203092), .CLK(I2702), .RSTB(I202891), .Q(I202859) );
nor I_11787 (I203123,I2391,I1319);
DFFARX1 I_11788  ( .D(I203123), .CLK(I2702), .RSTB(I202891), .Q(I203140) );
and I_11789 (I202856,I202956,I203140);
DFFARX1 I_11790  ( .D(I1687), .CLK(I2702), .RSTB(I202891), .Q(I203171) );
and I_11791 (I203188,I203171,I1999);
DFFARX1 I_11792  ( .D(I203188), .CLK(I2702), .RSTB(I202891), .Q(I203205) );
not I_11793 (I202868,I203205);
DFFARX1 I_11794  ( .D(I203188), .CLK(I2702), .RSTB(I202891), .Q(I202853) );
DFFARX1 I_11795  ( .D(I1895), .CLK(I2702), .RSTB(I202891), .Q(I203250) );
not I_11796 (I203267,I203250);
nor I_11797 (I203284,I202925,I203267);
and I_11798 (I203301,I203188,I203284);
or I_11799 (I203318,I202908,I203301);
DFFARX1 I_11800  ( .D(I203318), .CLK(I2702), .RSTB(I202891), .Q(I202874) );
nor I_11801 (I203349,I203250,I203058);
nand I_11802 (I202883,I203024,I203349);
nor I_11803 (I203380,I203250,I202973);
nand I_11804 (I202877,I203123,I203380);
not I_11805 (I202880,I203250);
nand I_11806 (I202871,I203250,I202973);
DFFARX1 I_11807  ( .D(I203250), .CLK(I2702), .RSTB(I202891), .Q(I202862) );
not I_11808 (I203486,I2709);
or I_11809 (I203503,I99514,I99508);
or I_11810 (I203520,I99502,I99514);
DFFARX1 I_11811  ( .D(I203520), .CLK(I2702), .RSTB(I203486), .Q(I203460) );
nor I_11812 (I203551,I99520,I99511);
not I_11813 (I203568,I203551);
not I_11814 (I203585,I99520);
and I_11815 (I203602,I203585,I99517);
nor I_11816 (I203619,I203602,I99508);
nor I_11817 (I203636,I99493,I99499);
DFFARX1 I_11818  ( .D(I203636), .CLK(I2702), .RSTB(I203486), .Q(I203653) );
nand I_11819 (I203670,I203653,I203503);
and I_11820 (I203687,I203619,I203670);
DFFARX1 I_11821  ( .D(I203687), .CLK(I2702), .RSTB(I203486), .Q(I203454) );
nor I_11822 (I203718,I99493,I99502);
DFFARX1 I_11823  ( .D(I203718), .CLK(I2702), .RSTB(I203486), .Q(I203735) );
and I_11824 (I203451,I203551,I203735);
DFFARX1 I_11825  ( .D(I99505), .CLK(I2702), .RSTB(I203486), .Q(I203766) );
and I_11826 (I203783,I203766,I99523);
DFFARX1 I_11827  ( .D(I203783), .CLK(I2702), .RSTB(I203486), .Q(I203800) );
not I_11828 (I203463,I203800);
DFFARX1 I_11829  ( .D(I203783), .CLK(I2702), .RSTB(I203486), .Q(I203448) );
DFFARX1 I_11830  ( .D(I99496), .CLK(I2702), .RSTB(I203486), .Q(I203845) );
not I_11831 (I203862,I203845);
nor I_11832 (I203879,I203520,I203862);
and I_11833 (I203896,I203783,I203879);
or I_11834 (I203913,I203503,I203896);
DFFARX1 I_11835  ( .D(I203913), .CLK(I2702), .RSTB(I203486), .Q(I203469) );
nor I_11836 (I203944,I203845,I203653);
nand I_11837 (I203478,I203619,I203944);
nor I_11838 (I203975,I203845,I203568);
nand I_11839 (I203472,I203718,I203975);
not I_11840 (I203475,I203845);
nand I_11841 (I203466,I203845,I203568);
DFFARX1 I_11842  ( .D(I203845), .CLK(I2702), .RSTB(I203486), .Q(I203457) );
not I_11843 (I204081,I2709);
or I_11844 (I204098,I40320,I40329);
or I_11845 (I204115,I40323,I40320);
DFFARX1 I_11846  ( .D(I204115), .CLK(I2702), .RSTB(I204081), .Q(I204055) );
nor I_11847 (I204146,I40299,I40302);
not I_11848 (I204163,I204146);
not I_11849 (I204180,I40299);
and I_11850 (I204197,I204180,I40311);
nor I_11851 (I204214,I204197,I40329);
nor I_11852 (I204231,I40317,I40308);
DFFARX1 I_11853  ( .D(I204231), .CLK(I2702), .RSTB(I204081), .Q(I204248) );
nand I_11854 (I204265,I204248,I204098);
and I_11855 (I204282,I204214,I204265);
DFFARX1 I_11856  ( .D(I204282), .CLK(I2702), .RSTB(I204081), .Q(I204049) );
nor I_11857 (I204313,I40317,I40323);
DFFARX1 I_11858  ( .D(I204313), .CLK(I2702), .RSTB(I204081), .Q(I204330) );
and I_11859 (I204046,I204146,I204330);
DFFARX1 I_11860  ( .D(I40314), .CLK(I2702), .RSTB(I204081), .Q(I204361) );
and I_11861 (I204378,I204361,I40305);
DFFARX1 I_11862  ( .D(I204378), .CLK(I2702), .RSTB(I204081), .Q(I204395) );
not I_11863 (I204058,I204395);
DFFARX1 I_11864  ( .D(I204378), .CLK(I2702), .RSTB(I204081), .Q(I204043) );
DFFARX1 I_11865  ( .D(I40326), .CLK(I2702), .RSTB(I204081), .Q(I204440) );
not I_11866 (I204457,I204440);
nor I_11867 (I204474,I204115,I204457);
and I_11868 (I204491,I204378,I204474);
or I_11869 (I204508,I204098,I204491);
DFFARX1 I_11870  ( .D(I204508), .CLK(I2702), .RSTB(I204081), .Q(I204064) );
nor I_11871 (I204539,I204440,I204248);
nand I_11872 (I204073,I204214,I204539);
nor I_11873 (I204570,I204440,I204163);
nand I_11874 (I204067,I204313,I204570);
not I_11875 (I204070,I204440);
nand I_11876 (I204061,I204440,I204163);
DFFARX1 I_11877  ( .D(I204440), .CLK(I2702), .RSTB(I204081), .Q(I204052) );
not I_11878 (I204676,I2709);
or I_11879 (I204693,I77550,I77544);
or I_11880 (I204710,I77538,I77550);
DFFARX1 I_11881  ( .D(I204710), .CLK(I2702), .RSTB(I204676), .Q(I204650) );
nor I_11882 (I204741,I77556,I77547);
not I_11883 (I204758,I204741);
not I_11884 (I204775,I77556);
and I_11885 (I204792,I204775,I77553);
nor I_11886 (I204809,I204792,I77544);
nor I_11887 (I204826,I77529,I77535);
DFFARX1 I_11888  ( .D(I204826), .CLK(I2702), .RSTB(I204676), .Q(I204843) );
nand I_11889 (I204860,I204843,I204693);
and I_11890 (I204877,I204809,I204860);
DFFARX1 I_11891  ( .D(I204877), .CLK(I2702), .RSTB(I204676), .Q(I204644) );
nor I_11892 (I204908,I77529,I77538);
DFFARX1 I_11893  ( .D(I204908), .CLK(I2702), .RSTB(I204676), .Q(I204925) );
and I_11894 (I204641,I204741,I204925);
DFFARX1 I_11895  ( .D(I77541), .CLK(I2702), .RSTB(I204676), .Q(I204956) );
and I_11896 (I204973,I204956,I77559);
DFFARX1 I_11897  ( .D(I204973), .CLK(I2702), .RSTB(I204676), .Q(I204990) );
not I_11898 (I204653,I204990);
DFFARX1 I_11899  ( .D(I204973), .CLK(I2702), .RSTB(I204676), .Q(I204638) );
DFFARX1 I_11900  ( .D(I77532), .CLK(I2702), .RSTB(I204676), .Q(I205035) );
not I_11901 (I205052,I205035);
nor I_11902 (I205069,I204710,I205052);
and I_11903 (I205086,I204973,I205069);
or I_11904 (I205103,I204693,I205086);
DFFARX1 I_11905  ( .D(I205103), .CLK(I2702), .RSTB(I204676), .Q(I204659) );
nor I_11906 (I205134,I205035,I204843);
nand I_11907 (I204668,I204809,I205134);
nor I_11908 (I205165,I205035,I204758);
nand I_11909 (I204662,I204908,I205165);
not I_11910 (I204665,I205035);
nand I_11911 (I204656,I205035,I204758);
DFFARX1 I_11912  ( .D(I205035), .CLK(I2702), .RSTB(I204676), .Q(I204647) );
not I_11913 (I205271,I2709);
or I_11914 (I205288,I266841,I266856);
or I_11915 (I205305,I266844,I266841);
DFFARX1 I_11916  ( .D(I205305), .CLK(I2702), .RSTB(I205271), .Q(I205245) );
nor I_11917 (I205336,I266847,I266862);
not I_11918 (I205353,I205336);
not I_11919 (I205370,I266847);
and I_11920 (I205387,I205370,I266850);
nor I_11921 (I205404,I205387,I266856);
nor I_11922 (I205421,I266853,I266871);
DFFARX1 I_11923  ( .D(I205421), .CLK(I2702), .RSTB(I205271), .Q(I205438) );
nand I_11924 (I205455,I205438,I205288);
and I_11925 (I205472,I205404,I205455);
DFFARX1 I_11926  ( .D(I205472), .CLK(I2702), .RSTB(I205271), .Q(I205239) );
nor I_11927 (I205503,I266853,I266844);
DFFARX1 I_11928  ( .D(I205503), .CLK(I2702), .RSTB(I205271), .Q(I205520) );
and I_11929 (I205236,I205336,I205520);
DFFARX1 I_11930  ( .D(I266868), .CLK(I2702), .RSTB(I205271), .Q(I205551) );
and I_11931 (I205568,I205551,I266859);
DFFARX1 I_11932  ( .D(I205568), .CLK(I2702), .RSTB(I205271), .Q(I205585) );
not I_11933 (I205248,I205585);
DFFARX1 I_11934  ( .D(I205568), .CLK(I2702), .RSTB(I205271), .Q(I205233) );
DFFARX1 I_11935  ( .D(I266865), .CLK(I2702), .RSTB(I205271), .Q(I205630) );
not I_11936 (I205647,I205630);
nor I_11937 (I205664,I205305,I205647);
and I_11938 (I205681,I205568,I205664);
or I_11939 (I205698,I205288,I205681);
DFFARX1 I_11940  ( .D(I205698), .CLK(I2702), .RSTB(I205271), .Q(I205254) );
nor I_11941 (I205729,I205630,I205438);
nand I_11942 (I205263,I205404,I205729);
nor I_11943 (I205760,I205630,I205353);
nand I_11944 (I205257,I205503,I205760);
not I_11945 (I205260,I205630);
nand I_11946 (I205251,I205630,I205353);
DFFARX1 I_11947  ( .D(I205630), .CLK(I2702), .RSTB(I205271), .Q(I205242) );
not I_11948 (I205866,I2709);
or I_11949 (I205883,I325185,I325200);
or I_11950 (I205900,I325188,I325185);
DFFARX1 I_11951  ( .D(I205900), .CLK(I2702), .RSTB(I205866), .Q(I205840) );
nor I_11952 (I205931,I325191,I325206);
not I_11953 (I205948,I205931);
not I_11954 (I205965,I325191);
and I_11955 (I205982,I205965,I325194);
nor I_11956 (I205999,I205982,I325200);
nor I_11957 (I206016,I325197,I325215);
DFFARX1 I_11958  ( .D(I206016), .CLK(I2702), .RSTB(I205866), .Q(I206033) );
nand I_11959 (I206050,I206033,I205883);
and I_11960 (I206067,I205999,I206050);
DFFARX1 I_11961  ( .D(I206067), .CLK(I2702), .RSTB(I205866), .Q(I205834) );
nor I_11962 (I206098,I325197,I325188);
DFFARX1 I_11963  ( .D(I206098), .CLK(I2702), .RSTB(I205866), .Q(I206115) );
and I_11964 (I205831,I205931,I206115);
DFFARX1 I_11965  ( .D(I325212), .CLK(I2702), .RSTB(I205866), .Q(I206146) );
and I_11966 (I206163,I206146,I325203);
DFFARX1 I_11967  ( .D(I206163), .CLK(I2702), .RSTB(I205866), .Q(I206180) );
not I_11968 (I205843,I206180);
DFFARX1 I_11969  ( .D(I206163), .CLK(I2702), .RSTB(I205866), .Q(I205828) );
DFFARX1 I_11970  ( .D(I325209), .CLK(I2702), .RSTB(I205866), .Q(I206225) );
not I_11971 (I206242,I206225);
nor I_11972 (I206259,I205900,I206242);
and I_11973 (I206276,I206163,I206259);
or I_11974 (I206293,I205883,I206276);
DFFARX1 I_11975  ( .D(I206293), .CLK(I2702), .RSTB(I205866), .Q(I205849) );
nor I_11976 (I206324,I206225,I206033);
nand I_11977 (I205858,I205999,I206324);
nor I_11978 (I206355,I206225,I205948);
nand I_11979 (I205852,I206098,I206355);
not I_11980 (I205855,I206225);
nand I_11981 (I205846,I206225,I205948);
DFFARX1 I_11982  ( .D(I206225), .CLK(I2702), .RSTB(I205866), .Q(I205837) );
not I_11983 (I206461,I2709);
or I_11984 (I206478,I230833,I230824);
or I_11985 (I206495,I230845,I230833);
DFFARX1 I_11986  ( .D(I206495), .CLK(I2702), .RSTB(I206461), .Q(I206435) );
nor I_11987 (I206526,I230848,I230827);
not I_11988 (I206543,I206526);
not I_11989 (I206560,I230848);
and I_11990 (I206577,I206560,I230836);
nor I_11991 (I206594,I206577,I230824);
nor I_11992 (I206611,I230821,I230839);
DFFARX1 I_11993  ( .D(I206611), .CLK(I2702), .RSTB(I206461), .Q(I206628) );
nand I_11994 (I206645,I206628,I206478);
and I_11995 (I206662,I206594,I206645);
DFFARX1 I_11996  ( .D(I206662), .CLK(I2702), .RSTB(I206461), .Q(I206429) );
nor I_11997 (I206693,I230821,I230845);
DFFARX1 I_11998  ( .D(I206693), .CLK(I2702), .RSTB(I206461), .Q(I206710) );
and I_11999 (I206426,I206526,I206710);
DFFARX1 I_12000  ( .D(I230842), .CLK(I2702), .RSTB(I206461), .Q(I206741) );
and I_12001 (I206758,I206741,I230818);
DFFARX1 I_12002  ( .D(I206758), .CLK(I2702), .RSTB(I206461), .Q(I206775) );
not I_12003 (I206438,I206775);
DFFARX1 I_12004  ( .D(I206758), .CLK(I2702), .RSTB(I206461), .Q(I206423) );
DFFARX1 I_12005  ( .D(I230830), .CLK(I2702), .RSTB(I206461), .Q(I206820) );
not I_12006 (I206837,I206820);
nor I_12007 (I206854,I206495,I206837);
and I_12008 (I206871,I206758,I206854);
or I_12009 (I206888,I206478,I206871);
DFFARX1 I_12010  ( .D(I206888), .CLK(I2702), .RSTB(I206461), .Q(I206444) );
nor I_12011 (I206919,I206820,I206628);
nand I_12012 (I206453,I206594,I206919);
nor I_12013 (I206950,I206820,I206543);
nand I_12014 (I206447,I206693,I206950);
not I_12015 (I206450,I206820);
nand I_12016 (I206441,I206820,I206543);
DFFARX1 I_12017  ( .D(I206820), .CLK(I2702), .RSTB(I206461), .Q(I206432) );
not I_12018 (I207056,I2709);
or I_12019 (I207073,I345433,I345430);
or I_12020 (I207090,I345415,I345433);
DFFARX1 I_12021  ( .D(I207090), .CLK(I2702), .RSTB(I207056), .Q(I207030) );
nor I_12022 (I207121,I345424,I345427);
not I_12023 (I207138,I207121);
not I_12024 (I207155,I345424);
and I_12025 (I207172,I207155,I345439);
nor I_12026 (I207189,I207172,I345430);
nor I_12027 (I207206,I345445,I345421);
DFFARX1 I_12028  ( .D(I207206), .CLK(I2702), .RSTB(I207056), .Q(I207223) );
nand I_12029 (I207240,I207223,I207073);
and I_12030 (I207257,I207189,I207240);
DFFARX1 I_12031  ( .D(I207257), .CLK(I2702), .RSTB(I207056), .Q(I207024) );
nor I_12032 (I207288,I345445,I345415);
DFFARX1 I_12033  ( .D(I207288), .CLK(I2702), .RSTB(I207056), .Q(I207305) );
and I_12034 (I207021,I207121,I207305);
DFFARX1 I_12035  ( .D(I345436), .CLK(I2702), .RSTB(I207056), .Q(I207336) );
and I_12036 (I207353,I207336,I345442);
DFFARX1 I_12037  ( .D(I207353), .CLK(I2702), .RSTB(I207056), .Q(I207370) );
not I_12038 (I207033,I207370);
DFFARX1 I_12039  ( .D(I207353), .CLK(I2702), .RSTB(I207056), .Q(I207018) );
DFFARX1 I_12040  ( .D(I345418), .CLK(I2702), .RSTB(I207056), .Q(I207415) );
not I_12041 (I207432,I207415);
nor I_12042 (I207449,I207090,I207432);
and I_12043 (I207466,I207353,I207449);
or I_12044 (I207483,I207073,I207466);
DFFARX1 I_12045  ( .D(I207483), .CLK(I2702), .RSTB(I207056), .Q(I207039) );
nor I_12046 (I207514,I207415,I207223);
nand I_12047 (I207048,I207189,I207514);
nor I_12048 (I207545,I207415,I207138);
nand I_12049 (I207042,I207288,I207545);
not I_12050 (I207045,I207415);
nand I_12051 (I207036,I207415,I207138);
DFFARX1 I_12052  ( .D(I207415), .CLK(I2702), .RSTB(I207056), .Q(I207027) );
not I_12053 (I207651,I2709);
or I_12054 (I207668,I546489,I546474);
or I_12055 (I207685,I546495,I546489);
DFFARX1 I_12056  ( .D(I207685), .CLK(I2702), .RSTB(I207651), .Q(I207625) );
nor I_12057 (I207716,I546501,I546483);
not I_12058 (I207733,I207716);
not I_12059 (I207750,I546501);
and I_12060 (I207767,I207750,I546480);
nor I_12061 (I207784,I207767,I546474);
nor I_12062 (I207801,I546477,I546486);
DFFARX1 I_12063  ( .D(I207801), .CLK(I2702), .RSTB(I207651), .Q(I207818) );
nand I_12064 (I207835,I207818,I207668);
and I_12065 (I207852,I207784,I207835);
DFFARX1 I_12066  ( .D(I207852), .CLK(I2702), .RSTB(I207651), .Q(I207619) );
nor I_12067 (I207883,I546477,I546495);
DFFARX1 I_12068  ( .D(I207883), .CLK(I2702), .RSTB(I207651), .Q(I207900) );
and I_12069 (I207616,I207716,I207900);
DFFARX1 I_12070  ( .D(I546504), .CLK(I2702), .RSTB(I207651), .Q(I207931) );
and I_12071 (I207948,I207931,I546492);
DFFARX1 I_12072  ( .D(I207948), .CLK(I2702), .RSTB(I207651), .Q(I207965) );
not I_12073 (I207628,I207965);
DFFARX1 I_12074  ( .D(I207948), .CLK(I2702), .RSTB(I207651), .Q(I207613) );
DFFARX1 I_12075  ( .D(I546498), .CLK(I2702), .RSTB(I207651), .Q(I208010) );
not I_12076 (I208027,I208010);
nor I_12077 (I208044,I207685,I208027);
and I_12078 (I208061,I207948,I208044);
or I_12079 (I208078,I207668,I208061);
DFFARX1 I_12080  ( .D(I208078), .CLK(I2702), .RSTB(I207651), .Q(I207634) );
nor I_12081 (I208109,I208010,I207818);
nand I_12082 (I207643,I207784,I208109);
nor I_12083 (I208140,I208010,I207733);
nand I_12084 (I207637,I207883,I208140);
not I_12085 (I207640,I208010);
nand I_12086 (I207631,I208010,I207733);
DFFARX1 I_12087  ( .D(I208010), .CLK(I2702), .RSTB(I207651), .Q(I207622) );
not I_12088 (I208246,I2709);
or I_12089 (I208263,I594681,I594675);
or I_12090 (I208280,I594669,I594681);
DFFARX1 I_12091  ( .D(I208280), .CLK(I2702), .RSTB(I208246), .Q(I208220) );
nor I_12092 (I208311,I594672,I594678);
not I_12093 (I208328,I208311);
not I_12094 (I208345,I594672);
and I_12095 (I208362,I208345,I594696);
nor I_12096 (I208379,I208362,I594675);
nor I_12097 (I208396,I594699,I594690);
DFFARX1 I_12098  ( .D(I208396), .CLK(I2702), .RSTB(I208246), .Q(I208413) );
nand I_12099 (I208430,I208413,I208263);
and I_12100 (I208447,I208379,I208430);
DFFARX1 I_12101  ( .D(I208447), .CLK(I2702), .RSTB(I208246), .Q(I208214) );
nor I_12102 (I208478,I594699,I594669);
DFFARX1 I_12103  ( .D(I208478), .CLK(I2702), .RSTB(I208246), .Q(I208495) );
and I_12104 (I208211,I208311,I208495);
DFFARX1 I_12105  ( .D(I594687), .CLK(I2702), .RSTB(I208246), .Q(I208526) );
and I_12106 (I208543,I208526,I594684);
DFFARX1 I_12107  ( .D(I208543), .CLK(I2702), .RSTB(I208246), .Q(I208560) );
not I_12108 (I208223,I208560);
DFFARX1 I_12109  ( .D(I208543), .CLK(I2702), .RSTB(I208246), .Q(I208208) );
DFFARX1 I_12110  ( .D(I594693), .CLK(I2702), .RSTB(I208246), .Q(I208605) );
not I_12111 (I208622,I208605);
nor I_12112 (I208639,I208280,I208622);
and I_12113 (I208656,I208543,I208639);
or I_12114 (I208673,I208263,I208656);
DFFARX1 I_12115  ( .D(I208673), .CLK(I2702), .RSTB(I208246), .Q(I208229) );
nor I_12116 (I208704,I208605,I208413);
nand I_12117 (I208238,I208379,I208704);
nor I_12118 (I208735,I208605,I208328);
nand I_12119 (I208232,I208478,I208735);
not I_12120 (I208235,I208605);
nand I_12121 (I208226,I208605,I208328);
DFFARX1 I_12122  ( .D(I208605), .CLK(I2702), .RSTB(I208246), .Q(I208217) );
not I_12123 (I208841,I2709);
or I_12124 (I208858,I7782,I7791);
or I_12125 (I208875,I7785,I7782);
DFFARX1 I_12126  ( .D(I208875), .CLK(I2702), .RSTB(I208841), .Q(I208815) );
nor I_12127 (I208906,I7761,I7764);
not I_12128 (I208923,I208906);
not I_12129 (I208940,I7761);
and I_12130 (I208957,I208940,I7773);
nor I_12131 (I208974,I208957,I7791);
nor I_12132 (I208991,I7779,I7770);
DFFARX1 I_12133  ( .D(I208991), .CLK(I2702), .RSTB(I208841), .Q(I209008) );
nand I_12134 (I209025,I209008,I208858);
and I_12135 (I209042,I208974,I209025);
DFFARX1 I_12136  ( .D(I209042), .CLK(I2702), .RSTB(I208841), .Q(I208809) );
nor I_12137 (I209073,I7779,I7785);
DFFARX1 I_12138  ( .D(I209073), .CLK(I2702), .RSTB(I208841), .Q(I209090) );
and I_12139 (I208806,I208906,I209090);
DFFARX1 I_12140  ( .D(I7776), .CLK(I2702), .RSTB(I208841), .Q(I209121) );
and I_12141 (I209138,I209121,I7767);
DFFARX1 I_12142  ( .D(I209138), .CLK(I2702), .RSTB(I208841), .Q(I209155) );
not I_12143 (I208818,I209155);
DFFARX1 I_12144  ( .D(I209138), .CLK(I2702), .RSTB(I208841), .Q(I208803) );
DFFARX1 I_12145  ( .D(I7788), .CLK(I2702), .RSTB(I208841), .Q(I209200) );
not I_12146 (I209217,I209200);
nor I_12147 (I209234,I208875,I209217);
and I_12148 (I209251,I209138,I209234);
or I_12149 (I209268,I208858,I209251);
DFFARX1 I_12150  ( .D(I209268), .CLK(I2702), .RSTB(I208841), .Q(I208824) );
nor I_12151 (I209299,I209200,I209008);
nand I_12152 (I208833,I208974,I209299);
nor I_12153 (I209330,I209200,I208923);
nand I_12154 (I208827,I209073,I209330);
not I_12155 (I208830,I209200);
nand I_12156 (I208821,I209200,I208923);
DFFARX1 I_12157  ( .D(I209200), .CLK(I2702), .RSTB(I208841), .Q(I208812) );
not I_12158 (I209436,I2709);
or I_12159 (I209453,I195267,I195252);
or I_12160 (I209470,I195249,I195267);
DFFARX1 I_12161  ( .D(I209470), .CLK(I2702), .RSTB(I209436), .Q(I209410) );
nor I_12162 (I209501,I195237,I195246);
not I_12163 (I209518,I209501);
not I_12164 (I209535,I195237);
and I_12165 (I209552,I209535,I195261);
nor I_12166 (I209569,I209552,I195252);
nor I_12167 (I209586,I195240,I195255);
DFFARX1 I_12168  ( .D(I209586), .CLK(I2702), .RSTB(I209436), .Q(I209603) );
nand I_12169 (I209620,I209603,I209453);
and I_12170 (I209637,I209569,I209620);
DFFARX1 I_12171  ( .D(I209637), .CLK(I2702), .RSTB(I209436), .Q(I209404) );
nor I_12172 (I209668,I195240,I195249);
DFFARX1 I_12173  ( .D(I209668), .CLK(I2702), .RSTB(I209436), .Q(I209685) );
and I_12174 (I209401,I209501,I209685);
DFFARX1 I_12175  ( .D(I195243), .CLK(I2702), .RSTB(I209436), .Q(I209716) );
and I_12176 (I209733,I209716,I195264);
DFFARX1 I_12177  ( .D(I209733), .CLK(I2702), .RSTB(I209436), .Q(I209750) );
not I_12178 (I209413,I209750);
DFFARX1 I_12179  ( .D(I209733), .CLK(I2702), .RSTB(I209436), .Q(I209398) );
DFFARX1 I_12180  ( .D(I195258), .CLK(I2702), .RSTB(I209436), .Q(I209795) );
not I_12181 (I209812,I209795);
nor I_12182 (I209829,I209470,I209812);
and I_12183 (I209846,I209733,I209829);
or I_12184 (I209863,I209453,I209846);
DFFARX1 I_12185  ( .D(I209863), .CLK(I2702), .RSTB(I209436), .Q(I209419) );
nor I_12186 (I209894,I209795,I209603);
nand I_12187 (I209428,I209569,I209894);
nor I_12188 (I209925,I209795,I209518);
nand I_12189 (I209422,I209668,I209925);
not I_12190 (I209425,I209795);
nand I_12191 (I209416,I209795,I209518);
DFFARX1 I_12192  ( .D(I209795), .CLK(I2702), .RSTB(I209436), .Q(I209407) );
not I_12193 (I210031,I2709);
or I_12194 (I210048,I76904,I76898);
or I_12195 (I210065,I76892,I76904);
DFFARX1 I_12196  ( .D(I210065), .CLK(I2702), .RSTB(I210031), .Q(I210005) );
nor I_12197 (I210096,I76910,I76901);
not I_12198 (I210113,I210096);
not I_12199 (I210130,I76910);
and I_12200 (I210147,I210130,I76907);
nor I_12201 (I210164,I210147,I76898);
nor I_12202 (I210181,I76883,I76889);
DFFARX1 I_12203  ( .D(I210181), .CLK(I2702), .RSTB(I210031), .Q(I210198) );
nand I_12204 (I210215,I210198,I210048);
and I_12205 (I210232,I210164,I210215);
DFFARX1 I_12206  ( .D(I210232), .CLK(I2702), .RSTB(I210031), .Q(I209999) );
nor I_12207 (I210263,I76883,I76892);
DFFARX1 I_12208  ( .D(I210263), .CLK(I2702), .RSTB(I210031), .Q(I210280) );
and I_12209 (I209996,I210096,I210280);
DFFARX1 I_12210  ( .D(I76895), .CLK(I2702), .RSTB(I210031), .Q(I210311) );
and I_12211 (I210328,I210311,I76913);
DFFARX1 I_12212  ( .D(I210328), .CLK(I2702), .RSTB(I210031), .Q(I210345) );
not I_12213 (I210008,I210345);
DFFARX1 I_12214  ( .D(I210328), .CLK(I2702), .RSTB(I210031), .Q(I209993) );
DFFARX1 I_12215  ( .D(I76886), .CLK(I2702), .RSTB(I210031), .Q(I210390) );
not I_12216 (I210407,I210390);
nor I_12217 (I210424,I210065,I210407);
and I_12218 (I210441,I210328,I210424);
or I_12219 (I210458,I210048,I210441);
DFFARX1 I_12220  ( .D(I210458), .CLK(I2702), .RSTB(I210031), .Q(I210014) );
nor I_12221 (I210489,I210390,I210198);
nand I_12222 (I210023,I210164,I210489);
nor I_12223 (I210520,I210390,I210113);
nand I_12224 (I210017,I210263,I210520);
not I_12225 (I210020,I210390);
nand I_12226 (I210011,I210390,I210113);
DFFARX1 I_12227  ( .D(I210390), .CLK(I2702), .RSTB(I210031), .Q(I210002) );
not I_12228 (I210626,I2709);
or I_12229 (I210643,I601821,I601815);
or I_12230 (I210660,I601809,I601821);
DFFARX1 I_12231  ( .D(I210660), .CLK(I2702), .RSTB(I210626), .Q(I210600) );
nor I_12232 (I210691,I601812,I601818);
not I_12233 (I210708,I210691);
not I_12234 (I210725,I601812);
and I_12235 (I210742,I210725,I601836);
nor I_12236 (I210759,I210742,I601815);
nor I_12237 (I210776,I601839,I601830);
DFFARX1 I_12238  ( .D(I210776), .CLK(I2702), .RSTB(I210626), .Q(I210793) );
nand I_12239 (I210810,I210793,I210643);
and I_12240 (I210827,I210759,I210810);
DFFARX1 I_12241  ( .D(I210827), .CLK(I2702), .RSTB(I210626), .Q(I210594) );
nor I_12242 (I210858,I601839,I601809);
DFFARX1 I_12243  ( .D(I210858), .CLK(I2702), .RSTB(I210626), .Q(I210875) );
and I_12244 (I210591,I210691,I210875);
DFFARX1 I_12245  ( .D(I601827), .CLK(I2702), .RSTB(I210626), .Q(I210906) );
and I_12246 (I210923,I210906,I601824);
DFFARX1 I_12247  ( .D(I210923), .CLK(I2702), .RSTB(I210626), .Q(I210940) );
not I_12248 (I210603,I210940);
DFFARX1 I_12249  ( .D(I210923), .CLK(I2702), .RSTB(I210626), .Q(I210588) );
DFFARX1 I_12250  ( .D(I601833), .CLK(I2702), .RSTB(I210626), .Q(I210985) );
not I_12251 (I211002,I210985);
nor I_12252 (I211019,I210660,I211002);
and I_12253 (I211036,I210923,I211019);
or I_12254 (I211053,I210643,I211036);
DFFARX1 I_12255  ( .D(I211053), .CLK(I2702), .RSTB(I210626), .Q(I210609) );
nor I_12256 (I211084,I210985,I210793);
nand I_12257 (I210618,I210759,I211084);
nor I_12258 (I211115,I210985,I210708);
nand I_12259 (I210612,I210858,I211115);
not I_12260 (I210615,I210985);
nand I_12261 (I210606,I210985,I210708);
DFFARX1 I_12262  ( .D(I210985), .CLK(I2702), .RSTB(I210626), .Q(I210597) );
not I_12263 (I211221,I2709);
or I_12264 (I211238,I555414,I555399);
or I_12265 (I211255,I555420,I555414);
DFFARX1 I_12266  ( .D(I211255), .CLK(I2702), .RSTB(I211221), .Q(I211195) );
nor I_12267 (I211286,I555426,I555408);
not I_12268 (I211303,I211286);
not I_12269 (I211320,I555426);
and I_12270 (I211337,I211320,I555405);
nor I_12271 (I211354,I211337,I555399);
nor I_12272 (I211371,I555402,I555411);
DFFARX1 I_12273  ( .D(I211371), .CLK(I2702), .RSTB(I211221), .Q(I211388) );
nand I_12274 (I211405,I211388,I211238);
and I_12275 (I211422,I211354,I211405);
DFFARX1 I_12276  ( .D(I211422), .CLK(I2702), .RSTB(I211221), .Q(I211189) );
nor I_12277 (I211453,I555402,I555420);
DFFARX1 I_12278  ( .D(I211453), .CLK(I2702), .RSTB(I211221), .Q(I211470) );
and I_12279 (I211186,I211286,I211470);
DFFARX1 I_12280  ( .D(I555429), .CLK(I2702), .RSTB(I211221), .Q(I211501) );
and I_12281 (I211518,I211501,I555417);
DFFARX1 I_12282  ( .D(I211518), .CLK(I2702), .RSTB(I211221), .Q(I211535) );
not I_12283 (I211198,I211535);
DFFARX1 I_12284  ( .D(I211518), .CLK(I2702), .RSTB(I211221), .Q(I211183) );
DFFARX1 I_12285  ( .D(I555423), .CLK(I2702), .RSTB(I211221), .Q(I211580) );
not I_12286 (I211597,I211580);
nor I_12287 (I211614,I211255,I211597);
and I_12288 (I211631,I211518,I211614);
or I_12289 (I211648,I211238,I211631);
DFFARX1 I_12290  ( .D(I211648), .CLK(I2702), .RSTB(I211221), .Q(I211204) );
nor I_12291 (I211679,I211580,I211388);
nand I_12292 (I211213,I211354,I211679);
nor I_12293 (I211710,I211580,I211303);
nand I_12294 (I211207,I211453,I211710);
not I_12295 (I211210,I211580);
nand I_12296 (I211201,I211580,I211303);
DFFARX1 I_12297  ( .D(I211580), .CLK(I2702), .RSTB(I211221), .Q(I211192) );
not I_12298 (I211816,I2709);
or I_12299 (I211833,I425432,I425417);
or I_12300 (I211850,I425426,I425432);
DFFARX1 I_12301  ( .D(I211850), .CLK(I2702), .RSTB(I211816), .Q(I211790) );
nor I_12302 (I211881,I425438,I425447);
not I_12303 (I211898,I211881);
not I_12304 (I211915,I425438);
and I_12305 (I211932,I211915,I425435);
nor I_12306 (I211949,I211932,I425417);
nor I_12307 (I211966,I425444,I425420);
DFFARX1 I_12308  ( .D(I211966), .CLK(I2702), .RSTB(I211816), .Q(I211983) );
nand I_12309 (I212000,I211983,I211833);
and I_12310 (I212017,I211949,I212000);
DFFARX1 I_12311  ( .D(I212017), .CLK(I2702), .RSTB(I211816), .Q(I211784) );
nor I_12312 (I212048,I425444,I425426);
DFFARX1 I_12313  ( .D(I212048), .CLK(I2702), .RSTB(I211816), .Q(I212065) );
and I_12314 (I211781,I211881,I212065);
DFFARX1 I_12315  ( .D(I425429), .CLK(I2702), .RSTB(I211816), .Q(I212096) );
and I_12316 (I212113,I212096,I425423);
DFFARX1 I_12317  ( .D(I212113), .CLK(I2702), .RSTB(I211816), .Q(I212130) );
not I_12318 (I211793,I212130);
DFFARX1 I_12319  ( .D(I212113), .CLK(I2702), .RSTB(I211816), .Q(I211778) );
DFFARX1 I_12320  ( .D(I425441), .CLK(I2702), .RSTB(I211816), .Q(I212175) );
not I_12321 (I212192,I212175);
nor I_12322 (I212209,I211850,I212192);
and I_12323 (I212226,I212113,I212209);
or I_12324 (I212243,I211833,I212226);
DFFARX1 I_12325  ( .D(I212243), .CLK(I2702), .RSTB(I211816), .Q(I211799) );
nor I_12326 (I212274,I212175,I211983);
nand I_12327 (I211808,I211949,I212274);
nor I_12328 (I212305,I212175,I211898);
nand I_12329 (I211802,I212048,I212305);
not I_12330 (I211805,I212175);
nand I_12331 (I211796,I212175,I211898);
DFFARX1 I_12332  ( .D(I212175), .CLK(I2702), .RSTB(I211816), .Q(I211787) );
not I_12333 (I212411,I2709);
or I_12334 (I212428,I403573,I403570);
or I_12335 (I212445,I403555,I403573);
DFFARX1 I_12336  ( .D(I212445), .CLK(I2702), .RSTB(I212411), .Q(I212385) );
nor I_12337 (I212476,I403564,I403567);
not I_12338 (I212493,I212476);
not I_12339 (I212510,I403564);
and I_12340 (I212527,I212510,I403579);
nor I_12341 (I212544,I212527,I403570);
nor I_12342 (I212561,I403585,I403561);
DFFARX1 I_12343  ( .D(I212561), .CLK(I2702), .RSTB(I212411), .Q(I212578) );
nand I_12344 (I212595,I212578,I212428);
and I_12345 (I212612,I212544,I212595);
DFFARX1 I_12346  ( .D(I212612), .CLK(I2702), .RSTB(I212411), .Q(I212379) );
nor I_12347 (I212643,I403585,I403555);
DFFARX1 I_12348  ( .D(I212643), .CLK(I2702), .RSTB(I212411), .Q(I212660) );
and I_12349 (I212376,I212476,I212660);
DFFARX1 I_12350  ( .D(I403576), .CLK(I2702), .RSTB(I212411), .Q(I212691) );
and I_12351 (I212708,I212691,I403582);
DFFARX1 I_12352  ( .D(I212708), .CLK(I2702), .RSTB(I212411), .Q(I212725) );
not I_12353 (I212388,I212725);
DFFARX1 I_12354  ( .D(I212708), .CLK(I2702), .RSTB(I212411), .Q(I212373) );
DFFARX1 I_12355  ( .D(I403558), .CLK(I2702), .RSTB(I212411), .Q(I212770) );
not I_12356 (I212787,I212770);
nor I_12357 (I212804,I212445,I212787);
and I_12358 (I212821,I212708,I212804);
or I_12359 (I212838,I212428,I212821);
DFFARX1 I_12360  ( .D(I212838), .CLK(I2702), .RSTB(I212411), .Q(I212394) );
nor I_12361 (I212869,I212770,I212578);
nand I_12362 (I212403,I212544,I212869);
nor I_12363 (I212900,I212770,I212493);
nand I_12364 (I212397,I212643,I212900);
not I_12365 (I212400,I212770);
nand I_12366 (I212391,I212770,I212493);
DFFARX1 I_12367  ( .D(I212770), .CLK(I2702), .RSTB(I212411), .Q(I212382) );
not I_12368 (I213006,I2709);
or I_12369 (I213023,I391299,I391296);
or I_12370 (I213040,I391281,I391299);
DFFARX1 I_12371  ( .D(I213040), .CLK(I2702), .RSTB(I213006), .Q(I212980) );
nor I_12372 (I213071,I391290,I391293);
not I_12373 (I213088,I213071);
not I_12374 (I213105,I391290);
and I_12375 (I213122,I213105,I391305);
nor I_12376 (I213139,I213122,I391296);
nor I_12377 (I213156,I391311,I391287);
DFFARX1 I_12378  ( .D(I213156), .CLK(I2702), .RSTB(I213006), .Q(I213173) );
nand I_12379 (I213190,I213173,I213023);
and I_12380 (I213207,I213139,I213190);
DFFARX1 I_12381  ( .D(I213207), .CLK(I2702), .RSTB(I213006), .Q(I212974) );
nor I_12382 (I213238,I391311,I391281);
DFFARX1 I_12383  ( .D(I213238), .CLK(I2702), .RSTB(I213006), .Q(I213255) );
and I_12384 (I212971,I213071,I213255);
DFFARX1 I_12385  ( .D(I391302), .CLK(I2702), .RSTB(I213006), .Q(I213286) );
and I_12386 (I213303,I213286,I391308);
DFFARX1 I_12387  ( .D(I213303), .CLK(I2702), .RSTB(I213006), .Q(I213320) );
not I_12388 (I212983,I213320);
DFFARX1 I_12389  ( .D(I213303), .CLK(I2702), .RSTB(I213006), .Q(I212968) );
DFFARX1 I_12390  ( .D(I391284), .CLK(I2702), .RSTB(I213006), .Q(I213365) );
not I_12391 (I213382,I213365);
nor I_12392 (I213399,I213040,I213382);
and I_12393 (I213416,I213303,I213399);
or I_12394 (I213433,I213023,I213416);
DFFARX1 I_12395  ( .D(I213433), .CLK(I2702), .RSTB(I213006), .Q(I212989) );
nor I_12396 (I213464,I213365,I213173);
nand I_12397 (I212998,I213139,I213464);
nor I_12398 (I213495,I213365,I213088);
nand I_12399 (I212992,I213238,I213495);
not I_12400 (I212995,I213365);
nand I_12401 (I212986,I213365,I213088);
DFFARX1 I_12402  ( .D(I213365), .CLK(I2702), .RSTB(I213006), .Q(I212977) );
not I_12403 (I213601,I2709);
or I_12404 (I213618,I496749,I496770);
or I_12405 (I213635,I496761,I496749);
DFFARX1 I_12406  ( .D(I213635), .CLK(I2702), .RSTB(I213601), .Q(I213575) );
nor I_12407 (I213666,I496779,I496773);
not I_12408 (I213683,I213666);
not I_12409 (I213700,I496779);
and I_12410 (I213717,I213700,I496758);
nor I_12411 (I213734,I213717,I496770);
nor I_12412 (I213751,I496767,I496752);
DFFARX1 I_12413  ( .D(I213751), .CLK(I2702), .RSTB(I213601), .Q(I213768) );
nand I_12414 (I213785,I213768,I213618);
and I_12415 (I213802,I213734,I213785);
DFFARX1 I_12416  ( .D(I213802), .CLK(I2702), .RSTB(I213601), .Q(I213569) );
nor I_12417 (I213833,I496767,I496761);
DFFARX1 I_12418  ( .D(I213833), .CLK(I2702), .RSTB(I213601), .Q(I213850) );
and I_12419 (I213566,I213666,I213850);
DFFARX1 I_12420  ( .D(I496764), .CLK(I2702), .RSTB(I213601), .Q(I213881) );
and I_12421 (I213898,I213881,I496755);
DFFARX1 I_12422  ( .D(I213898), .CLK(I2702), .RSTB(I213601), .Q(I213915) );
not I_12423 (I213578,I213915);
DFFARX1 I_12424  ( .D(I213898), .CLK(I2702), .RSTB(I213601), .Q(I213563) );
DFFARX1 I_12425  ( .D(I496776), .CLK(I2702), .RSTB(I213601), .Q(I213960) );
not I_12426 (I213977,I213960);
nor I_12427 (I213994,I213635,I213977);
and I_12428 (I214011,I213898,I213994);
or I_12429 (I214028,I213618,I214011);
DFFARX1 I_12430  ( .D(I214028), .CLK(I2702), .RSTB(I213601), .Q(I213584) );
nor I_12431 (I214059,I213960,I213768);
nand I_12432 (I213593,I213734,I214059);
nor I_12433 (I214090,I213960,I213683);
nand I_12434 (I213587,I213833,I214090);
not I_12435 (I213590,I213960);
nand I_12436 (I213581,I213960,I213683);
DFFARX1 I_12437  ( .D(I213960), .CLK(I2702), .RSTB(I213601), .Q(I213572) );
not I_12438 (I214196,I2709);
or I_12439 (I214213,I638838,I638835);
or I_12440 (I214230,I638865,I638838);
DFFARX1 I_12441  ( .D(I214230), .CLK(I2702), .RSTB(I214196), .Q(I214170) );
nor I_12442 (I214261,I638844,I638850);
not I_12443 (I214278,I214261);
not I_12444 (I214295,I638844);
and I_12445 (I214312,I214295,I638841);
nor I_12446 (I214329,I214312,I638835);
nor I_12447 (I214346,I638853,I638862);
DFFARX1 I_12448  ( .D(I214346), .CLK(I2702), .RSTB(I214196), .Q(I214363) );
nand I_12449 (I214380,I214363,I214213);
and I_12450 (I214397,I214329,I214380);
DFFARX1 I_12451  ( .D(I214397), .CLK(I2702), .RSTB(I214196), .Q(I214164) );
nor I_12452 (I214428,I638853,I638865);
DFFARX1 I_12453  ( .D(I214428), .CLK(I2702), .RSTB(I214196), .Q(I214445) );
and I_12454 (I214161,I214261,I214445);
DFFARX1 I_12455  ( .D(I638856), .CLK(I2702), .RSTB(I214196), .Q(I214476) );
and I_12456 (I214493,I214476,I638847);
DFFARX1 I_12457  ( .D(I214493), .CLK(I2702), .RSTB(I214196), .Q(I214510) );
not I_12458 (I214173,I214510);
DFFARX1 I_12459  ( .D(I214493), .CLK(I2702), .RSTB(I214196), .Q(I214158) );
DFFARX1 I_12460  ( .D(I638859), .CLK(I2702), .RSTB(I214196), .Q(I214555) );
not I_12461 (I214572,I214555);
nor I_12462 (I214589,I214230,I214572);
and I_12463 (I214606,I214493,I214589);
or I_12464 (I214623,I214213,I214606);
DFFARX1 I_12465  ( .D(I214623), .CLK(I2702), .RSTB(I214196), .Q(I214179) );
nor I_12466 (I214654,I214555,I214363);
nand I_12467 (I214188,I214329,I214654);
nor I_12468 (I214685,I214555,I214278);
nand I_12469 (I214182,I214428,I214685);
not I_12470 (I214185,I214555);
nand I_12471 (I214176,I214555,I214278);
DFFARX1 I_12472  ( .D(I214555), .CLK(I2702), .RSTB(I214196), .Q(I214167) );
not I_12473 (I214791,I2709);
or I_12474 (I214808,I186648,I186633);
or I_12475 (I214825,I186630,I186648);
DFFARX1 I_12476  ( .D(I214825), .CLK(I2702), .RSTB(I214791), .Q(I214765) );
nor I_12477 (I214856,I186618,I186627);
not I_12478 (I214873,I214856);
not I_12479 (I214890,I186618);
and I_12480 (I214907,I214890,I186642);
nor I_12481 (I214924,I214907,I186633);
nor I_12482 (I214941,I186621,I186636);
DFFARX1 I_12483  ( .D(I214941), .CLK(I2702), .RSTB(I214791), .Q(I214958) );
nand I_12484 (I214975,I214958,I214808);
and I_12485 (I214992,I214924,I214975);
DFFARX1 I_12486  ( .D(I214992), .CLK(I2702), .RSTB(I214791), .Q(I214759) );
nor I_12487 (I215023,I186621,I186630);
DFFARX1 I_12488  ( .D(I215023), .CLK(I2702), .RSTB(I214791), .Q(I215040) );
and I_12489 (I214756,I214856,I215040);
DFFARX1 I_12490  ( .D(I186624), .CLK(I2702), .RSTB(I214791), .Q(I215071) );
and I_12491 (I215088,I215071,I186645);
DFFARX1 I_12492  ( .D(I215088), .CLK(I2702), .RSTB(I214791), .Q(I215105) );
not I_12493 (I214768,I215105);
DFFARX1 I_12494  ( .D(I215088), .CLK(I2702), .RSTB(I214791), .Q(I214753) );
DFFARX1 I_12495  ( .D(I186639), .CLK(I2702), .RSTB(I214791), .Q(I215150) );
not I_12496 (I215167,I215150);
nor I_12497 (I215184,I214825,I215167);
and I_12498 (I215201,I215088,I215184);
or I_12499 (I215218,I214808,I215201);
DFFARX1 I_12500  ( .D(I215218), .CLK(I2702), .RSTB(I214791), .Q(I214774) );
nor I_12501 (I215249,I215150,I214958);
nand I_12502 (I214783,I214924,I215249);
nor I_12503 (I215280,I215150,I214873);
nand I_12504 (I214777,I215023,I215280);
not I_12505 (I214780,I215150);
nand I_12506 (I214771,I215150,I214873);
DFFARX1 I_12507  ( .D(I215150), .CLK(I2702), .RSTB(I214791), .Q(I214762) );
not I_12508 (I215386,I2709);
or I_12509 (I215403,I648273,I648270);
or I_12510 (I215420,I648300,I648273);
DFFARX1 I_12511  ( .D(I215420), .CLK(I2702), .RSTB(I215386), .Q(I215360) );
nor I_12512 (I215451,I648279,I648285);
not I_12513 (I215468,I215451);
not I_12514 (I215485,I648279);
and I_12515 (I215502,I215485,I648276);
nor I_12516 (I215519,I215502,I648270);
nor I_12517 (I215536,I648288,I648297);
DFFARX1 I_12518  ( .D(I215536), .CLK(I2702), .RSTB(I215386), .Q(I215553) );
nand I_12519 (I215570,I215553,I215403);
and I_12520 (I215587,I215519,I215570);
DFFARX1 I_12521  ( .D(I215587), .CLK(I2702), .RSTB(I215386), .Q(I215354) );
nor I_12522 (I215618,I648288,I648300);
DFFARX1 I_12523  ( .D(I215618), .CLK(I2702), .RSTB(I215386), .Q(I215635) );
and I_12524 (I215351,I215451,I215635);
DFFARX1 I_12525  ( .D(I648291), .CLK(I2702), .RSTB(I215386), .Q(I215666) );
and I_12526 (I215683,I215666,I648282);
DFFARX1 I_12527  ( .D(I215683), .CLK(I2702), .RSTB(I215386), .Q(I215700) );
not I_12528 (I215363,I215700);
DFFARX1 I_12529  ( .D(I215683), .CLK(I2702), .RSTB(I215386), .Q(I215348) );
DFFARX1 I_12530  ( .D(I648294), .CLK(I2702), .RSTB(I215386), .Q(I215745) );
not I_12531 (I215762,I215745);
nor I_12532 (I215779,I215420,I215762);
and I_12533 (I215796,I215683,I215779);
or I_12534 (I215813,I215403,I215796);
DFFARX1 I_12535  ( .D(I215813), .CLK(I2702), .RSTB(I215386), .Q(I215369) );
nor I_12536 (I215844,I215745,I215553);
nand I_12537 (I215378,I215519,I215844);
nor I_12538 (I215875,I215745,I215468);
nand I_12539 (I215372,I215618,I215875);
not I_12540 (I215375,I215745);
nand I_12541 (I215366,I215745,I215468);
DFFARX1 I_12542  ( .D(I215745), .CLK(I2702), .RSTB(I215386), .Q(I215357) );
not I_12543 (I215981,I2709);
or I_12544 (I215998,I378379,I378376);
or I_12545 (I216015,I378361,I378379);
DFFARX1 I_12546  ( .D(I216015), .CLK(I2702), .RSTB(I215981), .Q(I215955) );
nor I_12547 (I216046,I378370,I378373);
not I_12548 (I216063,I216046);
not I_12549 (I216080,I378370);
and I_12550 (I216097,I216080,I378385);
nor I_12551 (I216114,I216097,I378376);
nor I_12552 (I216131,I378391,I378367);
DFFARX1 I_12553  ( .D(I216131), .CLK(I2702), .RSTB(I215981), .Q(I216148) );
nand I_12554 (I216165,I216148,I215998);
and I_12555 (I216182,I216114,I216165);
DFFARX1 I_12556  ( .D(I216182), .CLK(I2702), .RSTB(I215981), .Q(I215949) );
nor I_12557 (I216213,I378391,I378361);
DFFARX1 I_12558  ( .D(I216213), .CLK(I2702), .RSTB(I215981), .Q(I216230) );
and I_12559 (I215946,I216046,I216230);
DFFARX1 I_12560  ( .D(I378382), .CLK(I2702), .RSTB(I215981), .Q(I216261) );
and I_12561 (I216278,I216261,I378388);
DFFARX1 I_12562  ( .D(I216278), .CLK(I2702), .RSTB(I215981), .Q(I216295) );
not I_12563 (I215958,I216295);
DFFARX1 I_12564  ( .D(I216278), .CLK(I2702), .RSTB(I215981), .Q(I215943) );
DFFARX1 I_12565  ( .D(I378364), .CLK(I2702), .RSTB(I215981), .Q(I216340) );
not I_12566 (I216357,I216340);
nor I_12567 (I216374,I216015,I216357);
and I_12568 (I216391,I216278,I216374);
or I_12569 (I216408,I215998,I216391);
DFFARX1 I_12570  ( .D(I216408), .CLK(I2702), .RSTB(I215981), .Q(I215964) );
nor I_12571 (I216439,I216340,I216148);
nand I_12572 (I215973,I216114,I216439);
nor I_12573 (I216470,I216340,I216063);
nand I_12574 (I215967,I216213,I216470);
not I_12575 (I215970,I216340);
nand I_12576 (I215961,I216340,I216063);
DFFARX1 I_12577  ( .D(I216340), .CLK(I2702), .RSTB(I215981), .Q(I215952) );
not I_12578 (I216576,I2709);
or I_12579 (I216593,I26295,I26304);
or I_12580 (I216610,I26298,I26295);
DFFARX1 I_12581  ( .D(I216610), .CLK(I2702), .RSTB(I216576), .Q(I216550) );
nor I_12582 (I216641,I26274,I26277);
not I_12583 (I216658,I216641);
not I_12584 (I216675,I26274);
and I_12585 (I216692,I216675,I26286);
nor I_12586 (I216709,I216692,I26304);
nor I_12587 (I216726,I26292,I26283);
DFFARX1 I_12588  ( .D(I216726), .CLK(I2702), .RSTB(I216576), .Q(I216743) );
nand I_12589 (I216760,I216743,I216593);
and I_12590 (I216777,I216709,I216760);
DFFARX1 I_12591  ( .D(I216777), .CLK(I2702), .RSTB(I216576), .Q(I216544) );
nor I_12592 (I216808,I26292,I26298);
DFFARX1 I_12593  ( .D(I216808), .CLK(I2702), .RSTB(I216576), .Q(I216825) );
and I_12594 (I216541,I216641,I216825);
DFFARX1 I_12595  ( .D(I26289), .CLK(I2702), .RSTB(I216576), .Q(I216856) );
and I_12596 (I216873,I216856,I26280);
DFFARX1 I_12597  ( .D(I216873), .CLK(I2702), .RSTB(I216576), .Q(I216890) );
not I_12598 (I216553,I216890);
DFFARX1 I_12599  ( .D(I216873), .CLK(I2702), .RSTB(I216576), .Q(I216538) );
DFFARX1 I_12600  ( .D(I26301), .CLK(I2702), .RSTB(I216576), .Q(I216935) );
not I_12601 (I216952,I216935);
nor I_12602 (I216969,I216610,I216952);
and I_12603 (I216986,I216873,I216969);
or I_12604 (I217003,I216593,I216986);
DFFARX1 I_12605  ( .D(I217003), .CLK(I2702), .RSTB(I216576), .Q(I216559) );
nor I_12606 (I217034,I216935,I216743);
nand I_12607 (I216568,I216709,I217034);
nor I_12608 (I217065,I216935,I216658);
nand I_12609 (I216562,I216808,I217065);
not I_12610 (I216565,I216935);
nand I_12611 (I216556,I216935,I216658);
DFFARX1 I_12612  ( .D(I216935), .CLK(I2702), .RSTB(I216576), .Q(I216547) );
not I_12613 (I217171,I2709);
or I_12614 (I217188,I459311,I459296);
or I_12615 (I217205,I459308,I459311);
DFFARX1 I_12616  ( .D(I217205), .CLK(I2702), .RSTB(I217171), .Q(I217145) );
nor I_12617 (I217236,I459290,I459281);
not I_12618 (I217253,I217236);
not I_12619 (I217270,I459290);
and I_12620 (I217287,I217270,I459305);
nor I_12621 (I217304,I217287,I459296);
nor I_12622 (I217321,I459284,I459302);
DFFARX1 I_12623  ( .D(I217321), .CLK(I2702), .RSTB(I217171), .Q(I217338) );
nand I_12624 (I217355,I217338,I217188);
and I_12625 (I217372,I217304,I217355);
DFFARX1 I_12626  ( .D(I217372), .CLK(I2702), .RSTB(I217171), .Q(I217139) );
nor I_12627 (I217403,I459284,I459308);
DFFARX1 I_12628  ( .D(I217403), .CLK(I2702), .RSTB(I217171), .Q(I217420) );
and I_12629 (I217136,I217236,I217420);
DFFARX1 I_12630  ( .D(I459293), .CLK(I2702), .RSTB(I217171), .Q(I217451) );
and I_12631 (I217468,I217451,I459287);
DFFARX1 I_12632  ( .D(I217468), .CLK(I2702), .RSTB(I217171), .Q(I217485) );
not I_12633 (I217148,I217485);
DFFARX1 I_12634  ( .D(I217468), .CLK(I2702), .RSTB(I217171), .Q(I217133) );
DFFARX1 I_12635  ( .D(I459299), .CLK(I2702), .RSTB(I217171), .Q(I217530) );
not I_12636 (I217547,I217530);
nor I_12637 (I217564,I217205,I217547);
and I_12638 (I217581,I217468,I217564);
or I_12639 (I217598,I217188,I217581);
DFFARX1 I_12640  ( .D(I217598), .CLK(I2702), .RSTB(I217171), .Q(I217154) );
nor I_12641 (I217629,I217530,I217338);
nand I_12642 (I217163,I217304,I217629);
nor I_12643 (I217660,I217530,I217253);
nand I_12644 (I217157,I217403,I217660);
not I_12645 (I217160,I217530);
nand I_12646 (I217151,I217530,I217253);
DFFARX1 I_12647  ( .D(I217530), .CLK(I2702), .RSTB(I217171), .Q(I217142) );
not I_12648 (I217766,I2709);
or I_12649 (I217783,I695564,I695582);
or I_12650 (I217800,I695567,I695564);
DFFARX1 I_12651  ( .D(I217800), .CLK(I2702), .RSTB(I217766), .Q(I217740) );
nor I_12652 (I217831,I695576,I695579);
not I_12653 (I217848,I217831);
not I_12654 (I217865,I695576);
and I_12655 (I217882,I217865,I695585);
nor I_12656 (I217899,I217882,I695582);
nor I_12657 (I217916,I695591,I695570);
DFFARX1 I_12658  ( .D(I217916), .CLK(I2702), .RSTB(I217766), .Q(I217933) );
nand I_12659 (I217950,I217933,I217783);
and I_12660 (I217967,I217899,I217950);
DFFARX1 I_12661  ( .D(I217967), .CLK(I2702), .RSTB(I217766), .Q(I217734) );
nor I_12662 (I217998,I695591,I695567);
DFFARX1 I_12663  ( .D(I217998), .CLK(I2702), .RSTB(I217766), .Q(I218015) );
and I_12664 (I217731,I217831,I218015);
DFFARX1 I_12665  ( .D(I695594), .CLK(I2702), .RSTB(I217766), .Q(I218046) );
and I_12666 (I218063,I218046,I695588);
DFFARX1 I_12667  ( .D(I218063), .CLK(I2702), .RSTB(I217766), .Q(I218080) );
not I_12668 (I217743,I218080);
DFFARX1 I_12669  ( .D(I218063), .CLK(I2702), .RSTB(I217766), .Q(I217728) );
DFFARX1 I_12670  ( .D(I695573), .CLK(I2702), .RSTB(I217766), .Q(I218125) );
not I_12671 (I218142,I218125);
nor I_12672 (I218159,I217800,I218142);
and I_12673 (I218176,I218063,I218159);
or I_12674 (I218193,I217783,I218176);
DFFARX1 I_12675  ( .D(I218193), .CLK(I2702), .RSTB(I217766), .Q(I217749) );
nor I_12676 (I218224,I218125,I217933);
nand I_12677 (I217758,I217899,I218224);
nor I_12678 (I218255,I218125,I217848);
nand I_12679 (I217752,I217998,I218255);
not I_12680 (I217755,I218125);
nand I_12681 (I217746,I218125,I217848);
DFFARX1 I_12682  ( .D(I218125), .CLK(I2702), .RSTB(I217766), .Q(I217737) );
not I_12683 (I218361,I2709);
or I_12684 (I218378,I106620,I106614);
or I_12685 (I218395,I106608,I106620);
DFFARX1 I_12686  ( .D(I218395), .CLK(I2702), .RSTB(I218361), .Q(I218335) );
nor I_12687 (I218426,I106626,I106617);
not I_12688 (I218443,I218426);
not I_12689 (I218460,I106626);
and I_12690 (I218477,I218460,I106623);
nor I_12691 (I218494,I218477,I106614);
nor I_12692 (I218511,I106599,I106605);
DFFARX1 I_12693  ( .D(I218511), .CLK(I2702), .RSTB(I218361), .Q(I218528) );
nand I_12694 (I218545,I218528,I218378);
and I_12695 (I218562,I218494,I218545);
DFFARX1 I_12696  ( .D(I218562), .CLK(I2702), .RSTB(I218361), .Q(I218329) );
nor I_12697 (I218593,I106599,I106608);
DFFARX1 I_12698  ( .D(I218593), .CLK(I2702), .RSTB(I218361), .Q(I218610) );
and I_12699 (I218326,I218426,I218610);
DFFARX1 I_12700  ( .D(I106611), .CLK(I2702), .RSTB(I218361), .Q(I218641) );
and I_12701 (I218658,I218641,I106629);
DFFARX1 I_12702  ( .D(I218658), .CLK(I2702), .RSTB(I218361), .Q(I218675) );
not I_12703 (I218338,I218675);
DFFARX1 I_12704  ( .D(I218658), .CLK(I2702), .RSTB(I218361), .Q(I218323) );
DFFARX1 I_12705  ( .D(I106602), .CLK(I2702), .RSTB(I218361), .Q(I218720) );
not I_12706 (I218737,I218720);
nor I_12707 (I218754,I218395,I218737);
and I_12708 (I218771,I218658,I218754);
or I_12709 (I218788,I218378,I218771);
DFFARX1 I_12710  ( .D(I218788), .CLK(I2702), .RSTB(I218361), .Q(I218344) );
nor I_12711 (I218819,I218720,I218528);
nand I_12712 (I218353,I218494,I218819);
nor I_12713 (I218850,I218720,I218443);
nand I_12714 (I218347,I218593,I218850);
not I_12715 (I218350,I218720);
nand I_12716 (I218341,I218720,I218443);
DFFARX1 I_12717  ( .D(I218720), .CLK(I2702), .RSTB(I218361), .Q(I218332) );
not I_12718 (I218956,I2709);
or I_12719 (I218973,I464513,I464498);
or I_12720 (I218990,I464510,I464513);
DFFARX1 I_12721  ( .D(I218990), .CLK(I2702), .RSTB(I218956), .Q(I218930) );
nor I_12722 (I219021,I464492,I464483);
not I_12723 (I219038,I219021);
not I_12724 (I219055,I464492);
and I_12725 (I219072,I219055,I464507);
nor I_12726 (I219089,I219072,I464498);
nor I_12727 (I219106,I464486,I464504);
DFFARX1 I_12728  ( .D(I219106), .CLK(I2702), .RSTB(I218956), .Q(I219123) );
nand I_12729 (I219140,I219123,I218973);
and I_12730 (I219157,I219089,I219140);
DFFARX1 I_12731  ( .D(I219157), .CLK(I2702), .RSTB(I218956), .Q(I218924) );
nor I_12732 (I219188,I464486,I464510);
DFFARX1 I_12733  ( .D(I219188), .CLK(I2702), .RSTB(I218956), .Q(I219205) );
and I_12734 (I218921,I219021,I219205);
DFFARX1 I_12735  ( .D(I464495), .CLK(I2702), .RSTB(I218956), .Q(I219236) );
and I_12736 (I219253,I219236,I464489);
DFFARX1 I_12737  ( .D(I219253), .CLK(I2702), .RSTB(I218956), .Q(I219270) );
not I_12738 (I218933,I219270);
DFFARX1 I_12739  ( .D(I219253), .CLK(I2702), .RSTB(I218956), .Q(I218918) );
DFFARX1 I_12740  ( .D(I464501), .CLK(I2702), .RSTB(I218956), .Q(I219315) );
not I_12741 (I219332,I219315);
nor I_12742 (I219349,I218990,I219332);
and I_12743 (I219366,I219253,I219349);
or I_12744 (I219383,I218973,I219366);
DFFARX1 I_12745  ( .D(I219383), .CLK(I2702), .RSTB(I218956), .Q(I218939) );
nor I_12746 (I219414,I219315,I219123);
nand I_12747 (I218948,I219089,I219414);
nor I_12748 (I219445,I219315,I219038);
nand I_12749 (I218942,I219188,I219445);
not I_12750 (I218945,I219315);
nand I_12751 (I218936,I219315,I219038);
DFFARX1 I_12752  ( .D(I219315), .CLK(I2702), .RSTB(I218956), .Q(I218927) );
not I_12753 (I219551,I2709);
or I_12754 (I219568,I632548,I632545);
or I_12755 (I219585,I632575,I632548);
DFFARX1 I_12756  ( .D(I219585), .CLK(I2702), .RSTB(I219551), .Q(I219525) );
nor I_12757 (I219616,I632554,I632560);
not I_12758 (I219633,I219616);
not I_12759 (I219650,I632554);
and I_12760 (I219667,I219650,I632551);
nor I_12761 (I219684,I219667,I632545);
nor I_12762 (I219701,I632563,I632572);
DFFARX1 I_12763  ( .D(I219701), .CLK(I2702), .RSTB(I219551), .Q(I219718) );
nand I_12764 (I219735,I219718,I219568);
and I_12765 (I219752,I219684,I219735);
DFFARX1 I_12766  ( .D(I219752), .CLK(I2702), .RSTB(I219551), .Q(I219519) );
nor I_12767 (I219783,I632563,I632575);
DFFARX1 I_12768  ( .D(I219783), .CLK(I2702), .RSTB(I219551), .Q(I219800) );
and I_12769 (I219516,I219616,I219800);
DFFARX1 I_12770  ( .D(I632566), .CLK(I2702), .RSTB(I219551), .Q(I219831) );
and I_12771 (I219848,I219831,I632557);
DFFARX1 I_12772  ( .D(I219848), .CLK(I2702), .RSTB(I219551), .Q(I219865) );
not I_12773 (I219528,I219865);
DFFARX1 I_12774  ( .D(I219848), .CLK(I2702), .RSTB(I219551), .Q(I219513) );
DFFARX1 I_12775  ( .D(I632569), .CLK(I2702), .RSTB(I219551), .Q(I219910) );
not I_12776 (I219927,I219910);
nor I_12777 (I219944,I219585,I219927);
and I_12778 (I219961,I219848,I219944);
or I_12779 (I219978,I219568,I219961);
DFFARX1 I_12780  ( .D(I219978), .CLK(I2702), .RSTB(I219551), .Q(I219534) );
nor I_12781 (I220009,I219910,I219718);
nand I_12782 (I219543,I219684,I220009);
nor I_12783 (I220040,I219910,I219633);
nand I_12784 (I219537,I219783,I220040);
not I_12785 (I219540,I219910);
nand I_12786 (I219531,I219910,I219633);
DFFARX1 I_12787  ( .D(I219910), .CLK(I2702), .RSTB(I219551), .Q(I219522) );
not I_12788 (I220146,I2709);
or I_12789 (I220163,I73028,I73022);
or I_12790 (I220180,I73016,I73028);
DFFARX1 I_12791  ( .D(I220180), .CLK(I2702), .RSTB(I220146), .Q(I220120) );
nor I_12792 (I220211,I73034,I73025);
not I_12793 (I220228,I220211);
not I_12794 (I220245,I73034);
and I_12795 (I220262,I220245,I73031);
nor I_12796 (I220279,I220262,I73022);
nor I_12797 (I220296,I73007,I73013);
DFFARX1 I_12798  ( .D(I220296), .CLK(I2702), .RSTB(I220146), .Q(I220313) );
nand I_12799 (I220330,I220313,I220163);
and I_12800 (I220347,I220279,I220330);
DFFARX1 I_12801  ( .D(I220347), .CLK(I2702), .RSTB(I220146), .Q(I220114) );
nor I_12802 (I220378,I73007,I73016);
DFFARX1 I_12803  ( .D(I220378), .CLK(I2702), .RSTB(I220146), .Q(I220395) );
and I_12804 (I220111,I220211,I220395);
DFFARX1 I_12805  ( .D(I73019), .CLK(I2702), .RSTB(I220146), .Q(I220426) );
and I_12806 (I220443,I220426,I73037);
DFFARX1 I_12807  ( .D(I220443), .CLK(I2702), .RSTB(I220146), .Q(I220460) );
not I_12808 (I220123,I220460);
DFFARX1 I_12809  ( .D(I220443), .CLK(I2702), .RSTB(I220146), .Q(I220108) );
DFFARX1 I_12810  ( .D(I73010), .CLK(I2702), .RSTB(I220146), .Q(I220505) );
not I_12811 (I220522,I220505);
nor I_12812 (I220539,I220180,I220522);
and I_12813 (I220556,I220443,I220539);
or I_12814 (I220573,I220163,I220556);
DFFARX1 I_12815  ( .D(I220573), .CLK(I2702), .RSTB(I220146), .Q(I220129) );
nor I_12816 (I220604,I220505,I220313);
nand I_12817 (I220138,I220279,I220604);
nor I_12818 (I220635,I220505,I220228);
nand I_12819 (I220132,I220378,I220635);
not I_12820 (I220135,I220505);
nand I_12821 (I220126,I220505,I220228);
DFFARX1 I_12822  ( .D(I220505), .CLK(I2702), .RSTB(I220146), .Q(I220117) );
not I_12823 (I220741,I2709);
or I_12824 (I220758,I232023,I232014);
or I_12825 (I220775,I232035,I232023);
DFFARX1 I_12826  ( .D(I220775), .CLK(I2702), .RSTB(I220741), .Q(I220715) );
nor I_12827 (I220806,I232038,I232017);
not I_12828 (I220823,I220806);
not I_12829 (I220840,I232038);
and I_12830 (I220857,I220840,I232026);
nor I_12831 (I220874,I220857,I232014);
nor I_12832 (I220891,I232011,I232029);
DFFARX1 I_12833  ( .D(I220891), .CLK(I2702), .RSTB(I220741), .Q(I220908) );
nand I_12834 (I220925,I220908,I220758);
and I_12835 (I220942,I220874,I220925);
DFFARX1 I_12836  ( .D(I220942), .CLK(I2702), .RSTB(I220741), .Q(I220709) );
nor I_12837 (I220973,I232011,I232035);
DFFARX1 I_12838  ( .D(I220973), .CLK(I2702), .RSTB(I220741), .Q(I220990) );
and I_12839 (I220706,I220806,I220990);
DFFARX1 I_12840  ( .D(I232032), .CLK(I2702), .RSTB(I220741), .Q(I221021) );
and I_12841 (I221038,I221021,I232008);
DFFARX1 I_12842  ( .D(I221038), .CLK(I2702), .RSTB(I220741), .Q(I221055) );
not I_12843 (I220718,I221055);
DFFARX1 I_12844  ( .D(I221038), .CLK(I2702), .RSTB(I220741), .Q(I220703) );
DFFARX1 I_12845  ( .D(I232020), .CLK(I2702), .RSTB(I220741), .Q(I221100) );
not I_12846 (I221117,I221100);
nor I_12847 (I221134,I220775,I221117);
and I_12848 (I221151,I221038,I221134);
or I_12849 (I221168,I220758,I221151);
DFFARX1 I_12850  ( .D(I221168), .CLK(I2702), .RSTB(I220741), .Q(I220724) );
nor I_12851 (I221199,I221100,I220908);
nand I_12852 (I220733,I220874,I221199);
nor I_12853 (I221230,I221100,I220823);
nand I_12854 (I220727,I220973,I221230);
not I_12855 (I220730,I221100);
nand I_12856 (I220721,I221100,I220823);
DFFARX1 I_12857  ( .D(I221100), .CLK(I2702), .RSTB(I220741), .Q(I220712) );
not I_12858 (I221336,I2709);
or I_12859 (I221353,I562554,I562539);
or I_12860 (I221370,I562560,I562554);
DFFARX1 I_12861  ( .D(I221370), .CLK(I2702), .RSTB(I221336), .Q(I221310) );
nor I_12862 (I221401,I562566,I562548);
not I_12863 (I221418,I221401);
not I_12864 (I221435,I562566);
and I_12865 (I221452,I221435,I562545);
nor I_12866 (I221469,I221452,I562539);
nor I_12867 (I221486,I562542,I562551);
DFFARX1 I_12868  ( .D(I221486), .CLK(I2702), .RSTB(I221336), .Q(I221503) );
nand I_12869 (I221520,I221503,I221353);
and I_12870 (I221537,I221469,I221520);
DFFARX1 I_12871  ( .D(I221537), .CLK(I2702), .RSTB(I221336), .Q(I221304) );
nor I_12872 (I221568,I562542,I562560);
DFFARX1 I_12873  ( .D(I221568), .CLK(I2702), .RSTB(I221336), .Q(I221585) );
and I_12874 (I221301,I221401,I221585);
DFFARX1 I_12875  ( .D(I562569), .CLK(I2702), .RSTB(I221336), .Q(I221616) );
and I_12876 (I221633,I221616,I562557);
DFFARX1 I_12877  ( .D(I221633), .CLK(I2702), .RSTB(I221336), .Q(I221650) );
not I_12878 (I221313,I221650);
DFFARX1 I_12879  ( .D(I221633), .CLK(I2702), .RSTB(I221336), .Q(I221298) );
DFFARX1 I_12880  ( .D(I562563), .CLK(I2702), .RSTB(I221336), .Q(I221695) );
not I_12881 (I221712,I221695);
nor I_12882 (I221729,I221370,I221712);
and I_12883 (I221746,I221633,I221729);
or I_12884 (I221763,I221353,I221746);
DFFARX1 I_12885  ( .D(I221763), .CLK(I2702), .RSTB(I221336), .Q(I221319) );
nor I_12886 (I221794,I221695,I221503);
nand I_12887 (I221328,I221469,I221794);
nor I_12888 (I221825,I221695,I221418);
nand I_12889 (I221322,I221568,I221825);
not I_12890 (I221325,I221695);
nand I_12891 (I221316,I221695,I221418);
DFFARX1 I_12892  ( .D(I221695), .CLK(I2702), .RSTB(I221336), .Q(I221307) );
not I_12893 (I221931,I2709);
or I_12894 (I221948,I87240,I87234);
or I_12895 (I221965,I87228,I87240);
DFFARX1 I_12896  ( .D(I221965), .CLK(I2702), .RSTB(I221931), .Q(I221905) );
nor I_12897 (I221996,I87246,I87237);
not I_12898 (I222013,I221996);
not I_12899 (I222030,I87246);
and I_12900 (I222047,I222030,I87243);
nor I_12901 (I222064,I222047,I87234);
nor I_12902 (I222081,I87219,I87225);
DFFARX1 I_12903  ( .D(I222081), .CLK(I2702), .RSTB(I221931), .Q(I222098) );
nand I_12904 (I222115,I222098,I221948);
and I_12905 (I222132,I222064,I222115);
DFFARX1 I_12906  ( .D(I222132), .CLK(I2702), .RSTB(I221931), .Q(I221899) );
nor I_12907 (I222163,I87219,I87228);
DFFARX1 I_12908  ( .D(I222163), .CLK(I2702), .RSTB(I221931), .Q(I222180) );
and I_12909 (I221896,I221996,I222180);
DFFARX1 I_12910  ( .D(I87231), .CLK(I2702), .RSTB(I221931), .Q(I222211) );
and I_12911 (I222228,I222211,I87249);
DFFARX1 I_12912  ( .D(I222228), .CLK(I2702), .RSTB(I221931), .Q(I222245) );
not I_12913 (I221908,I222245);
DFFARX1 I_12914  ( .D(I222228), .CLK(I2702), .RSTB(I221931), .Q(I221893) );
DFFARX1 I_12915  ( .D(I87222), .CLK(I2702), .RSTB(I221931), .Q(I222290) );
not I_12916 (I222307,I222290);
nor I_12917 (I222324,I221965,I222307);
and I_12918 (I222341,I222228,I222324);
or I_12919 (I222358,I221948,I222341);
DFFARX1 I_12920  ( .D(I222358), .CLK(I2702), .RSTB(I221931), .Q(I221914) );
nor I_12921 (I222389,I222290,I222098);
nand I_12922 (I221923,I222064,I222389);
nor I_12923 (I222420,I222290,I222013);
nand I_12924 (I221917,I222163,I222420);
not I_12925 (I221920,I222290);
nand I_12926 (I221911,I222290,I222013);
DFFARX1 I_12927  ( .D(I222290), .CLK(I2702), .RSTB(I221931), .Q(I221902) );
not I_12928 (I222526,I2709);
or I_12929 (I222543,I294687,I294702);
or I_12930 (I222560,I294690,I294687);
DFFARX1 I_12931  ( .D(I222560), .CLK(I2702), .RSTB(I222526), .Q(I222500) );
nor I_12932 (I222591,I294693,I294708);
not I_12933 (I222608,I222591);
not I_12934 (I222625,I294693);
and I_12935 (I222642,I222625,I294696);
nor I_12936 (I222659,I222642,I294702);
nor I_12937 (I222676,I294699,I294717);
DFFARX1 I_12938  ( .D(I222676), .CLK(I2702), .RSTB(I222526), .Q(I222693) );
nand I_12939 (I222710,I222693,I222543);
and I_12940 (I222727,I222659,I222710);
DFFARX1 I_12941  ( .D(I222727), .CLK(I2702), .RSTB(I222526), .Q(I222494) );
nor I_12942 (I222758,I294699,I294690);
DFFARX1 I_12943  ( .D(I222758), .CLK(I2702), .RSTB(I222526), .Q(I222775) );
and I_12944 (I222491,I222591,I222775);
DFFARX1 I_12945  ( .D(I294714), .CLK(I2702), .RSTB(I222526), .Q(I222806) );
and I_12946 (I222823,I222806,I294705);
DFFARX1 I_12947  ( .D(I222823), .CLK(I2702), .RSTB(I222526), .Q(I222840) );
not I_12948 (I222503,I222840);
DFFARX1 I_12949  ( .D(I222823), .CLK(I2702), .RSTB(I222526), .Q(I222488) );
DFFARX1 I_12950  ( .D(I294711), .CLK(I2702), .RSTB(I222526), .Q(I222885) );
not I_12951 (I222902,I222885);
nor I_12952 (I222919,I222560,I222902);
and I_12953 (I222936,I222823,I222919);
or I_12954 (I222953,I222543,I222936);
DFFARX1 I_12955  ( .D(I222953), .CLK(I2702), .RSTB(I222526), .Q(I222509) );
nor I_12956 (I222984,I222885,I222693);
nand I_12957 (I222518,I222659,I222984);
nor I_12958 (I223015,I222885,I222608);
nand I_12959 (I222512,I222758,I223015);
not I_12960 (I222515,I222885);
nand I_12961 (I222506,I222885,I222608);
DFFARX1 I_12962  ( .D(I222885), .CLK(I2702), .RSTB(I222526), .Q(I222497) );
not I_12963 (I223121,I2709);
or I_12964 (I223138,I590516,I590510);
or I_12965 (I223155,I590504,I590516);
DFFARX1 I_12966  ( .D(I223155), .CLK(I2702), .RSTB(I223121), .Q(I223095) );
nor I_12967 (I223186,I590507,I590513);
not I_12968 (I223203,I223186);
not I_12969 (I223220,I590507);
and I_12970 (I223237,I223220,I590531);
nor I_12971 (I223254,I223237,I590510);
nor I_12972 (I223271,I590534,I590525);
DFFARX1 I_12973  ( .D(I223271), .CLK(I2702), .RSTB(I223121), .Q(I223288) );
nand I_12974 (I223305,I223288,I223138);
and I_12975 (I223322,I223254,I223305);
DFFARX1 I_12976  ( .D(I223322), .CLK(I2702), .RSTB(I223121), .Q(I223089) );
nor I_12977 (I223353,I590534,I590504);
DFFARX1 I_12978  ( .D(I223353), .CLK(I2702), .RSTB(I223121), .Q(I223370) );
and I_12979 (I223086,I223186,I223370);
DFFARX1 I_12980  ( .D(I590522), .CLK(I2702), .RSTB(I223121), .Q(I223401) );
and I_12981 (I223418,I223401,I590519);
DFFARX1 I_12982  ( .D(I223418), .CLK(I2702), .RSTB(I223121), .Q(I223435) );
not I_12983 (I223098,I223435);
DFFARX1 I_12984  ( .D(I223418), .CLK(I2702), .RSTB(I223121), .Q(I223083) );
DFFARX1 I_12985  ( .D(I590528), .CLK(I2702), .RSTB(I223121), .Q(I223480) );
not I_12986 (I223497,I223480);
nor I_12987 (I223514,I223155,I223497);
and I_12988 (I223531,I223418,I223514);
or I_12989 (I223548,I223138,I223531);
DFFARX1 I_12990  ( .D(I223548), .CLK(I2702), .RSTB(I223121), .Q(I223104) );
nor I_12991 (I223579,I223480,I223288);
nand I_12992 (I223113,I223254,I223579);
nor I_12993 (I223610,I223480,I223203);
nand I_12994 (I223107,I223353,I223610);
not I_12995 (I223110,I223480);
nand I_12996 (I223101,I223480,I223203);
DFFARX1 I_12997  ( .D(I223480), .CLK(I2702), .RSTB(I223121), .Q(I223092) );
not I_12998 (I223716,I2709);
or I_12999 (I223733,I388715,I388712);
or I_13000 (I223750,I388697,I388715);
DFFARX1 I_13001  ( .D(I223750), .CLK(I2702), .RSTB(I223716), .Q(I223690) );
nor I_13002 (I223781,I388706,I388709);
not I_13003 (I223798,I223781);
not I_13004 (I223815,I388706);
and I_13005 (I223832,I223815,I388721);
nor I_13006 (I223849,I223832,I388712);
nor I_13007 (I223866,I388727,I388703);
DFFARX1 I_13008  ( .D(I223866), .CLK(I2702), .RSTB(I223716), .Q(I223883) );
nand I_13009 (I223900,I223883,I223733);
and I_13010 (I223917,I223849,I223900);
DFFARX1 I_13011  ( .D(I223917), .CLK(I2702), .RSTB(I223716), .Q(I223684) );
nor I_13012 (I223948,I388727,I388697);
DFFARX1 I_13013  ( .D(I223948), .CLK(I2702), .RSTB(I223716), .Q(I223965) );
and I_13014 (I223681,I223781,I223965);
DFFARX1 I_13015  ( .D(I388718), .CLK(I2702), .RSTB(I223716), .Q(I223996) );
and I_13016 (I224013,I223996,I388724);
DFFARX1 I_13017  ( .D(I224013), .CLK(I2702), .RSTB(I223716), .Q(I224030) );
not I_13018 (I223693,I224030);
DFFARX1 I_13019  ( .D(I224013), .CLK(I2702), .RSTB(I223716), .Q(I223678) );
DFFARX1 I_13020  ( .D(I388700), .CLK(I2702), .RSTB(I223716), .Q(I224075) );
not I_13021 (I224092,I224075);
nor I_13022 (I224109,I223750,I224092);
and I_13023 (I224126,I224013,I224109);
or I_13024 (I224143,I223733,I224126);
DFFARX1 I_13025  ( .D(I224143), .CLK(I2702), .RSTB(I223716), .Q(I223699) );
nor I_13026 (I224174,I224075,I223883);
nand I_13027 (I223708,I223849,I224174);
nor I_13028 (I224205,I224075,I223798);
nand I_13029 (I223702,I223948,I224205);
not I_13030 (I223705,I224075);
nand I_13031 (I223696,I224075,I223798);
DFFARX1 I_13032  ( .D(I224075), .CLK(I2702), .RSTB(I223716), .Q(I223687) );
not I_13033 (I224311,I2709);
or I_13034 (I224328,I400989,I400986);
or I_13035 (I224345,I400971,I400989);
DFFARX1 I_13036  ( .D(I224345), .CLK(I2702), .RSTB(I224311), .Q(I224285) );
nor I_13037 (I224376,I400980,I400983);
not I_13038 (I224393,I224376);
not I_13039 (I224410,I400980);
and I_13040 (I224427,I224410,I400995);
nor I_13041 (I224444,I224427,I400986);
nor I_13042 (I224461,I401001,I400977);
DFFARX1 I_13043  ( .D(I224461), .CLK(I2702), .RSTB(I224311), .Q(I224478) );
nand I_13044 (I224495,I224478,I224328);
and I_13045 (I224512,I224444,I224495);
DFFARX1 I_13046  ( .D(I224512), .CLK(I2702), .RSTB(I224311), .Q(I224279) );
nor I_13047 (I224543,I401001,I400971);
DFFARX1 I_13048  ( .D(I224543), .CLK(I2702), .RSTB(I224311), .Q(I224560) );
and I_13049 (I224276,I224376,I224560);
DFFARX1 I_13050  ( .D(I400992), .CLK(I2702), .RSTB(I224311), .Q(I224591) );
and I_13051 (I224608,I224591,I400998);
DFFARX1 I_13052  ( .D(I224608), .CLK(I2702), .RSTB(I224311), .Q(I224625) );
not I_13053 (I224288,I224625);
DFFARX1 I_13054  ( .D(I224608), .CLK(I2702), .RSTB(I224311), .Q(I224273) );
DFFARX1 I_13055  ( .D(I400974), .CLK(I2702), .RSTB(I224311), .Q(I224670) );
not I_13056 (I224687,I224670);
nor I_13057 (I224704,I224345,I224687);
and I_13058 (I224721,I224608,I224704);
or I_13059 (I224738,I224328,I224721);
DFFARX1 I_13060  ( .D(I224738), .CLK(I2702), .RSTB(I224311), .Q(I224294) );
nor I_13061 (I224769,I224670,I224478);
nand I_13062 (I224303,I224444,I224769);
nor I_13063 (I224800,I224670,I224393);
nand I_13064 (I224297,I224543,I224800);
not I_13065 (I224300,I224670);
nand I_13066 (I224291,I224670,I224393);
DFFARX1 I_13067  ( .D(I224670), .CLK(I2702), .RSTB(I224311), .Q(I224282) );
not I_13068 (I224906,I2709);
or I_13069 (I224923,I265515,I265530);
or I_13070 (I224940,I265518,I265515);
DFFARX1 I_13071  ( .D(I224940), .CLK(I2702), .RSTB(I224906), .Q(I224880) );
nor I_13072 (I224971,I265521,I265536);
not I_13073 (I224988,I224971);
not I_13074 (I225005,I265521);
and I_13075 (I225022,I225005,I265524);
nor I_13076 (I225039,I225022,I265530);
nor I_13077 (I225056,I265527,I265545);
DFFARX1 I_13078  ( .D(I225056), .CLK(I2702), .RSTB(I224906), .Q(I225073) );
nand I_13079 (I225090,I225073,I224923);
and I_13080 (I225107,I225039,I225090);
DFFARX1 I_13081  ( .D(I225107), .CLK(I2702), .RSTB(I224906), .Q(I224874) );
nor I_13082 (I225138,I265527,I265518);
DFFARX1 I_13083  ( .D(I225138), .CLK(I2702), .RSTB(I224906), .Q(I225155) );
and I_13084 (I224871,I224971,I225155);
DFFARX1 I_13085  ( .D(I265542), .CLK(I2702), .RSTB(I224906), .Q(I225186) );
and I_13086 (I225203,I225186,I265533);
DFFARX1 I_13087  ( .D(I225203), .CLK(I2702), .RSTB(I224906), .Q(I225220) );
not I_13088 (I224883,I225220);
DFFARX1 I_13089  ( .D(I225203), .CLK(I2702), .RSTB(I224906), .Q(I224868) );
DFFARX1 I_13090  ( .D(I265539), .CLK(I2702), .RSTB(I224906), .Q(I225265) );
not I_13091 (I225282,I225265);
nor I_13092 (I225299,I224940,I225282);
and I_13093 (I225316,I225203,I225299);
or I_13094 (I225333,I224923,I225316);
DFFARX1 I_13095  ( .D(I225333), .CLK(I2702), .RSTB(I224906), .Q(I224889) );
nor I_13096 (I225364,I225265,I225073);
nand I_13097 (I224898,I225039,I225364);
nor I_13098 (I225395,I225265,I224988);
nand I_13099 (I224892,I225138,I225395);
not I_13100 (I224895,I225265);
nand I_13101 (I224886,I225265,I224988);
DFFARX1 I_13102  ( .D(I225265), .CLK(I2702), .RSTB(I224906), .Q(I224877) );
not I_13103 (I225501,I2709);
or I_13104 (I225518,I288057,I288072);
or I_13105 (I225535,I288060,I288057);
DFFARX1 I_13106  ( .D(I225535), .CLK(I2702), .RSTB(I225501), .Q(I225475) );
nor I_13107 (I225566,I288063,I288078);
not I_13108 (I225583,I225566);
not I_13109 (I225600,I288063);
and I_13110 (I225617,I225600,I288066);
nor I_13111 (I225634,I225617,I288072);
nor I_13112 (I225651,I288069,I288087);
DFFARX1 I_13113  ( .D(I225651), .CLK(I2702), .RSTB(I225501), .Q(I225668) );
nand I_13114 (I225685,I225668,I225518);
and I_13115 (I225702,I225634,I225685);
DFFARX1 I_13116  ( .D(I225702), .CLK(I2702), .RSTB(I225501), .Q(I225469) );
nor I_13117 (I225733,I288069,I288060);
DFFARX1 I_13118  ( .D(I225733), .CLK(I2702), .RSTB(I225501), .Q(I225750) );
and I_13119 (I225466,I225566,I225750);
DFFARX1 I_13120  ( .D(I288084), .CLK(I2702), .RSTB(I225501), .Q(I225781) );
and I_13121 (I225798,I225781,I288075);
DFFARX1 I_13122  ( .D(I225798), .CLK(I2702), .RSTB(I225501), .Q(I225815) );
not I_13123 (I225478,I225815);
DFFARX1 I_13124  ( .D(I225798), .CLK(I2702), .RSTB(I225501), .Q(I225463) );
DFFARX1 I_13125  ( .D(I288081), .CLK(I2702), .RSTB(I225501), .Q(I225860) );
not I_13126 (I225877,I225860);
nor I_13127 (I225894,I225535,I225877);
and I_13128 (I225911,I225798,I225894);
or I_13129 (I225928,I225518,I225911);
DFFARX1 I_13130  ( .D(I225928), .CLK(I2702), .RSTB(I225501), .Q(I225484) );
nor I_13131 (I225959,I225860,I225668);
nand I_13132 (I225493,I225634,I225959);
nor I_13133 (I225990,I225860,I225583);
nand I_13134 (I225487,I225733,I225990);
not I_13135 (I225490,I225860);
nand I_13136 (I225481,I225860,I225583);
DFFARX1 I_13137  ( .D(I225860), .CLK(I2702), .RSTB(I225501), .Q(I225472) );
not I_13138 (I226096,I2709);
or I_13139 (I226113,I241543,I241534);
or I_13140 (I226130,I241555,I241543);
DFFARX1 I_13141  ( .D(I226130), .CLK(I2702), .RSTB(I226096), .Q(I226070) );
nor I_13142 (I226161,I241558,I241537);
not I_13143 (I226178,I226161);
not I_13144 (I226195,I241558);
and I_13145 (I226212,I226195,I241546);
nor I_13146 (I226229,I226212,I241534);
nor I_13147 (I226246,I241531,I241549);
DFFARX1 I_13148  ( .D(I226246), .CLK(I2702), .RSTB(I226096), .Q(I226263) );
nand I_13149 (I226280,I226263,I226113);
and I_13150 (I226297,I226229,I226280);
DFFARX1 I_13151  ( .D(I226297), .CLK(I2702), .RSTB(I226096), .Q(I226064) );
nor I_13152 (I226328,I241531,I241555);
DFFARX1 I_13153  ( .D(I226328), .CLK(I2702), .RSTB(I226096), .Q(I226345) );
and I_13154 (I226061,I226161,I226345);
DFFARX1 I_13155  ( .D(I241552), .CLK(I2702), .RSTB(I226096), .Q(I226376) );
and I_13156 (I226393,I226376,I241528);
DFFARX1 I_13157  ( .D(I226393), .CLK(I2702), .RSTB(I226096), .Q(I226410) );
not I_13158 (I226073,I226410);
DFFARX1 I_13159  ( .D(I226393), .CLK(I2702), .RSTB(I226096), .Q(I226058) );
DFFARX1 I_13160  ( .D(I241540), .CLK(I2702), .RSTB(I226096), .Q(I226455) );
not I_13161 (I226472,I226455);
nor I_13162 (I226489,I226130,I226472);
and I_13163 (I226506,I226393,I226489);
or I_13164 (I226523,I226113,I226506);
DFFARX1 I_13165  ( .D(I226523), .CLK(I2702), .RSTB(I226096), .Q(I226079) );
nor I_13166 (I226554,I226455,I226263);
nand I_13167 (I226088,I226229,I226554);
nor I_13168 (I226585,I226455,I226178);
nand I_13169 (I226082,I226328,I226585);
not I_13170 (I226085,I226455);
nand I_13171 (I226076,I226455,I226178);
DFFARX1 I_13172  ( .D(I226455), .CLK(I2702), .RSTB(I226096), .Q(I226067) );
not I_13173 (I226691,I2709);
or I_13174 (I226708,I104036,I104030);
or I_13175 (I226725,I104024,I104036);
DFFARX1 I_13176  ( .D(I226725), .CLK(I2702), .RSTB(I226691), .Q(I226665) );
nor I_13177 (I226756,I104042,I104033);
not I_13178 (I226773,I226756);
not I_13179 (I226790,I104042);
and I_13180 (I226807,I226790,I104039);
nor I_13181 (I226824,I226807,I104030);
nor I_13182 (I226841,I104015,I104021);
DFFARX1 I_13183  ( .D(I226841), .CLK(I2702), .RSTB(I226691), .Q(I226858) );
nand I_13184 (I226875,I226858,I226708);
and I_13185 (I226892,I226824,I226875);
DFFARX1 I_13186  ( .D(I226892), .CLK(I2702), .RSTB(I226691), .Q(I226659) );
nor I_13187 (I226923,I104015,I104024);
DFFARX1 I_13188  ( .D(I226923), .CLK(I2702), .RSTB(I226691), .Q(I226940) );
and I_13189 (I226656,I226756,I226940);
DFFARX1 I_13190  ( .D(I104027), .CLK(I2702), .RSTB(I226691), .Q(I226971) );
and I_13191 (I226988,I226971,I104045);
DFFARX1 I_13192  ( .D(I226988), .CLK(I2702), .RSTB(I226691), .Q(I227005) );
not I_13193 (I226668,I227005);
DFFARX1 I_13194  ( .D(I226988), .CLK(I2702), .RSTB(I226691), .Q(I226653) );
DFFARX1 I_13195  ( .D(I104018), .CLK(I2702), .RSTB(I226691), .Q(I227050) );
not I_13196 (I227067,I227050);
nor I_13197 (I227084,I226725,I227067);
and I_13198 (I227101,I226988,I227084);
or I_13199 (I227118,I226708,I227101);
DFFARX1 I_13200  ( .D(I227118), .CLK(I2702), .RSTB(I226691), .Q(I226674) );
nor I_13201 (I227149,I227050,I226858);
nand I_13202 (I226683,I226824,I227149);
nor I_13203 (I227180,I227050,I226773);
nand I_13204 (I226677,I226923,I227180);
not I_13205 (I226680,I227050);
nand I_13206 (I226671,I227050,I226773);
DFFARX1 I_13207  ( .D(I227050), .CLK(I2702), .RSTB(I226691), .Q(I226662) );
not I_13208 (I227286,I2709);
or I_13209 (I227303,I326511,I326526);
or I_13210 (I227320,I326514,I326511);
DFFARX1 I_13211  ( .D(I227320), .CLK(I2702), .RSTB(I227286), .Q(I227260) );
nor I_13212 (I227351,I326517,I326532);
not I_13213 (I227368,I227351);
not I_13214 (I227385,I326517);
and I_13215 (I227402,I227385,I326520);
nor I_13216 (I227419,I227402,I326526);
nor I_13217 (I227436,I326523,I326541);
DFFARX1 I_13218  ( .D(I227436), .CLK(I2702), .RSTB(I227286), .Q(I227453) );
nand I_13219 (I227470,I227453,I227303);
and I_13220 (I227487,I227419,I227470);
DFFARX1 I_13221  ( .D(I227487), .CLK(I2702), .RSTB(I227286), .Q(I227254) );
nor I_13222 (I227518,I326523,I326514);
DFFARX1 I_13223  ( .D(I227518), .CLK(I2702), .RSTB(I227286), .Q(I227535) );
and I_13224 (I227251,I227351,I227535);
DFFARX1 I_13225  ( .D(I326538), .CLK(I2702), .RSTB(I227286), .Q(I227566) );
and I_13226 (I227583,I227566,I326529);
DFFARX1 I_13227  ( .D(I227583), .CLK(I2702), .RSTB(I227286), .Q(I227600) );
not I_13228 (I227263,I227600);
DFFARX1 I_13229  ( .D(I227583), .CLK(I2702), .RSTB(I227286), .Q(I227248) );
DFFARX1 I_13230  ( .D(I326535), .CLK(I2702), .RSTB(I227286), .Q(I227645) );
not I_13231 (I227662,I227645);
nor I_13232 (I227679,I227320,I227662);
and I_13233 (I227696,I227583,I227679);
or I_13234 (I227713,I227303,I227696);
DFFARX1 I_13235  ( .D(I227713), .CLK(I2702), .RSTB(I227286), .Q(I227269) );
nor I_13236 (I227744,I227645,I227453);
nand I_13237 (I227278,I227419,I227744);
nor I_13238 (I227775,I227645,I227368);
nand I_13239 (I227272,I227518,I227775);
not I_13240 (I227275,I227645);
nand I_13241 (I227266,I227645,I227368);
DFFARX1 I_13242  ( .D(I227645), .CLK(I2702), .RSTB(I227286), .Q(I227257) );
not I_13243 (I227881,I2709);
or I_13244 (I227898,I135041,I135038);
not I_13245 (I227864,I227898);
DFFARX1 I_13246  ( .D(I227898), .CLK(I2702), .RSTB(I227881), .Q(I227843) );
or I_13247 (I227943,I135032,I135041);
nor I_13248 (I227960,I135050,I135023);
nor I_13249 (I227977,I227960,I227898);
not I_13250 (I227994,I135050);
and I_13251 (I228011,I227994,I135044);
nor I_13252 (I228028,I228011,I135038);
DFFARX1 I_13253  ( .D(I228028), .CLK(I2702), .RSTB(I227881), .Q(I228045) );
nor I_13254 (I228062,I135026,I135053);
DFFARX1 I_13255  ( .D(I228062), .CLK(I2702), .RSTB(I227881), .Q(I228079) );
nor I_13256 (I227870,I228079,I228028);
not I_13257 (I228110,I228079);
nor I_13258 (I228127,I135026,I135032);
nand I_13259 (I228144,I228028,I228127);
and I_13260 (I228161,I227943,I228144);
DFFARX1 I_13261  ( .D(I228161), .CLK(I2702), .RSTB(I227881), .Q(I227873) );
DFFARX1 I_13262  ( .D(I135029), .CLK(I2702), .RSTB(I227881), .Q(I228192) );
and I_13263 (I228209,I228192,I135035);
nor I_13264 (I228226,I228209,I228110);
and I_13265 (I228243,I228127,I228226);
or I_13266 (I228260,I227960,I228243);
DFFARX1 I_13267  ( .D(I228260), .CLK(I2702), .RSTB(I227881), .Q(I227858) );
not I_13268 (I228291,I228209);
nor I_13269 (I228308,I227898,I228291);
nand I_13270 (I227861,I227943,I228308);
nand I_13271 (I227855,I228079,I228291);
DFFARX1 I_13272  ( .D(I228209), .CLK(I2702), .RSTB(I227881), .Q(I227849) );
DFFARX1 I_13273  ( .D(I135047), .CLK(I2702), .RSTB(I227881), .Q(I228367) );
nand I_13274 (I227867,I228367,I227977);
DFFARX1 I_13275  ( .D(I228367), .CLK(I2702), .RSTB(I227881), .Q(I228398) );
not I_13276 (I227852,I228398);
and I_13277 (I227846,I228367,I228045);
not I_13278 (I228476,I2709);
or I_13279 (I228493,I193920,I193917);
not I_13280 (I228459,I228493);
DFFARX1 I_13281  ( .D(I228493), .CLK(I2702), .RSTB(I228476), .Q(I228438) );
or I_13282 (I228538,I193935,I193920);
nor I_13283 (I228555,I193926,I193911);
nor I_13284 (I228572,I228555,I228493);
not I_13285 (I228589,I193926);
and I_13286 (I228606,I228589,I193929);
nor I_13287 (I228623,I228606,I193917);
DFFARX1 I_13288  ( .D(I228623), .CLK(I2702), .RSTB(I228476), .Q(I228640) );
nor I_13289 (I228657,I193914,I193923);
DFFARX1 I_13290  ( .D(I228657), .CLK(I2702), .RSTB(I228476), .Q(I228674) );
nor I_13291 (I228465,I228674,I228623);
not I_13292 (I228705,I228674);
nor I_13293 (I228722,I193914,I193935);
nand I_13294 (I228739,I228623,I228722);
and I_13295 (I228756,I228538,I228739);
DFFARX1 I_13296  ( .D(I228756), .CLK(I2702), .RSTB(I228476), .Q(I228468) );
DFFARX1 I_13297  ( .D(I193932), .CLK(I2702), .RSTB(I228476), .Q(I228787) );
and I_13298 (I228804,I228787,I193941);
nor I_13299 (I228821,I228804,I228705);
and I_13300 (I228838,I228722,I228821);
or I_13301 (I228855,I228555,I228838);
DFFARX1 I_13302  ( .D(I228855), .CLK(I2702), .RSTB(I228476), .Q(I228453) );
not I_13303 (I228886,I228804);
nor I_13304 (I228903,I228493,I228886);
nand I_13305 (I228456,I228538,I228903);
nand I_13306 (I228450,I228674,I228886);
DFFARX1 I_13307  ( .D(I228804), .CLK(I2702), .RSTB(I228476), .Q(I228444) );
DFFARX1 I_13308  ( .D(I193938), .CLK(I2702), .RSTB(I228476), .Q(I228962) );
nand I_13309 (I228462,I228962,I228572);
DFFARX1 I_13310  ( .D(I228962), .CLK(I2702), .RSTB(I228476), .Q(I228993) );
not I_13311 (I228447,I228993);
and I_13312 (I228441,I228962,I228640);
not I_13313 (I229071,I2709);
or I_13314 (I229088,I189279,I189276);
not I_13315 (I229054,I229088);
DFFARX1 I_13316  ( .D(I229088), .CLK(I2702), .RSTB(I229071), .Q(I229033) );
or I_13317 (I229133,I189294,I189279);
nor I_13318 (I229150,I189285,I189270);
nor I_13319 (I229167,I229150,I229088);
not I_13320 (I229184,I189285);
and I_13321 (I229201,I229184,I189288);
nor I_13322 (I229218,I229201,I189276);
DFFARX1 I_13323  ( .D(I229218), .CLK(I2702), .RSTB(I229071), .Q(I229235) );
nor I_13324 (I229252,I189273,I189282);
DFFARX1 I_13325  ( .D(I229252), .CLK(I2702), .RSTB(I229071), .Q(I229269) );
nor I_13326 (I229060,I229269,I229218);
not I_13327 (I229300,I229269);
nor I_13328 (I229317,I189273,I189294);
nand I_13329 (I229334,I229218,I229317);
and I_13330 (I229351,I229133,I229334);
DFFARX1 I_13331  ( .D(I229351), .CLK(I2702), .RSTB(I229071), .Q(I229063) );
DFFARX1 I_13332  ( .D(I189291), .CLK(I2702), .RSTB(I229071), .Q(I229382) );
and I_13333 (I229399,I229382,I189300);
nor I_13334 (I229416,I229399,I229300);
and I_13335 (I229433,I229317,I229416);
or I_13336 (I229450,I229150,I229433);
DFFARX1 I_13337  ( .D(I229450), .CLK(I2702), .RSTB(I229071), .Q(I229048) );
not I_13338 (I229481,I229399);
nor I_13339 (I229498,I229088,I229481);
nand I_13340 (I229051,I229133,I229498);
nand I_13341 (I229045,I229269,I229481);
DFFARX1 I_13342  ( .D(I229399), .CLK(I2702), .RSTB(I229071), .Q(I229039) );
DFFARX1 I_13343  ( .D(I189297), .CLK(I2702), .RSTB(I229071), .Q(I229557) );
nand I_13344 (I229057,I229557,I229167);
DFFARX1 I_13345  ( .D(I229557), .CLK(I2702), .RSTB(I229071), .Q(I229588) );
not I_13346 (I229042,I229588);
and I_13347 (I229036,I229557,I229235);
not I_13348 (I229666,I2709);
or I_13349 (I229683,I2543,I2199);
not I_13350 (I229649,I229683);
DFFARX1 I_13351  ( .D(I229683), .CLK(I2702), .RSTB(I229666), .Q(I229628) );
or I_13352 (I229728,I1975,I2543);
nor I_13353 (I229745,I1231,I2239);
nor I_13354 (I229762,I229745,I229683);
not I_13355 (I229779,I1231);
and I_13356 (I229796,I229779,I1487);
nor I_13357 (I229813,I229796,I2199);
DFFARX1 I_13358  ( .D(I229813), .CLK(I2702), .RSTB(I229666), .Q(I229830) );
nor I_13359 (I229847,I2551,I2351);
DFFARX1 I_13360  ( .D(I229847), .CLK(I2702), .RSTB(I229666), .Q(I229864) );
nor I_13361 (I229655,I229864,I229813);
not I_13362 (I229895,I229864);
nor I_13363 (I229912,I2551,I1975);
nand I_13364 (I229929,I229813,I229912);
and I_13365 (I229946,I229728,I229929);
DFFARX1 I_13366  ( .D(I229946), .CLK(I2702), .RSTB(I229666), .Q(I229658) );
DFFARX1 I_13367  ( .D(I1479), .CLK(I2702), .RSTB(I229666), .Q(I229977) );
and I_13368 (I229994,I229977,I1959);
nor I_13369 (I230011,I229994,I229895);
and I_13370 (I230028,I229912,I230011);
or I_13371 (I230045,I229745,I230028);
DFFARX1 I_13372  ( .D(I230045), .CLK(I2702), .RSTB(I229666), .Q(I229643) );
not I_13373 (I230076,I229994);
nor I_13374 (I230093,I229683,I230076);
nand I_13375 (I229646,I229728,I230093);
nand I_13376 (I229640,I229864,I230076);
DFFARX1 I_13377  ( .D(I229994), .CLK(I2702), .RSTB(I229666), .Q(I229634) );
DFFARX1 I_13378  ( .D(I1359), .CLK(I2702), .RSTB(I229666), .Q(I230152) );
nand I_13379 (I229652,I230152,I229762);
DFFARX1 I_13380  ( .D(I230152), .CLK(I2702), .RSTB(I229666), .Q(I230183) );
not I_13381 (I229637,I230183);
and I_13382 (I229631,I230152,I229830);
not I_13383 (I230261,I2709);
or I_13384 (I230278,I645131,I645140);
not I_13385 (I230244,I230278);
DFFARX1 I_13386  ( .D(I230278), .CLK(I2702), .RSTB(I230261), .Q(I230223) );
or I_13387 (I230323,I645149,I645131);
nor I_13388 (I230340,I645143,I645137);
nor I_13389 (I230357,I230340,I230278);
not I_13390 (I230374,I645143);
and I_13391 (I230391,I230374,I645146);
nor I_13392 (I230408,I230391,I645140);
DFFARX1 I_13393  ( .D(I230408), .CLK(I2702), .RSTB(I230261), .Q(I230425) );
nor I_13394 (I230442,I645134,I645152);
DFFARX1 I_13395  ( .D(I230442), .CLK(I2702), .RSTB(I230261), .Q(I230459) );
nor I_13396 (I230250,I230459,I230408);
not I_13397 (I230490,I230459);
nor I_13398 (I230507,I645134,I645149);
nand I_13399 (I230524,I230408,I230507);
and I_13400 (I230541,I230323,I230524);
DFFARX1 I_13401  ( .D(I230541), .CLK(I2702), .RSTB(I230261), .Q(I230253) );
DFFARX1 I_13402  ( .D(I645155), .CLK(I2702), .RSTB(I230261), .Q(I230572) );
and I_13403 (I230589,I230572,I645128);
nor I_13404 (I230606,I230589,I230490);
and I_13405 (I230623,I230507,I230606);
or I_13406 (I230640,I230340,I230623);
DFFARX1 I_13407  ( .D(I230640), .CLK(I2702), .RSTB(I230261), .Q(I230238) );
not I_13408 (I230671,I230589);
nor I_13409 (I230688,I230278,I230671);
nand I_13410 (I230241,I230323,I230688);
nand I_13411 (I230235,I230459,I230671);
DFFARX1 I_13412  ( .D(I230589), .CLK(I2702), .RSTB(I230261), .Q(I230229) );
DFFARX1 I_13413  ( .D(I645125), .CLK(I2702), .RSTB(I230261), .Q(I230747) );
nand I_13414 (I230247,I230747,I230357);
DFFARX1 I_13415  ( .D(I230747), .CLK(I2702), .RSTB(I230261), .Q(I230778) );
not I_13416 (I230232,I230778);
and I_13417 (I230226,I230747,I230425);
not I_13418 (I230856,I2709);
or I_13419 (I230873,I380948,I380945);
not I_13420 (I230839,I230873);
DFFARX1 I_13421  ( .D(I230873), .CLK(I2702), .RSTB(I230856), .Q(I230818) );
or I_13422 (I230918,I380954,I380948);
nor I_13423 (I230935,I380969,I380960);
nor I_13424 (I230952,I230935,I230873);
not I_13425 (I230969,I380969);
and I_13426 (I230986,I230969,I380963);
nor I_13427 (I231003,I230986,I380945);
DFFARX1 I_13428  ( .D(I231003), .CLK(I2702), .RSTB(I230856), .Q(I231020) );
nor I_13429 (I231037,I380975,I380972);
DFFARX1 I_13430  ( .D(I231037), .CLK(I2702), .RSTB(I230856), .Q(I231054) );
nor I_13431 (I230845,I231054,I231003);
not I_13432 (I231085,I231054);
nor I_13433 (I231102,I380975,I380954);
nand I_13434 (I231119,I231003,I231102);
and I_13435 (I231136,I230918,I231119);
DFFARX1 I_13436  ( .D(I231136), .CLK(I2702), .RSTB(I230856), .Q(I230848) );
DFFARX1 I_13437  ( .D(I380951), .CLK(I2702), .RSTB(I230856), .Q(I231167) );
and I_13438 (I231184,I231167,I380966);
nor I_13439 (I231201,I231184,I231085);
and I_13440 (I231218,I231102,I231201);
or I_13441 (I231235,I230935,I231218);
DFFARX1 I_13442  ( .D(I231235), .CLK(I2702), .RSTB(I230856), .Q(I230833) );
not I_13443 (I231266,I231184);
nor I_13444 (I231283,I230873,I231266);
nand I_13445 (I230836,I230918,I231283);
nand I_13446 (I230830,I231054,I231266);
DFFARX1 I_13447  ( .D(I231184), .CLK(I2702), .RSTB(I230856), .Q(I230824) );
DFFARX1 I_13448  ( .D(I380957), .CLK(I2702), .RSTB(I230856), .Q(I231342) );
nand I_13449 (I230842,I231342,I230952);
DFFARX1 I_13450  ( .D(I231342), .CLK(I2702), .RSTB(I230856), .Q(I231373) );
not I_13451 (I230827,I231373);
and I_13452 (I230821,I231342,I231020);
not I_13453 (I231451,I2709);
or I_13454 (I231468,I684129,I684138);
not I_13455 (I231434,I231468);
DFFARX1 I_13456  ( .D(I231468), .CLK(I2702), .RSTB(I231451), .Q(I231413) );
or I_13457 (I231513,I684147,I684129);
nor I_13458 (I231530,I684141,I684135);
nor I_13459 (I231547,I231530,I231468);
not I_13460 (I231564,I684141);
and I_13461 (I231581,I231564,I684144);
nor I_13462 (I231598,I231581,I684138);
DFFARX1 I_13463  ( .D(I231598), .CLK(I2702), .RSTB(I231451), .Q(I231615) );
nor I_13464 (I231632,I684132,I684150);
DFFARX1 I_13465  ( .D(I231632), .CLK(I2702), .RSTB(I231451), .Q(I231649) );
nor I_13466 (I231440,I231649,I231598);
not I_13467 (I231680,I231649);
nor I_13468 (I231697,I684132,I684147);
nand I_13469 (I231714,I231598,I231697);
and I_13470 (I231731,I231513,I231714);
DFFARX1 I_13471  ( .D(I231731), .CLK(I2702), .RSTB(I231451), .Q(I231443) );
DFFARX1 I_13472  ( .D(I684153), .CLK(I2702), .RSTB(I231451), .Q(I231762) );
and I_13473 (I231779,I231762,I684126);
nor I_13474 (I231796,I231779,I231680);
and I_13475 (I231813,I231697,I231796);
or I_13476 (I231830,I231530,I231813);
DFFARX1 I_13477  ( .D(I231830), .CLK(I2702), .RSTB(I231451), .Q(I231428) );
not I_13478 (I231861,I231779);
nor I_13479 (I231878,I231468,I231861);
nand I_13480 (I231431,I231513,I231878);
nand I_13481 (I231425,I231649,I231861);
DFFARX1 I_13482  ( .D(I231779), .CLK(I2702), .RSTB(I231451), .Q(I231419) );
DFFARX1 I_13483  ( .D(I684123), .CLK(I2702), .RSTB(I231451), .Q(I231937) );
nand I_13484 (I231437,I231937,I231547);
DFFARX1 I_13485  ( .D(I231937), .CLK(I2702), .RSTB(I231451), .Q(I231968) );
not I_13486 (I231422,I231968);
and I_13487 (I231416,I231937,I231615);
not I_13488 (I232046,I2709);
or I_13489 (I232063,I548265,I548277);
not I_13490 (I232029,I232063);
DFFARX1 I_13491  ( .D(I232063), .CLK(I2702), .RSTB(I232046), .Q(I232008) );
or I_13492 (I232108,I548289,I548265);
nor I_13493 (I232125,I548283,I548268);
nor I_13494 (I232142,I232125,I232063);
not I_13495 (I232159,I548283);
and I_13496 (I232176,I232159,I548280);
nor I_13497 (I232193,I232176,I548277);
DFFARX1 I_13498  ( .D(I232193), .CLK(I2702), .RSTB(I232046), .Q(I232210) );
nor I_13499 (I232227,I548274,I548271);
DFFARX1 I_13500  ( .D(I232227), .CLK(I2702), .RSTB(I232046), .Q(I232244) );
nor I_13501 (I232035,I232244,I232193);
not I_13502 (I232275,I232244);
nor I_13503 (I232292,I548274,I548289);
nand I_13504 (I232309,I232193,I232292);
and I_13505 (I232326,I232108,I232309);
DFFARX1 I_13506  ( .D(I232326), .CLK(I2702), .RSTB(I232046), .Q(I232038) );
DFFARX1 I_13507  ( .D(I548286), .CLK(I2702), .RSTB(I232046), .Q(I232357) );
and I_13508 (I232374,I232357,I548259);
nor I_13509 (I232391,I232374,I232275);
and I_13510 (I232408,I232292,I232391);
or I_13511 (I232425,I232125,I232408);
DFFARX1 I_13512  ( .D(I232425), .CLK(I2702), .RSTB(I232046), .Q(I232023) );
not I_13513 (I232456,I232374);
nor I_13514 (I232473,I232063,I232456);
nand I_13515 (I232026,I232108,I232473);
nand I_13516 (I232020,I232244,I232456);
DFFARX1 I_13517  ( .D(I232374), .CLK(I2702), .RSTB(I232046), .Q(I232014) );
DFFARX1 I_13518  ( .D(I548262), .CLK(I2702), .RSTB(I232046), .Q(I232532) );
nand I_13519 (I232032,I232532,I232142);
DFFARX1 I_13520  ( .D(I232532), .CLK(I2702), .RSTB(I232046), .Q(I232563) );
not I_13521 (I232017,I232563);
and I_13522 (I232011,I232532,I232210);
not I_13523 (I232641,I2709);
or I_13524 (I232658,I468529,I468559);
not I_13525 (I232624,I232658);
DFFARX1 I_13526  ( .D(I232658), .CLK(I2702), .RSTB(I232641), .Q(I232603) );
or I_13527 (I232703,I468538,I468529);
nor I_13528 (I232720,I468544,I468541);
nor I_13529 (I232737,I232720,I232658);
not I_13530 (I232754,I468544);
and I_13531 (I232771,I232754,I468550);
nor I_13532 (I232788,I232771,I468559);
DFFARX1 I_13533  ( .D(I232788), .CLK(I2702), .RSTB(I232641), .Q(I232805) );
nor I_13534 (I232822,I468535,I468553);
DFFARX1 I_13535  ( .D(I232822), .CLK(I2702), .RSTB(I232641), .Q(I232839) );
nor I_13536 (I232630,I232839,I232788);
not I_13537 (I232870,I232839);
nor I_13538 (I232887,I468535,I468538);
nand I_13539 (I232904,I232788,I232887);
and I_13540 (I232921,I232703,I232904);
DFFARX1 I_13541  ( .D(I232921), .CLK(I2702), .RSTB(I232641), .Q(I232633) );
DFFARX1 I_13542  ( .D(I468556), .CLK(I2702), .RSTB(I232641), .Q(I232952) );
and I_13543 (I232969,I232952,I468547);
nor I_13544 (I232986,I232969,I232870);
and I_13545 (I233003,I232887,I232986);
or I_13546 (I233020,I232720,I233003);
DFFARX1 I_13547  ( .D(I233020), .CLK(I2702), .RSTB(I232641), .Q(I232618) );
not I_13548 (I233051,I232969);
nor I_13549 (I233068,I232658,I233051);
nand I_13550 (I232621,I232703,I233068);
nand I_13551 (I232615,I232839,I233051);
DFFARX1 I_13552  ( .D(I232969), .CLK(I2702), .RSTB(I232641), .Q(I232609) );
DFFARX1 I_13553  ( .D(I468532), .CLK(I2702), .RSTB(I232641), .Q(I233127) );
nand I_13554 (I232627,I233127,I232737);
DFFARX1 I_13555  ( .D(I233127), .CLK(I2702), .RSTB(I232641), .Q(I233158) );
not I_13556 (I232612,I233158);
and I_13557 (I232606,I233127,I232805);
not I_13558 (I233236,I2709);
or I_13559 (I233253,I222500,I222497);
not I_13560 (I233219,I233253);
DFFARX1 I_13561  ( .D(I233253), .CLK(I2702), .RSTB(I233236), .Q(I233198) );
or I_13562 (I233298,I222488,I222500);
nor I_13563 (I233315,I222515,I222494);
nor I_13564 (I233332,I233315,I233253);
not I_13565 (I233349,I222515);
and I_13566 (I233366,I233349,I222503);
nor I_13567 (I233383,I233366,I222497);
DFFARX1 I_13568  ( .D(I233383), .CLK(I2702), .RSTB(I233236), .Q(I233400) );
nor I_13569 (I233417,I222491,I222509);
DFFARX1 I_13570  ( .D(I233417), .CLK(I2702), .RSTB(I233236), .Q(I233434) );
nor I_13571 (I233225,I233434,I233383);
not I_13572 (I233465,I233434);
nor I_13573 (I233482,I222491,I222488);
nand I_13574 (I233499,I233383,I233482);
and I_13575 (I233516,I233298,I233499);
DFFARX1 I_13576  ( .D(I233516), .CLK(I2702), .RSTB(I233236), .Q(I233228) );
DFFARX1 I_13577  ( .D(I222506), .CLK(I2702), .RSTB(I233236), .Q(I233547) );
and I_13578 (I233564,I233547,I222518);
nor I_13579 (I233581,I233564,I233465);
and I_13580 (I233598,I233482,I233581);
or I_13581 (I233615,I233315,I233598);
DFFARX1 I_13582  ( .D(I233615), .CLK(I2702), .RSTB(I233236), .Q(I233213) );
not I_13583 (I233646,I233564);
nor I_13584 (I233663,I233253,I233646);
nand I_13585 (I233216,I233298,I233663);
nand I_13586 (I233210,I233434,I233646);
DFFARX1 I_13587  ( .D(I233564), .CLK(I2702), .RSTB(I233236), .Q(I233204) );
DFFARX1 I_13588  ( .D(I222512), .CLK(I2702), .RSTB(I233236), .Q(I233722) );
nand I_13589 (I233222,I233722,I233332);
DFFARX1 I_13590  ( .D(I233722), .CLK(I2702), .RSTB(I233236), .Q(I233753) );
not I_13591 (I233207,I233753);
and I_13592 (I233201,I233722,I233400);
not I_13593 (I233831,I2709);
or I_13594 (I233848,I105971,I105968);
not I_13595 (I233814,I233848);
DFFARX1 I_13596  ( .D(I233848), .CLK(I2702), .RSTB(I233831), .Q(I233793) );
or I_13597 (I233893,I105962,I105971);
nor I_13598 (I233910,I105980,I105953);
nor I_13599 (I233927,I233910,I233848);
not I_13600 (I233944,I105980);
and I_13601 (I233961,I233944,I105974);
nor I_13602 (I233978,I233961,I105968);
DFFARX1 I_13603  ( .D(I233978), .CLK(I2702), .RSTB(I233831), .Q(I233995) );
nor I_13604 (I234012,I105956,I105983);
DFFARX1 I_13605  ( .D(I234012), .CLK(I2702), .RSTB(I233831), .Q(I234029) );
nor I_13606 (I233820,I234029,I233978);
not I_13607 (I234060,I234029);
nor I_13608 (I234077,I105956,I105962);
nand I_13609 (I234094,I233978,I234077);
and I_13610 (I234111,I233893,I234094);
DFFARX1 I_13611  ( .D(I234111), .CLK(I2702), .RSTB(I233831), .Q(I233823) );
DFFARX1 I_13612  ( .D(I105959), .CLK(I2702), .RSTB(I233831), .Q(I234142) );
and I_13613 (I234159,I234142,I105965);
nor I_13614 (I234176,I234159,I234060);
and I_13615 (I234193,I234077,I234176);
or I_13616 (I234210,I233910,I234193);
DFFARX1 I_13617  ( .D(I234210), .CLK(I2702), .RSTB(I233831), .Q(I233808) );
not I_13618 (I234241,I234159);
nor I_13619 (I234258,I233848,I234241);
nand I_13620 (I233811,I233893,I234258);
nand I_13621 (I233805,I234029,I234241);
DFFARX1 I_13622  ( .D(I234159), .CLK(I2702), .RSTB(I233831), .Q(I233799) );
DFFARX1 I_13623  ( .D(I105977), .CLK(I2702), .RSTB(I233831), .Q(I234317) );
nand I_13624 (I233817,I234317,I233927);
DFFARX1 I_13625  ( .D(I234317), .CLK(I2702), .RSTB(I233831), .Q(I234348) );
not I_13626 (I233802,I234348);
and I_13627 (I233796,I234317,I233995);
not I_13628 (I234426,I2709);
or I_13629 (I234443,I643873,I643882);
not I_13630 (I234409,I234443);
DFFARX1 I_13631  ( .D(I234443), .CLK(I2702), .RSTB(I234426), .Q(I234388) );
or I_13632 (I234488,I643891,I643873);
nor I_13633 (I234505,I643885,I643879);
nor I_13634 (I234522,I234505,I234443);
not I_13635 (I234539,I643885);
and I_13636 (I234556,I234539,I643888);
nor I_13637 (I234573,I234556,I643882);
DFFARX1 I_13638  ( .D(I234573), .CLK(I2702), .RSTB(I234426), .Q(I234590) );
nor I_13639 (I234607,I643876,I643894);
DFFARX1 I_13640  ( .D(I234607), .CLK(I2702), .RSTB(I234426), .Q(I234624) );
nor I_13641 (I234415,I234624,I234573);
not I_13642 (I234655,I234624);
nor I_13643 (I234672,I643876,I643891);
nand I_13644 (I234689,I234573,I234672);
and I_13645 (I234706,I234488,I234689);
DFFARX1 I_13646  ( .D(I234706), .CLK(I2702), .RSTB(I234426), .Q(I234418) );
DFFARX1 I_13647  ( .D(I643897), .CLK(I2702), .RSTB(I234426), .Q(I234737) );
and I_13648 (I234754,I234737,I643870);
nor I_13649 (I234771,I234754,I234655);
and I_13650 (I234788,I234672,I234771);
or I_13651 (I234805,I234505,I234788);
DFFARX1 I_13652  ( .D(I234805), .CLK(I2702), .RSTB(I234426), .Q(I234403) );
not I_13653 (I234836,I234754);
nor I_13654 (I234853,I234443,I234836);
nand I_13655 (I234406,I234488,I234853);
nand I_13656 (I234400,I234624,I234836);
DFFARX1 I_13657  ( .D(I234754), .CLK(I2702), .RSTB(I234426), .Q(I234394) );
DFFARX1 I_13658  ( .D(I643867), .CLK(I2702), .RSTB(I234426), .Q(I234912) );
nand I_13659 (I234412,I234912,I234522);
DFFARX1 I_13660  ( .D(I234912), .CLK(I2702), .RSTB(I234426), .Q(I234943) );
not I_13661 (I234397,I234943);
and I_13662 (I234391,I234912,I234590);
not I_13663 (I235021,I2709);
or I_13664 (I235038,I384178,I384175);
not I_13665 (I235004,I235038);
DFFARX1 I_13666  ( .D(I235038), .CLK(I2702), .RSTB(I235021), .Q(I234983) );
or I_13667 (I235083,I384184,I384178);
nor I_13668 (I235100,I384199,I384190);
nor I_13669 (I235117,I235100,I235038);
not I_13670 (I235134,I384199);
and I_13671 (I235151,I235134,I384193);
nor I_13672 (I235168,I235151,I384175);
DFFARX1 I_13673  ( .D(I235168), .CLK(I2702), .RSTB(I235021), .Q(I235185) );
nor I_13674 (I235202,I384205,I384202);
DFFARX1 I_13675  ( .D(I235202), .CLK(I2702), .RSTB(I235021), .Q(I235219) );
nor I_13676 (I235010,I235219,I235168);
not I_13677 (I235250,I235219);
nor I_13678 (I235267,I384205,I384184);
nand I_13679 (I235284,I235168,I235267);
and I_13680 (I235301,I235083,I235284);
DFFARX1 I_13681  ( .D(I235301), .CLK(I2702), .RSTB(I235021), .Q(I235013) );
DFFARX1 I_13682  ( .D(I384181), .CLK(I2702), .RSTB(I235021), .Q(I235332) );
and I_13683 (I235349,I235332,I384196);
nor I_13684 (I235366,I235349,I235250);
and I_13685 (I235383,I235267,I235366);
or I_13686 (I235400,I235100,I235383);
DFFARX1 I_13687  ( .D(I235400), .CLK(I2702), .RSTB(I235021), .Q(I234998) );
not I_13688 (I235431,I235349);
nor I_13689 (I235448,I235038,I235431);
nand I_13690 (I235001,I235083,I235448);
nand I_13691 (I234995,I235219,I235431);
DFFARX1 I_13692  ( .D(I235349), .CLK(I2702), .RSTB(I235021), .Q(I234989) );
DFFARX1 I_13693  ( .D(I384187), .CLK(I2702), .RSTB(I235021), .Q(I235507) );
nand I_13694 (I235007,I235507,I235117);
DFFARX1 I_13695  ( .D(I235507), .CLK(I2702), .RSTB(I235021), .Q(I235538) );
not I_13696 (I234992,I235538);
and I_13697 (I234986,I235507,I235185);
not I_13698 (I235616,I2709);
or I_13699 (I235633,I598245,I598239);
not I_13700 (I235599,I235633);
DFFARX1 I_13701  ( .D(I235633), .CLK(I2702), .RSTB(I235616), .Q(I235578) );
or I_13702 (I235678,I598266,I598245);
nor I_13703 (I235695,I598269,I598254);
nor I_13704 (I235712,I235695,I235633);
not I_13705 (I235729,I598269);
and I_13706 (I235746,I235729,I598263);
nor I_13707 (I235763,I235746,I598239);
DFFARX1 I_13708  ( .D(I235763), .CLK(I2702), .RSTB(I235616), .Q(I235780) );
nor I_13709 (I235797,I598248,I598251);
DFFARX1 I_13710  ( .D(I235797), .CLK(I2702), .RSTB(I235616), .Q(I235814) );
nor I_13711 (I235605,I235814,I235763);
not I_13712 (I235845,I235814);
nor I_13713 (I235862,I598248,I598266);
nand I_13714 (I235879,I235763,I235862);
and I_13715 (I235896,I235678,I235879);
DFFARX1 I_13716  ( .D(I235896), .CLK(I2702), .RSTB(I235616), .Q(I235608) );
DFFARX1 I_13717  ( .D(I598260), .CLK(I2702), .RSTB(I235616), .Q(I235927) );
and I_13718 (I235944,I235927,I598242);
nor I_13719 (I235961,I235944,I235845);
and I_13720 (I235978,I235862,I235961);
or I_13721 (I235995,I235695,I235978);
DFFARX1 I_13722  ( .D(I235995), .CLK(I2702), .RSTB(I235616), .Q(I235593) );
not I_13723 (I236026,I235944);
nor I_13724 (I236043,I235633,I236026);
nand I_13725 (I235596,I235678,I236043);
nand I_13726 (I235590,I235814,I236026);
DFFARX1 I_13727  ( .D(I235944), .CLK(I2702), .RSTB(I235616), .Q(I235584) );
DFFARX1 I_13728  ( .D(I598257), .CLK(I2702), .RSTB(I235616), .Q(I236102) );
nand I_13729 (I235602,I236102,I235712);
DFFARX1 I_13730  ( .D(I236102), .CLK(I2702), .RSTB(I235616), .Q(I236133) );
not I_13731 (I235587,I236133);
and I_13732 (I235581,I236102,I235780);
not I_13733 (I236211,I2709);
or I_13734 (I236228,I572660,I572672);
not I_13735 (I236194,I236228);
DFFARX1 I_13736  ( .D(I236228), .CLK(I2702), .RSTB(I236211), .Q(I236173) );
or I_13737 (I236273,I572684,I572660);
nor I_13738 (I236290,I572678,I572663);
nor I_13739 (I236307,I236290,I236228);
not I_13740 (I236324,I572678);
and I_13741 (I236341,I236324,I572675);
nor I_13742 (I236358,I236341,I572672);
DFFARX1 I_13743  ( .D(I236358), .CLK(I2702), .RSTB(I236211), .Q(I236375) );
nor I_13744 (I236392,I572669,I572666);
DFFARX1 I_13745  ( .D(I236392), .CLK(I2702), .RSTB(I236211), .Q(I236409) );
nor I_13746 (I236200,I236409,I236358);
not I_13747 (I236440,I236409);
nor I_13748 (I236457,I572669,I572684);
nand I_13749 (I236474,I236358,I236457);
and I_13750 (I236491,I236273,I236474);
DFFARX1 I_13751  ( .D(I236491), .CLK(I2702), .RSTB(I236211), .Q(I236203) );
DFFARX1 I_13752  ( .D(I572681), .CLK(I2702), .RSTB(I236211), .Q(I236522) );
and I_13753 (I236539,I236522,I572654);
nor I_13754 (I236556,I236539,I236440);
and I_13755 (I236573,I236457,I236556);
or I_13756 (I236590,I236290,I236573);
DFFARX1 I_13757  ( .D(I236590), .CLK(I2702), .RSTB(I236211), .Q(I236188) );
not I_13758 (I236621,I236539);
nor I_13759 (I236638,I236228,I236621);
nand I_13760 (I236191,I236273,I236638);
nand I_13761 (I236185,I236409,I236621);
DFFARX1 I_13762  ( .D(I236539), .CLK(I2702), .RSTB(I236211), .Q(I236179) );
DFFARX1 I_13763  ( .D(I572657), .CLK(I2702), .RSTB(I236211), .Q(I236697) );
nand I_13764 (I236197,I236697,I236307);
DFFARX1 I_13765  ( .D(I236697), .CLK(I2702), .RSTB(I236211), .Q(I236728) );
not I_13766 (I236182,I236728);
and I_13767 (I236176,I236697,I236375);
not I_13768 (I236806,I2709);
or I_13769 (I236823,I259563,I259551);
not I_13770 (I236789,I236823);
DFFARX1 I_13771  ( .D(I236823), .CLK(I2702), .RSTB(I236806), .Q(I236768) );
or I_13772 (I236868,I259548,I259563);
nor I_13773 (I236885,I259578,I259569);
nor I_13774 (I236902,I236885,I236823);
not I_13775 (I236919,I259578);
and I_13776 (I236936,I236919,I259557);
nor I_13777 (I236953,I236936,I259551);
DFFARX1 I_13778  ( .D(I236953), .CLK(I2702), .RSTB(I236806), .Q(I236970) );
nor I_13779 (I236987,I259560,I259554);
DFFARX1 I_13780  ( .D(I236987), .CLK(I2702), .RSTB(I236806), .Q(I237004) );
nor I_13781 (I236795,I237004,I236953);
not I_13782 (I237035,I237004);
nor I_13783 (I237052,I259560,I259548);
nand I_13784 (I237069,I236953,I237052);
and I_13785 (I237086,I236868,I237069);
DFFARX1 I_13786  ( .D(I237086), .CLK(I2702), .RSTB(I236806), .Q(I236798) );
DFFARX1 I_13787  ( .D(I259575), .CLK(I2702), .RSTB(I236806), .Q(I237117) );
and I_13788 (I237134,I237117,I259572);
nor I_13789 (I237151,I237134,I237035);
and I_13790 (I237168,I237052,I237151);
or I_13791 (I237185,I236885,I237168);
DFFARX1 I_13792  ( .D(I237185), .CLK(I2702), .RSTB(I236806), .Q(I236783) );
not I_13793 (I237216,I237134);
nor I_13794 (I237233,I236823,I237216);
nand I_13795 (I236786,I236868,I237233);
nand I_13796 (I236780,I237004,I237216);
DFFARX1 I_13797  ( .D(I237134), .CLK(I2702), .RSTB(I236806), .Q(I236774) );
DFFARX1 I_13798  ( .D(I259566), .CLK(I2702), .RSTB(I236806), .Q(I237292) );
nand I_13799 (I236792,I237292,I236902);
DFFARX1 I_13800  ( .D(I237292), .CLK(I2702), .RSTB(I236806), .Q(I237323) );
not I_13801 (I236777,I237323);
and I_13802 (I236771,I237292,I236970);
not I_13803 (I237401,I2709);
or I_13804 (I237418,I522085,I522097);
not I_13805 (I237384,I237418);
DFFARX1 I_13806  ( .D(I237418), .CLK(I2702), .RSTB(I237401), .Q(I237363) );
or I_13807 (I237463,I522109,I522085);
nor I_13808 (I237480,I522103,I522088);
nor I_13809 (I237497,I237480,I237418);
not I_13810 (I237514,I522103);
and I_13811 (I237531,I237514,I522100);
nor I_13812 (I237548,I237531,I522097);
DFFARX1 I_13813  ( .D(I237548), .CLK(I2702), .RSTB(I237401), .Q(I237565) );
nor I_13814 (I237582,I522094,I522091);
DFFARX1 I_13815  ( .D(I237582), .CLK(I2702), .RSTB(I237401), .Q(I237599) );
nor I_13816 (I237390,I237599,I237548);
not I_13817 (I237630,I237599);
nor I_13818 (I237647,I522094,I522109);
nand I_13819 (I237664,I237548,I237647);
and I_13820 (I237681,I237463,I237664);
DFFARX1 I_13821  ( .D(I237681), .CLK(I2702), .RSTB(I237401), .Q(I237393) );
DFFARX1 I_13822  ( .D(I522106), .CLK(I2702), .RSTB(I237401), .Q(I237712) );
and I_13823 (I237729,I237712,I522079);
nor I_13824 (I237746,I237729,I237630);
and I_13825 (I237763,I237647,I237746);
or I_13826 (I237780,I237480,I237763);
DFFARX1 I_13827  ( .D(I237780), .CLK(I2702), .RSTB(I237401), .Q(I237378) );
not I_13828 (I237811,I237729);
nor I_13829 (I237828,I237418,I237811);
nand I_13830 (I237381,I237463,I237828);
nand I_13831 (I237375,I237599,I237811);
DFFARX1 I_13832  ( .D(I237729), .CLK(I2702), .RSTB(I237401), .Q(I237369) );
DFFARX1 I_13833  ( .D(I522082), .CLK(I2702), .RSTB(I237401), .Q(I237887) );
nand I_13834 (I237387,I237887,I237497);
DFFARX1 I_13835  ( .D(I237887), .CLK(I2702), .RSTB(I237401), .Q(I237918) );
not I_13836 (I237372,I237918);
and I_13837 (I237366,I237887,I237565);
not I_13838 (I237996,I2709);
or I_13839 (I238013,I509590,I509602);
not I_13840 (I237979,I238013);
DFFARX1 I_13841  ( .D(I238013), .CLK(I2702), .RSTB(I237996), .Q(I237958) );
or I_13842 (I238058,I509614,I509590);
nor I_13843 (I238075,I509608,I509593);
nor I_13844 (I238092,I238075,I238013);
not I_13845 (I238109,I509608);
and I_13846 (I238126,I238109,I509605);
nor I_13847 (I238143,I238126,I509602);
DFFARX1 I_13848  ( .D(I238143), .CLK(I2702), .RSTB(I237996), .Q(I238160) );
nor I_13849 (I238177,I509599,I509596);
DFFARX1 I_13850  ( .D(I238177), .CLK(I2702), .RSTB(I237996), .Q(I238194) );
nor I_13851 (I237985,I238194,I238143);
not I_13852 (I238225,I238194);
nor I_13853 (I238242,I509599,I509614);
nand I_13854 (I238259,I238143,I238242);
and I_13855 (I238276,I238058,I238259);
DFFARX1 I_13856  ( .D(I238276), .CLK(I2702), .RSTB(I237996), .Q(I237988) );
DFFARX1 I_13857  ( .D(I509611), .CLK(I2702), .RSTB(I237996), .Q(I238307) );
and I_13858 (I238324,I238307,I509584);
nor I_13859 (I238341,I238324,I238225);
and I_13860 (I238358,I238242,I238341);
or I_13861 (I238375,I238075,I238358);
DFFARX1 I_13862  ( .D(I238375), .CLK(I2702), .RSTB(I237996), .Q(I237973) );
not I_13863 (I238406,I238324);
nor I_13864 (I238423,I238013,I238406);
nand I_13865 (I237976,I238058,I238423);
nand I_13866 (I237970,I238194,I238406);
DFFARX1 I_13867  ( .D(I238324), .CLK(I2702), .RSTB(I237996), .Q(I237964) );
DFFARX1 I_13868  ( .D(I509587), .CLK(I2702), .RSTB(I237996), .Q(I238482) );
nand I_13869 (I237982,I238482,I238092);
DFFARX1 I_13870  ( .D(I238482), .CLK(I2702), .RSTB(I237996), .Q(I238513) );
not I_13871 (I237967,I238513);
and I_13872 (I237961,I238482,I238160);
not I_13873 (I238591,I2709);
or I_13874 (I238608,I580395,I580389);
not I_13875 (I238574,I238608);
DFFARX1 I_13876  ( .D(I238608), .CLK(I2702), .RSTB(I238591), .Q(I238553) );
or I_13877 (I238653,I580416,I580395);
nor I_13878 (I238670,I580419,I580404);
nor I_13879 (I238687,I238670,I238608);
not I_13880 (I238704,I580419);
and I_13881 (I238721,I238704,I580413);
nor I_13882 (I238738,I238721,I580389);
DFFARX1 I_13883  ( .D(I238738), .CLK(I2702), .RSTB(I238591), .Q(I238755) );
nor I_13884 (I238772,I580398,I580401);
DFFARX1 I_13885  ( .D(I238772), .CLK(I2702), .RSTB(I238591), .Q(I238789) );
nor I_13886 (I238580,I238789,I238738);
not I_13887 (I238820,I238789);
nor I_13888 (I238837,I580398,I580416);
nand I_13889 (I238854,I238738,I238837);
and I_13890 (I238871,I238653,I238854);
DFFARX1 I_13891  ( .D(I238871), .CLK(I2702), .RSTB(I238591), .Q(I238583) );
DFFARX1 I_13892  ( .D(I580410), .CLK(I2702), .RSTB(I238591), .Q(I238902) );
and I_13893 (I238919,I238902,I580392);
nor I_13894 (I238936,I238919,I238820);
and I_13895 (I238953,I238837,I238936);
or I_13896 (I238970,I238670,I238953);
DFFARX1 I_13897  ( .D(I238970), .CLK(I2702), .RSTB(I238591), .Q(I238568) );
not I_13898 (I239001,I238919);
nor I_13899 (I239018,I238608,I239001);
nand I_13900 (I238571,I238653,I239018);
nand I_13901 (I238565,I238789,I239001);
DFFARX1 I_13902  ( .D(I238919), .CLK(I2702), .RSTB(I238591), .Q(I238559) );
DFFARX1 I_13903  ( .D(I580407), .CLK(I2702), .RSTB(I238591), .Q(I239077) );
nand I_13904 (I238577,I239077,I238687);
DFFARX1 I_13905  ( .D(I239077), .CLK(I2702), .RSTB(I238591), .Q(I239108) );
not I_13906 (I238562,I239108);
and I_13907 (I238556,I239077,I238755);
not I_13908 (I239186,I2709);
or I_13909 (I239203,I107909,I107906);
not I_13910 (I239169,I239203);
DFFARX1 I_13911  ( .D(I239203), .CLK(I2702), .RSTB(I239186), .Q(I239148) );
or I_13912 (I239248,I107900,I107909);
nor I_13913 (I239265,I107918,I107891);
nor I_13914 (I239282,I239265,I239203);
not I_13915 (I239299,I107918);
and I_13916 (I239316,I239299,I107912);
nor I_13917 (I239333,I239316,I107906);
DFFARX1 I_13918  ( .D(I239333), .CLK(I2702), .RSTB(I239186), .Q(I239350) );
nor I_13919 (I239367,I107894,I107921);
DFFARX1 I_13920  ( .D(I239367), .CLK(I2702), .RSTB(I239186), .Q(I239384) );
nor I_13921 (I239175,I239384,I239333);
not I_13922 (I239415,I239384);
nor I_13923 (I239432,I107894,I107900);
nand I_13924 (I239449,I239333,I239432);
and I_13925 (I239466,I239248,I239449);
DFFARX1 I_13926  ( .D(I239466), .CLK(I2702), .RSTB(I239186), .Q(I239178) );
DFFARX1 I_13927  ( .D(I107897), .CLK(I2702), .RSTB(I239186), .Q(I239497) );
and I_13928 (I239514,I239497,I107903);
nor I_13929 (I239531,I239514,I239415);
and I_13930 (I239548,I239432,I239531);
or I_13931 (I239565,I239265,I239548);
DFFARX1 I_13932  ( .D(I239565), .CLK(I2702), .RSTB(I239186), .Q(I239163) );
not I_13933 (I239596,I239514);
nor I_13934 (I239613,I239203,I239596);
nand I_13935 (I239166,I239248,I239613);
nand I_13936 (I239160,I239384,I239596);
DFFARX1 I_13937  ( .D(I239514), .CLK(I2702), .RSTB(I239186), .Q(I239154) );
DFFARX1 I_13938  ( .D(I107915), .CLK(I2702), .RSTB(I239186), .Q(I239672) );
nand I_13939 (I239172,I239672,I239282);
DFFARX1 I_13940  ( .D(I239672), .CLK(I2702), .RSTB(I239186), .Q(I239703) );
not I_13941 (I239157,I239703);
and I_13942 (I239151,I239672,I239350);
not I_13943 (I239781,I2709);
or I_13944 (I239798,I205840,I205837);
not I_13945 (I239764,I239798);
DFFARX1 I_13946  ( .D(I239798), .CLK(I2702), .RSTB(I239781), .Q(I239743) );
or I_13947 (I239843,I205828,I205840);
nor I_13948 (I239860,I205855,I205834);
nor I_13949 (I239877,I239860,I239798);
not I_13950 (I239894,I205855);
and I_13951 (I239911,I239894,I205843);
nor I_13952 (I239928,I239911,I205837);
DFFARX1 I_13953  ( .D(I239928), .CLK(I2702), .RSTB(I239781), .Q(I239945) );
nor I_13954 (I239962,I205831,I205849);
DFFARX1 I_13955  ( .D(I239962), .CLK(I2702), .RSTB(I239781), .Q(I239979) );
nor I_13956 (I239770,I239979,I239928);
not I_13957 (I240010,I239979);
nor I_13958 (I240027,I205831,I205828);
nand I_13959 (I240044,I239928,I240027);
and I_13960 (I240061,I239843,I240044);
DFFARX1 I_13961  ( .D(I240061), .CLK(I2702), .RSTB(I239781), .Q(I239773) );
DFFARX1 I_13962  ( .D(I205846), .CLK(I2702), .RSTB(I239781), .Q(I240092) );
and I_13963 (I240109,I240092,I205858);
nor I_13964 (I240126,I240109,I240010);
and I_13965 (I240143,I240027,I240126);
or I_13966 (I240160,I239860,I240143);
DFFARX1 I_13967  ( .D(I240160), .CLK(I2702), .RSTB(I239781), .Q(I239758) );
not I_13968 (I240191,I240109);
nor I_13969 (I240208,I239798,I240191);
nand I_13970 (I239761,I239843,I240208);
nand I_13971 (I239755,I239979,I240191);
DFFARX1 I_13972  ( .D(I240109), .CLK(I2702), .RSTB(I239781), .Q(I239749) );
DFFARX1 I_13973  ( .D(I205852), .CLK(I2702), .RSTB(I239781), .Q(I240267) );
nand I_13974 (I239767,I240267,I239877);
DFFARX1 I_13975  ( .D(I240267), .CLK(I2702), .RSTB(I239781), .Q(I240298) );
not I_13976 (I239752,I240298);
and I_13977 (I239746,I240267,I239945);
not I_13978 (I240376,I2709);
or I_13979 (I240393,I703099,I703081);
not I_13980 (I240359,I240393);
DFFARX1 I_13981  ( .D(I240393), .CLK(I2702), .RSTB(I240376), .Q(I240338) );
or I_13982 (I240438,I703108,I703099);
nor I_13983 (I240455,I703090,I703105);
nor I_13984 (I240472,I240455,I240393);
not I_13985 (I240489,I703090);
and I_13986 (I240506,I240489,I703087);
nor I_13987 (I240523,I240506,I703081);
DFFARX1 I_13988  ( .D(I240523), .CLK(I2702), .RSTB(I240376), .Q(I240540) );
nor I_13989 (I240557,I703102,I703078);
DFFARX1 I_13990  ( .D(I240557), .CLK(I2702), .RSTB(I240376), .Q(I240574) );
nor I_13991 (I240365,I240574,I240523);
not I_13992 (I240605,I240574);
nor I_13993 (I240622,I703102,I703108);
nand I_13994 (I240639,I240523,I240622);
and I_13995 (I240656,I240438,I240639);
DFFARX1 I_13996  ( .D(I240656), .CLK(I2702), .RSTB(I240376), .Q(I240368) );
DFFARX1 I_13997  ( .D(I703096), .CLK(I2702), .RSTB(I240376), .Q(I240687) );
and I_13998 (I240704,I240687,I703084);
nor I_13999 (I240721,I240704,I240605);
and I_14000 (I240738,I240622,I240721);
or I_14001 (I240755,I240455,I240738);
DFFARX1 I_14002  ( .D(I240755), .CLK(I2702), .RSTB(I240376), .Q(I240353) );
not I_14003 (I240786,I240704);
nor I_14004 (I240803,I240393,I240786);
nand I_14005 (I240356,I240438,I240803);
nand I_14006 (I240350,I240574,I240786);
DFFARX1 I_14007  ( .D(I240704), .CLK(I2702), .RSTB(I240376), .Q(I240344) );
DFFARX1 I_14008  ( .D(I703093), .CLK(I2702), .RSTB(I240376), .Q(I240862) );
nand I_14009 (I240362,I240862,I240472);
DFFARX1 I_14010  ( .D(I240862), .CLK(I2702), .RSTB(I240376), .Q(I240893) );
not I_14011 (I240347,I240893);
and I_14012 (I240341,I240862,I240540);
not I_14013 (I240971,I2709);
or I_14014 (I240988,I69149,I69146);
not I_14015 (I240954,I240988);
DFFARX1 I_14016  ( .D(I240988), .CLK(I2702), .RSTB(I240971), .Q(I240933) );
or I_14017 (I241033,I69140,I69149);
nor I_14018 (I241050,I69158,I69131);
nor I_14019 (I241067,I241050,I240988);
not I_14020 (I241084,I69158);
and I_14021 (I241101,I241084,I69152);
nor I_14022 (I241118,I241101,I69146);
DFFARX1 I_14023  ( .D(I241118), .CLK(I2702), .RSTB(I240971), .Q(I241135) );
nor I_14024 (I241152,I69134,I69161);
DFFARX1 I_14025  ( .D(I241152), .CLK(I2702), .RSTB(I240971), .Q(I241169) );
nor I_14026 (I240960,I241169,I241118);
not I_14027 (I241200,I241169);
nor I_14028 (I241217,I69134,I69140);
nand I_14029 (I241234,I241118,I241217);
and I_14030 (I241251,I241033,I241234);
DFFARX1 I_14031  ( .D(I241251), .CLK(I2702), .RSTB(I240971), .Q(I240963) );
DFFARX1 I_14032  ( .D(I69137), .CLK(I2702), .RSTB(I240971), .Q(I241282) );
and I_14033 (I241299,I241282,I69143);
nor I_14034 (I241316,I241299,I241200);
and I_14035 (I241333,I241217,I241316);
or I_14036 (I241350,I241050,I241333);
DFFARX1 I_14037  ( .D(I241350), .CLK(I2702), .RSTB(I240971), .Q(I240948) );
not I_14038 (I241381,I241299);
nor I_14039 (I241398,I240988,I241381);
nand I_14040 (I240951,I241033,I241398);
nand I_14041 (I240945,I241169,I241381);
DFFARX1 I_14042  ( .D(I241299), .CLK(I2702), .RSTB(I240971), .Q(I240939) );
DFFARX1 I_14043  ( .D(I69155), .CLK(I2702), .RSTB(I240971), .Q(I241457) );
nand I_14044 (I240957,I241457,I241067);
DFFARX1 I_14045  ( .D(I241457), .CLK(I2702), .RSTB(I240971), .Q(I241488) );
not I_14046 (I240942,I241488);
and I_14047 (I240936,I241457,I241135);
not I_14048 (I241566,I2709);
or I_14049 (I241583,I348002,I347999);
not I_14050 (I241549,I241583);
DFFARX1 I_14051  ( .D(I241583), .CLK(I2702), .RSTB(I241566), .Q(I241528) );
or I_14052 (I241628,I348008,I348002);
nor I_14053 (I241645,I348023,I348014);
nor I_14054 (I241662,I241645,I241583);
not I_14055 (I241679,I348023);
and I_14056 (I241696,I241679,I348017);
nor I_14057 (I241713,I241696,I347999);
DFFARX1 I_14058  ( .D(I241713), .CLK(I2702), .RSTB(I241566), .Q(I241730) );
nor I_14059 (I241747,I348029,I348026);
DFFARX1 I_14060  ( .D(I241747), .CLK(I2702), .RSTB(I241566), .Q(I241764) );
nor I_14061 (I241555,I241764,I241713);
not I_14062 (I241795,I241764);
nor I_14063 (I241812,I348029,I348008);
nand I_14064 (I241829,I241713,I241812);
and I_14065 (I241846,I241628,I241829);
DFFARX1 I_14066  ( .D(I241846), .CLK(I2702), .RSTB(I241566), .Q(I241558) );
DFFARX1 I_14067  ( .D(I348005), .CLK(I2702), .RSTB(I241566), .Q(I241877) );
and I_14068 (I241894,I241877,I348020);
nor I_14069 (I241911,I241894,I241795);
and I_14070 (I241928,I241812,I241911);
or I_14071 (I241945,I241645,I241928);
DFFARX1 I_14072  ( .D(I241945), .CLK(I2702), .RSTB(I241566), .Q(I241543) );
not I_14073 (I241976,I241894);
nor I_14074 (I241993,I241583,I241976);
nand I_14075 (I241546,I241628,I241993);
nand I_14076 (I241540,I241764,I241976);
DFFARX1 I_14077  ( .D(I241894), .CLK(I2702), .RSTB(I241566), .Q(I241534) );
DFFARX1 I_14078  ( .D(I348011), .CLK(I2702), .RSTB(I241566), .Q(I242052) );
nand I_14079 (I241552,I242052,I241662);
DFFARX1 I_14080  ( .D(I242052), .CLK(I2702), .RSTB(I241566), .Q(I242083) );
not I_14081 (I241537,I242083);
and I_14082 (I241531,I242052,I241730);
not I_14083 (I242161,I2709);
or I_14084 (I242178,I631922,I631931);
not I_14085 (I242144,I242178);
DFFARX1 I_14086  ( .D(I242178), .CLK(I2702), .RSTB(I242161), .Q(I242123) );
or I_14087 (I242223,I631940,I631922);
nor I_14088 (I242240,I631934,I631928);
nor I_14089 (I242257,I242240,I242178);
not I_14090 (I242274,I631934);
and I_14091 (I242291,I242274,I631937);
nor I_14092 (I242308,I242291,I631931);
DFFARX1 I_14093  ( .D(I242308), .CLK(I2702), .RSTB(I242161), .Q(I242325) );
nor I_14094 (I242342,I631925,I631943);
DFFARX1 I_14095  ( .D(I242342), .CLK(I2702), .RSTB(I242161), .Q(I242359) );
nor I_14096 (I242150,I242359,I242308);
not I_14097 (I242390,I242359);
nor I_14098 (I242407,I631925,I631940);
nand I_14099 (I242424,I242308,I242407);
and I_14100 (I242441,I242223,I242424);
DFFARX1 I_14101  ( .D(I242441), .CLK(I2702), .RSTB(I242161), .Q(I242153) );
DFFARX1 I_14102  ( .D(I631946), .CLK(I2702), .RSTB(I242161), .Q(I242472) );
and I_14103 (I242489,I242472,I631919);
nor I_14104 (I242506,I242489,I242390);
and I_14105 (I242523,I242407,I242506);
or I_14106 (I242540,I242240,I242523);
DFFARX1 I_14107  ( .D(I242540), .CLK(I2702), .RSTB(I242161), .Q(I242138) );
not I_14108 (I242571,I242489);
nor I_14109 (I242588,I242178,I242571);
nand I_14110 (I242141,I242223,I242588);
nand I_14111 (I242135,I242359,I242571);
DFFARX1 I_14112  ( .D(I242489), .CLK(I2702), .RSTB(I242161), .Q(I242129) );
DFFARX1 I_14113  ( .D(I631916), .CLK(I2702), .RSTB(I242161), .Q(I242647) );
nand I_14114 (I242147,I242647,I242257);
DFFARX1 I_14115  ( .D(I242647), .CLK(I2702), .RSTB(I242161), .Q(I242678) );
not I_14116 (I242132,I242678);
and I_14117 (I242126,I242647,I242325);
not I_14118 (I242756,I2709);
or I_14119 (I242773,I402266,I402263);
not I_14120 (I242739,I242773);
DFFARX1 I_14121  ( .D(I242773), .CLK(I2702), .RSTB(I242756), .Q(I242718) );
or I_14122 (I242818,I402272,I402266);
nor I_14123 (I242835,I402287,I402278);
nor I_14124 (I242852,I242835,I242773);
not I_14125 (I242869,I402287);
and I_14126 (I242886,I242869,I402281);
nor I_14127 (I242903,I242886,I402263);
DFFARX1 I_14128  ( .D(I242903), .CLK(I2702), .RSTB(I242756), .Q(I242920) );
nor I_14129 (I242937,I402293,I402290);
DFFARX1 I_14130  ( .D(I242937), .CLK(I2702), .RSTB(I242756), .Q(I242954) );
nor I_14131 (I242745,I242954,I242903);
not I_14132 (I242985,I242954);
nor I_14133 (I243002,I402293,I402272);
nand I_14134 (I243019,I242903,I243002);
and I_14135 (I243036,I242818,I243019);
DFFARX1 I_14136  ( .D(I243036), .CLK(I2702), .RSTB(I242756), .Q(I242748) );
DFFARX1 I_14137  ( .D(I402269), .CLK(I2702), .RSTB(I242756), .Q(I243067) );
and I_14138 (I243084,I243067,I402284);
nor I_14139 (I243101,I243084,I242985);
and I_14140 (I243118,I243002,I243101);
or I_14141 (I243135,I242835,I243118);
DFFARX1 I_14142  ( .D(I243135), .CLK(I2702), .RSTB(I242756), .Q(I242733) );
not I_14143 (I243166,I243084);
nor I_14144 (I243183,I242773,I243166);
nand I_14145 (I242736,I242818,I243183);
nand I_14146 (I242730,I242954,I243166);
DFFARX1 I_14147  ( .D(I243084), .CLK(I2702), .RSTB(I242756), .Q(I242724) );
DFFARX1 I_14148  ( .D(I402275), .CLK(I2702), .RSTB(I242756), .Q(I243242) );
nand I_14149 (I242742,I243242,I242852);
DFFARX1 I_14150  ( .D(I243242), .CLK(I2702), .RSTB(I242756), .Q(I243273) );
not I_14151 (I242727,I243273);
and I_14152 (I242721,I243242,I242920);
not I_14153 (I243351,I2709);
or I_14154 (I243368,I394514,I394511);
not I_14155 (I243334,I243368);
DFFARX1 I_14156  ( .D(I243368), .CLK(I2702), .RSTB(I243351), .Q(I243313) );
or I_14157 (I243413,I394520,I394514);
nor I_14158 (I243430,I394535,I394526);
nor I_14159 (I243447,I243430,I243368);
not I_14160 (I243464,I394535);
and I_14161 (I243481,I243464,I394529);
nor I_14162 (I243498,I243481,I394511);
DFFARX1 I_14163  ( .D(I243498), .CLK(I2702), .RSTB(I243351), .Q(I243515) );
nor I_14164 (I243532,I394541,I394538);
DFFARX1 I_14165  ( .D(I243532), .CLK(I2702), .RSTB(I243351), .Q(I243549) );
nor I_14166 (I243340,I243549,I243498);
not I_14167 (I243580,I243549);
nor I_14168 (I243597,I394541,I394520);
nand I_14169 (I243614,I243498,I243597);
and I_14170 (I243631,I243413,I243614);
DFFARX1 I_14171  ( .D(I243631), .CLK(I2702), .RSTB(I243351), .Q(I243343) );
DFFARX1 I_14172  ( .D(I394517), .CLK(I2702), .RSTB(I243351), .Q(I243662) );
and I_14173 (I243679,I243662,I394532);
nor I_14174 (I243696,I243679,I243580);
and I_14175 (I243713,I243597,I243696);
or I_14176 (I243730,I243430,I243713);
DFFARX1 I_14177  ( .D(I243730), .CLK(I2702), .RSTB(I243351), .Q(I243328) );
not I_14178 (I243761,I243679);
nor I_14179 (I243778,I243368,I243761);
nand I_14180 (I243331,I243413,I243778);
nand I_14181 (I243325,I243549,I243761);
DFFARX1 I_14182  ( .D(I243679), .CLK(I2702), .RSTB(I243351), .Q(I243319) );
DFFARX1 I_14183  ( .D(I394523), .CLK(I2702), .RSTB(I243351), .Q(I243837) );
nand I_14184 (I243337,I243837,I243447);
DFFARX1 I_14185  ( .D(I243837), .CLK(I2702), .RSTB(I243351), .Q(I243868) );
not I_14186 (I243322,I243868);
and I_14187 (I243316,I243837,I243515);
not I_14188 (I243946,I2709);
or I_14189 (I243963,I129227,I129224);
not I_14190 (I243929,I243963);
DFFARX1 I_14191  ( .D(I243963), .CLK(I2702), .RSTB(I243946), .Q(I243908) );
or I_14192 (I244008,I129218,I129227);
nor I_14193 (I244025,I129236,I129209);
nor I_14194 (I244042,I244025,I243963);
not I_14195 (I244059,I129236);
and I_14196 (I244076,I244059,I129230);
nor I_14197 (I244093,I244076,I129224);
DFFARX1 I_14198  ( .D(I244093), .CLK(I2702), .RSTB(I243946), .Q(I244110) );
nor I_14199 (I244127,I129212,I129239);
DFFARX1 I_14200  ( .D(I244127), .CLK(I2702), .RSTB(I243946), .Q(I244144) );
nor I_14201 (I243935,I244144,I244093);
not I_14202 (I244175,I244144);
nor I_14203 (I244192,I129212,I129218);
nand I_14204 (I244209,I244093,I244192);
and I_14205 (I244226,I244008,I244209);
DFFARX1 I_14206  ( .D(I244226), .CLK(I2702), .RSTB(I243946), .Q(I243938) );
DFFARX1 I_14207  ( .D(I129215), .CLK(I2702), .RSTB(I243946), .Q(I244257) );
and I_14208 (I244274,I244257,I129221);
nor I_14209 (I244291,I244274,I244175);
and I_14210 (I244308,I244192,I244291);
or I_14211 (I244325,I244025,I244308);
DFFARX1 I_14212  ( .D(I244325), .CLK(I2702), .RSTB(I243946), .Q(I243923) );
not I_14213 (I244356,I244274);
nor I_14214 (I244373,I243963,I244356);
nand I_14215 (I243926,I244008,I244373);
nand I_14216 (I243920,I244144,I244356);
DFFARX1 I_14217  ( .D(I244274), .CLK(I2702), .RSTB(I243946), .Q(I243914) );
DFFARX1 I_14218  ( .D(I129233), .CLK(I2702), .RSTB(I243946), .Q(I244432) );
nand I_14219 (I243932,I244432,I244042);
DFFARX1 I_14220  ( .D(I244432), .CLK(I2702), .RSTB(I243946), .Q(I244463) );
not I_14221 (I243917,I244463);
and I_14222 (I243911,I244432,I244110);
not I_14223 (I244541,I2709);
or I_14224 (I244558,I65919,I65916);
not I_14225 (I244524,I244558);
DFFARX1 I_14226  ( .D(I244558), .CLK(I2702), .RSTB(I244541), .Q(I244503) );
or I_14227 (I244603,I65910,I65919);
nor I_14228 (I244620,I65928,I65901);
nor I_14229 (I244637,I244620,I244558);
not I_14230 (I244654,I65928);
and I_14231 (I244671,I244654,I65922);
nor I_14232 (I244688,I244671,I65916);
DFFARX1 I_14233  ( .D(I244688), .CLK(I2702), .RSTB(I244541), .Q(I244705) );
nor I_14234 (I244722,I65904,I65931);
DFFARX1 I_14235  ( .D(I244722), .CLK(I2702), .RSTB(I244541), .Q(I244739) );
nor I_14236 (I244530,I244739,I244688);
not I_14237 (I244770,I244739);
nor I_14238 (I244787,I65904,I65910);
nand I_14239 (I244804,I244688,I244787);
and I_14240 (I244821,I244603,I244804);
DFFARX1 I_14241  ( .D(I244821), .CLK(I2702), .RSTB(I244541), .Q(I244533) );
DFFARX1 I_14242  ( .D(I65907), .CLK(I2702), .RSTB(I244541), .Q(I244852) );
and I_14243 (I244869,I244852,I65913);
nor I_14244 (I244886,I244869,I244770);
and I_14245 (I244903,I244787,I244886);
or I_14246 (I244920,I244620,I244903);
DFFARX1 I_14247  ( .D(I244920), .CLK(I2702), .RSTB(I244541), .Q(I244518) );
not I_14248 (I244951,I244869);
nor I_14249 (I244968,I244558,I244951);
nand I_14250 (I244521,I244603,I244968);
nand I_14251 (I244515,I244739,I244951);
DFFARX1 I_14252  ( .D(I244869), .CLK(I2702), .RSTB(I244541), .Q(I244509) );
DFFARX1 I_14253  ( .D(I65925), .CLK(I2702), .RSTB(I244541), .Q(I245027) );
nand I_14254 (I244527,I245027,I244637);
DFFARX1 I_14255  ( .D(I245027), .CLK(I2702), .RSTB(I244541), .Q(I245058) );
not I_14256 (I244512,I245058);
and I_14257 (I244506,I245027,I244705);
not I_14258 (I245136,I2709);
or I_14259 (I245153,I543505,I543517);
not I_14260 (I245119,I245153);
DFFARX1 I_14261  ( .D(I245153), .CLK(I2702), .RSTB(I245136), .Q(I245098) );
or I_14262 (I245198,I543529,I543505);
nor I_14263 (I245215,I543523,I543508);
nor I_14264 (I245232,I245215,I245153);
not I_14265 (I245249,I543523);
and I_14266 (I245266,I245249,I543520);
nor I_14267 (I245283,I245266,I543517);
DFFARX1 I_14268  ( .D(I245283), .CLK(I2702), .RSTB(I245136), .Q(I245300) );
nor I_14269 (I245317,I543514,I543511);
DFFARX1 I_14270  ( .D(I245317), .CLK(I2702), .RSTB(I245136), .Q(I245334) );
nor I_14271 (I245125,I245334,I245283);
not I_14272 (I245365,I245334);
nor I_14273 (I245382,I543514,I543529);
nand I_14274 (I245399,I245283,I245382);
and I_14275 (I245416,I245198,I245399);
DFFARX1 I_14276  ( .D(I245416), .CLK(I2702), .RSTB(I245136), .Q(I245128) );
DFFARX1 I_14277  ( .D(I543526), .CLK(I2702), .RSTB(I245136), .Q(I245447) );
and I_14278 (I245464,I245447,I543499);
nor I_14279 (I245481,I245464,I245365);
and I_14280 (I245498,I245382,I245481);
or I_14281 (I245515,I245215,I245498);
DFFARX1 I_14282  ( .D(I245515), .CLK(I2702), .RSTB(I245136), .Q(I245113) );
not I_14283 (I245546,I245464);
nor I_14284 (I245563,I245153,I245546);
nand I_14285 (I245116,I245198,I245563);
nand I_14286 (I245110,I245334,I245546);
DFFARX1 I_14287  ( .D(I245464), .CLK(I2702), .RSTB(I245136), .Q(I245104) );
DFFARX1 I_14288  ( .D(I543502), .CLK(I2702), .RSTB(I245136), .Q(I245622) );
nand I_14289 (I245122,I245622,I245232);
DFFARX1 I_14290  ( .D(I245622), .CLK(I2702), .RSTB(I245136), .Q(I245653) );
not I_14291 (I245107,I245653);
and I_14292 (I245101,I245622,I245300);
not I_14293 (I245731,I2709);
or I_14294 (I245748,I36957,I36933);
not I_14295 (I245714,I245748);
DFFARX1 I_14296  ( .D(I245748), .CLK(I2702), .RSTB(I245731), .Q(I245693) );
or I_14297 (I245793,I36960,I36957);
nor I_14298 (I245810,I36942,I36948);
nor I_14299 (I245827,I245810,I245748);
not I_14300 (I245844,I36942);
and I_14301 (I245861,I245844,I36936);
nor I_14302 (I245878,I245861,I36933);
DFFARX1 I_14303  ( .D(I245878), .CLK(I2702), .RSTB(I245731), .Q(I245895) );
nor I_14304 (I245912,I36963,I36954);
DFFARX1 I_14305  ( .D(I245912), .CLK(I2702), .RSTB(I245731), .Q(I245929) );
nor I_14306 (I245720,I245929,I245878);
not I_14307 (I245960,I245929);
nor I_14308 (I245977,I36963,I36960);
nand I_14309 (I245994,I245878,I245977);
and I_14310 (I246011,I245793,I245994);
DFFARX1 I_14311  ( .D(I246011), .CLK(I2702), .RSTB(I245731), .Q(I245723) );
DFFARX1 I_14312  ( .D(I36939), .CLK(I2702), .RSTB(I245731), .Q(I246042) );
and I_14313 (I246059,I246042,I36951);
nor I_14314 (I246076,I246059,I245960);
and I_14315 (I246093,I245977,I246076);
or I_14316 (I246110,I245810,I246093);
DFFARX1 I_14317  ( .D(I246110), .CLK(I2702), .RSTB(I245731), .Q(I245708) );
not I_14318 (I246141,I246059);
nor I_14319 (I246158,I245748,I246141);
nand I_14320 (I245711,I245793,I246158);
nand I_14321 (I245705,I245929,I246141);
DFFARX1 I_14322  ( .D(I246059), .CLK(I2702), .RSTB(I245731), .Q(I245699) );
DFFARX1 I_14323  ( .D(I36945), .CLK(I2702), .RSTB(I245731), .Q(I246217) );
nand I_14324 (I245717,I246217,I245827);
DFFARX1 I_14325  ( .D(I246217), .CLK(I2702), .RSTB(I245731), .Q(I246248) );
not I_14326 (I245702,I246248);
and I_14327 (I245696,I246217,I245895);
not I_14328 (I246326,I2709);
not I_14329 (I246343,I520312);
nor I_14330 (I246360,I520321,I520303);
nand I_14331 (I246377,I246360,I520324);
nor I_14332 (I246394,I246343,I520321);
nand I_14333 (I246411,I246394,I520315);
not I_14334 (I246428,I246411);
not I_14335 (I246445,I520321);
nor I_14336 (I246315,I246411,I246445);
not I_14337 (I246476,I246445);
nand I_14338 (I246300,I246411,I246476);
not I_14339 (I246507,I520309);
nor I_14340 (I246524,I246507,I520300);
and I_14341 (I246541,I246524,I520297);
or I_14342 (I246558,I246541,I520294);
DFFARX1 I_14343  ( .D(I246558), .CLK(I2702), .RSTB(I246326), .Q(I246575) );
nor I_14344 (I246592,I246575,I246428);
DFFARX1 I_14345  ( .D(I246575), .CLK(I2702), .RSTB(I246326), .Q(I246609) );
not I_14346 (I246297,I246609);
nand I_14347 (I246640,I246343,I520309);
and I_14348 (I246657,I246640,I246592);
DFFARX1 I_14349  ( .D(I246640), .CLK(I2702), .RSTB(I246326), .Q(I246294) );
DFFARX1 I_14350  ( .D(I520318), .CLK(I2702), .RSTB(I246326), .Q(I246688) );
nor I_14351 (I246705,I246688,I246411);
nand I_14352 (I246312,I246575,I246705);
nor I_14353 (I246736,I246688,I246476);
not I_14354 (I246309,I246688);
nand I_14355 (I246767,I246688,I246377);
and I_14356 (I246784,I246445,I246767);
DFFARX1 I_14357  ( .D(I246784), .CLK(I2702), .RSTB(I246326), .Q(I246288) );
DFFARX1 I_14358  ( .D(I246688), .CLK(I2702), .RSTB(I246326), .Q(I246291) );
DFFARX1 I_14359  ( .D(I520306), .CLK(I2702), .RSTB(I246326), .Q(I246829) );
not I_14360 (I246846,I246829);
nand I_14361 (I246863,I246846,I246411);
and I_14362 (I246880,I246640,I246863);
DFFARX1 I_14363  ( .D(I246880), .CLK(I2702), .RSTB(I246326), .Q(I246318) );
or I_14364 (I246911,I246846,I246657);
DFFARX1 I_14365  ( .D(I246911), .CLK(I2702), .RSTB(I246326), .Q(I246303) );
nand I_14366 (I246306,I246846,I246736);
not I_14367 (I246989,I2709);
not I_14368 (I247006,I166731);
nor I_14369 (I247023,I166737,I166743);
nand I_14370 (I247040,I247023,I166746);
nor I_14371 (I247057,I247006,I166737);
nand I_14372 (I247074,I247057,I166728);
not I_14373 (I247091,I247074);
not I_14374 (I247108,I166737);
nor I_14375 (I246978,I247074,I247108);
not I_14376 (I247139,I247108);
nand I_14377 (I246963,I247074,I247139);
not I_14378 (I247170,I166740);
nor I_14379 (I247187,I247170,I166734);
and I_14380 (I247204,I247187,I166749);
or I_14381 (I247221,I247204,I166755);
DFFARX1 I_14382  ( .D(I247221), .CLK(I2702), .RSTB(I246989), .Q(I247238) );
nor I_14383 (I247255,I247238,I247091);
DFFARX1 I_14384  ( .D(I247238), .CLK(I2702), .RSTB(I246989), .Q(I247272) );
not I_14385 (I246960,I247272);
nand I_14386 (I247303,I247006,I166740);
and I_14387 (I247320,I247303,I247255);
DFFARX1 I_14388  ( .D(I247303), .CLK(I2702), .RSTB(I246989), .Q(I246957) );
DFFARX1 I_14389  ( .D(I166752), .CLK(I2702), .RSTB(I246989), .Q(I247351) );
nor I_14390 (I247368,I247351,I247074);
nand I_14391 (I246975,I247238,I247368);
nor I_14392 (I247399,I247351,I247139);
not I_14393 (I246972,I247351);
nand I_14394 (I247430,I247351,I247040);
and I_14395 (I247447,I247108,I247430);
DFFARX1 I_14396  ( .D(I247447), .CLK(I2702), .RSTB(I246989), .Q(I246951) );
DFFARX1 I_14397  ( .D(I247351), .CLK(I2702), .RSTB(I246989), .Q(I246954) );
DFFARX1 I_14398  ( .D(I166758), .CLK(I2702), .RSTB(I246989), .Q(I247492) );
not I_14399 (I247509,I247492);
nand I_14400 (I247526,I247509,I247074);
and I_14401 (I247543,I247303,I247526);
DFFARX1 I_14402  ( .D(I247543), .CLK(I2702), .RSTB(I246989), .Q(I246981) );
or I_14403 (I247574,I247509,I247320);
DFFARX1 I_14404  ( .D(I247574), .CLK(I2702), .RSTB(I246989), .Q(I246966) );
nand I_14405 (I246969,I247509,I247399);
not I_14406 (I247652,I2709);
not I_14407 (I247669,I412571);
nor I_14408 (I247686,I412574,I412580);
nand I_14409 (I247703,I247686,I412586);
nor I_14410 (I247720,I247669,I412574);
nand I_14411 (I247737,I247720,I412565);
not I_14412 (I247754,I247737);
not I_14413 (I247771,I412574);
nor I_14414 (I247641,I247737,I247771);
not I_14415 (I247802,I247771);
nand I_14416 (I247626,I247737,I247802);
not I_14417 (I247833,I412577);
nor I_14418 (I247850,I247833,I412592);
and I_14419 (I247867,I247850,I412595);
or I_14420 (I247884,I247867,I412568);
DFFARX1 I_14421  ( .D(I247884), .CLK(I2702), .RSTB(I247652), .Q(I247901) );
nor I_14422 (I247918,I247901,I247754);
DFFARX1 I_14423  ( .D(I247901), .CLK(I2702), .RSTB(I247652), .Q(I247935) );
not I_14424 (I247623,I247935);
nand I_14425 (I247966,I247669,I412577);
and I_14426 (I247983,I247966,I247918);
DFFARX1 I_14427  ( .D(I247966), .CLK(I2702), .RSTB(I247652), .Q(I247620) );
DFFARX1 I_14428  ( .D(I412589), .CLK(I2702), .RSTB(I247652), .Q(I248014) );
nor I_14429 (I248031,I248014,I247737);
nand I_14430 (I247638,I247901,I248031);
nor I_14431 (I248062,I248014,I247802);
not I_14432 (I247635,I248014);
nand I_14433 (I248093,I248014,I247703);
and I_14434 (I248110,I247771,I248093);
DFFARX1 I_14435  ( .D(I248110), .CLK(I2702), .RSTB(I247652), .Q(I247614) );
DFFARX1 I_14436  ( .D(I248014), .CLK(I2702), .RSTB(I247652), .Q(I247617) );
DFFARX1 I_14437  ( .D(I412583), .CLK(I2702), .RSTB(I247652), .Q(I248155) );
not I_14438 (I248172,I248155);
nand I_14439 (I248189,I248172,I247737);
and I_14440 (I248206,I247966,I248189);
DFFARX1 I_14441  ( .D(I248206), .CLK(I2702), .RSTB(I247652), .Q(I247644) );
or I_14442 (I248237,I248172,I247983);
DFFARX1 I_14443  ( .D(I248237), .CLK(I2702), .RSTB(I247652), .Q(I247629) );
nand I_14444 (I247632,I248172,I248062);
not I_14445 (I248315,I2709);
not I_14446 (I248332,I154797);
nor I_14447 (I248349,I154803,I154809);
nand I_14448 (I248366,I248349,I154812);
nor I_14449 (I248383,I248332,I154803);
nand I_14450 (I248400,I248383,I154794);
not I_14451 (I248417,I248400);
not I_14452 (I248434,I154803);
nor I_14453 (I248304,I248400,I248434);
not I_14454 (I248465,I248434);
nand I_14455 (I248289,I248400,I248465);
not I_14456 (I248496,I154806);
nor I_14457 (I248513,I248496,I154800);
and I_14458 (I248530,I248513,I154815);
or I_14459 (I248547,I248530,I154821);
DFFARX1 I_14460  ( .D(I248547), .CLK(I2702), .RSTB(I248315), .Q(I248564) );
nor I_14461 (I248581,I248564,I248417);
DFFARX1 I_14462  ( .D(I248564), .CLK(I2702), .RSTB(I248315), .Q(I248598) );
not I_14463 (I248286,I248598);
nand I_14464 (I248629,I248332,I154806);
and I_14465 (I248646,I248629,I248581);
DFFARX1 I_14466  ( .D(I248629), .CLK(I2702), .RSTB(I248315), .Q(I248283) );
DFFARX1 I_14467  ( .D(I154818), .CLK(I2702), .RSTB(I248315), .Q(I248677) );
nor I_14468 (I248694,I248677,I248400);
nand I_14469 (I248301,I248564,I248694);
nor I_14470 (I248725,I248677,I248465);
not I_14471 (I248298,I248677);
nand I_14472 (I248756,I248677,I248366);
and I_14473 (I248773,I248434,I248756);
DFFARX1 I_14474  ( .D(I248773), .CLK(I2702), .RSTB(I248315), .Q(I248277) );
DFFARX1 I_14475  ( .D(I248677), .CLK(I2702), .RSTB(I248315), .Q(I248280) );
DFFARX1 I_14476  ( .D(I154824), .CLK(I2702), .RSTB(I248315), .Q(I248818) );
not I_14477 (I248835,I248818);
nand I_14478 (I248852,I248835,I248400);
and I_14479 (I248869,I248629,I248852);
DFFARX1 I_14480  ( .D(I248869), .CLK(I2702), .RSTB(I248315), .Q(I248307) );
or I_14481 (I248900,I248835,I248646);
DFFARX1 I_14482  ( .D(I248900), .CLK(I2702), .RSTB(I248315), .Q(I248292) );
nand I_14483 (I248295,I248835,I248725);
not I_14484 (I248978,I2709);
not I_14485 (I248995,I435598);
nor I_14486 (I249012,I435610,I435592);
nand I_14487 (I249029,I249012,I435613);
nor I_14488 (I249046,I248995,I435610);
nand I_14489 (I249063,I249046,I435604);
not I_14490 (I249080,I249063);
not I_14491 (I249097,I435610);
nor I_14492 (I248967,I249063,I249097);
not I_14493 (I249128,I249097);
nand I_14494 (I248952,I249063,I249128);
not I_14495 (I249159,I435595);
nor I_14496 (I249176,I249159,I435589);
and I_14497 (I249193,I249176,I435601);
or I_14498 (I249210,I249193,I435586);
DFFARX1 I_14499  ( .D(I249210), .CLK(I2702), .RSTB(I248978), .Q(I249227) );
nor I_14500 (I249244,I249227,I249080);
DFFARX1 I_14501  ( .D(I249227), .CLK(I2702), .RSTB(I248978), .Q(I249261) );
not I_14502 (I248949,I249261);
nand I_14503 (I249292,I248995,I435595);
and I_14504 (I249309,I249292,I249244);
DFFARX1 I_14505  ( .D(I249292), .CLK(I2702), .RSTB(I248978), .Q(I248946) );
DFFARX1 I_14506  ( .D(I435583), .CLK(I2702), .RSTB(I248978), .Q(I249340) );
nor I_14507 (I249357,I249340,I249063);
nand I_14508 (I248964,I249227,I249357);
nor I_14509 (I249388,I249340,I249128);
not I_14510 (I248961,I249340);
nand I_14511 (I249419,I249340,I249029);
and I_14512 (I249436,I249097,I249419);
DFFARX1 I_14513  ( .D(I249436), .CLK(I2702), .RSTB(I248978), .Q(I248940) );
DFFARX1 I_14514  ( .D(I249340), .CLK(I2702), .RSTB(I248978), .Q(I248943) );
DFFARX1 I_14515  ( .D(I435607), .CLK(I2702), .RSTB(I248978), .Q(I249481) );
not I_14516 (I249498,I249481);
nand I_14517 (I249515,I249498,I249063);
and I_14518 (I249532,I249292,I249515);
DFFARX1 I_14519  ( .D(I249532), .CLK(I2702), .RSTB(I248978), .Q(I248970) );
or I_14520 (I249563,I249498,I249309);
DFFARX1 I_14521  ( .D(I249563), .CLK(I2702), .RSTB(I248978), .Q(I248955) );
nand I_14522 (I248958,I249498,I249388);
not I_14523 (I249641,I2709);
not I_14524 (I249658,I507817);
nor I_14525 (I249675,I507826,I507808);
nand I_14526 (I249692,I249675,I507829);
nor I_14527 (I249709,I249658,I507826);
nand I_14528 (I249726,I249709,I507820);
not I_14529 (I249743,I249726);
not I_14530 (I249760,I507826);
nor I_14531 (I249630,I249726,I249760);
not I_14532 (I249791,I249760);
nand I_14533 (I249615,I249726,I249791);
not I_14534 (I249822,I507814);
nor I_14535 (I249839,I249822,I507805);
and I_14536 (I249856,I249839,I507802);
or I_14537 (I249873,I249856,I507799);
DFFARX1 I_14538  ( .D(I249873), .CLK(I2702), .RSTB(I249641), .Q(I249890) );
nor I_14539 (I249907,I249890,I249743);
DFFARX1 I_14540  ( .D(I249890), .CLK(I2702), .RSTB(I249641), .Q(I249924) );
not I_14541 (I249612,I249924);
nand I_14542 (I249955,I249658,I507814);
and I_14543 (I249972,I249955,I249907);
DFFARX1 I_14544  ( .D(I249955), .CLK(I2702), .RSTB(I249641), .Q(I249609) );
DFFARX1 I_14545  ( .D(I507823), .CLK(I2702), .RSTB(I249641), .Q(I250003) );
nor I_14546 (I250020,I250003,I249726);
nand I_14547 (I249627,I249890,I250020);
nor I_14548 (I250051,I250003,I249791);
not I_14549 (I249624,I250003);
nand I_14550 (I250082,I250003,I249692);
and I_14551 (I250099,I249760,I250082);
DFFARX1 I_14552  ( .D(I250099), .CLK(I2702), .RSTB(I249641), .Q(I249603) );
DFFARX1 I_14553  ( .D(I250003), .CLK(I2702), .RSTB(I249641), .Q(I249606) );
DFFARX1 I_14554  ( .D(I507811), .CLK(I2702), .RSTB(I249641), .Q(I250144) );
not I_14555 (I250161,I250144);
nand I_14556 (I250178,I250161,I249726);
and I_14557 (I250195,I249955,I250178);
DFFARX1 I_14558  ( .D(I250195), .CLK(I2702), .RSTB(I249641), .Q(I249633) );
or I_14559 (I250226,I250161,I249972);
DFFARX1 I_14560  ( .D(I250226), .CLK(I2702), .RSTB(I249641), .Q(I249618) );
nand I_14561 (I249621,I250161,I250051);
not I_14562 (I250304,I2709);
not I_14563 (I250321,I592902);
nor I_14564 (I250338,I592899,I592890);
nand I_14565 (I250355,I250338,I592893);
nor I_14566 (I250372,I250321,I592899);
nand I_14567 (I250389,I250372,I592887);
not I_14568 (I250406,I250389);
not I_14569 (I250423,I592899);
nor I_14570 (I250293,I250389,I250423);
not I_14571 (I250454,I250423);
nand I_14572 (I250278,I250389,I250454);
not I_14573 (I250485,I592908);
nor I_14574 (I250502,I250485,I592911);
and I_14575 (I250519,I250502,I592896);
or I_14576 (I250536,I250519,I592884);
DFFARX1 I_14577  ( .D(I250536), .CLK(I2702), .RSTB(I250304), .Q(I250553) );
nor I_14578 (I250570,I250553,I250406);
DFFARX1 I_14579  ( .D(I250553), .CLK(I2702), .RSTB(I250304), .Q(I250587) );
not I_14580 (I250275,I250587);
nand I_14581 (I250618,I250321,I592908);
and I_14582 (I250635,I250618,I250570);
DFFARX1 I_14583  ( .D(I250618), .CLK(I2702), .RSTB(I250304), .Q(I250272) );
DFFARX1 I_14584  ( .D(I592905), .CLK(I2702), .RSTB(I250304), .Q(I250666) );
nor I_14585 (I250683,I250666,I250389);
nand I_14586 (I250290,I250553,I250683);
nor I_14587 (I250714,I250666,I250454);
not I_14588 (I250287,I250666);
nand I_14589 (I250745,I250666,I250355);
and I_14590 (I250762,I250423,I250745);
DFFARX1 I_14591  ( .D(I250762), .CLK(I2702), .RSTB(I250304), .Q(I250266) );
DFFARX1 I_14592  ( .D(I250666), .CLK(I2702), .RSTB(I250304), .Q(I250269) );
DFFARX1 I_14593  ( .D(I592914), .CLK(I2702), .RSTB(I250304), .Q(I250807) );
not I_14594 (I250824,I250807);
nand I_14595 (I250841,I250824,I250389);
and I_14596 (I250858,I250618,I250841);
DFFARX1 I_14597  ( .D(I250858), .CLK(I2702), .RSTB(I250304), .Q(I250296) );
or I_14598 (I250889,I250824,I250635);
DFFARX1 I_14599  ( .D(I250889), .CLK(I2702), .RSTB(I250304), .Q(I250281) );
nand I_14600 (I250284,I250824,I250714);
not I_14601 (I250967,I2709);
not I_14602 (I250984,I187947);
nor I_14603 (I251001,I187953,I187959);
nand I_14604 (I251018,I251001,I187962);
nor I_14605 (I251035,I250984,I187953);
nand I_14606 (I251052,I251035,I187944);
not I_14607 (I251069,I251052);
not I_14608 (I251086,I187953);
nor I_14609 (I250956,I251052,I251086);
not I_14610 (I251117,I251086);
nand I_14611 (I250941,I251052,I251117);
not I_14612 (I251148,I187956);
nor I_14613 (I251165,I251148,I187950);
and I_14614 (I251182,I251165,I187965);
or I_14615 (I251199,I251182,I187971);
DFFARX1 I_14616  ( .D(I251199), .CLK(I2702), .RSTB(I250967), .Q(I251216) );
nor I_14617 (I251233,I251216,I251069);
DFFARX1 I_14618  ( .D(I251216), .CLK(I2702), .RSTB(I250967), .Q(I251250) );
not I_14619 (I250938,I251250);
nand I_14620 (I251281,I250984,I187956);
and I_14621 (I251298,I251281,I251233);
DFFARX1 I_14622  ( .D(I251281), .CLK(I2702), .RSTB(I250967), .Q(I250935) );
DFFARX1 I_14623  ( .D(I187968), .CLK(I2702), .RSTB(I250967), .Q(I251329) );
nor I_14624 (I251346,I251329,I251052);
nand I_14625 (I250953,I251216,I251346);
nor I_14626 (I251377,I251329,I251117);
not I_14627 (I250950,I251329);
nand I_14628 (I251408,I251329,I251018);
and I_14629 (I251425,I251086,I251408);
DFFARX1 I_14630  ( .D(I251425), .CLK(I2702), .RSTB(I250967), .Q(I250929) );
DFFARX1 I_14631  ( .D(I251329), .CLK(I2702), .RSTB(I250967), .Q(I250932) );
DFFARX1 I_14632  ( .D(I187974), .CLK(I2702), .RSTB(I250967), .Q(I251470) );
not I_14633 (I251487,I251470);
nand I_14634 (I251504,I251487,I251052);
and I_14635 (I251521,I251281,I251504);
DFFARX1 I_14636  ( .D(I251521), .CLK(I2702), .RSTB(I250967), .Q(I250959) );
or I_14637 (I251552,I251487,I251298);
DFFARX1 I_14638  ( .D(I251552), .CLK(I2702), .RSTB(I250967), .Q(I250944) );
nand I_14639 (I250947,I251487,I251377);
not I_14640 (I251630,I2709);
not I_14641 (I251647,I40878);
nor I_14642 (I251664,I40884,I40887);
nand I_14643 (I251681,I251664,I40863);
nor I_14644 (I251698,I251647,I40884);
nand I_14645 (I251715,I251698,I40872);
not I_14646 (I251732,I251715);
not I_14647 (I251749,I40884);
nor I_14648 (I251619,I251715,I251749);
not I_14649 (I251780,I251749);
nand I_14650 (I251604,I251715,I251780);
not I_14651 (I251811,I40866);
nor I_14652 (I251828,I251811,I40890);
and I_14653 (I251845,I251828,I40860);
or I_14654 (I251862,I251845,I40869);
DFFARX1 I_14655  ( .D(I251862), .CLK(I2702), .RSTB(I251630), .Q(I251879) );
nor I_14656 (I251896,I251879,I251732);
DFFARX1 I_14657  ( .D(I251879), .CLK(I2702), .RSTB(I251630), .Q(I251913) );
not I_14658 (I251601,I251913);
nand I_14659 (I251944,I251647,I40866);
and I_14660 (I251961,I251944,I251896);
DFFARX1 I_14661  ( .D(I251944), .CLK(I2702), .RSTB(I251630), .Q(I251598) );
DFFARX1 I_14662  ( .D(I40875), .CLK(I2702), .RSTB(I251630), .Q(I251992) );
nor I_14663 (I252009,I251992,I251715);
nand I_14664 (I251616,I251879,I252009);
nor I_14665 (I252040,I251992,I251780);
not I_14666 (I251613,I251992);
nand I_14667 (I252071,I251992,I251681);
and I_14668 (I252088,I251749,I252071);
DFFARX1 I_14669  ( .D(I252088), .CLK(I2702), .RSTB(I251630), .Q(I251592) );
DFFARX1 I_14670  ( .D(I251992), .CLK(I2702), .RSTB(I251630), .Q(I251595) );
DFFARX1 I_14671  ( .D(I40881), .CLK(I2702), .RSTB(I251630), .Q(I252133) );
not I_14672 (I252150,I252133);
nand I_14673 (I252167,I252150,I251715);
and I_14674 (I252184,I251944,I252167);
DFFARX1 I_14675  ( .D(I252184), .CLK(I2702), .RSTB(I251630), .Q(I251622) );
or I_14676 (I252215,I252150,I251961);
DFFARX1 I_14677  ( .D(I252215), .CLK(I2702), .RSTB(I251630), .Q(I251607) );
nand I_14678 (I251610,I252150,I252040);
not I_14679 (I252293,I2709);
not I_14680 (I252310,I707714);
nor I_14681 (I252327,I707705,I707711);
nand I_14682 (I252344,I252327,I707723);
nor I_14683 (I252361,I252310,I707705);
nand I_14684 (I252378,I252361,I707708);
not I_14685 (I252395,I252378);
not I_14686 (I252412,I707705);
nor I_14687 (I252282,I252378,I252412);
not I_14688 (I252443,I252412);
nand I_14689 (I252267,I252378,I252443);
not I_14690 (I252474,I707732);
nor I_14691 (I252491,I252474,I707726);
and I_14692 (I252508,I252491,I707717);
or I_14693 (I252525,I252508,I707702);
DFFARX1 I_14694  ( .D(I252525), .CLK(I2702), .RSTB(I252293), .Q(I252542) );
nor I_14695 (I252559,I252542,I252395);
DFFARX1 I_14696  ( .D(I252542), .CLK(I2702), .RSTB(I252293), .Q(I252576) );
not I_14697 (I252264,I252576);
nand I_14698 (I252607,I252310,I707732);
and I_14699 (I252624,I252607,I252559);
DFFARX1 I_14700  ( .D(I252607), .CLK(I2702), .RSTB(I252293), .Q(I252261) );
DFFARX1 I_14701  ( .D(I707720), .CLK(I2702), .RSTB(I252293), .Q(I252655) );
nor I_14702 (I252672,I252655,I252378);
nand I_14703 (I252279,I252542,I252672);
nor I_14704 (I252703,I252655,I252443);
not I_14705 (I252276,I252655);
nand I_14706 (I252734,I252655,I252344);
and I_14707 (I252751,I252412,I252734);
DFFARX1 I_14708  ( .D(I252751), .CLK(I2702), .RSTB(I252293), .Q(I252255) );
DFFARX1 I_14709  ( .D(I252655), .CLK(I2702), .RSTB(I252293), .Q(I252258) );
DFFARX1 I_14710  ( .D(I707729), .CLK(I2702), .RSTB(I252293), .Q(I252796) );
not I_14711 (I252813,I252796);
nand I_14712 (I252830,I252813,I252378);
and I_14713 (I252847,I252607,I252830);
DFFARX1 I_14714  ( .D(I252847), .CLK(I2702), .RSTB(I252293), .Q(I252285) );
or I_14715 (I252878,I252813,I252624);
DFFARX1 I_14716  ( .D(I252878), .CLK(I2702), .RSTB(I252293), .Q(I252270) );
nand I_14717 (I252273,I252813,I252703);
not I_14718 (I252956,I2709);
not I_14719 (I252973,I477214);
nor I_14720 (I252990,I477226,I477208);
nand I_14721 (I253007,I252990,I477229);
nor I_14722 (I253024,I252973,I477226);
nand I_14723 (I253041,I253024,I477220);
not I_14724 (I253058,I253041);
not I_14725 (I253075,I477226);
nor I_14726 (I252945,I253041,I253075);
not I_14727 (I253106,I253075);
nand I_14728 (I252930,I253041,I253106);
not I_14729 (I253137,I477211);
nor I_14730 (I253154,I253137,I477205);
and I_14731 (I253171,I253154,I477217);
or I_14732 (I253188,I253171,I477202);
DFFARX1 I_14733  ( .D(I253188), .CLK(I2702), .RSTB(I252956), .Q(I253205) );
nor I_14734 (I253222,I253205,I253058);
DFFARX1 I_14735  ( .D(I253205), .CLK(I2702), .RSTB(I252956), .Q(I253239) );
not I_14736 (I252927,I253239);
nand I_14737 (I253270,I252973,I477211);
and I_14738 (I253287,I253270,I253222);
DFFARX1 I_14739  ( .D(I253270), .CLK(I2702), .RSTB(I252956), .Q(I252924) );
DFFARX1 I_14740  ( .D(I477199), .CLK(I2702), .RSTB(I252956), .Q(I253318) );
nor I_14741 (I253335,I253318,I253041);
nand I_14742 (I252942,I253205,I253335);
nor I_14743 (I253366,I253318,I253106);
not I_14744 (I252939,I253318);
nand I_14745 (I253397,I253318,I253007);
and I_14746 (I253414,I253075,I253397);
DFFARX1 I_14747  ( .D(I253414), .CLK(I2702), .RSTB(I252956), .Q(I252918) );
DFFARX1 I_14748  ( .D(I253318), .CLK(I2702), .RSTB(I252956), .Q(I252921) );
DFFARX1 I_14749  ( .D(I477223), .CLK(I2702), .RSTB(I252956), .Q(I253459) );
not I_14750 (I253476,I253459);
nand I_14751 (I253493,I253476,I253041);
and I_14752 (I253510,I253270,I253493);
DFFARX1 I_14753  ( .D(I253510), .CLK(I2702), .RSTB(I252956), .Q(I252948) );
or I_14754 (I253541,I253476,I253287);
DFFARX1 I_14755  ( .D(I253541), .CLK(I2702), .RSTB(I252956), .Q(I252933) );
nand I_14756 (I252936,I253476,I253366);
not I_14757 (I253619,I2709);
not I_14758 (I253636,I688532);
nor I_14759 (I253653,I688550,I688541);
nand I_14760 (I253670,I253653,I688547);
nor I_14761 (I253687,I253636,I688550);
nand I_14762 (I253704,I253687,I688553);
not I_14763 (I253721,I253704);
not I_14764 (I253738,I688550);
nor I_14765 (I253608,I253704,I253738);
not I_14766 (I253769,I253738);
nand I_14767 (I253593,I253704,I253769);
not I_14768 (I253800,I688529);
nor I_14769 (I253817,I253800,I688544);
and I_14770 (I253834,I253817,I688526);
or I_14771 (I253851,I253834,I688535);
DFFARX1 I_14772  ( .D(I253851), .CLK(I2702), .RSTB(I253619), .Q(I253868) );
nor I_14773 (I253885,I253868,I253721);
DFFARX1 I_14774  ( .D(I253868), .CLK(I2702), .RSTB(I253619), .Q(I253902) );
not I_14775 (I253590,I253902);
nand I_14776 (I253933,I253636,I688529);
and I_14777 (I253950,I253933,I253885);
DFFARX1 I_14778  ( .D(I253933), .CLK(I2702), .RSTB(I253619), .Q(I253587) );
DFFARX1 I_14779  ( .D(I688538), .CLK(I2702), .RSTB(I253619), .Q(I253981) );
nor I_14780 (I253998,I253981,I253704);
nand I_14781 (I253605,I253868,I253998);
nor I_14782 (I254029,I253981,I253769);
not I_14783 (I253602,I253981);
nand I_14784 (I254060,I253981,I253670);
and I_14785 (I254077,I253738,I254060);
DFFARX1 I_14786  ( .D(I254077), .CLK(I2702), .RSTB(I253619), .Q(I253581) );
DFFARX1 I_14787  ( .D(I253981), .CLK(I2702), .RSTB(I253619), .Q(I253584) );
DFFARX1 I_14788  ( .D(I688556), .CLK(I2702), .RSTB(I253619), .Q(I254122) );
not I_14789 (I254139,I254122);
nand I_14790 (I254156,I254139,I253704);
and I_14791 (I254173,I253933,I254156);
DFFARX1 I_14792  ( .D(I254173), .CLK(I2702), .RSTB(I253619), .Q(I253611) );
or I_14793 (I254204,I254139,I253950);
DFFARX1 I_14794  ( .D(I254204), .CLK(I2702), .RSTB(I253619), .Q(I253596) );
nand I_14795 (I253599,I254139,I254029);
not I_14796 (I254282,I2709);
not I_14797 (I254299,I544112);
nor I_14798 (I254316,I544121,I544103);
nand I_14799 (I254333,I254316,I544124);
nor I_14800 (I254350,I254299,I544121);
nand I_14801 (I254367,I254350,I544115);
not I_14802 (I254384,I254367);
not I_14803 (I254401,I544121);
nor I_14804 (I254271,I254367,I254401);
not I_14805 (I254432,I254401);
nand I_14806 (I254256,I254367,I254432);
not I_14807 (I254463,I544109);
nor I_14808 (I254480,I254463,I544100);
and I_14809 (I254497,I254480,I544097);
or I_14810 (I254514,I254497,I544094);
DFFARX1 I_14811  ( .D(I254514), .CLK(I2702), .RSTB(I254282), .Q(I254531) );
nor I_14812 (I254548,I254531,I254384);
DFFARX1 I_14813  ( .D(I254531), .CLK(I2702), .RSTB(I254282), .Q(I254565) );
not I_14814 (I254253,I254565);
nand I_14815 (I254596,I254299,I544109);
and I_14816 (I254613,I254596,I254548);
DFFARX1 I_14817  ( .D(I254596), .CLK(I2702), .RSTB(I254282), .Q(I254250) );
DFFARX1 I_14818  ( .D(I544118), .CLK(I2702), .RSTB(I254282), .Q(I254644) );
nor I_14819 (I254661,I254644,I254367);
nand I_14820 (I254268,I254531,I254661);
nor I_14821 (I254692,I254644,I254432);
not I_14822 (I254265,I254644);
nand I_14823 (I254723,I254644,I254333);
and I_14824 (I254740,I254401,I254723);
DFFARX1 I_14825  ( .D(I254740), .CLK(I2702), .RSTB(I254282), .Q(I254244) );
DFFARX1 I_14826  ( .D(I254644), .CLK(I2702), .RSTB(I254282), .Q(I254247) );
DFFARX1 I_14827  ( .D(I544106), .CLK(I2702), .RSTB(I254282), .Q(I254785) );
not I_14828 (I254802,I254785);
nand I_14829 (I254819,I254802,I254367);
and I_14830 (I254836,I254596,I254819);
DFFARX1 I_14831  ( .D(I254836), .CLK(I2702), .RSTB(I254282), .Q(I254274) );
or I_14832 (I254867,I254802,I254613);
DFFARX1 I_14833  ( .D(I254867), .CLK(I2702), .RSTB(I254282), .Q(I254259) );
nand I_14834 (I254262,I254802,I254692);
not I_14835 (I254945,I2709);
not I_14836 (I254962,I371267);
nor I_14837 (I254979,I371264,I371282);
nand I_14838 (I254996,I254979,I371285);
nor I_14839 (I255013,I254962,I371264);
nand I_14840 (I255030,I255013,I371270);
not I_14841 (I255047,I255030);
not I_14842 (I255064,I371264);
nor I_14843 (I254934,I255030,I255064);
not I_14844 (I255095,I255064);
nand I_14845 (I254919,I255030,I255095);
not I_14846 (I255126,I371279);
nor I_14847 (I255143,I255126,I371261);
and I_14848 (I255160,I255143,I371255);
or I_14849 (I255177,I255160,I371273);
DFFARX1 I_14850  ( .D(I255177), .CLK(I2702), .RSTB(I254945), .Q(I255194) );
nor I_14851 (I255211,I255194,I255047);
DFFARX1 I_14852  ( .D(I255194), .CLK(I2702), .RSTB(I254945), .Q(I255228) );
not I_14853 (I254916,I255228);
nand I_14854 (I255259,I254962,I371279);
and I_14855 (I255276,I255259,I255211);
DFFARX1 I_14856  ( .D(I255259), .CLK(I2702), .RSTB(I254945), .Q(I254913) );
DFFARX1 I_14857  ( .D(I371258), .CLK(I2702), .RSTB(I254945), .Q(I255307) );
nor I_14858 (I255324,I255307,I255030);
nand I_14859 (I254931,I255194,I255324);
nor I_14860 (I255355,I255307,I255095);
not I_14861 (I254928,I255307);
nand I_14862 (I255386,I255307,I254996);
and I_14863 (I255403,I255064,I255386);
DFFARX1 I_14864  ( .D(I255403), .CLK(I2702), .RSTB(I254945), .Q(I254907) );
DFFARX1 I_14865  ( .D(I255307), .CLK(I2702), .RSTB(I254945), .Q(I254910) );
DFFARX1 I_14866  ( .D(I371276), .CLK(I2702), .RSTB(I254945), .Q(I255448) );
not I_14867 (I255465,I255448);
nand I_14868 (I255482,I255465,I255030);
and I_14869 (I255499,I255259,I255482);
DFFARX1 I_14870  ( .D(I255499), .CLK(I2702), .RSTB(I254945), .Q(I254937) );
or I_14871 (I255530,I255465,I255276);
DFFARX1 I_14872  ( .D(I255530), .CLK(I2702), .RSTB(I254945), .Q(I254922) );
nand I_14873 (I254925,I255465,I255355);
not I_14874 (I255608,I2709);
not I_14875 (I255625,I553632);
nor I_14876 (I255642,I553641,I553623);
nand I_14877 (I255659,I255642,I553644);
nor I_14878 (I255676,I255625,I553641);
nand I_14879 (I255693,I255676,I553635);
not I_14880 (I255710,I255693);
not I_14881 (I255727,I553641);
nor I_14882 (I255597,I255693,I255727);
not I_14883 (I255758,I255727);
nand I_14884 (I255582,I255693,I255758);
not I_14885 (I255789,I553629);
nor I_14886 (I255806,I255789,I553620);
and I_14887 (I255823,I255806,I553617);
or I_14888 (I255840,I255823,I553614);
DFFARX1 I_14889  ( .D(I255840), .CLK(I2702), .RSTB(I255608), .Q(I255857) );
nor I_14890 (I255874,I255857,I255710);
DFFARX1 I_14891  ( .D(I255857), .CLK(I2702), .RSTB(I255608), .Q(I255891) );
not I_14892 (I255579,I255891);
nand I_14893 (I255922,I255625,I553629);
and I_14894 (I255939,I255922,I255874);
DFFARX1 I_14895  ( .D(I255922), .CLK(I2702), .RSTB(I255608), .Q(I255576) );
DFFARX1 I_14896  ( .D(I553638), .CLK(I2702), .RSTB(I255608), .Q(I255970) );
nor I_14897 (I255987,I255970,I255693);
nand I_14898 (I255594,I255857,I255987);
nor I_14899 (I256018,I255970,I255758);
not I_14900 (I255591,I255970);
nand I_14901 (I256049,I255970,I255659);
and I_14902 (I256066,I255727,I256049);
DFFARX1 I_14903  ( .D(I256066), .CLK(I2702), .RSTB(I255608), .Q(I255570) );
DFFARX1 I_14904  ( .D(I255970), .CLK(I2702), .RSTB(I255608), .Q(I255573) );
DFFARX1 I_14905  ( .D(I553626), .CLK(I2702), .RSTB(I255608), .Q(I256111) );
not I_14906 (I256128,I256111);
nand I_14907 (I256145,I256128,I255693);
and I_14908 (I256162,I255922,I256145);
DFFARX1 I_14909  ( .D(I256162), .CLK(I2702), .RSTB(I255608), .Q(I255600) );
or I_14910 (I256193,I256128,I255939);
DFFARX1 I_14911  ( .D(I256193), .CLK(I2702), .RSTB(I255608), .Q(I255585) );
nand I_14912 (I255588,I256128,I256018);
not I_14913 (I256271,I2709);
not I_14914 (I256288,I348657);
nor I_14915 (I256305,I348654,I348672);
nand I_14916 (I256322,I256305,I348675);
nor I_14917 (I256339,I256288,I348654);
nand I_14918 (I256356,I256339,I348660);
not I_14919 (I256373,I256356);
not I_14920 (I256390,I348654);
nor I_14921 (I256260,I256356,I256390);
not I_14922 (I256421,I256390);
nand I_14923 (I256245,I256356,I256421);
not I_14924 (I256452,I348669);
nor I_14925 (I256469,I256452,I348651);
and I_14926 (I256486,I256469,I348645);
or I_14927 (I256503,I256486,I348663);
DFFARX1 I_14928  ( .D(I256503), .CLK(I2702), .RSTB(I256271), .Q(I256520) );
nor I_14929 (I256537,I256520,I256373);
DFFARX1 I_14930  ( .D(I256520), .CLK(I2702), .RSTB(I256271), .Q(I256554) );
not I_14931 (I256242,I256554);
nand I_14932 (I256585,I256288,I348669);
and I_14933 (I256602,I256585,I256537);
DFFARX1 I_14934  ( .D(I256585), .CLK(I2702), .RSTB(I256271), .Q(I256239) );
DFFARX1 I_14935  ( .D(I348648), .CLK(I2702), .RSTB(I256271), .Q(I256633) );
nor I_14936 (I256650,I256633,I256356);
nand I_14937 (I256257,I256520,I256650);
nor I_14938 (I256681,I256633,I256421);
not I_14939 (I256254,I256633);
nand I_14940 (I256712,I256633,I256322);
and I_14941 (I256729,I256390,I256712);
DFFARX1 I_14942  ( .D(I256729), .CLK(I2702), .RSTB(I256271), .Q(I256233) );
DFFARX1 I_14943  ( .D(I256633), .CLK(I2702), .RSTB(I256271), .Q(I256236) );
DFFARX1 I_14944  ( .D(I348666), .CLK(I2702), .RSTB(I256271), .Q(I256774) );
not I_14945 (I256791,I256774);
nand I_14946 (I256808,I256791,I256356);
and I_14947 (I256825,I256585,I256808);
DFFARX1 I_14948  ( .D(I256825), .CLK(I2702), .RSTB(I256271), .Q(I256263) );
or I_14949 (I256856,I256791,I256602);
DFFARX1 I_14950  ( .D(I256856), .CLK(I2702), .RSTB(I256271), .Q(I256248) );
nand I_14951 (I256251,I256791,I256681);
not I_14952 (I256934,I2709);
not I_14953 (I256951,I113065);
nor I_14954 (I256968,I113062,I113086);
nand I_14955 (I256985,I256968,I113083);
nor I_14956 (I257002,I256951,I113062);
nand I_14957 (I257019,I257002,I113089);
not I_14958 (I257036,I257019);
not I_14959 (I257053,I113062);
nor I_14960 (I256923,I257019,I257053);
not I_14961 (I257084,I257053);
nand I_14962 (I256908,I257019,I257084);
not I_14963 (I257115,I113080);
nor I_14964 (I257132,I257115,I113071);
and I_14965 (I257149,I257132,I113068);
or I_14966 (I257166,I257149,I113077);
DFFARX1 I_14967  ( .D(I257166), .CLK(I2702), .RSTB(I256934), .Q(I257183) );
nor I_14968 (I257200,I257183,I257036);
DFFARX1 I_14969  ( .D(I257183), .CLK(I2702), .RSTB(I256934), .Q(I257217) );
not I_14970 (I256905,I257217);
nand I_14971 (I257248,I256951,I113080);
and I_14972 (I257265,I257248,I257200);
DFFARX1 I_14973  ( .D(I257248), .CLK(I2702), .RSTB(I256934), .Q(I256902) );
DFFARX1 I_14974  ( .D(I113059), .CLK(I2702), .RSTB(I256934), .Q(I257296) );
nor I_14975 (I257313,I257296,I257019);
nand I_14976 (I256920,I257183,I257313);
nor I_14977 (I257344,I257296,I257084);
not I_14978 (I256917,I257296);
nand I_14979 (I257375,I257296,I256985);
and I_14980 (I257392,I257053,I257375);
DFFARX1 I_14981  ( .D(I257392), .CLK(I2702), .RSTB(I256934), .Q(I256896) );
DFFARX1 I_14982  ( .D(I257296), .CLK(I2702), .RSTB(I256934), .Q(I256899) );
DFFARX1 I_14983  ( .D(I113074), .CLK(I2702), .RSTB(I256934), .Q(I257437) );
not I_14984 (I257454,I257437);
nand I_14985 (I257471,I257454,I257019);
and I_14986 (I257488,I257248,I257471);
DFFARX1 I_14987  ( .D(I257488), .CLK(I2702), .RSTB(I256934), .Q(I256926) );
or I_14988 (I257519,I257454,I257265);
DFFARX1 I_14989  ( .D(I257519), .CLK(I2702), .RSTB(I256934), .Q(I256911) );
nand I_14990 (I256914,I257454,I257344);
not I_14991 (I257597,I2709);
not I_14992 (I257614,I242150);
nor I_14993 (I257631,I242123,I242126);
nand I_14994 (I257648,I257631,I242138);
nor I_14995 (I257665,I257614,I242123);
nand I_14996 (I257682,I257665,I242144);
not I_14997 (I257699,I257682);
not I_14998 (I257716,I242123);
nor I_14999 (I257586,I257682,I257716);
not I_15000 (I257747,I257716);
nand I_15001 (I257571,I257682,I257747);
not I_15002 (I257778,I242147);
nor I_15003 (I257795,I257778,I242129);
and I_15004 (I257812,I257795,I242132);
or I_15005 (I257829,I257812,I242153);
DFFARX1 I_15006  ( .D(I257829), .CLK(I2702), .RSTB(I257597), .Q(I257846) );
nor I_15007 (I257863,I257846,I257699);
DFFARX1 I_15008  ( .D(I257846), .CLK(I2702), .RSTB(I257597), .Q(I257880) );
not I_15009 (I257568,I257880);
nand I_15010 (I257911,I257614,I242147);
and I_15011 (I257928,I257911,I257863);
DFFARX1 I_15012  ( .D(I257911), .CLK(I2702), .RSTB(I257597), .Q(I257565) );
DFFARX1 I_15013  ( .D(I242135), .CLK(I2702), .RSTB(I257597), .Q(I257959) );
nor I_15014 (I257976,I257959,I257682);
nand I_15015 (I257583,I257846,I257976);
nor I_15016 (I258007,I257959,I257747);
not I_15017 (I257580,I257959);
nand I_15018 (I258038,I257959,I257648);
and I_15019 (I258055,I257716,I258038);
DFFARX1 I_15020  ( .D(I258055), .CLK(I2702), .RSTB(I257597), .Q(I257559) );
DFFARX1 I_15021  ( .D(I257959), .CLK(I2702), .RSTB(I257597), .Q(I257562) );
DFFARX1 I_15022  ( .D(I242141), .CLK(I2702), .RSTB(I257597), .Q(I258100) );
not I_15023 (I258117,I258100);
nand I_15024 (I258134,I258117,I257682);
and I_15025 (I258151,I257911,I258134);
DFFARX1 I_15026  ( .D(I258151), .CLK(I2702), .RSTB(I257597), .Q(I257589) );
or I_15027 (I258182,I258117,I257928);
DFFARX1 I_15028  ( .D(I258182), .CLK(I2702), .RSTB(I257597), .Q(I257574) );
nand I_15029 (I257577,I258117,I258007);
not I_15030 (I258260,I2709);
not I_15031 (I258277,I636954);
nor I_15032 (I258294,I636972,I636963);
nand I_15033 (I258311,I258294,I636969);
nor I_15034 (I258328,I258277,I636972);
nand I_15035 (I258345,I258328,I636975);
not I_15036 (I258362,I258345);
not I_15037 (I258379,I636972);
nor I_15038 (I258249,I258345,I258379);
not I_15039 (I258410,I258379);
nand I_15040 (I258234,I258345,I258410);
not I_15041 (I258441,I636951);
nor I_15042 (I258458,I258441,I636966);
and I_15043 (I258475,I258458,I636948);
or I_15044 (I258492,I258475,I636957);
DFFARX1 I_15045  ( .D(I258492), .CLK(I2702), .RSTB(I258260), .Q(I258509) );
nor I_15046 (I258526,I258509,I258362);
DFFARX1 I_15047  ( .D(I258509), .CLK(I2702), .RSTB(I258260), .Q(I258543) );
not I_15048 (I258231,I258543);
nand I_15049 (I258574,I258277,I636951);
and I_15050 (I258591,I258574,I258526);
DFFARX1 I_15051  ( .D(I258574), .CLK(I2702), .RSTB(I258260), .Q(I258228) );
DFFARX1 I_15052  ( .D(I636960), .CLK(I2702), .RSTB(I258260), .Q(I258622) );
nor I_15053 (I258639,I258622,I258345);
nand I_15054 (I258246,I258509,I258639);
nor I_15055 (I258670,I258622,I258410);
not I_15056 (I258243,I258622);
nand I_15057 (I258701,I258622,I258311);
and I_15058 (I258718,I258379,I258701);
DFFARX1 I_15059  ( .D(I258718), .CLK(I2702), .RSTB(I258260), .Q(I258222) );
DFFARX1 I_15060  ( .D(I258622), .CLK(I2702), .RSTB(I258260), .Q(I258225) );
DFFARX1 I_15061  ( .D(I636978), .CLK(I2702), .RSTB(I258260), .Q(I258763) );
not I_15062 (I258780,I258763);
nand I_15063 (I258797,I258780,I258345);
and I_15064 (I258814,I258574,I258797);
DFFARX1 I_15065  ( .D(I258814), .CLK(I2702), .RSTB(I258260), .Q(I258252) );
or I_15066 (I258845,I258780,I258591);
DFFARX1 I_15067  ( .D(I258845), .CLK(I2702), .RSTB(I258260), .Q(I258237) );
nand I_15068 (I258240,I258780,I258670);
not I_15069 (I258923,I2709);
not I_15070 (I258940,I22365);
nor I_15071 (I258957,I22371,I22374);
nand I_15072 (I258974,I258957,I22350);
nor I_15073 (I258991,I258940,I22371);
nand I_15074 (I259008,I258991,I22359);
not I_15075 (I259025,I259008);
not I_15076 (I259042,I22371);
nor I_15077 (I258912,I259008,I259042);
not I_15078 (I259073,I259042);
nand I_15079 (I258897,I259008,I259073);
not I_15080 (I259104,I22353);
nor I_15081 (I259121,I259104,I22377);
and I_15082 (I259138,I259121,I22347);
or I_15083 (I259155,I259138,I22356);
DFFARX1 I_15084  ( .D(I259155), .CLK(I2702), .RSTB(I258923), .Q(I259172) );
nor I_15085 (I259189,I259172,I259025);
DFFARX1 I_15086  ( .D(I259172), .CLK(I2702), .RSTB(I258923), .Q(I259206) );
not I_15087 (I258894,I259206);
nand I_15088 (I259237,I258940,I22353);
and I_15089 (I259254,I259237,I259189);
DFFARX1 I_15090  ( .D(I259237), .CLK(I2702), .RSTB(I258923), .Q(I258891) );
DFFARX1 I_15091  ( .D(I22362), .CLK(I2702), .RSTB(I258923), .Q(I259285) );
nor I_15092 (I259302,I259285,I259008);
nand I_15093 (I258909,I259172,I259302);
nor I_15094 (I259333,I259285,I259073);
not I_15095 (I258906,I259285);
nand I_15096 (I259364,I259285,I258974);
and I_15097 (I259381,I259042,I259364);
DFFARX1 I_15098  ( .D(I259381), .CLK(I2702), .RSTB(I258923), .Q(I258885) );
DFFARX1 I_15099  ( .D(I259285), .CLK(I2702), .RSTB(I258923), .Q(I258888) );
DFFARX1 I_15100  ( .D(I22368), .CLK(I2702), .RSTB(I258923), .Q(I259426) );
not I_15101 (I259443,I259426);
nand I_15102 (I259460,I259443,I259008);
and I_15103 (I259477,I259237,I259460);
DFFARX1 I_15104  ( .D(I259477), .CLK(I2702), .RSTB(I258923), .Q(I258915) );
or I_15105 (I259508,I259443,I259254);
DFFARX1 I_15106  ( .D(I259508), .CLK(I2702), .RSTB(I258923), .Q(I258900) );
nand I_15107 (I258903,I259443,I259333);
not I_15108 (I259586,I2709);
not I_15109 (I259603,I510197);
nor I_15110 (I259620,I510206,I510188);
nand I_15111 (I259637,I259620,I510209);
nor I_15112 (I259654,I259603,I510206);
nand I_15113 (I259671,I259654,I510200);
not I_15114 (I259688,I259671);
not I_15115 (I259705,I510206);
nor I_15116 (I259575,I259671,I259705);
not I_15117 (I259736,I259705);
nand I_15118 (I259560,I259671,I259736);
not I_15119 (I259767,I510194);
nor I_15120 (I259784,I259767,I510185);
and I_15121 (I259801,I259784,I510182);
or I_15122 (I259818,I259801,I510179);
DFFARX1 I_15123  ( .D(I259818), .CLK(I2702), .RSTB(I259586), .Q(I259835) );
nor I_15124 (I259852,I259835,I259688);
DFFARX1 I_15125  ( .D(I259835), .CLK(I2702), .RSTB(I259586), .Q(I259869) );
not I_15126 (I259557,I259869);
nand I_15127 (I259900,I259603,I510194);
and I_15128 (I259917,I259900,I259852);
DFFARX1 I_15129  ( .D(I259900), .CLK(I2702), .RSTB(I259586), .Q(I259554) );
DFFARX1 I_15130  ( .D(I510203), .CLK(I2702), .RSTB(I259586), .Q(I259948) );
nor I_15131 (I259965,I259948,I259671);
nand I_15132 (I259572,I259835,I259965);
nor I_15133 (I259996,I259948,I259736);
not I_15134 (I259569,I259948);
nand I_15135 (I260027,I259948,I259637);
and I_15136 (I260044,I259705,I260027);
DFFARX1 I_15137  ( .D(I260044), .CLK(I2702), .RSTB(I259586), .Q(I259548) );
DFFARX1 I_15138  ( .D(I259948), .CLK(I2702), .RSTB(I259586), .Q(I259551) );
DFFARX1 I_15139  ( .D(I510191), .CLK(I2702), .RSTB(I259586), .Q(I260089) );
not I_15140 (I260106,I260089);
nand I_15141 (I260123,I260106,I259671);
and I_15142 (I260140,I259900,I260123);
DFFARX1 I_15143  ( .D(I260140), .CLK(I2702), .RSTB(I259586), .Q(I259578) );
or I_15144 (I260171,I260106,I259917);
DFFARX1 I_15145  ( .D(I260171), .CLK(I2702), .RSTB(I259586), .Q(I259563) );
nand I_15146 (I259566,I260106,I259996);
not I_15147 (I260249,I2709);
not I_15148 (I260266,I13950);
nor I_15149 (I260283,I13956,I13959);
nand I_15150 (I260300,I260283,I13935);
nor I_15151 (I260317,I260266,I13956);
nand I_15152 (I260334,I260317,I13944);
not I_15153 (I260351,I260334);
not I_15154 (I260368,I13956);
nor I_15155 (I260238,I260334,I260368);
not I_15156 (I260399,I260368);
nand I_15157 (I260223,I260334,I260399);
not I_15158 (I260430,I13938);
nor I_15159 (I260447,I260430,I13962);
and I_15160 (I260464,I260447,I13932);
or I_15161 (I260481,I260464,I13941);
DFFARX1 I_15162  ( .D(I260481), .CLK(I2702), .RSTB(I260249), .Q(I260498) );
nor I_15163 (I260515,I260498,I260351);
DFFARX1 I_15164  ( .D(I260498), .CLK(I2702), .RSTB(I260249), .Q(I260532) );
not I_15165 (I260220,I260532);
nand I_15166 (I260563,I260266,I13938);
and I_15167 (I260580,I260563,I260515);
DFFARX1 I_15168  ( .D(I260563), .CLK(I2702), .RSTB(I260249), .Q(I260217) );
DFFARX1 I_15169  ( .D(I13947), .CLK(I2702), .RSTB(I260249), .Q(I260611) );
nor I_15170 (I260628,I260611,I260334);
nand I_15171 (I260235,I260498,I260628);
nor I_15172 (I260659,I260611,I260399);
not I_15173 (I260232,I260611);
nand I_15174 (I260690,I260611,I260300);
and I_15175 (I260707,I260368,I260690);
DFFARX1 I_15176  ( .D(I260707), .CLK(I2702), .RSTB(I260249), .Q(I260211) );
DFFARX1 I_15177  ( .D(I260611), .CLK(I2702), .RSTB(I260249), .Q(I260214) );
DFFARX1 I_15178  ( .D(I13953), .CLK(I2702), .RSTB(I260249), .Q(I260752) );
not I_15179 (I260769,I260752);
nand I_15180 (I260786,I260769,I260334);
and I_15181 (I260803,I260563,I260786);
DFFARX1 I_15182  ( .D(I260803), .CLK(I2702), .RSTB(I260249), .Q(I260241) );
or I_15183 (I260834,I260769,I260580);
DFFARX1 I_15184  ( .D(I260834), .CLK(I2702), .RSTB(I260249), .Q(I260226) );
nand I_15185 (I260229,I260769,I260659);
not I_15186 (I260912,I2709);
not I_15187 (I260929,I163416);
nor I_15188 (I260946,I163422,I163428);
nand I_15189 (I260963,I260946,I163431);
nor I_15190 (I260980,I260929,I163422);
nand I_15191 (I260997,I260980,I163413);
not I_15192 (I261014,I260997);
not I_15193 (I261031,I163422);
nor I_15194 (I260901,I260997,I261031);
not I_15195 (I261062,I261031);
nand I_15196 (I260886,I260997,I261062);
not I_15197 (I261093,I163425);
nor I_15198 (I261110,I261093,I163419);
and I_15199 (I261127,I261110,I163434);
or I_15200 (I261144,I261127,I163440);
DFFARX1 I_15201  ( .D(I261144), .CLK(I2702), .RSTB(I260912), .Q(I261161) );
nor I_15202 (I261178,I261161,I261014);
DFFARX1 I_15203  ( .D(I261161), .CLK(I2702), .RSTB(I260912), .Q(I261195) );
not I_15204 (I260883,I261195);
nand I_15205 (I261226,I260929,I163425);
and I_15206 (I261243,I261226,I261178);
DFFARX1 I_15207  ( .D(I261226), .CLK(I2702), .RSTB(I260912), .Q(I260880) );
DFFARX1 I_15208  ( .D(I163437), .CLK(I2702), .RSTB(I260912), .Q(I261274) );
nor I_15209 (I261291,I261274,I260997);
nand I_15210 (I260898,I261161,I261291);
nor I_15211 (I261322,I261274,I261062);
not I_15212 (I260895,I261274);
nand I_15213 (I261353,I261274,I260963);
and I_15214 (I261370,I261031,I261353);
DFFARX1 I_15215  ( .D(I261370), .CLK(I2702), .RSTB(I260912), .Q(I260874) );
DFFARX1 I_15216  ( .D(I261274), .CLK(I2702), .RSTB(I260912), .Q(I260877) );
DFFARX1 I_15217  ( .D(I163443), .CLK(I2702), .RSTB(I260912), .Q(I261415) );
not I_15218 (I261432,I261415);
nand I_15219 (I261449,I261432,I260997);
and I_15220 (I261466,I261226,I261449);
DFFARX1 I_15221  ( .D(I261466), .CLK(I2702), .RSTB(I260912), .Q(I260904) );
or I_15222 (I261497,I261432,I261243);
DFFARX1 I_15223  ( .D(I261497), .CLK(I2702), .RSTB(I260912), .Q(I260889) );
nand I_15224 (I260892,I261432,I261322);
not I_15225 (I261575,I2709);
not I_15226 (I261592,I1279);
nor I_15227 (I261609,I1799,I1991);
nand I_15228 (I261626,I261609,I2487);
nor I_15229 (I261643,I261592,I1799);
nand I_15230 (I261660,I261643,I1807);
not I_15231 (I261677,I261660);
not I_15232 (I261694,I1799);
nor I_15233 (I261564,I261660,I261694);
not I_15234 (I261725,I261694);
nand I_15235 (I261549,I261660,I261725);
not I_15236 (I261756,I1503);
nor I_15237 (I261773,I261756,I2327);
and I_15238 (I261790,I261773,I1727);
or I_15239 (I261807,I261790,I1839);
DFFARX1 I_15240  ( .D(I261807), .CLK(I2702), .RSTB(I261575), .Q(I261824) );
nor I_15241 (I261841,I261824,I261677);
DFFARX1 I_15242  ( .D(I261824), .CLK(I2702), .RSTB(I261575), .Q(I261858) );
not I_15243 (I261546,I261858);
nand I_15244 (I261889,I261592,I1503);
and I_15245 (I261906,I261889,I261841);
DFFARX1 I_15246  ( .D(I261889), .CLK(I2702), .RSTB(I261575), .Q(I261543) );
DFFARX1 I_15247  ( .D(I1439), .CLK(I2702), .RSTB(I261575), .Q(I261937) );
nor I_15248 (I261954,I261937,I261660);
nand I_15249 (I261561,I261824,I261954);
nor I_15250 (I261985,I261937,I261725);
not I_15251 (I261558,I261937);
nand I_15252 (I262016,I261937,I261626);
and I_15253 (I262033,I261694,I262016);
DFFARX1 I_15254  ( .D(I262033), .CLK(I2702), .RSTB(I261575), .Q(I261537) );
DFFARX1 I_15255  ( .D(I261937), .CLK(I2702), .RSTB(I261575), .Q(I261540) );
DFFARX1 I_15256  ( .D(I1567), .CLK(I2702), .RSTB(I261575), .Q(I262078) );
not I_15257 (I262095,I262078);
nand I_15258 (I262112,I262095,I261660);
and I_15259 (I262129,I261889,I262112);
DFFARX1 I_15260  ( .D(I262129), .CLK(I2702), .RSTB(I261575), .Q(I261567) );
or I_15261 (I262160,I262095,I261906);
DFFARX1 I_15262  ( .D(I262160), .CLK(I2702), .RSTB(I261575), .Q(I261552) );
nand I_15263 (I261555,I262095,I261985);
not I_15264 (I262238,I2709);
not I_15265 (I262255,I507222);
nor I_15266 (I262272,I507231,I507213);
nand I_15267 (I262289,I262272,I507234);
nor I_15268 (I262306,I262255,I507231);
nand I_15269 (I262323,I262306,I507225);
not I_15270 (I262340,I262323);
not I_15271 (I262357,I507231);
nor I_15272 (I262227,I262323,I262357);
not I_15273 (I262388,I262357);
nand I_15274 (I262212,I262323,I262388);
not I_15275 (I262419,I507219);
nor I_15276 (I262436,I262419,I507210);
and I_15277 (I262453,I262436,I507207);
or I_15278 (I262470,I262453,I507204);
DFFARX1 I_15279  ( .D(I262470), .CLK(I2702), .RSTB(I262238), .Q(I262487) );
nor I_15280 (I262504,I262487,I262340);
DFFARX1 I_15281  ( .D(I262487), .CLK(I2702), .RSTB(I262238), .Q(I262521) );
not I_15282 (I262209,I262521);
nand I_15283 (I262552,I262255,I507219);
and I_15284 (I262569,I262552,I262504);
DFFARX1 I_15285  ( .D(I262552), .CLK(I2702), .RSTB(I262238), .Q(I262206) );
DFFARX1 I_15286  ( .D(I507228), .CLK(I2702), .RSTB(I262238), .Q(I262600) );
nor I_15287 (I262617,I262600,I262323);
nand I_15288 (I262224,I262487,I262617);
nor I_15289 (I262648,I262600,I262388);
not I_15290 (I262221,I262600);
nand I_15291 (I262679,I262600,I262289);
and I_15292 (I262696,I262357,I262679);
DFFARX1 I_15293  ( .D(I262696), .CLK(I2702), .RSTB(I262238), .Q(I262200) );
DFFARX1 I_15294  ( .D(I262600), .CLK(I2702), .RSTB(I262238), .Q(I262203) );
DFFARX1 I_15295  ( .D(I507216), .CLK(I2702), .RSTB(I262238), .Q(I262741) );
not I_15296 (I262758,I262741);
nand I_15297 (I262775,I262758,I262323);
and I_15298 (I262792,I262552,I262775);
DFFARX1 I_15299  ( .D(I262792), .CLK(I2702), .RSTB(I262238), .Q(I262230) );
or I_15300 (I262823,I262758,I262569);
DFFARX1 I_15301  ( .D(I262823), .CLK(I2702), .RSTB(I262238), .Q(I262215) );
nand I_15302 (I262218,I262758,I262648);
not I_15303 (I262901,I2709);
not I_15304 (I262918,I105313);
nor I_15305 (I262935,I105310,I105334);
nand I_15306 (I262952,I262935,I105331);
nor I_15307 (I262969,I262918,I105310);
nand I_15308 (I262986,I262969,I105337);
not I_15309 (I263003,I262986);
not I_15310 (I263020,I105310);
nor I_15311 (I262890,I262986,I263020);
not I_15312 (I263051,I263020);
nand I_15313 (I262875,I262986,I263051);
not I_15314 (I263082,I105328);
nor I_15315 (I263099,I263082,I105319);
and I_15316 (I263116,I263099,I105316);
or I_15317 (I263133,I263116,I105325);
DFFARX1 I_15318  ( .D(I263133), .CLK(I2702), .RSTB(I262901), .Q(I263150) );
nor I_15319 (I263167,I263150,I263003);
DFFARX1 I_15320  ( .D(I263150), .CLK(I2702), .RSTB(I262901), .Q(I263184) );
not I_15321 (I262872,I263184);
nand I_15322 (I263215,I262918,I105328);
and I_15323 (I263232,I263215,I263167);
DFFARX1 I_15324  ( .D(I263215), .CLK(I2702), .RSTB(I262901), .Q(I262869) );
DFFARX1 I_15325  ( .D(I105307), .CLK(I2702), .RSTB(I262901), .Q(I263263) );
nor I_15326 (I263280,I263263,I262986);
nand I_15327 (I262887,I263150,I263280);
nor I_15328 (I263311,I263263,I263051);
not I_15329 (I262884,I263263);
nand I_15330 (I263342,I263263,I262952);
and I_15331 (I263359,I263020,I263342);
DFFARX1 I_15332  ( .D(I263359), .CLK(I2702), .RSTB(I262901), .Q(I262863) );
DFFARX1 I_15333  ( .D(I263263), .CLK(I2702), .RSTB(I262901), .Q(I262866) );
DFFARX1 I_15334  ( .D(I105322), .CLK(I2702), .RSTB(I262901), .Q(I263404) );
not I_15335 (I263421,I263404);
nand I_15336 (I263438,I263421,I262986);
and I_15337 (I263455,I263215,I263438);
DFFARX1 I_15338  ( .D(I263455), .CLK(I2702), .RSTB(I262901), .Q(I262893) );
or I_15339 (I263486,I263421,I263232);
DFFARX1 I_15340  ( .D(I263486), .CLK(I2702), .RSTB(I262901), .Q(I262878) );
nand I_15341 (I262881,I263421,I263311);
not I_15342 (I263564,I2709);
not I_15343 (I263581,I528642);
nor I_15344 (I263598,I528651,I528633);
nand I_15345 (I263615,I263598,I528654);
nor I_15346 (I263632,I263581,I528651);
nand I_15347 (I263649,I263632,I528645);
not I_15348 (I263666,I263649);
not I_15349 (I263683,I528651);
nor I_15350 (I263553,I263649,I263683);
not I_15351 (I263714,I263683);
nand I_15352 (I263538,I263649,I263714);
not I_15353 (I263745,I528639);
nor I_15354 (I263762,I263745,I528630);
and I_15355 (I263779,I263762,I528627);
or I_15356 (I263796,I263779,I528624);
DFFARX1 I_15357  ( .D(I263796), .CLK(I2702), .RSTB(I263564), .Q(I263813) );
nor I_15358 (I263830,I263813,I263666);
DFFARX1 I_15359  ( .D(I263813), .CLK(I2702), .RSTB(I263564), .Q(I263847) );
not I_15360 (I263535,I263847);
nand I_15361 (I263878,I263581,I528639);
and I_15362 (I263895,I263878,I263830);
DFFARX1 I_15363  ( .D(I263878), .CLK(I2702), .RSTB(I263564), .Q(I263532) );
DFFARX1 I_15364  ( .D(I528648), .CLK(I2702), .RSTB(I263564), .Q(I263926) );
nor I_15365 (I263943,I263926,I263649);
nand I_15366 (I263550,I263813,I263943);
nor I_15367 (I263974,I263926,I263714);
not I_15368 (I263547,I263926);
nand I_15369 (I264005,I263926,I263615);
and I_15370 (I264022,I263683,I264005);
DFFARX1 I_15371  ( .D(I264022), .CLK(I2702), .RSTB(I263564), .Q(I263526) );
DFFARX1 I_15372  ( .D(I263926), .CLK(I2702), .RSTB(I263564), .Q(I263529) );
DFFARX1 I_15373  ( .D(I528636), .CLK(I2702), .RSTB(I263564), .Q(I264067) );
not I_15374 (I264084,I264067);
nand I_15375 (I264101,I264084,I263649);
and I_15376 (I264118,I263878,I264101);
DFFARX1 I_15377  ( .D(I264118), .CLK(I2702), .RSTB(I263564), .Q(I263556) );
or I_15378 (I264149,I264084,I263895);
DFFARX1 I_15379  ( .D(I264149), .CLK(I2702), .RSTB(I263564), .Q(I263541) );
nand I_15380 (I263544,I264084,I263974);
not I_15381 (I264227,I2709);
not I_15382 (I264244,I559582);
nor I_15383 (I264261,I559591,I559573);
nand I_15384 (I264278,I264261,I559594);
nor I_15385 (I264295,I264244,I559591);
nand I_15386 (I264312,I264295,I559585);
not I_15387 (I264329,I264312);
not I_15388 (I264346,I559591);
nor I_15389 (I264216,I264312,I264346);
not I_15390 (I264377,I264346);
nand I_15391 (I264201,I264312,I264377);
not I_15392 (I264408,I559579);
nor I_15393 (I264425,I264408,I559570);
and I_15394 (I264442,I264425,I559567);
or I_15395 (I264459,I264442,I559564);
DFFARX1 I_15396  ( .D(I264459), .CLK(I2702), .RSTB(I264227), .Q(I264476) );
nor I_15397 (I264493,I264476,I264329);
DFFARX1 I_15398  ( .D(I264476), .CLK(I2702), .RSTB(I264227), .Q(I264510) );
not I_15399 (I264198,I264510);
nand I_15400 (I264541,I264244,I559579);
and I_15401 (I264558,I264541,I264493);
DFFARX1 I_15402  ( .D(I264541), .CLK(I2702), .RSTB(I264227), .Q(I264195) );
DFFARX1 I_15403  ( .D(I559588), .CLK(I2702), .RSTB(I264227), .Q(I264589) );
nor I_15404 (I264606,I264589,I264312);
nand I_15405 (I264213,I264476,I264606);
nor I_15406 (I264637,I264589,I264377);
not I_15407 (I264210,I264589);
nand I_15408 (I264668,I264589,I264278);
and I_15409 (I264685,I264346,I264668);
DFFARX1 I_15410  ( .D(I264685), .CLK(I2702), .RSTB(I264227), .Q(I264189) );
DFFARX1 I_15411  ( .D(I264589), .CLK(I2702), .RSTB(I264227), .Q(I264192) );
DFFARX1 I_15412  ( .D(I559576), .CLK(I2702), .RSTB(I264227), .Q(I264730) );
not I_15413 (I264747,I264730);
nand I_15414 (I264764,I264747,I264312);
and I_15415 (I264781,I264541,I264764);
DFFARX1 I_15416  ( .D(I264781), .CLK(I2702), .RSTB(I264227), .Q(I264219) );
or I_15417 (I264812,I264747,I264558);
DFFARX1 I_15418  ( .D(I264812), .CLK(I2702), .RSTB(I264227), .Q(I264204) );
nand I_15419 (I264207,I264747,I264637);
not I_15420 (I264890,I2709);
not I_15421 (I264907,I429095);
nor I_15422 (I264924,I429098,I429104);
nand I_15423 (I264941,I264924,I429110);
nor I_15424 (I264958,I264907,I429098);
nand I_15425 (I264975,I264958,I429089);
not I_15426 (I264992,I264975);
not I_15427 (I265009,I429098);
nor I_15428 (I264879,I264975,I265009);
not I_15429 (I265040,I265009);
nand I_15430 (I264864,I264975,I265040);
not I_15431 (I265071,I429101);
nor I_15432 (I265088,I265071,I429116);
and I_15433 (I265105,I265088,I429119);
or I_15434 (I265122,I265105,I429092);
DFFARX1 I_15435  ( .D(I265122), .CLK(I2702), .RSTB(I264890), .Q(I265139) );
nor I_15436 (I265156,I265139,I264992);
DFFARX1 I_15437  ( .D(I265139), .CLK(I2702), .RSTB(I264890), .Q(I265173) );
not I_15438 (I264861,I265173);
nand I_15439 (I265204,I264907,I429101);
and I_15440 (I265221,I265204,I265156);
DFFARX1 I_15441  ( .D(I265204), .CLK(I2702), .RSTB(I264890), .Q(I264858) );
DFFARX1 I_15442  ( .D(I429113), .CLK(I2702), .RSTB(I264890), .Q(I265252) );
nor I_15443 (I265269,I265252,I264975);
nand I_15444 (I264876,I265139,I265269);
nor I_15445 (I265300,I265252,I265040);
not I_15446 (I264873,I265252);
nand I_15447 (I265331,I265252,I264941);
and I_15448 (I265348,I265009,I265331);
DFFARX1 I_15449  ( .D(I265348), .CLK(I2702), .RSTB(I264890), .Q(I264852) );
DFFARX1 I_15450  ( .D(I265252), .CLK(I2702), .RSTB(I264890), .Q(I264855) );
DFFARX1 I_15451  ( .D(I429107), .CLK(I2702), .RSTB(I264890), .Q(I265393) );
not I_15452 (I265410,I265393);
nand I_15453 (I265427,I265410,I264975);
and I_15454 (I265444,I265204,I265427);
DFFARX1 I_15455  ( .D(I265444), .CLK(I2702), .RSTB(I264890), .Q(I264882) );
or I_15456 (I265475,I265410,I265221);
DFFARX1 I_15457  ( .D(I265475), .CLK(I2702), .RSTB(I264890), .Q(I264867) );
nand I_15458 (I264870,I265410,I265300);
not I_15459 (I265553,I2709);
not I_15460 (I265570,I670920);
nor I_15461 (I265587,I670938,I670929);
nand I_15462 (I265604,I265587,I670935);
nor I_15463 (I265621,I265570,I670938);
nand I_15464 (I265638,I265621,I670941);
not I_15465 (I265655,I265638);
not I_15466 (I265672,I670938);
nor I_15467 (I265542,I265638,I265672);
not I_15468 (I265703,I265672);
nand I_15469 (I265527,I265638,I265703);
not I_15470 (I265734,I670917);
nor I_15471 (I265751,I265734,I670932);
and I_15472 (I265768,I265751,I670914);
or I_15473 (I265785,I265768,I670923);
DFFARX1 I_15474  ( .D(I265785), .CLK(I2702), .RSTB(I265553), .Q(I265802) );
nor I_15475 (I265819,I265802,I265655);
DFFARX1 I_15476  ( .D(I265802), .CLK(I2702), .RSTB(I265553), .Q(I265836) );
not I_15477 (I265524,I265836);
nand I_15478 (I265867,I265570,I670917);
and I_15479 (I265884,I265867,I265819);
DFFARX1 I_15480  ( .D(I265867), .CLK(I2702), .RSTB(I265553), .Q(I265521) );
DFFARX1 I_15481  ( .D(I670926), .CLK(I2702), .RSTB(I265553), .Q(I265915) );
nor I_15482 (I265932,I265915,I265638);
nand I_15483 (I265539,I265802,I265932);
nor I_15484 (I265963,I265915,I265703);
not I_15485 (I265536,I265915);
nand I_15486 (I265994,I265915,I265604);
and I_15487 (I266011,I265672,I265994);
DFFARX1 I_15488  ( .D(I266011), .CLK(I2702), .RSTB(I265553), .Q(I265515) );
DFFARX1 I_15489  ( .D(I265915), .CLK(I2702), .RSTB(I265553), .Q(I265518) );
DFFARX1 I_15490  ( .D(I670944), .CLK(I2702), .RSTB(I265553), .Q(I266056) );
not I_15491 (I266073,I266056);
nand I_15492 (I266090,I266073,I265638);
and I_15493 (I266107,I265867,I266090);
DFFARX1 I_15494  ( .D(I266107), .CLK(I2702), .RSTB(I265553), .Q(I265545) );
or I_15495 (I266138,I266073,I265884);
DFFARX1 I_15496  ( .D(I266138), .CLK(I2702), .RSTB(I265553), .Q(I265530) );
nand I_15497 (I265533,I266073,I265963);
not I_15498 (I266216,I2709);
not I_15499 (I266233,I93685);
nor I_15500 (I266250,I93682,I93706);
nand I_15501 (I266267,I266250,I93703);
nor I_15502 (I266284,I266233,I93682);
nand I_15503 (I266301,I266284,I93709);
not I_15504 (I266318,I266301);
not I_15505 (I266335,I93682);
nor I_15506 (I266205,I266301,I266335);
not I_15507 (I266366,I266335);
nand I_15508 (I266190,I266301,I266366);
not I_15509 (I266397,I93700);
nor I_15510 (I266414,I266397,I93691);
and I_15511 (I266431,I266414,I93688);
or I_15512 (I266448,I266431,I93697);
DFFARX1 I_15513  ( .D(I266448), .CLK(I2702), .RSTB(I266216), .Q(I266465) );
nor I_15514 (I266482,I266465,I266318);
DFFARX1 I_15515  ( .D(I266465), .CLK(I2702), .RSTB(I266216), .Q(I266499) );
not I_15516 (I266187,I266499);
nand I_15517 (I266530,I266233,I93700);
and I_15518 (I266547,I266530,I266482);
DFFARX1 I_15519  ( .D(I266530), .CLK(I2702), .RSTB(I266216), .Q(I266184) );
DFFARX1 I_15520  ( .D(I93679), .CLK(I2702), .RSTB(I266216), .Q(I266578) );
nor I_15521 (I266595,I266578,I266301);
nand I_15522 (I266202,I266465,I266595);
nor I_15523 (I266626,I266578,I266366);
not I_15524 (I266199,I266578);
nand I_15525 (I266657,I266578,I266267);
and I_15526 (I266674,I266335,I266657);
DFFARX1 I_15527  ( .D(I266674), .CLK(I2702), .RSTB(I266216), .Q(I266178) );
DFFARX1 I_15528  ( .D(I266578), .CLK(I2702), .RSTB(I266216), .Q(I266181) );
DFFARX1 I_15529  ( .D(I93694), .CLK(I2702), .RSTB(I266216), .Q(I266719) );
not I_15530 (I266736,I266719);
nand I_15531 (I266753,I266736,I266301);
and I_15532 (I266770,I266530,I266753);
DFFARX1 I_15533  ( .D(I266770), .CLK(I2702), .RSTB(I266216), .Q(I266208) );
or I_15534 (I266801,I266736,I266547);
DFFARX1 I_15535  ( .D(I266801), .CLK(I2702), .RSTB(I266216), .Q(I266193) );
nand I_15536 (I266196,I266736,I266626);
not I_15537 (I266879,I2709);
not I_15538 (I266896,I664001);
nor I_15539 (I266913,I664019,I664010);
nand I_15540 (I266930,I266913,I664016);
nor I_15541 (I266947,I266896,I664019);
nand I_15542 (I266964,I266947,I664022);
not I_15543 (I266981,I266964);
not I_15544 (I266998,I664019);
nor I_15545 (I266868,I266964,I266998);
not I_15546 (I267029,I266998);
nand I_15547 (I266853,I266964,I267029);
not I_15548 (I267060,I663998);
nor I_15549 (I267077,I267060,I664013);
and I_15550 (I267094,I267077,I663995);
or I_15551 (I267111,I267094,I664004);
DFFARX1 I_15552  ( .D(I267111), .CLK(I2702), .RSTB(I266879), .Q(I267128) );
nor I_15553 (I267145,I267128,I266981);
DFFARX1 I_15554  ( .D(I267128), .CLK(I2702), .RSTB(I266879), .Q(I267162) );
not I_15555 (I266850,I267162);
nand I_15556 (I267193,I266896,I663998);
and I_15557 (I267210,I267193,I267145);
DFFARX1 I_15558  ( .D(I267193), .CLK(I2702), .RSTB(I266879), .Q(I266847) );
DFFARX1 I_15559  ( .D(I664007), .CLK(I2702), .RSTB(I266879), .Q(I267241) );
nor I_15560 (I267258,I267241,I266964);
nand I_15561 (I266865,I267128,I267258);
nor I_15562 (I267289,I267241,I267029);
not I_15563 (I266862,I267241);
nand I_15564 (I267320,I267241,I266930);
and I_15565 (I267337,I266998,I267320);
DFFARX1 I_15566  ( .D(I267337), .CLK(I2702), .RSTB(I266879), .Q(I266841) );
DFFARX1 I_15567  ( .D(I267241), .CLK(I2702), .RSTB(I266879), .Q(I266844) );
DFFARX1 I_15568  ( .D(I664025), .CLK(I2702), .RSTB(I266879), .Q(I267382) );
not I_15569 (I267399,I267382);
nand I_15570 (I267416,I267399,I266964);
and I_15571 (I267433,I267193,I267416);
DFFARX1 I_15572  ( .D(I267433), .CLK(I2702), .RSTB(I266879), .Q(I266871) );
or I_15573 (I267464,I267399,I267210);
DFFARX1 I_15574  ( .D(I267464), .CLK(I2702), .RSTB(I266879), .Q(I266856) );
nand I_15575 (I266859,I267399,I267289);
not I_15576 (I267542,I2709);
not I_15577 (I267559,I463342);
nor I_15578 (I267576,I463354,I463336);
nand I_15579 (I267593,I267576,I463357);
nor I_15580 (I267610,I267559,I463354);
nand I_15581 (I267627,I267610,I463348);
not I_15582 (I267644,I267627);
not I_15583 (I267661,I463354);
nor I_15584 (I267531,I267627,I267661);
not I_15585 (I267692,I267661);
nand I_15586 (I267516,I267627,I267692);
not I_15587 (I267723,I463339);
nor I_15588 (I267740,I267723,I463333);
and I_15589 (I267757,I267740,I463345);
or I_15590 (I267774,I267757,I463330);
DFFARX1 I_15591  ( .D(I267774), .CLK(I2702), .RSTB(I267542), .Q(I267791) );
nor I_15592 (I267808,I267791,I267644);
DFFARX1 I_15593  ( .D(I267791), .CLK(I2702), .RSTB(I267542), .Q(I267825) );
not I_15594 (I267513,I267825);
nand I_15595 (I267856,I267559,I463339);
and I_15596 (I267873,I267856,I267808);
DFFARX1 I_15597  ( .D(I267856), .CLK(I2702), .RSTB(I267542), .Q(I267510) );
DFFARX1 I_15598  ( .D(I463327), .CLK(I2702), .RSTB(I267542), .Q(I267904) );
nor I_15599 (I267921,I267904,I267627);
nand I_15600 (I267528,I267791,I267921);
nor I_15601 (I267952,I267904,I267692);
not I_15602 (I267525,I267904);
nand I_15603 (I267983,I267904,I267593);
and I_15604 (I268000,I267661,I267983);
DFFARX1 I_15605  ( .D(I268000), .CLK(I2702), .RSTB(I267542), .Q(I267504) );
DFFARX1 I_15606  ( .D(I267904), .CLK(I2702), .RSTB(I267542), .Q(I267507) );
DFFARX1 I_15607  ( .D(I463351), .CLK(I2702), .RSTB(I267542), .Q(I268045) );
not I_15608 (I268062,I268045);
nand I_15609 (I268079,I268062,I267627);
and I_15610 (I268096,I267856,I268079);
DFFARX1 I_15611  ( .D(I268096), .CLK(I2702), .RSTB(I267542), .Q(I267534) );
or I_15612 (I268127,I268062,I267873);
DFFARX1 I_15613  ( .D(I268127), .CLK(I2702), .RSTB(I267542), .Q(I267519) );
nand I_15614 (I267522,I268062,I267952);
not I_15615 (I268205,I2709);
not I_15616 (I268222,I550657);
nor I_15617 (I268239,I550666,I550648);
nand I_15618 (I268256,I268239,I550669);
nor I_15619 (I268273,I268222,I550666);
nand I_15620 (I268290,I268273,I550660);
not I_15621 (I268307,I268290);
not I_15622 (I268324,I550666);
nor I_15623 (I268194,I268290,I268324);
not I_15624 (I268355,I268324);
nand I_15625 (I268179,I268290,I268355);
not I_15626 (I268386,I550654);
nor I_15627 (I268403,I268386,I550645);
and I_15628 (I268420,I268403,I550642);
or I_15629 (I268437,I268420,I550639);
DFFARX1 I_15630  ( .D(I268437), .CLK(I2702), .RSTB(I268205), .Q(I268454) );
nor I_15631 (I268471,I268454,I268307);
DFFARX1 I_15632  ( .D(I268454), .CLK(I2702), .RSTB(I268205), .Q(I268488) );
not I_15633 (I268176,I268488);
nand I_15634 (I268519,I268222,I550654);
and I_15635 (I268536,I268519,I268471);
DFFARX1 I_15636  ( .D(I268519), .CLK(I2702), .RSTB(I268205), .Q(I268173) );
DFFARX1 I_15637  ( .D(I550663), .CLK(I2702), .RSTB(I268205), .Q(I268567) );
nor I_15638 (I268584,I268567,I268290);
nand I_15639 (I268191,I268454,I268584);
nor I_15640 (I268615,I268567,I268355);
not I_15641 (I268188,I268567);
nand I_15642 (I268646,I268567,I268256);
and I_15643 (I268663,I268324,I268646);
DFFARX1 I_15644  ( .D(I268663), .CLK(I2702), .RSTB(I268205), .Q(I268167) );
DFFARX1 I_15645  ( .D(I268567), .CLK(I2702), .RSTB(I268205), .Q(I268170) );
DFFARX1 I_15646  ( .D(I550651), .CLK(I2702), .RSTB(I268205), .Q(I268708) );
not I_15647 (I268725,I268708);
nand I_15648 (I268742,I268725,I268290);
and I_15649 (I268759,I268519,I268742);
DFFARX1 I_15650  ( .D(I268759), .CLK(I2702), .RSTB(I268205), .Q(I268197) );
or I_15651 (I268790,I268725,I268536);
DFFARX1 I_15652  ( .D(I268790), .CLK(I2702), .RSTB(I268205), .Q(I268182) );
nand I_15653 (I268185,I268725,I268615);
not I_15654 (I268868,I2709);
not I_15655 (I268885,I722742);
nor I_15656 (I268902,I722733,I722739);
nand I_15657 (I268919,I268902,I722751);
nor I_15658 (I268936,I268885,I722733);
nand I_15659 (I268953,I268936,I722736);
not I_15660 (I268970,I268953);
not I_15661 (I268987,I722733);
nor I_15662 (I268857,I268953,I268987);
not I_15663 (I269018,I268987);
nand I_15664 (I268842,I268953,I269018);
not I_15665 (I269049,I722760);
nor I_15666 (I269066,I269049,I722754);
and I_15667 (I269083,I269066,I722745);
or I_15668 (I269100,I269083,I722730);
DFFARX1 I_15669  ( .D(I269100), .CLK(I2702), .RSTB(I268868), .Q(I269117) );
nor I_15670 (I269134,I269117,I268970);
DFFARX1 I_15671  ( .D(I269117), .CLK(I2702), .RSTB(I268868), .Q(I269151) );
not I_15672 (I268839,I269151);
nand I_15673 (I269182,I268885,I722760);
and I_15674 (I269199,I269182,I269134);
DFFARX1 I_15675  ( .D(I269182), .CLK(I2702), .RSTB(I268868), .Q(I268836) );
DFFARX1 I_15676  ( .D(I722748), .CLK(I2702), .RSTB(I268868), .Q(I269230) );
nor I_15677 (I269247,I269230,I268953);
nand I_15678 (I268854,I269117,I269247);
nor I_15679 (I269278,I269230,I269018);
not I_15680 (I268851,I269230);
nand I_15681 (I269309,I269230,I268919);
and I_15682 (I269326,I268987,I269309);
DFFARX1 I_15683  ( .D(I269326), .CLK(I2702), .RSTB(I268868), .Q(I268830) );
DFFARX1 I_15684  ( .D(I269230), .CLK(I2702), .RSTB(I268868), .Q(I268833) );
DFFARX1 I_15685  ( .D(I722757), .CLK(I2702), .RSTB(I268868), .Q(I269371) );
not I_15686 (I269388,I269371);
nand I_15687 (I269405,I269388,I268953);
and I_15688 (I269422,I269182,I269405);
DFFARX1 I_15689  ( .D(I269422), .CLK(I2702), .RSTB(I268868), .Q(I268860) );
or I_15690 (I269453,I269388,I269199);
DFFARX1 I_15691  ( .D(I269453), .CLK(I2702), .RSTB(I268868), .Q(I268845) );
nand I_15692 (I268848,I269388,I269278);
not I_15693 (I269531,I2709);
not I_15694 (I269548,I579217);
nor I_15695 (I269565,I579214,I579205);
nand I_15696 (I269582,I269565,I579208);
nor I_15697 (I269599,I269548,I579214);
nand I_15698 (I269616,I269599,I579202);
not I_15699 (I269633,I269616);
not I_15700 (I269650,I579214);
nor I_15701 (I269520,I269616,I269650);
not I_15702 (I269681,I269650);
nand I_15703 (I269505,I269616,I269681);
not I_15704 (I269712,I579223);
nor I_15705 (I269729,I269712,I579226);
and I_15706 (I269746,I269729,I579211);
or I_15707 (I269763,I269746,I579199);
DFFARX1 I_15708  ( .D(I269763), .CLK(I2702), .RSTB(I269531), .Q(I269780) );
nor I_15709 (I269797,I269780,I269633);
DFFARX1 I_15710  ( .D(I269780), .CLK(I2702), .RSTB(I269531), .Q(I269814) );
not I_15711 (I269502,I269814);
nand I_15712 (I269845,I269548,I579223);
and I_15713 (I269862,I269845,I269797);
DFFARX1 I_15714  ( .D(I269845), .CLK(I2702), .RSTB(I269531), .Q(I269499) );
DFFARX1 I_15715  ( .D(I579220), .CLK(I2702), .RSTB(I269531), .Q(I269893) );
nor I_15716 (I269910,I269893,I269616);
nand I_15717 (I269517,I269780,I269910);
nor I_15718 (I269941,I269893,I269681);
not I_15719 (I269514,I269893);
nand I_15720 (I269972,I269893,I269582);
and I_15721 (I269989,I269650,I269972);
DFFARX1 I_15722  ( .D(I269989), .CLK(I2702), .RSTB(I269531), .Q(I269493) );
DFFARX1 I_15723  ( .D(I269893), .CLK(I2702), .RSTB(I269531), .Q(I269496) );
DFFARX1 I_15724  ( .D(I579229), .CLK(I2702), .RSTB(I269531), .Q(I270034) );
not I_15725 (I270051,I270034);
nand I_15726 (I270068,I270051,I269616);
and I_15727 (I270085,I269845,I270068);
DFFARX1 I_15728  ( .D(I270085), .CLK(I2702), .RSTB(I269531), .Q(I269523) );
or I_15729 (I270116,I270051,I269862);
DFFARX1 I_15730  ( .D(I270116), .CLK(I2702), .RSTB(I269531), .Q(I269508) );
nand I_15731 (I269511,I270051,I269941);
not I_15732 (I270194,I2709);
not I_15733 (I270211,I78827);
nor I_15734 (I270228,I78824,I78848);
nand I_15735 (I270245,I270228,I78845);
nor I_15736 (I270262,I270211,I78824);
nand I_15737 (I270279,I270262,I78851);
not I_15738 (I270296,I270279);
not I_15739 (I270313,I78824);
nor I_15740 (I270183,I270279,I270313);
not I_15741 (I270344,I270313);
nand I_15742 (I270168,I270279,I270344);
not I_15743 (I270375,I78842);
nor I_15744 (I270392,I270375,I78833);
and I_15745 (I270409,I270392,I78830);
or I_15746 (I270426,I270409,I78839);
DFFARX1 I_15747  ( .D(I270426), .CLK(I2702), .RSTB(I270194), .Q(I270443) );
nor I_15748 (I270460,I270443,I270296);
DFFARX1 I_15749  ( .D(I270443), .CLK(I2702), .RSTB(I270194), .Q(I270477) );
not I_15750 (I270165,I270477);
nand I_15751 (I270508,I270211,I78842);
and I_15752 (I270525,I270508,I270460);
DFFARX1 I_15753  ( .D(I270508), .CLK(I2702), .RSTB(I270194), .Q(I270162) );
DFFARX1 I_15754  ( .D(I78821), .CLK(I2702), .RSTB(I270194), .Q(I270556) );
nor I_15755 (I270573,I270556,I270279);
nand I_15756 (I270180,I270443,I270573);
nor I_15757 (I270604,I270556,I270344);
not I_15758 (I270177,I270556);
nand I_15759 (I270635,I270556,I270245);
and I_15760 (I270652,I270313,I270635);
DFFARX1 I_15761  ( .D(I270652), .CLK(I2702), .RSTB(I270194), .Q(I270156) );
DFFARX1 I_15762  ( .D(I270556), .CLK(I2702), .RSTB(I270194), .Q(I270159) );
DFFARX1 I_15763  ( .D(I78836), .CLK(I2702), .RSTB(I270194), .Q(I270697) );
not I_15764 (I270714,I270697);
nand I_15765 (I270731,I270714,I270279);
and I_15766 (I270748,I270508,I270731);
DFFARX1 I_15767  ( .D(I270748), .CLK(I2702), .RSTB(I270194), .Q(I270186) );
or I_15768 (I270779,I270714,I270525);
DFFARX1 I_15769  ( .D(I270779), .CLK(I2702), .RSTB(I270194), .Q(I270171) );
nand I_15770 (I270174,I270714,I270604);
not I_15771 (I270857,I2709);
not I_15772 (I270874,I43683);
nor I_15773 (I270891,I43689,I43692);
nand I_15774 (I270908,I270891,I43668);
nor I_15775 (I270925,I270874,I43689);
nand I_15776 (I270942,I270925,I43677);
not I_15777 (I270959,I270942);
not I_15778 (I270976,I43689);
nor I_15779 (I270846,I270942,I270976);
not I_15780 (I271007,I270976);
nand I_15781 (I270831,I270942,I271007);
not I_15782 (I271038,I43671);
nor I_15783 (I271055,I271038,I43695);
and I_15784 (I271072,I271055,I43665);
or I_15785 (I271089,I271072,I43674);
DFFARX1 I_15786  ( .D(I271089), .CLK(I2702), .RSTB(I270857), .Q(I271106) );
nor I_15787 (I271123,I271106,I270959);
DFFARX1 I_15788  ( .D(I271106), .CLK(I2702), .RSTB(I270857), .Q(I271140) );
not I_15789 (I270828,I271140);
nand I_15790 (I271171,I270874,I43671);
and I_15791 (I271188,I271171,I271123);
DFFARX1 I_15792  ( .D(I271171), .CLK(I2702), .RSTB(I270857), .Q(I270825) );
DFFARX1 I_15793  ( .D(I43680), .CLK(I2702), .RSTB(I270857), .Q(I271219) );
nor I_15794 (I271236,I271219,I270942);
nand I_15795 (I270843,I271106,I271236);
nor I_15796 (I271267,I271219,I271007);
not I_15797 (I270840,I271219);
nand I_15798 (I271298,I271219,I270908);
and I_15799 (I271315,I270976,I271298);
DFFARX1 I_15800  ( .D(I271315), .CLK(I2702), .RSTB(I270857), .Q(I270819) );
DFFARX1 I_15801  ( .D(I271219), .CLK(I2702), .RSTB(I270857), .Q(I270822) );
DFFARX1 I_15802  ( .D(I43686), .CLK(I2702), .RSTB(I270857), .Q(I271360) );
not I_15803 (I271377,I271360);
nand I_15804 (I271394,I271377,I270942);
and I_15805 (I271411,I271171,I271394);
DFFARX1 I_15806  ( .D(I271411), .CLK(I2702), .RSTB(I270857), .Q(I270849) );
or I_15807 (I271442,I271377,I271188);
DFFARX1 I_15808  ( .D(I271442), .CLK(I2702), .RSTB(I270857), .Q(I270834) );
nand I_15809 (I270837,I271377,I271267);
not I_15810 (I271520,I2709);
not I_15811 (I271537,I3852);
nor I_15812 (I271554,I3858,I3861);
nand I_15813 (I271571,I271554,I3837);
nor I_15814 (I271588,I271537,I3858);
nand I_15815 (I271605,I271588,I3846);
not I_15816 (I271622,I271605);
not I_15817 (I271639,I3858);
nor I_15818 (I271509,I271605,I271639);
not I_15819 (I271670,I271639);
nand I_15820 (I271494,I271605,I271670);
not I_15821 (I271701,I3840);
nor I_15822 (I271718,I271701,I3864);
and I_15823 (I271735,I271718,I3834);
or I_15824 (I271752,I271735,I3843);
DFFARX1 I_15825  ( .D(I271752), .CLK(I2702), .RSTB(I271520), .Q(I271769) );
nor I_15826 (I271786,I271769,I271622);
DFFARX1 I_15827  ( .D(I271769), .CLK(I2702), .RSTB(I271520), .Q(I271803) );
not I_15828 (I271491,I271803);
nand I_15829 (I271834,I271537,I3840);
and I_15830 (I271851,I271834,I271786);
DFFARX1 I_15831  ( .D(I271834), .CLK(I2702), .RSTB(I271520), .Q(I271488) );
DFFARX1 I_15832  ( .D(I3849), .CLK(I2702), .RSTB(I271520), .Q(I271882) );
nor I_15833 (I271899,I271882,I271605);
nand I_15834 (I271506,I271769,I271899);
nor I_15835 (I271930,I271882,I271670);
not I_15836 (I271503,I271882);
nand I_15837 (I271961,I271882,I271571);
and I_15838 (I271978,I271639,I271961);
DFFARX1 I_15839  ( .D(I271978), .CLK(I2702), .RSTB(I271520), .Q(I271482) );
DFFARX1 I_15840  ( .D(I271882), .CLK(I2702), .RSTB(I271520), .Q(I271485) );
DFFARX1 I_15841  ( .D(I3855), .CLK(I2702), .RSTB(I271520), .Q(I272023) );
not I_15842 (I272040,I272023);
nand I_15843 (I272057,I272040,I271605);
and I_15844 (I272074,I271834,I272057);
DFFARX1 I_15845  ( .D(I272074), .CLK(I2702), .RSTB(I271520), .Q(I271512) );
or I_15846 (I272105,I272040,I271851);
DFFARX1 I_15847  ( .D(I272105), .CLK(I2702), .RSTB(I271520), .Q(I271497) );
nand I_15848 (I271500,I272040,I271930);
not I_15849 (I272183,I2709);
not I_15850 (I272200,I86579);
nor I_15851 (I272217,I86576,I86600);
nand I_15852 (I272234,I272217,I86597);
nor I_15853 (I272251,I272200,I86576);
nand I_15854 (I272268,I272251,I86603);
not I_15855 (I272285,I272268);
not I_15856 (I272302,I86576);
nor I_15857 (I272172,I272268,I272302);
not I_15858 (I272333,I272302);
nand I_15859 (I272157,I272268,I272333);
not I_15860 (I272364,I86594);
nor I_15861 (I272381,I272364,I86585);
and I_15862 (I272398,I272381,I86582);
or I_15863 (I272415,I272398,I86591);
DFFARX1 I_15864  ( .D(I272415), .CLK(I2702), .RSTB(I272183), .Q(I272432) );
nor I_15865 (I272449,I272432,I272285);
DFFARX1 I_15866  ( .D(I272432), .CLK(I2702), .RSTB(I272183), .Q(I272466) );
not I_15867 (I272154,I272466);
nand I_15868 (I272497,I272200,I86594);
and I_15869 (I272514,I272497,I272449);
DFFARX1 I_15870  ( .D(I272497), .CLK(I2702), .RSTB(I272183), .Q(I272151) );
DFFARX1 I_15871  ( .D(I86573), .CLK(I2702), .RSTB(I272183), .Q(I272545) );
nor I_15872 (I272562,I272545,I272268);
nand I_15873 (I272169,I272432,I272562);
nor I_15874 (I272593,I272545,I272333);
not I_15875 (I272166,I272545);
nand I_15876 (I272624,I272545,I272234);
and I_15877 (I272641,I272302,I272624);
DFFARX1 I_15878  ( .D(I272641), .CLK(I2702), .RSTB(I272183), .Q(I272145) );
DFFARX1 I_15879  ( .D(I272545), .CLK(I2702), .RSTB(I272183), .Q(I272148) );
DFFARX1 I_15880  ( .D(I86588), .CLK(I2702), .RSTB(I272183), .Q(I272686) );
not I_15881 (I272703,I272686);
nand I_15882 (I272720,I272703,I272268);
and I_15883 (I272737,I272497,I272720);
DFFARX1 I_15884  ( .D(I272737), .CLK(I2702), .RSTB(I272183), .Q(I272175) );
or I_15885 (I272768,I272703,I272514);
DFFARX1 I_15886  ( .D(I272768), .CLK(I2702), .RSTB(I272183), .Q(I272160) );
nand I_15887 (I272163,I272703,I272593);
not I_15888 (I272846,I2709);
not I_15889 (I272863,I527452);
nor I_15890 (I272880,I527461,I527443);
nand I_15891 (I272897,I272880,I527464);
nor I_15892 (I272914,I272863,I527461);
nand I_15893 (I272931,I272914,I527455);
not I_15894 (I272948,I272931);
not I_15895 (I272965,I527461);
nor I_15896 (I272835,I272931,I272965);
not I_15897 (I272996,I272965);
nand I_15898 (I272820,I272931,I272996);
not I_15899 (I273027,I527449);
nor I_15900 (I273044,I273027,I527440);
and I_15901 (I273061,I273044,I527437);
or I_15902 (I273078,I273061,I527434);
DFFARX1 I_15903  ( .D(I273078), .CLK(I2702), .RSTB(I272846), .Q(I273095) );
nor I_15904 (I273112,I273095,I272948);
DFFARX1 I_15905  ( .D(I273095), .CLK(I2702), .RSTB(I272846), .Q(I273129) );
not I_15906 (I272817,I273129);
nand I_15907 (I273160,I272863,I527449);
and I_15908 (I273177,I273160,I273112);
DFFARX1 I_15909  ( .D(I273160), .CLK(I2702), .RSTB(I272846), .Q(I272814) );
DFFARX1 I_15910  ( .D(I527458), .CLK(I2702), .RSTB(I272846), .Q(I273208) );
nor I_15911 (I273225,I273208,I272931);
nand I_15912 (I272832,I273095,I273225);
nor I_15913 (I273256,I273208,I272996);
not I_15914 (I272829,I273208);
nand I_15915 (I273287,I273208,I272897);
and I_15916 (I273304,I272965,I273287);
DFFARX1 I_15917  ( .D(I273304), .CLK(I2702), .RSTB(I272846), .Q(I272808) );
DFFARX1 I_15918  ( .D(I273208), .CLK(I2702), .RSTB(I272846), .Q(I272811) );
DFFARX1 I_15919  ( .D(I527446), .CLK(I2702), .RSTB(I272846), .Q(I273349) );
not I_15920 (I273366,I273349);
nand I_15921 (I273383,I273366,I272931);
and I_15922 (I273400,I273160,I273383);
DFFARX1 I_15923  ( .D(I273400), .CLK(I2702), .RSTB(I272846), .Q(I272838) );
or I_15924 (I273431,I273366,I273177);
DFFARX1 I_15925  ( .D(I273431), .CLK(I2702), .RSTB(I272846), .Q(I272823) );
nand I_15926 (I272826,I273366,I273256);
not I_15927 (I273509,I2709);
not I_15928 (I273526,I25731);
nor I_15929 (I273543,I25737,I25740);
nand I_15930 (I273560,I273543,I25716);
nor I_15931 (I273577,I273526,I25737);
nand I_15932 (I273594,I273577,I25725);
not I_15933 (I273611,I273594);
not I_15934 (I273628,I25737);
nor I_15935 (I273498,I273594,I273628);
not I_15936 (I273659,I273628);
nand I_15937 (I273483,I273594,I273659);
not I_15938 (I273690,I25719);
nor I_15939 (I273707,I273690,I25743);
and I_15940 (I273724,I273707,I25713);
or I_15941 (I273741,I273724,I25722);
DFFARX1 I_15942  ( .D(I273741), .CLK(I2702), .RSTB(I273509), .Q(I273758) );
nor I_15943 (I273775,I273758,I273611);
DFFARX1 I_15944  ( .D(I273758), .CLK(I2702), .RSTB(I273509), .Q(I273792) );
not I_15945 (I273480,I273792);
nand I_15946 (I273823,I273526,I25719);
and I_15947 (I273840,I273823,I273775);
DFFARX1 I_15948  ( .D(I273823), .CLK(I2702), .RSTB(I273509), .Q(I273477) );
DFFARX1 I_15949  ( .D(I25728), .CLK(I2702), .RSTB(I273509), .Q(I273871) );
nor I_15950 (I273888,I273871,I273594);
nand I_15951 (I273495,I273758,I273888);
nor I_15952 (I273919,I273871,I273659);
not I_15953 (I273492,I273871);
nand I_15954 (I273950,I273871,I273560);
and I_15955 (I273967,I273628,I273950);
DFFARX1 I_15956  ( .D(I273967), .CLK(I2702), .RSTB(I273509), .Q(I273471) );
DFFARX1 I_15957  ( .D(I273871), .CLK(I2702), .RSTB(I273509), .Q(I273474) );
DFFARX1 I_15958  ( .D(I25734), .CLK(I2702), .RSTB(I273509), .Q(I274012) );
not I_15959 (I274029,I274012);
nand I_15960 (I274046,I274029,I273594);
and I_15961 (I274063,I273823,I274046);
DFFARX1 I_15962  ( .D(I274063), .CLK(I2702), .RSTB(I273509), .Q(I273501) );
or I_15963 (I274094,I274029,I273840);
DFFARX1 I_15964  ( .D(I274094), .CLK(I2702), .RSTB(I273509), .Q(I273486) );
nand I_15965 (I273489,I274029,I273919);
not I_15966 (I274172,I2709);
not I_15967 (I274189,I454672);
nor I_15968 (I274206,I454684,I454666);
nand I_15969 (I274223,I274206,I454687);
nor I_15970 (I274240,I274189,I454684);
nand I_15971 (I274257,I274240,I454678);
not I_15972 (I274274,I274257);
not I_15973 (I274291,I454684);
nor I_15974 (I274161,I274257,I274291);
not I_15975 (I274322,I274291);
nand I_15976 (I274146,I274257,I274322);
not I_15977 (I274353,I454669);
nor I_15978 (I274370,I274353,I454663);
and I_15979 (I274387,I274370,I454675);
or I_15980 (I274404,I274387,I454660);
DFFARX1 I_15981  ( .D(I274404), .CLK(I2702), .RSTB(I274172), .Q(I274421) );
nor I_15982 (I274438,I274421,I274274);
DFFARX1 I_15983  ( .D(I274421), .CLK(I2702), .RSTB(I274172), .Q(I274455) );
not I_15984 (I274143,I274455);
nand I_15985 (I274486,I274189,I454669);
and I_15986 (I274503,I274486,I274438);
DFFARX1 I_15987  ( .D(I274486), .CLK(I2702), .RSTB(I274172), .Q(I274140) );
DFFARX1 I_15988  ( .D(I454657), .CLK(I2702), .RSTB(I274172), .Q(I274534) );
nor I_15989 (I274551,I274534,I274257);
nand I_15990 (I274158,I274421,I274551);
nor I_15991 (I274582,I274534,I274322);
not I_15992 (I274155,I274534);
nand I_15993 (I274613,I274534,I274223);
and I_15994 (I274630,I274291,I274613);
DFFARX1 I_15995  ( .D(I274630), .CLK(I2702), .RSTB(I274172), .Q(I274134) );
DFFARX1 I_15996  ( .D(I274534), .CLK(I2702), .RSTB(I274172), .Q(I274137) );
DFFARX1 I_15997  ( .D(I454681), .CLK(I2702), .RSTB(I274172), .Q(I274675) );
not I_15998 (I274692,I274675);
nand I_15999 (I274709,I274692,I274257);
and I_16000 (I274726,I274486,I274709);
DFFARX1 I_16001  ( .D(I274726), .CLK(I2702), .RSTB(I274172), .Q(I274164) );
or I_16002 (I274757,I274692,I274503);
DFFARX1 I_16003  ( .D(I274757), .CLK(I2702), .RSTB(I274172), .Q(I274149) );
nand I_16004 (I274152,I274692,I274582);
not I_16005 (I274835,I2709);
not I_16006 (I274852,I467966);
nor I_16007 (I274869,I467978,I467960);
nand I_16008 (I274886,I274869,I467981);
nor I_16009 (I274903,I274852,I467978);
nand I_16010 (I274920,I274903,I467972);
not I_16011 (I274937,I274920);
not I_16012 (I274954,I467978);
nor I_16013 (I274824,I274920,I274954);
not I_16014 (I274985,I274954);
nand I_16015 (I274809,I274920,I274985);
not I_16016 (I275016,I467963);
nor I_16017 (I275033,I275016,I467957);
and I_16018 (I275050,I275033,I467969);
or I_16019 (I275067,I275050,I467954);
DFFARX1 I_16020  ( .D(I275067), .CLK(I2702), .RSTB(I274835), .Q(I275084) );
nor I_16021 (I275101,I275084,I274937);
DFFARX1 I_16022  ( .D(I275084), .CLK(I2702), .RSTB(I274835), .Q(I275118) );
not I_16023 (I274806,I275118);
nand I_16024 (I275149,I274852,I467963);
and I_16025 (I275166,I275149,I275101);
DFFARX1 I_16026  ( .D(I275149), .CLK(I2702), .RSTB(I274835), .Q(I274803) );
DFFARX1 I_16027  ( .D(I467951), .CLK(I2702), .RSTB(I274835), .Q(I275197) );
nor I_16028 (I275214,I275197,I274920);
nand I_16029 (I274821,I275084,I275214);
nor I_16030 (I275245,I275197,I274985);
not I_16031 (I274818,I275197);
nand I_16032 (I275276,I275197,I274886);
and I_16033 (I275293,I274954,I275276);
DFFARX1 I_16034  ( .D(I275293), .CLK(I2702), .RSTB(I274835), .Q(I274797) );
DFFARX1 I_16035  ( .D(I275197), .CLK(I2702), .RSTB(I274835), .Q(I274800) );
DFFARX1 I_16036  ( .D(I467975), .CLK(I2702), .RSTB(I274835), .Q(I275338) );
not I_16037 (I275355,I275338);
nand I_16038 (I275372,I275355,I274920);
and I_16039 (I275389,I275149,I275372);
DFFARX1 I_16040  ( .D(I275389), .CLK(I2702), .RSTB(I274835), .Q(I274827) );
or I_16041 (I275420,I275355,I275166);
DFFARX1 I_16042  ( .D(I275420), .CLK(I2702), .RSTB(I274835), .Q(I274812) );
nand I_16043 (I274815,I275355,I275245);
not I_16044 (I275498,I2709);
not I_16045 (I275515,I127277);
nor I_16046 (I275532,I127274,I127298);
nand I_16047 (I275549,I275532,I127295);
nor I_16048 (I275566,I275515,I127274);
nand I_16049 (I275583,I275566,I127301);
not I_16050 (I275600,I275583);
not I_16051 (I275617,I127274);
nor I_16052 (I275487,I275583,I275617);
not I_16053 (I275648,I275617);
nand I_16054 (I275472,I275583,I275648);
not I_16055 (I275679,I127292);
nor I_16056 (I275696,I275679,I127283);
and I_16057 (I275713,I275696,I127280);
or I_16058 (I275730,I275713,I127289);
DFFARX1 I_16059  ( .D(I275730), .CLK(I2702), .RSTB(I275498), .Q(I275747) );
nor I_16060 (I275764,I275747,I275600);
DFFARX1 I_16061  ( .D(I275747), .CLK(I2702), .RSTB(I275498), .Q(I275781) );
not I_16062 (I275469,I275781);
nand I_16063 (I275812,I275515,I127292);
and I_16064 (I275829,I275812,I275764);
DFFARX1 I_16065  ( .D(I275812), .CLK(I2702), .RSTB(I275498), .Q(I275466) );
DFFARX1 I_16066  ( .D(I127271), .CLK(I2702), .RSTB(I275498), .Q(I275860) );
nor I_16067 (I275877,I275860,I275583);
nand I_16068 (I275484,I275747,I275877);
nor I_16069 (I275908,I275860,I275648);
not I_16070 (I275481,I275860);
nand I_16071 (I275939,I275860,I275549);
and I_16072 (I275956,I275617,I275939);
DFFARX1 I_16073  ( .D(I275956), .CLK(I2702), .RSTB(I275498), .Q(I275460) );
DFFARX1 I_16074  ( .D(I275860), .CLK(I2702), .RSTB(I275498), .Q(I275463) );
DFFARX1 I_16075  ( .D(I127286), .CLK(I2702), .RSTB(I275498), .Q(I276001) );
not I_16076 (I276018,I276001);
nand I_16077 (I276035,I276018,I275583);
and I_16078 (I276052,I275812,I276035);
DFFARX1 I_16079  ( .D(I276052), .CLK(I2702), .RSTB(I275498), .Q(I275490) );
or I_16080 (I276083,I276018,I275829);
DFFARX1 I_16081  ( .D(I276083), .CLK(I2702), .RSTB(I275498), .Q(I275475) );
nand I_16082 (I275478,I276018,I275908);
not I_16083 (I276161,I2709);
not I_16084 (I276178,I484728);
nor I_16085 (I276195,I484740,I484722);
nand I_16086 (I276212,I276195,I484743);
nor I_16087 (I276229,I276178,I484740);
nand I_16088 (I276246,I276229,I484734);
not I_16089 (I276263,I276246);
not I_16090 (I276280,I484740);
nor I_16091 (I276150,I276246,I276280);
not I_16092 (I276311,I276280);
nand I_16093 (I276135,I276246,I276311);
not I_16094 (I276342,I484725);
nor I_16095 (I276359,I276342,I484719);
and I_16096 (I276376,I276359,I484731);
or I_16097 (I276393,I276376,I484716);
DFFARX1 I_16098  ( .D(I276393), .CLK(I2702), .RSTB(I276161), .Q(I276410) );
nor I_16099 (I276427,I276410,I276263);
DFFARX1 I_16100  ( .D(I276410), .CLK(I2702), .RSTB(I276161), .Q(I276444) );
not I_16101 (I276132,I276444);
nand I_16102 (I276475,I276178,I484725);
and I_16103 (I276492,I276475,I276427);
DFFARX1 I_16104  ( .D(I276475), .CLK(I2702), .RSTB(I276161), .Q(I276129) );
DFFARX1 I_16105  ( .D(I484713), .CLK(I2702), .RSTB(I276161), .Q(I276523) );
nor I_16106 (I276540,I276523,I276246);
nand I_16107 (I276147,I276410,I276540);
nor I_16108 (I276571,I276523,I276311);
not I_16109 (I276144,I276523);
nand I_16110 (I276602,I276523,I276212);
and I_16111 (I276619,I276280,I276602);
DFFARX1 I_16112  ( .D(I276619), .CLK(I2702), .RSTB(I276161), .Q(I276123) );
DFFARX1 I_16113  ( .D(I276523), .CLK(I2702), .RSTB(I276161), .Q(I276126) );
DFFARX1 I_16114  ( .D(I484737), .CLK(I2702), .RSTB(I276161), .Q(I276664) );
not I_16115 (I276681,I276664);
nand I_16116 (I276698,I276681,I276246);
and I_16117 (I276715,I276475,I276698);
DFFARX1 I_16118  ( .D(I276715), .CLK(I2702), .RSTB(I276161), .Q(I276153) );
or I_16119 (I276746,I276681,I276492);
DFFARX1 I_16120  ( .D(I276746), .CLK(I2702), .RSTB(I276161), .Q(I276138) );
nand I_16121 (I276141,I276681,I276571);
not I_16122 (I276824,I2709);
not I_16123 (I276841,I193251);
nor I_16124 (I276858,I193257,I193263);
nand I_16125 (I276875,I276858,I193266);
nor I_16126 (I276892,I276841,I193257);
nand I_16127 (I276909,I276892,I193248);
not I_16128 (I276926,I276909);
not I_16129 (I276943,I193257);
nor I_16130 (I276813,I276909,I276943);
not I_16131 (I276974,I276943);
nand I_16132 (I276798,I276909,I276974);
not I_16133 (I277005,I193260);
nor I_16134 (I277022,I277005,I193254);
and I_16135 (I277039,I277022,I193269);
or I_16136 (I277056,I277039,I193275);
DFFARX1 I_16137  ( .D(I277056), .CLK(I2702), .RSTB(I276824), .Q(I277073) );
nor I_16138 (I277090,I277073,I276926);
DFFARX1 I_16139  ( .D(I277073), .CLK(I2702), .RSTB(I276824), .Q(I277107) );
not I_16140 (I276795,I277107);
nand I_16141 (I277138,I276841,I193260);
and I_16142 (I277155,I277138,I277090);
DFFARX1 I_16143  ( .D(I277138), .CLK(I2702), .RSTB(I276824), .Q(I276792) );
DFFARX1 I_16144  ( .D(I193272), .CLK(I2702), .RSTB(I276824), .Q(I277186) );
nor I_16145 (I277203,I277186,I276909);
nand I_16146 (I276810,I277073,I277203);
nor I_16147 (I277234,I277186,I276974);
not I_16148 (I276807,I277186);
nand I_16149 (I277265,I277186,I276875);
and I_16150 (I277282,I276943,I277265);
DFFARX1 I_16151  ( .D(I277282), .CLK(I2702), .RSTB(I276824), .Q(I276786) );
DFFARX1 I_16152  ( .D(I277186), .CLK(I2702), .RSTB(I276824), .Q(I276789) );
DFFARX1 I_16153  ( .D(I193278), .CLK(I2702), .RSTB(I276824), .Q(I277327) );
not I_16154 (I277344,I277327);
nand I_16155 (I277361,I277344,I276909);
and I_16156 (I277378,I277138,I277361);
DFFARX1 I_16157  ( .D(I277378), .CLK(I2702), .RSTB(I276824), .Q(I276816) );
or I_16158 (I277409,I277344,I277155);
DFFARX1 I_16159  ( .D(I277409), .CLK(I2702), .RSTB(I276824), .Q(I276801) );
nand I_16160 (I276804,I277344,I277234);
not I_16161 (I277487,I2709);
not I_16162 (I277504,I682242);
nor I_16163 (I277521,I682260,I682251);
nand I_16164 (I277538,I277521,I682257);
nor I_16165 (I277555,I277504,I682260);
nand I_16166 (I277572,I277555,I682263);
not I_16167 (I277589,I277572);
not I_16168 (I277606,I682260);
nor I_16169 (I277476,I277572,I277606);
not I_16170 (I277637,I277606);
nand I_16171 (I277461,I277572,I277637);
not I_16172 (I277668,I682239);
nor I_16173 (I277685,I277668,I682254);
and I_16174 (I277702,I277685,I682236);
or I_16175 (I277719,I277702,I682245);
DFFARX1 I_16176  ( .D(I277719), .CLK(I2702), .RSTB(I277487), .Q(I277736) );
nor I_16177 (I277753,I277736,I277589);
DFFARX1 I_16178  ( .D(I277736), .CLK(I2702), .RSTB(I277487), .Q(I277770) );
not I_16179 (I277458,I277770);
nand I_16180 (I277801,I277504,I682239);
and I_16181 (I277818,I277801,I277753);
DFFARX1 I_16182  ( .D(I277801), .CLK(I2702), .RSTB(I277487), .Q(I277455) );
DFFARX1 I_16183  ( .D(I682248), .CLK(I2702), .RSTB(I277487), .Q(I277849) );
nor I_16184 (I277866,I277849,I277572);
nand I_16185 (I277473,I277736,I277866);
nor I_16186 (I277897,I277849,I277637);
not I_16187 (I277470,I277849);
nand I_16188 (I277928,I277849,I277538);
and I_16189 (I277945,I277606,I277928);
DFFARX1 I_16190  ( .D(I277945), .CLK(I2702), .RSTB(I277487), .Q(I277449) );
DFFARX1 I_16191  ( .D(I277849), .CLK(I2702), .RSTB(I277487), .Q(I277452) );
DFFARX1 I_16192  ( .D(I682266), .CLK(I2702), .RSTB(I277487), .Q(I277990) );
not I_16193 (I278007,I277990);
nand I_16194 (I278024,I278007,I277572);
and I_16195 (I278041,I277801,I278024);
DFFARX1 I_16196  ( .D(I278041), .CLK(I2702), .RSTB(I277487), .Q(I277479) );
or I_16197 (I278072,I278007,I277818);
DFFARX1 I_16198  ( .D(I278072), .CLK(I2702), .RSTB(I277487), .Q(I277464) );
nand I_16199 (I277467,I278007,I277897);
not I_16200 (I278150,I2709);
not I_16201 (I278167,I335091);
nor I_16202 (I278184,I335088,I335106);
nand I_16203 (I278201,I278184,I335109);
nor I_16204 (I278218,I278167,I335088);
nand I_16205 (I278235,I278218,I335094);
not I_16206 (I278252,I278235);
not I_16207 (I278269,I335088);
nor I_16208 (I278139,I278235,I278269);
not I_16209 (I278300,I278269);
nand I_16210 (I278124,I278235,I278300);
not I_16211 (I278331,I335103);
nor I_16212 (I278348,I278331,I335085);
and I_16213 (I278365,I278348,I335079);
or I_16214 (I278382,I278365,I335097);
DFFARX1 I_16215  ( .D(I278382), .CLK(I2702), .RSTB(I278150), .Q(I278399) );
nor I_16216 (I278416,I278399,I278252);
DFFARX1 I_16217  ( .D(I278399), .CLK(I2702), .RSTB(I278150), .Q(I278433) );
not I_16218 (I278121,I278433);
nand I_16219 (I278464,I278167,I335103);
and I_16220 (I278481,I278464,I278416);
DFFARX1 I_16221  ( .D(I278464), .CLK(I2702), .RSTB(I278150), .Q(I278118) );
DFFARX1 I_16222  ( .D(I335082), .CLK(I2702), .RSTB(I278150), .Q(I278512) );
nor I_16223 (I278529,I278512,I278235);
nand I_16224 (I278136,I278399,I278529);
nor I_16225 (I278560,I278512,I278300);
not I_16226 (I278133,I278512);
nand I_16227 (I278591,I278512,I278201);
and I_16228 (I278608,I278269,I278591);
DFFARX1 I_16229  ( .D(I278608), .CLK(I2702), .RSTB(I278150), .Q(I278112) );
DFFARX1 I_16230  ( .D(I278512), .CLK(I2702), .RSTB(I278150), .Q(I278115) );
DFFARX1 I_16231  ( .D(I335100), .CLK(I2702), .RSTB(I278150), .Q(I278653) );
not I_16232 (I278670,I278653);
nand I_16233 (I278687,I278670,I278235);
and I_16234 (I278704,I278464,I278687);
DFFARX1 I_16235  ( .D(I278704), .CLK(I2702), .RSTB(I278150), .Q(I278142) );
or I_16236 (I278735,I278670,I278481);
DFFARX1 I_16237  ( .D(I278735), .CLK(I2702), .RSTB(I278150), .Q(I278127) );
nand I_16238 (I278130,I278670,I278560);
not I_16239 (I278813,I2709);
not I_16240 (I278830,I439644);
nor I_16241 (I278847,I439656,I439638);
nand I_16242 (I278864,I278847,I439659);
nor I_16243 (I278881,I278830,I439656);
nand I_16244 (I278898,I278881,I439650);
not I_16245 (I278915,I278898);
not I_16246 (I278932,I439656);
nor I_16247 (I278802,I278898,I278932);
not I_16248 (I278963,I278932);
nand I_16249 (I278787,I278898,I278963);
not I_16250 (I278994,I439641);
nor I_16251 (I279011,I278994,I439635);
and I_16252 (I279028,I279011,I439647);
or I_16253 (I279045,I279028,I439632);
DFFARX1 I_16254  ( .D(I279045), .CLK(I2702), .RSTB(I278813), .Q(I279062) );
nor I_16255 (I279079,I279062,I278915);
DFFARX1 I_16256  ( .D(I279062), .CLK(I2702), .RSTB(I278813), .Q(I279096) );
not I_16257 (I278784,I279096);
nand I_16258 (I279127,I278830,I439641);
and I_16259 (I279144,I279127,I279079);
DFFARX1 I_16260  ( .D(I279127), .CLK(I2702), .RSTB(I278813), .Q(I278781) );
DFFARX1 I_16261  ( .D(I439629), .CLK(I2702), .RSTB(I278813), .Q(I279175) );
nor I_16262 (I279192,I279175,I278898);
nand I_16263 (I278799,I279062,I279192);
nor I_16264 (I279223,I279175,I278963);
not I_16265 (I278796,I279175);
nand I_16266 (I279254,I279175,I278864);
and I_16267 (I279271,I278932,I279254);
DFFARX1 I_16268  ( .D(I279271), .CLK(I2702), .RSTB(I278813), .Q(I278775) );
DFFARX1 I_16269  ( .D(I279175), .CLK(I2702), .RSTB(I278813), .Q(I278778) );
DFFARX1 I_16270  ( .D(I439653), .CLK(I2702), .RSTB(I278813), .Q(I279316) );
not I_16271 (I279333,I279316);
nand I_16272 (I279350,I279333,I278898);
and I_16273 (I279367,I279127,I279350);
DFFARX1 I_16274  ( .D(I279367), .CLK(I2702), .RSTB(I278813), .Q(I278805) );
or I_16275 (I279398,I279333,I279144);
DFFARX1 I_16276  ( .D(I279398), .CLK(I2702), .RSTB(I278813), .Q(I278790) );
nand I_16277 (I278793,I279333,I279223);
not I_16278 (I279476,I2709);
not I_16279 (I279493,I508412);
nor I_16280 (I279510,I508421,I508403);
nand I_16281 (I279527,I279510,I508424);
nor I_16282 (I279544,I279493,I508421);
nand I_16283 (I279561,I279544,I508415);
not I_16284 (I279578,I279561);
not I_16285 (I279595,I508421);
nor I_16286 (I279465,I279561,I279595);
not I_16287 (I279626,I279595);
nand I_16288 (I279450,I279561,I279626);
not I_16289 (I279657,I508409);
nor I_16290 (I279674,I279657,I508400);
and I_16291 (I279691,I279674,I508397);
or I_16292 (I279708,I279691,I508394);
DFFARX1 I_16293  ( .D(I279708), .CLK(I2702), .RSTB(I279476), .Q(I279725) );
nor I_16294 (I279742,I279725,I279578);
DFFARX1 I_16295  ( .D(I279725), .CLK(I2702), .RSTB(I279476), .Q(I279759) );
not I_16296 (I279447,I279759);
nand I_16297 (I279790,I279493,I508409);
and I_16298 (I279807,I279790,I279742);
DFFARX1 I_16299  ( .D(I279790), .CLK(I2702), .RSTB(I279476), .Q(I279444) );
DFFARX1 I_16300  ( .D(I508418), .CLK(I2702), .RSTB(I279476), .Q(I279838) );
nor I_16301 (I279855,I279838,I279561);
nand I_16302 (I279462,I279725,I279855);
nor I_16303 (I279886,I279838,I279626);
not I_16304 (I279459,I279838);
nand I_16305 (I279917,I279838,I279527);
and I_16306 (I279934,I279595,I279917);
DFFARX1 I_16307  ( .D(I279934), .CLK(I2702), .RSTB(I279476), .Q(I279438) );
DFFARX1 I_16308  ( .D(I279838), .CLK(I2702), .RSTB(I279476), .Q(I279441) );
DFFARX1 I_16309  ( .D(I508406), .CLK(I2702), .RSTB(I279476), .Q(I279979) );
not I_16310 (I279996,I279979);
nand I_16311 (I280013,I279996,I279561);
and I_16312 (I280030,I279790,I280013);
DFFARX1 I_16313  ( .D(I280030), .CLK(I2702), .RSTB(I279476), .Q(I279468) );
or I_16314 (I280061,I279996,I279807);
DFFARX1 I_16315  ( .D(I280061), .CLK(I2702), .RSTB(I279476), .Q(I279453) );
nand I_16316 (I279456,I279996,I279886);
not I_16317 (I280139,I2709);
not I_16318 (I280156,I552442);
nor I_16319 (I280173,I552451,I552433);
nand I_16320 (I280190,I280173,I552454);
nor I_16321 (I280207,I280156,I552451);
nand I_16322 (I280224,I280207,I552445);
not I_16323 (I280241,I280224);
not I_16324 (I280258,I552451);
nor I_16325 (I280128,I280224,I280258);
not I_16326 (I280289,I280258);
nand I_16327 (I280113,I280224,I280289);
not I_16328 (I280320,I552439);
nor I_16329 (I280337,I280320,I552430);
and I_16330 (I280354,I280337,I552427);
or I_16331 (I280371,I280354,I552424);
DFFARX1 I_16332  ( .D(I280371), .CLK(I2702), .RSTB(I280139), .Q(I280388) );
nor I_16333 (I280405,I280388,I280241);
DFFARX1 I_16334  ( .D(I280388), .CLK(I2702), .RSTB(I280139), .Q(I280422) );
not I_16335 (I280110,I280422);
nand I_16336 (I280453,I280156,I552439);
and I_16337 (I280470,I280453,I280405);
DFFARX1 I_16338  ( .D(I280453), .CLK(I2702), .RSTB(I280139), .Q(I280107) );
DFFARX1 I_16339  ( .D(I552448), .CLK(I2702), .RSTB(I280139), .Q(I280501) );
nor I_16340 (I280518,I280501,I280224);
nand I_16341 (I280125,I280388,I280518);
nor I_16342 (I280549,I280501,I280289);
not I_16343 (I280122,I280501);
nand I_16344 (I280580,I280501,I280190);
and I_16345 (I280597,I280258,I280580);
DFFARX1 I_16346  ( .D(I280597), .CLK(I2702), .RSTB(I280139), .Q(I280101) );
DFFARX1 I_16347  ( .D(I280501), .CLK(I2702), .RSTB(I280139), .Q(I280104) );
DFFARX1 I_16348  ( .D(I552436), .CLK(I2702), .RSTB(I280139), .Q(I280642) );
not I_16349 (I280659,I280642);
nand I_16350 (I280676,I280659,I280224);
and I_16351 (I280693,I280453,I280676);
DFFARX1 I_16352  ( .D(I280693), .CLK(I2702), .RSTB(I280139), .Q(I280131) );
or I_16353 (I280724,I280659,I280470);
DFFARX1 I_16354  ( .D(I280724), .CLK(I2702), .RSTB(I280139), .Q(I280116) );
nand I_16355 (I280119,I280659,I280549);
not I_16356 (I280802,I2709);
not I_16357 (I280819,I98853);
nor I_16358 (I280836,I98850,I98874);
nand I_16359 (I280853,I280836,I98871);
nor I_16360 (I280870,I280819,I98850);
nand I_16361 (I280887,I280870,I98877);
not I_16362 (I280904,I280887);
not I_16363 (I280921,I98850);
nor I_16364 (I280791,I280887,I280921);
not I_16365 (I280952,I280921);
nand I_16366 (I280776,I280887,I280952);
not I_16367 (I280983,I98868);
nor I_16368 (I281000,I280983,I98859);
and I_16369 (I281017,I281000,I98856);
or I_16370 (I281034,I281017,I98865);
DFFARX1 I_16371  ( .D(I281034), .CLK(I2702), .RSTB(I280802), .Q(I281051) );
nor I_16372 (I281068,I281051,I280904);
DFFARX1 I_16373  ( .D(I281051), .CLK(I2702), .RSTB(I280802), .Q(I281085) );
not I_16374 (I280773,I281085);
nand I_16375 (I281116,I280819,I98868);
and I_16376 (I281133,I281116,I281068);
DFFARX1 I_16377  ( .D(I281116), .CLK(I2702), .RSTB(I280802), .Q(I280770) );
DFFARX1 I_16378  ( .D(I98847), .CLK(I2702), .RSTB(I280802), .Q(I281164) );
nor I_16379 (I281181,I281164,I280887);
nand I_16380 (I280788,I281051,I281181);
nor I_16381 (I281212,I281164,I280952);
not I_16382 (I280785,I281164);
nand I_16383 (I281243,I281164,I280853);
and I_16384 (I281260,I280921,I281243);
DFFARX1 I_16385  ( .D(I281260), .CLK(I2702), .RSTB(I280802), .Q(I280764) );
DFFARX1 I_16386  ( .D(I281164), .CLK(I2702), .RSTB(I280802), .Q(I280767) );
DFFARX1 I_16387  ( .D(I98862), .CLK(I2702), .RSTB(I280802), .Q(I281305) );
not I_16388 (I281322,I281305);
nand I_16389 (I281339,I281322,I280887);
and I_16390 (I281356,I281116,I281339);
DFFARX1 I_16391  ( .D(I281356), .CLK(I2702), .RSTB(I280802), .Q(I280794) );
or I_16392 (I281387,I281322,I281133);
DFFARX1 I_16393  ( .D(I281387), .CLK(I2702), .RSTB(I280802), .Q(I280779) );
nand I_16394 (I280782,I281322,I281212);
not I_16395 (I281465,I2709);
not I_16396 (I281482,I158775);
nor I_16397 (I281499,I158781,I158787);
nand I_16398 (I281516,I281499,I158790);
nor I_16399 (I281533,I281482,I158781);
nand I_16400 (I281550,I281533,I158772);
not I_16401 (I281567,I281550);
not I_16402 (I281584,I158781);
nor I_16403 (I281454,I281550,I281584);
not I_16404 (I281615,I281584);
nand I_16405 (I281439,I281550,I281615);
not I_16406 (I281646,I158784);
nor I_16407 (I281663,I281646,I158778);
and I_16408 (I281680,I281663,I158793);
or I_16409 (I281697,I281680,I158799);
DFFARX1 I_16410  ( .D(I281697), .CLK(I2702), .RSTB(I281465), .Q(I281714) );
nor I_16411 (I281731,I281714,I281567);
DFFARX1 I_16412  ( .D(I281714), .CLK(I2702), .RSTB(I281465), .Q(I281748) );
not I_16413 (I281436,I281748);
nand I_16414 (I281779,I281482,I158784);
and I_16415 (I281796,I281779,I281731);
DFFARX1 I_16416  ( .D(I281779), .CLK(I2702), .RSTB(I281465), .Q(I281433) );
DFFARX1 I_16417  ( .D(I158796), .CLK(I2702), .RSTB(I281465), .Q(I281827) );
nor I_16418 (I281844,I281827,I281550);
nand I_16419 (I281451,I281714,I281844);
nor I_16420 (I281875,I281827,I281615);
not I_16421 (I281448,I281827);
nand I_16422 (I281906,I281827,I281516);
and I_16423 (I281923,I281584,I281906);
DFFARX1 I_16424  ( .D(I281923), .CLK(I2702), .RSTB(I281465), .Q(I281427) );
DFFARX1 I_16425  ( .D(I281827), .CLK(I2702), .RSTB(I281465), .Q(I281430) );
DFFARX1 I_16426  ( .D(I158802), .CLK(I2702), .RSTB(I281465), .Q(I281968) );
not I_16427 (I281985,I281968);
nand I_16428 (I282002,I281985,I281550);
and I_16429 (I282019,I281779,I282002);
DFFARX1 I_16430  ( .D(I282019), .CLK(I2702), .RSTB(I281465), .Q(I281457) );
or I_16431 (I282050,I281985,I281796);
DFFARX1 I_16432  ( .D(I282050), .CLK(I2702), .RSTB(I281465), .Q(I281442) );
nand I_16433 (I281445,I281985,I281875);
not I_16434 (I282128,I2709);
not I_16435 (I282145,I34707);
nor I_16436 (I282162,I34713,I34716);
nand I_16437 (I282179,I282162,I34692);
nor I_16438 (I282196,I282145,I34713);
nand I_16439 (I282213,I282196,I34701);
not I_16440 (I282230,I282213);
not I_16441 (I282247,I34713);
nor I_16442 (I282117,I282213,I282247);
not I_16443 (I282278,I282247);
nand I_16444 (I282102,I282213,I282278);
not I_16445 (I282309,I34695);
nor I_16446 (I282326,I282309,I34719);
and I_16447 (I282343,I282326,I34689);
or I_16448 (I282360,I282343,I34698);
DFFARX1 I_16449  ( .D(I282360), .CLK(I2702), .RSTB(I282128), .Q(I282377) );
nor I_16450 (I282394,I282377,I282230);
DFFARX1 I_16451  ( .D(I282377), .CLK(I2702), .RSTB(I282128), .Q(I282411) );
not I_16452 (I282099,I282411);
nand I_16453 (I282442,I282145,I34695);
and I_16454 (I282459,I282442,I282394);
DFFARX1 I_16455  ( .D(I282442), .CLK(I2702), .RSTB(I282128), .Q(I282096) );
DFFARX1 I_16456  ( .D(I34704), .CLK(I2702), .RSTB(I282128), .Q(I282490) );
nor I_16457 (I282507,I282490,I282213);
nand I_16458 (I282114,I282377,I282507);
nor I_16459 (I282538,I282490,I282278);
not I_16460 (I282111,I282490);
nand I_16461 (I282569,I282490,I282179);
and I_16462 (I282586,I282247,I282569);
DFFARX1 I_16463  ( .D(I282586), .CLK(I2702), .RSTB(I282128), .Q(I282090) );
DFFARX1 I_16464  ( .D(I282490), .CLK(I2702), .RSTB(I282128), .Q(I282093) );
DFFARX1 I_16465  ( .D(I34710), .CLK(I2702), .RSTB(I282128), .Q(I282631) );
not I_16466 (I282648,I282631);
nand I_16467 (I282665,I282648,I282213);
and I_16468 (I282682,I282442,I282665);
DFFARX1 I_16469  ( .D(I282682), .CLK(I2702), .RSTB(I282128), .Q(I282120) );
or I_16470 (I282713,I282648,I282459);
DFFARX1 I_16471  ( .D(I282713), .CLK(I2702), .RSTB(I282128), .Q(I282105) );
nand I_16472 (I282108,I282648,I282538);
not I_16473 (I282791,I2709);
not I_16474 (I282808,I485884);
nor I_16475 (I282825,I485896,I485878);
nand I_16476 (I282842,I282825,I485899);
nor I_16477 (I282859,I282808,I485896);
nand I_16478 (I282876,I282859,I485890);
not I_16479 (I282893,I282876);
not I_16480 (I282910,I485896);
nor I_16481 (I282780,I282876,I282910);
not I_16482 (I282941,I282910);
nand I_16483 (I282765,I282876,I282941);
not I_16484 (I282972,I485881);
nor I_16485 (I282989,I282972,I485875);
and I_16486 (I283006,I282989,I485887);
or I_16487 (I283023,I283006,I485872);
DFFARX1 I_16488  ( .D(I283023), .CLK(I2702), .RSTB(I282791), .Q(I283040) );
nor I_16489 (I283057,I283040,I282893);
DFFARX1 I_16490  ( .D(I283040), .CLK(I2702), .RSTB(I282791), .Q(I283074) );
not I_16491 (I282762,I283074);
nand I_16492 (I283105,I282808,I485881);
and I_16493 (I283122,I283105,I283057);
DFFARX1 I_16494  ( .D(I283105), .CLK(I2702), .RSTB(I282791), .Q(I282759) );
DFFARX1 I_16495  ( .D(I485869), .CLK(I2702), .RSTB(I282791), .Q(I283153) );
nor I_16496 (I283170,I283153,I282876);
nand I_16497 (I282777,I283040,I283170);
nor I_16498 (I283201,I283153,I282941);
not I_16499 (I282774,I283153);
nand I_16500 (I283232,I283153,I282842);
and I_16501 (I283249,I282910,I283232);
DFFARX1 I_16502  ( .D(I283249), .CLK(I2702), .RSTB(I282791), .Q(I282753) );
DFFARX1 I_16503  ( .D(I283153), .CLK(I2702), .RSTB(I282791), .Q(I282756) );
DFFARX1 I_16504  ( .D(I485893), .CLK(I2702), .RSTB(I282791), .Q(I283294) );
not I_16505 (I283311,I283294);
nand I_16506 (I283328,I283311,I282876);
and I_16507 (I283345,I283105,I283328);
DFFARX1 I_16508  ( .D(I283345), .CLK(I2702), .RSTB(I282791), .Q(I282783) );
or I_16509 (I283376,I283311,I283122);
DFFARX1 I_16510  ( .D(I283376), .CLK(I2702), .RSTB(I282791), .Q(I282768) );
nand I_16511 (I282771,I283311,I283201);
not I_16512 (I283454,I2709);
not I_16513 (I283471,I82057);
nor I_16514 (I283488,I82054,I82078);
nand I_16515 (I283505,I283488,I82075);
nor I_16516 (I283522,I283471,I82054);
nand I_16517 (I283539,I283522,I82081);
not I_16518 (I283556,I283539);
not I_16519 (I283573,I82054);
nor I_16520 (I283443,I283539,I283573);
not I_16521 (I283604,I283573);
nand I_16522 (I283428,I283539,I283604);
not I_16523 (I283635,I82072);
nor I_16524 (I283652,I283635,I82063);
and I_16525 (I283669,I283652,I82060);
or I_16526 (I283686,I283669,I82069);
DFFARX1 I_16527  ( .D(I283686), .CLK(I2702), .RSTB(I283454), .Q(I283703) );
nor I_16528 (I283720,I283703,I283556);
DFFARX1 I_16529  ( .D(I283703), .CLK(I2702), .RSTB(I283454), .Q(I283737) );
not I_16530 (I283425,I283737);
nand I_16531 (I283768,I283471,I82072);
and I_16532 (I283785,I283768,I283720);
DFFARX1 I_16533  ( .D(I283768), .CLK(I2702), .RSTB(I283454), .Q(I283422) );
DFFARX1 I_16534  ( .D(I82051), .CLK(I2702), .RSTB(I283454), .Q(I283816) );
nor I_16535 (I283833,I283816,I283539);
nand I_16536 (I283440,I283703,I283833);
nor I_16537 (I283864,I283816,I283604);
not I_16538 (I283437,I283816);
nand I_16539 (I283895,I283816,I283505);
and I_16540 (I283912,I283573,I283895);
DFFARX1 I_16541  ( .D(I283912), .CLK(I2702), .RSTB(I283454), .Q(I283416) );
DFFARX1 I_16542  ( .D(I283816), .CLK(I2702), .RSTB(I283454), .Q(I283419) );
DFFARX1 I_16543  ( .D(I82066), .CLK(I2702), .RSTB(I283454), .Q(I283957) );
not I_16544 (I283974,I283957);
nand I_16545 (I283991,I283974,I283539);
and I_16546 (I284008,I283768,I283991);
DFFARX1 I_16547  ( .D(I284008), .CLK(I2702), .RSTB(I283454), .Q(I283446) );
or I_16548 (I284039,I283974,I283785);
DFFARX1 I_16549  ( .D(I284039), .CLK(I2702), .RSTB(I283454), .Q(I283431) );
nand I_16550 (I283434,I283974,I283864);
not I_16551 (I284117,I2709);
not I_16552 (I284134,I373851);
nor I_16553 (I284151,I373848,I373866);
nand I_16554 (I284168,I284151,I373869);
nor I_16555 (I284185,I284134,I373848);
nand I_16556 (I284202,I284185,I373854);
not I_16557 (I284219,I284202);
not I_16558 (I284236,I373848);
nor I_16559 (I284106,I284202,I284236);
not I_16560 (I284267,I284236);
nand I_16561 (I284091,I284202,I284267);
not I_16562 (I284298,I373863);
nor I_16563 (I284315,I284298,I373845);
and I_16564 (I284332,I284315,I373839);
or I_16565 (I284349,I284332,I373857);
DFFARX1 I_16566  ( .D(I284349), .CLK(I2702), .RSTB(I284117), .Q(I284366) );
nor I_16567 (I284383,I284366,I284219);
DFFARX1 I_16568  ( .D(I284366), .CLK(I2702), .RSTB(I284117), .Q(I284400) );
not I_16569 (I284088,I284400);
nand I_16570 (I284431,I284134,I373863);
and I_16571 (I284448,I284431,I284383);
DFFARX1 I_16572  ( .D(I284431), .CLK(I2702), .RSTB(I284117), .Q(I284085) );
DFFARX1 I_16573  ( .D(I373842), .CLK(I2702), .RSTB(I284117), .Q(I284479) );
nor I_16574 (I284496,I284479,I284202);
nand I_16575 (I284103,I284366,I284496);
nor I_16576 (I284527,I284479,I284267);
not I_16577 (I284100,I284479);
nand I_16578 (I284558,I284479,I284168);
and I_16579 (I284575,I284236,I284558);
DFFARX1 I_16580  ( .D(I284575), .CLK(I2702), .RSTB(I284117), .Q(I284079) );
DFFARX1 I_16581  ( .D(I284479), .CLK(I2702), .RSTB(I284117), .Q(I284082) );
DFFARX1 I_16582  ( .D(I373860), .CLK(I2702), .RSTB(I284117), .Q(I284620) );
not I_16583 (I284637,I284620);
nand I_16584 (I284654,I284637,I284202);
and I_16585 (I284671,I284431,I284654);
DFFARX1 I_16586  ( .D(I284671), .CLK(I2702), .RSTB(I284117), .Q(I284109) );
or I_16587 (I284702,I284637,I284448);
DFFARX1 I_16588  ( .D(I284702), .CLK(I2702), .RSTB(I284117), .Q(I284094) );
nand I_16589 (I284097,I284637,I284527);
not I_16590 (I284780,I2709);
not I_16591 (I284797,I550062);
nor I_16592 (I284814,I550071,I550053);
nand I_16593 (I284831,I284814,I550074);
nor I_16594 (I284848,I284797,I550071);
nand I_16595 (I284865,I284848,I550065);
not I_16596 (I284882,I284865);
not I_16597 (I284899,I550071);
nor I_16598 (I284769,I284865,I284899);
not I_16599 (I284930,I284899);
nand I_16600 (I284754,I284865,I284930);
not I_16601 (I284961,I550059);
nor I_16602 (I284978,I284961,I550050);
and I_16603 (I284995,I284978,I550047);
or I_16604 (I285012,I284995,I550044);
DFFARX1 I_16605  ( .D(I285012), .CLK(I2702), .RSTB(I284780), .Q(I285029) );
nor I_16606 (I285046,I285029,I284882);
DFFARX1 I_16607  ( .D(I285029), .CLK(I2702), .RSTB(I284780), .Q(I285063) );
not I_16608 (I284751,I285063);
nand I_16609 (I285094,I284797,I550059);
and I_16610 (I285111,I285094,I285046);
DFFARX1 I_16611  ( .D(I285094), .CLK(I2702), .RSTB(I284780), .Q(I284748) );
DFFARX1 I_16612  ( .D(I550068), .CLK(I2702), .RSTB(I284780), .Q(I285142) );
nor I_16613 (I285159,I285142,I284865);
nand I_16614 (I284766,I285029,I285159);
nor I_16615 (I285190,I285142,I284930);
not I_16616 (I284763,I285142);
nand I_16617 (I285221,I285142,I284831);
and I_16618 (I285238,I284899,I285221);
DFFARX1 I_16619  ( .D(I285238), .CLK(I2702), .RSTB(I284780), .Q(I284742) );
DFFARX1 I_16620  ( .D(I285142), .CLK(I2702), .RSTB(I284780), .Q(I284745) );
DFFARX1 I_16621  ( .D(I550056), .CLK(I2702), .RSTB(I284780), .Q(I285283) );
not I_16622 (I285300,I285283);
nand I_16623 (I285317,I285300,I284865);
and I_16624 (I285334,I285094,I285317);
DFFARX1 I_16625  ( .D(I285334), .CLK(I2702), .RSTB(I284780), .Q(I284772) );
or I_16626 (I285365,I285300,I285111);
DFFARX1 I_16627  ( .D(I285365), .CLK(I2702), .RSTB(I284780), .Q(I284757) );
nand I_16628 (I284760,I285300,I285190);
not I_16629 (I285443,I2709);
not I_16630 (I285460,I584572);
nor I_16631 (I285477,I584569,I584560);
nand I_16632 (I285494,I285477,I584563);
nor I_16633 (I285511,I285460,I584569);
nand I_16634 (I285528,I285511,I584557);
not I_16635 (I285545,I285528);
not I_16636 (I285562,I584569);
nor I_16637 (I285432,I285528,I285562);
not I_16638 (I285593,I285562);
nand I_16639 (I285417,I285528,I285593);
not I_16640 (I285624,I584578);
nor I_16641 (I285641,I285624,I584581);
and I_16642 (I285658,I285641,I584566);
or I_16643 (I285675,I285658,I584554);
DFFARX1 I_16644  ( .D(I285675), .CLK(I2702), .RSTB(I285443), .Q(I285692) );
nor I_16645 (I285709,I285692,I285545);
DFFARX1 I_16646  ( .D(I285692), .CLK(I2702), .RSTB(I285443), .Q(I285726) );
not I_16647 (I285414,I285726);
nand I_16648 (I285757,I285460,I584578);
and I_16649 (I285774,I285757,I285709);
DFFARX1 I_16650  ( .D(I285757), .CLK(I2702), .RSTB(I285443), .Q(I285411) );
DFFARX1 I_16651  ( .D(I584575), .CLK(I2702), .RSTB(I285443), .Q(I285805) );
nor I_16652 (I285822,I285805,I285528);
nand I_16653 (I285429,I285692,I285822);
nor I_16654 (I285853,I285805,I285593);
not I_16655 (I285426,I285805);
nand I_16656 (I285884,I285805,I285494);
and I_16657 (I285901,I285562,I285884);
DFFARX1 I_16658  ( .D(I285901), .CLK(I2702), .RSTB(I285443), .Q(I285405) );
DFFARX1 I_16659  ( .D(I285805), .CLK(I2702), .RSTB(I285443), .Q(I285408) );
DFFARX1 I_16660  ( .D(I584584), .CLK(I2702), .RSTB(I285443), .Q(I285946) );
not I_16661 (I285963,I285946);
nand I_16662 (I285980,I285963,I285528);
and I_16663 (I285997,I285757,I285980);
DFFARX1 I_16664  ( .D(I285997), .CLK(I2702), .RSTB(I285443), .Q(I285435) );
or I_16665 (I286028,I285963,I285774);
DFFARX1 I_16666  ( .D(I286028), .CLK(I2702), .RSTB(I285443), .Q(I285420) );
nand I_16667 (I285423,I285963,I285853);
not I_16668 (I286106,I2709);
not I_16669 (I286123,I456984);
nor I_16670 (I286140,I456996,I456978);
nand I_16671 (I286157,I286140,I456999);
nor I_16672 (I286174,I286123,I456996);
nand I_16673 (I286191,I286174,I456990);
not I_16674 (I286208,I286191);
not I_16675 (I286225,I456996);
nor I_16676 (I286095,I286191,I286225);
not I_16677 (I286256,I286225);
nand I_16678 (I286080,I286191,I286256);
not I_16679 (I286287,I456981);
nor I_16680 (I286304,I286287,I456975);
and I_16681 (I286321,I286304,I456987);
or I_16682 (I286338,I286321,I456972);
DFFARX1 I_16683  ( .D(I286338), .CLK(I2702), .RSTB(I286106), .Q(I286355) );
nor I_16684 (I286372,I286355,I286208);
DFFARX1 I_16685  ( .D(I286355), .CLK(I2702), .RSTB(I286106), .Q(I286389) );
not I_16686 (I286077,I286389);
nand I_16687 (I286420,I286123,I456981);
and I_16688 (I286437,I286420,I286372);
DFFARX1 I_16689  ( .D(I286420), .CLK(I2702), .RSTB(I286106), .Q(I286074) );
DFFARX1 I_16690  ( .D(I456969), .CLK(I2702), .RSTB(I286106), .Q(I286468) );
nor I_16691 (I286485,I286468,I286191);
nand I_16692 (I286092,I286355,I286485);
nor I_16693 (I286516,I286468,I286256);
not I_16694 (I286089,I286468);
nand I_16695 (I286547,I286468,I286157);
and I_16696 (I286564,I286225,I286547);
DFFARX1 I_16697  ( .D(I286564), .CLK(I2702), .RSTB(I286106), .Q(I286068) );
DFFARX1 I_16698  ( .D(I286468), .CLK(I2702), .RSTB(I286106), .Q(I286071) );
DFFARX1 I_16699  ( .D(I456993), .CLK(I2702), .RSTB(I286106), .Q(I286609) );
not I_16700 (I286626,I286609);
nand I_16701 (I286643,I286626,I286191);
and I_16702 (I286660,I286420,I286643);
DFFARX1 I_16703  ( .D(I286660), .CLK(I2702), .RSTB(I286106), .Q(I286098) );
or I_16704 (I286691,I286626,I286437);
DFFARX1 I_16705  ( .D(I286691), .CLK(I2702), .RSTB(I286106), .Q(I286083) );
nand I_16706 (I286086,I286626,I286516);
not I_16707 (I286769,I2709);
not I_16708 (I286786,I451782);
nor I_16709 (I286803,I451794,I451776);
nand I_16710 (I286820,I286803,I451797);
nor I_16711 (I286837,I286786,I451794);
nand I_16712 (I286854,I286837,I451788);
not I_16713 (I286871,I286854);
not I_16714 (I286888,I451794);
nor I_16715 (I286758,I286854,I286888);
not I_16716 (I286919,I286888);
nand I_16717 (I286743,I286854,I286919);
not I_16718 (I286950,I451779);
nor I_16719 (I286967,I286950,I451773);
and I_16720 (I286984,I286967,I451785);
or I_16721 (I287001,I286984,I451770);
DFFARX1 I_16722  ( .D(I287001), .CLK(I2702), .RSTB(I286769), .Q(I287018) );
nor I_16723 (I287035,I287018,I286871);
DFFARX1 I_16724  ( .D(I287018), .CLK(I2702), .RSTB(I286769), .Q(I287052) );
not I_16725 (I286740,I287052);
nand I_16726 (I287083,I286786,I451779);
and I_16727 (I287100,I287083,I287035);
DFFARX1 I_16728  ( .D(I287083), .CLK(I2702), .RSTB(I286769), .Q(I286737) );
DFFARX1 I_16729  ( .D(I451767), .CLK(I2702), .RSTB(I286769), .Q(I287131) );
nor I_16730 (I287148,I287131,I286854);
nand I_16731 (I286755,I287018,I287148);
nor I_16732 (I287179,I287131,I286919);
not I_16733 (I286752,I287131);
nand I_16734 (I287210,I287131,I286820);
and I_16735 (I287227,I286888,I287210);
DFFARX1 I_16736  ( .D(I287227), .CLK(I2702), .RSTB(I286769), .Q(I286731) );
DFFARX1 I_16737  ( .D(I287131), .CLK(I2702), .RSTB(I286769), .Q(I286734) );
DFFARX1 I_16738  ( .D(I451791), .CLK(I2702), .RSTB(I286769), .Q(I287272) );
not I_16739 (I287289,I287272);
nand I_16740 (I287306,I287289,I286854);
and I_16741 (I287323,I287083,I287306);
DFFARX1 I_16742  ( .D(I287323), .CLK(I2702), .RSTB(I286769), .Q(I286761) );
or I_16743 (I287354,I287289,I287100);
DFFARX1 I_16744  ( .D(I287354), .CLK(I2702), .RSTB(I286769), .Q(I286746) );
nand I_16745 (I286749,I287289,I287179);
not I_16746 (I287432,I2709);
not I_16747 (I287449,I351241);
nor I_16748 (I287466,I351238,I351256);
nand I_16749 (I287483,I287466,I351259);
nor I_16750 (I287500,I287449,I351238);
nand I_16751 (I287517,I287500,I351244);
not I_16752 (I287534,I287517);
not I_16753 (I287551,I351238);
nor I_16754 (I287421,I287517,I287551);
not I_16755 (I287582,I287551);
nand I_16756 (I287406,I287517,I287582);
not I_16757 (I287613,I351253);
nor I_16758 (I287630,I287613,I351235);
and I_16759 (I287647,I287630,I351229);
or I_16760 (I287664,I287647,I351247);
DFFARX1 I_16761  ( .D(I287664), .CLK(I2702), .RSTB(I287432), .Q(I287681) );
nor I_16762 (I287698,I287681,I287534);
DFFARX1 I_16763  ( .D(I287681), .CLK(I2702), .RSTB(I287432), .Q(I287715) );
not I_16764 (I287403,I287715);
nand I_16765 (I287746,I287449,I351253);
and I_16766 (I287763,I287746,I287698);
DFFARX1 I_16767  ( .D(I287746), .CLK(I2702), .RSTB(I287432), .Q(I287400) );
DFFARX1 I_16768  ( .D(I351232), .CLK(I2702), .RSTB(I287432), .Q(I287794) );
nor I_16769 (I287811,I287794,I287517);
nand I_16770 (I287418,I287681,I287811);
nor I_16771 (I287842,I287794,I287582);
not I_16772 (I287415,I287794);
nand I_16773 (I287873,I287794,I287483);
and I_16774 (I287890,I287551,I287873);
DFFARX1 I_16775  ( .D(I287890), .CLK(I2702), .RSTB(I287432), .Q(I287394) );
DFFARX1 I_16776  ( .D(I287794), .CLK(I2702), .RSTB(I287432), .Q(I287397) );
DFFARX1 I_16777  ( .D(I351250), .CLK(I2702), .RSTB(I287432), .Q(I287935) );
not I_16778 (I287952,I287935);
nand I_16779 (I287969,I287952,I287517);
and I_16780 (I287986,I287746,I287969);
DFFARX1 I_16781  ( .D(I287986), .CLK(I2702), .RSTB(I287432), .Q(I287424) );
or I_16782 (I288017,I287952,I287763);
DFFARX1 I_16783  ( .D(I288017), .CLK(I2702), .RSTB(I287432), .Q(I287409) );
nand I_16784 (I287412,I287952,I287842);
not I_16785 (I288095,I2709);
not I_16786 (I288112,I338321);
nor I_16787 (I288129,I338318,I338336);
nand I_16788 (I288146,I288129,I338339);
nor I_16789 (I288163,I288112,I338318);
nand I_16790 (I288180,I288163,I338324);
not I_16791 (I288197,I288180);
not I_16792 (I288214,I338318);
nor I_16793 (I288084,I288180,I288214);
not I_16794 (I288245,I288214);
nand I_16795 (I288069,I288180,I288245);
not I_16796 (I288276,I338333);
nor I_16797 (I288293,I288276,I338315);
and I_16798 (I288310,I288293,I338309);
or I_16799 (I288327,I288310,I338327);
DFFARX1 I_16800  ( .D(I288327), .CLK(I2702), .RSTB(I288095), .Q(I288344) );
nor I_16801 (I288361,I288344,I288197);
DFFARX1 I_16802  ( .D(I288344), .CLK(I2702), .RSTB(I288095), .Q(I288378) );
not I_16803 (I288066,I288378);
nand I_16804 (I288409,I288112,I338333);
and I_16805 (I288426,I288409,I288361);
DFFARX1 I_16806  ( .D(I288409), .CLK(I2702), .RSTB(I288095), .Q(I288063) );
DFFARX1 I_16807  ( .D(I338312), .CLK(I2702), .RSTB(I288095), .Q(I288457) );
nor I_16808 (I288474,I288457,I288180);
nand I_16809 (I288081,I288344,I288474);
nor I_16810 (I288505,I288457,I288245);
not I_16811 (I288078,I288457);
nand I_16812 (I288536,I288457,I288146);
and I_16813 (I288553,I288214,I288536);
DFFARX1 I_16814  ( .D(I288553), .CLK(I2702), .RSTB(I288095), .Q(I288057) );
DFFARX1 I_16815  ( .D(I288457), .CLK(I2702), .RSTB(I288095), .Q(I288060) );
DFFARX1 I_16816  ( .D(I338330), .CLK(I2702), .RSTB(I288095), .Q(I288598) );
not I_16817 (I288615,I288598);
nand I_16818 (I288632,I288615,I288180);
and I_16819 (I288649,I288409,I288632);
DFFARX1 I_16820  ( .D(I288649), .CLK(I2702), .RSTB(I288095), .Q(I288087) );
or I_16821 (I288680,I288615,I288426);
DFFARX1 I_16822  ( .D(I288680), .CLK(I2702), .RSTB(I288095), .Q(I288072) );
nand I_16823 (I288075,I288615,I288505);
not I_16824 (I288758,I2709);
not I_16825 (I288775,I154134);
nor I_16826 (I288792,I154140,I154146);
nand I_16827 (I288809,I288792,I154149);
nor I_16828 (I288826,I288775,I154140);
nand I_16829 (I288843,I288826,I154131);
not I_16830 (I288860,I288843);
not I_16831 (I288877,I154140);
nor I_16832 (I288747,I288843,I288877);
not I_16833 (I288908,I288877);
nand I_16834 (I288732,I288843,I288908);
not I_16835 (I288939,I154143);
nor I_16836 (I288956,I288939,I154137);
and I_16837 (I288973,I288956,I154152);
or I_16838 (I288990,I288973,I154158);
DFFARX1 I_16839  ( .D(I288990), .CLK(I2702), .RSTB(I288758), .Q(I289007) );
nor I_16840 (I289024,I289007,I288860);
DFFARX1 I_16841  ( .D(I289007), .CLK(I2702), .RSTB(I288758), .Q(I289041) );
not I_16842 (I288729,I289041);
nand I_16843 (I289072,I288775,I154143);
and I_16844 (I289089,I289072,I289024);
DFFARX1 I_16845  ( .D(I289072), .CLK(I2702), .RSTB(I288758), .Q(I288726) );
DFFARX1 I_16846  ( .D(I154155), .CLK(I2702), .RSTB(I288758), .Q(I289120) );
nor I_16847 (I289137,I289120,I288843);
nand I_16848 (I288744,I289007,I289137);
nor I_16849 (I289168,I289120,I288908);
not I_16850 (I288741,I289120);
nand I_16851 (I289199,I289120,I288809);
and I_16852 (I289216,I288877,I289199);
DFFARX1 I_16853  ( .D(I289216), .CLK(I2702), .RSTB(I288758), .Q(I288720) );
DFFARX1 I_16854  ( .D(I289120), .CLK(I2702), .RSTB(I288758), .Q(I288723) );
DFFARX1 I_16855  ( .D(I154161), .CLK(I2702), .RSTB(I288758), .Q(I289261) );
not I_16856 (I289278,I289261);
nand I_16857 (I289295,I289278,I288843);
and I_16858 (I289312,I289072,I289295);
DFFARX1 I_16859  ( .D(I289312), .CLK(I2702), .RSTB(I288758), .Q(I288750) );
or I_16860 (I289343,I289278,I289089);
DFFARX1 I_16861  ( .D(I289343), .CLK(I2702), .RSTB(I288758), .Q(I288735) );
nand I_16862 (I288738,I289278,I289168);
not I_16863 (I289421,I2709);
not I_16864 (I289438,I487043);
nor I_16865 (I289455,I487040,I487037);
nand I_16866 (I289472,I289455,I487025);
nor I_16867 (I289489,I289438,I487040);
nand I_16868 (I289506,I289489,I487046);
not I_16869 (I289523,I289506);
not I_16870 (I289540,I487040);
nor I_16871 (I289410,I289506,I289540);
not I_16872 (I289571,I289540);
nand I_16873 (I289395,I289506,I289571);
not I_16874 (I289602,I487028);
nor I_16875 (I289619,I289602,I487034);
and I_16876 (I289636,I289619,I487031);
or I_16877 (I289653,I289636,I487055);
DFFARX1 I_16878  ( .D(I289653), .CLK(I2702), .RSTB(I289421), .Q(I289670) );
nor I_16879 (I289687,I289670,I289523);
DFFARX1 I_16880  ( .D(I289670), .CLK(I2702), .RSTB(I289421), .Q(I289704) );
not I_16881 (I289392,I289704);
nand I_16882 (I289735,I289438,I487028);
and I_16883 (I289752,I289735,I289687);
DFFARX1 I_16884  ( .D(I289735), .CLK(I2702), .RSTB(I289421), .Q(I289389) );
DFFARX1 I_16885  ( .D(I487052), .CLK(I2702), .RSTB(I289421), .Q(I289783) );
nor I_16886 (I289800,I289783,I289506);
nand I_16887 (I289407,I289670,I289800);
nor I_16888 (I289831,I289783,I289571);
not I_16889 (I289404,I289783);
nand I_16890 (I289862,I289783,I289472);
and I_16891 (I289879,I289540,I289862);
DFFARX1 I_16892  ( .D(I289879), .CLK(I2702), .RSTB(I289421), .Q(I289383) );
DFFARX1 I_16893  ( .D(I289783), .CLK(I2702), .RSTB(I289421), .Q(I289386) );
DFFARX1 I_16894  ( .D(I487049), .CLK(I2702), .RSTB(I289421), .Q(I289924) );
not I_16895 (I289941,I289924);
nand I_16896 (I289958,I289941,I289506);
and I_16897 (I289975,I289735,I289958);
DFFARX1 I_16898  ( .D(I289975), .CLK(I2702), .RSTB(I289421), .Q(I289413) );
or I_16899 (I290006,I289941,I289752);
DFFARX1 I_16900  ( .D(I290006), .CLK(I2702), .RSTB(I289421), .Q(I289398) );
nand I_16901 (I289401,I289941,I289831);
not I_16902 (I290084,I2709);
not I_16903 (I290101,I90455);
nor I_16904 (I290118,I90452,I90476);
nand I_16905 (I290135,I290118,I90473);
nor I_16906 (I290152,I290101,I90452);
nand I_16907 (I290169,I290152,I90479);
not I_16908 (I290186,I290169);
not I_16909 (I290203,I90452);
nor I_16910 (I290073,I290169,I290203);
not I_16911 (I290234,I290203);
nand I_16912 (I290058,I290169,I290234);
not I_16913 (I290265,I90470);
nor I_16914 (I290282,I290265,I90461);
and I_16915 (I290299,I290282,I90458);
or I_16916 (I290316,I290299,I90467);
DFFARX1 I_16917  ( .D(I290316), .CLK(I2702), .RSTB(I290084), .Q(I290333) );
nor I_16918 (I290350,I290333,I290186);
DFFARX1 I_16919  ( .D(I290333), .CLK(I2702), .RSTB(I290084), .Q(I290367) );
not I_16920 (I290055,I290367);
nand I_16921 (I290398,I290101,I90470);
and I_16922 (I290415,I290398,I290350);
DFFARX1 I_16923  ( .D(I290398), .CLK(I2702), .RSTB(I290084), .Q(I290052) );
DFFARX1 I_16924  ( .D(I90449), .CLK(I2702), .RSTB(I290084), .Q(I290446) );
nor I_16925 (I290463,I290446,I290169);
nand I_16926 (I290070,I290333,I290463);
nor I_16927 (I290494,I290446,I290234);
not I_16928 (I290067,I290446);
nand I_16929 (I290525,I290446,I290135);
and I_16930 (I290542,I290203,I290525);
DFFARX1 I_16931  ( .D(I290542), .CLK(I2702), .RSTB(I290084), .Q(I290046) );
DFFARX1 I_16932  ( .D(I290446), .CLK(I2702), .RSTB(I290084), .Q(I290049) );
DFFARX1 I_16933  ( .D(I90464), .CLK(I2702), .RSTB(I290084), .Q(I290587) );
not I_16934 (I290604,I290587);
nand I_16935 (I290621,I290604,I290169);
and I_16936 (I290638,I290398,I290621);
DFFARX1 I_16937  ( .D(I290638), .CLK(I2702), .RSTB(I290084), .Q(I290076) );
or I_16938 (I290669,I290604,I290415);
DFFARX1 I_16939  ( .D(I290669), .CLK(I2702), .RSTB(I290084), .Q(I290061) );
nand I_16940 (I290064,I290604,I290494);
not I_16941 (I290747,I2709);
not I_16942 (I290764,I663372);
nor I_16943 (I290781,I663390,I663381);
nand I_16944 (I290798,I290781,I663387);
nor I_16945 (I290815,I290764,I663390);
nand I_16946 (I290832,I290815,I663393);
not I_16947 (I290849,I290832);
not I_16948 (I290866,I663390);
nor I_16949 (I290736,I290832,I290866);
not I_16950 (I290897,I290866);
nand I_16951 (I290721,I290832,I290897);
not I_16952 (I290928,I663369);
nor I_16953 (I290945,I290928,I663384);
and I_16954 (I290962,I290945,I663366);
or I_16955 (I290979,I290962,I663375);
DFFARX1 I_16956  ( .D(I290979), .CLK(I2702), .RSTB(I290747), .Q(I290996) );
nor I_16957 (I291013,I290996,I290849);
DFFARX1 I_16958  ( .D(I290996), .CLK(I2702), .RSTB(I290747), .Q(I291030) );
not I_16959 (I290718,I291030);
nand I_16960 (I291061,I290764,I663369);
and I_16961 (I291078,I291061,I291013);
DFFARX1 I_16962  ( .D(I291061), .CLK(I2702), .RSTB(I290747), .Q(I290715) );
DFFARX1 I_16963  ( .D(I663378), .CLK(I2702), .RSTB(I290747), .Q(I291109) );
nor I_16964 (I291126,I291109,I290832);
nand I_16965 (I290733,I290996,I291126);
nor I_16966 (I291157,I291109,I290897);
not I_16967 (I290730,I291109);
nand I_16968 (I291188,I291109,I290798);
and I_16969 (I291205,I290866,I291188);
DFFARX1 I_16970  ( .D(I291205), .CLK(I2702), .RSTB(I290747), .Q(I290709) );
DFFARX1 I_16971  ( .D(I291109), .CLK(I2702), .RSTB(I290747), .Q(I290712) );
DFFARX1 I_16972  ( .D(I663396), .CLK(I2702), .RSTB(I290747), .Q(I291250) );
not I_16973 (I291267,I291250);
nand I_16974 (I291284,I291267,I290832);
and I_16975 (I291301,I291061,I291284);
DFFARX1 I_16976  ( .D(I291301), .CLK(I2702), .RSTB(I290747), .Q(I290739) );
or I_16977 (I291332,I291267,I291078);
DFFARX1 I_16978  ( .D(I291332), .CLK(I2702), .RSTB(I290747), .Q(I290724) );
nand I_16979 (I290727,I291267,I291157);
not I_16980 (I291410,I2709);
not I_16981 (I291427,I644502);
nor I_16982 (I291444,I644520,I644511);
nand I_16983 (I291461,I291444,I644517);
nor I_16984 (I291478,I291427,I644520);
nand I_16985 (I291495,I291478,I644523);
not I_16986 (I291512,I291495);
not I_16987 (I291529,I644520);
nor I_16988 (I291399,I291495,I291529);
not I_16989 (I291560,I291529);
nand I_16990 (I291384,I291495,I291560);
not I_16991 (I291591,I644499);
nor I_16992 (I291608,I291591,I644514);
and I_16993 (I291625,I291608,I644496);
or I_16994 (I291642,I291625,I644505);
DFFARX1 I_16995  ( .D(I291642), .CLK(I2702), .RSTB(I291410), .Q(I291659) );
nor I_16996 (I291676,I291659,I291512);
DFFARX1 I_16997  ( .D(I291659), .CLK(I2702), .RSTB(I291410), .Q(I291693) );
not I_16998 (I291381,I291693);
nand I_16999 (I291724,I291427,I644499);
and I_17000 (I291741,I291724,I291676);
DFFARX1 I_17001  ( .D(I291724), .CLK(I2702), .RSTB(I291410), .Q(I291378) );
DFFARX1 I_17002  ( .D(I644508), .CLK(I2702), .RSTB(I291410), .Q(I291772) );
nor I_17003 (I291789,I291772,I291495);
nand I_17004 (I291396,I291659,I291789);
nor I_17005 (I291820,I291772,I291560);
not I_17006 (I291393,I291772);
nand I_17007 (I291851,I291772,I291461);
and I_17008 (I291868,I291529,I291851);
DFFARX1 I_17009  ( .D(I291868), .CLK(I2702), .RSTB(I291410), .Q(I291372) );
DFFARX1 I_17010  ( .D(I291772), .CLK(I2702), .RSTB(I291410), .Q(I291375) );
DFFARX1 I_17011  ( .D(I644526), .CLK(I2702), .RSTB(I291410), .Q(I291913) );
not I_17012 (I291930,I291913);
nand I_17013 (I291947,I291930,I291495);
and I_17014 (I291964,I291724,I291947);
DFFARX1 I_17015  ( .D(I291964), .CLK(I2702), .RSTB(I291410), .Q(I291402) );
or I_17016 (I291995,I291930,I291741);
DFFARX1 I_17017  ( .D(I291995), .CLK(I2702), .RSTB(I291410), .Q(I291387) );
nand I_17018 (I291390,I291930,I291820);
not I_17019 (I292073,I2709);
not I_17020 (I292090,I96269);
nor I_17021 (I292107,I96266,I96290);
nand I_17022 (I292124,I292107,I96287);
nor I_17023 (I292141,I292090,I96266);
nand I_17024 (I292158,I292141,I96293);
not I_17025 (I292175,I292158);
not I_17026 (I292192,I96266);
nor I_17027 (I292062,I292158,I292192);
not I_17028 (I292223,I292192);
nand I_17029 (I292047,I292158,I292223);
not I_17030 (I292254,I96284);
nor I_17031 (I292271,I292254,I96275);
and I_17032 (I292288,I292271,I96272);
or I_17033 (I292305,I292288,I96281);
DFFARX1 I_17034  ( .D(I292305), .CLK(I2702), .RSTB(I292073), .Q(I292322) );
nor I_17035 (I292339,I292322,I292175);
DFFARX1 I_17036  ( .D(I292322), .CLK(I2702), .RSTB(I292073), .Q(I292356) );
not I_17037 (I292044,I292356);
nand I_17038 (I292387,I292090,I96284);
and I_17039 (I292404,I292387,I292339);
DFFARX1 I_17040  ( .D(I292387), .CLK(I2702), .RSTB(I292073), .Q(I292041) );
DFFARX1 I_17041  ( .D(I96263), .CLK(I2702), .RSTB(I292073), .Q(I292435) );
nor I_17042 (I292452,I292435,I292158);
nand I_17043 (I292059,I292322,I292452);
nor I_17044 (I292483,I292435,I292223);
not I_17045 (I292056,I292435);
nand I_17046 (I292514,I292435,I292124);
and I_17047 (I292531,I292192,I292514);
DFFARX1 I_17048  ( .D(I292531), .CLK(I2702), .RSTB(I292073), .Q(I292035) );
DFFARX1 I_17049  ( .D(I292435), .CLK(I2702), .RSTB(I292073), .Q(I292038) );
DFFARX1 I_17050  ( .D(I96278), .CLK(I2702), .RSTB(I292073), .Q(I292576) );
not I_17051 (I292593,I292576);
nand I_17052 (I292610,I292593,I292158);
and I_17053 (I292627,I292387,I292610);
DFFARX1 I_17054  ( .D(I292627), .CLK(I2702), .RSTB(I292073), .Q(I292065) );
or I_17055 (I292658,I292593,I292404);
DFFARX1 I_17056  ( .D(I292658), .CLK(I2702), .RSTB(I292073), .Q(I292050) );
nand I_17057 (I292053,I292593,I292483);
not I_17058 (I292736,I2709);
not I_17059 (I292753,I15072);
nor I_17060 (I292770,I15078,I15081);
nand I_17061 (I292787,I292770,I15057);
nor I_17062 (I292804,I292753,I15078);
nand I_17063 (I292821,I292804,I15066);
not I_17064 (I292838,I292821);
not I_17065 (I292855,I15078);
nor I_17066 (I292725,I292821,I292855);
not I_17067 (I292886,I292855);
nand I_17068 (I292710,I292821,I292886);
not I_17069 (I292917,I15060);
nor I_17070 (I292934,I292917,I15084);
and I_17071 (I292951,I292934,I15054);
or I_17072 (I292968,I292951,I15063);
DFFARX1 I_17073  ( .D(I292968), .CLK(I2702), .RSTB(I292736), .Q(I292985) );
nor I_17074 (I293002,I292985,I292838);
DFFARX1 I_17075  ( .D(I292985), .CLK(I2702), .RSTB(I292736), .Q(I293019) );
not I_17076 (I292707,I293019);
nand I_17077 (I293050,I292753,I15060);
and I_17078 (I293067,I293050,I293002);
DFFARX1 I_17079  ( .D(I293050), .CLK(I2702), .RSTB(I292736), .Q(I292704) );
DFFARX1 I_17080  ( .D(I15069), .CLK(I2702), .RSTB(I292736), .Q(I293098) );
nor I_17081 (I293115,I293098,I292821);
nand I_17082 (I292722,I292985,I293115);
nor I_17083 (I293146,I293098,I292886);
not I_17084 (I292719,I293098);
nand I_17085 (I293177,I293098,I292787);
and I_17086 (I293194,I292855,I293177);
DFFARX1 I_17087  ( .D(I293194), .CLK(I2702), .RSTB(I292736), .Q(I292698) );
DFFARX1 I_17088  ( .D(I293098), .CLK(I2702), .RSTB(I292736), .Q(I292701) );
DFFARX1 I_17089  ( .D(I15075), .CLK(I2702), .RSTB(I292736), .Q(I293239) );
not I_17090 (I293256,I293239);
nand I_17091 (I293273,I293256,I292821);
and I_17092 (I293290,I293050,I293273);
DFFARX1 I_17093  ( .D(I293290), .CLK(I2702), .RSTB(I292736), .Q(I292728) );
or I_17094 (I293321,I293256,I293067);
DFFARX1 I_17095  ( .D(I293321), .CLK(I2702), .RSTB(I292736), .Q(I292713) );
nand I_17096 (I292716,I293256,I293146);
not I_17097 (I293399,I2709);
not I_17098 (I293416,I399045);
nor I_17099 (I293433,I399042,I399060);
nand I_17100 (I293450,I293433,I399063);
nor I_17101 (I293467,I293416,I399042);
nand I_17102 (I293484,I293467,I399048);
not I_17103 (I293501,I293484);
not I_17104 (I293518,I399042);
nor I_17105 (I293388,I293484,I293518);
not I_17106 (I293549,I293518);
nand I_17107 (I293373,I293484,I293549);
not I_17108 (I293580,I399057);
nor I_17109 (I293597,I293580,I399039);
and I_17110 (I293614,I293597,I399033);
or I_17111 (I293631,I293614,I399051);
DFFARX1 I_17112  ( .D(I293631), .CLK(I2702), .RSTB(I293399), .Q(I293648) );
nor I_17113 (I293665,I293648,I293501);
DFFARX1 I_17114  ( .D(I293648), .CLK(I2702), .RSTB(I293399), .Q(I293682) );
not I_17115 (I293370,I293682);
nand I_17116 (I293713,I293416,I399057);
and I_17117 (I293730,I293713,I293665);
DFFARX1 I_17118  ( .D(I293713), .CLK(I2702), .RSTB(I293399), .Q(I293367) );
DFFARX1 I_17119  ( .D(I399036), .CLK(I2702), .RSTB(I293399), .Q(I293761) );
nor I_17120 (I293778,I293761,I293484);
nand I_17121 (I293385,I293648,I293778);
nor I_17122 (I293809,I293761,I293549);
not I_17123 (I293382,I293761);
nand I_17124 (I293840,I293761,I293450);
and I_17125 (I293857,I293518,I293840);
DFFARX1 I_17126  ( .D(I293857), .CLK(I2702), .RSTB(I293399), .Q(I293361) );
DFFARX1 I_17127  ( .D(I293761), .CLK(I2702), .RSTB(I293399), .Q(I293364) );
DFFARX1 I_17128  ( .D(I399054), .CLK(I2702), .RSTB(I293399), .Q(I293902) );
not I_17129 (I293919,I293902);
nand I_17130 (I293936,I293919,I293484);
and I_17131 (I293953,I293713,I293936);
DFFARX1 I_17132  ( .D(I293953), .CLK(I2702), .RSTB(I293399), .Q(I293391) );
or I_17133 (I293984,I293919,I293730);
DFFARX1 I_17134  ( .D(I293984), .CLK(I2702), .RSTB(I293399), .Q(I293376) );
nand I_17135 (I293379,I293919,I293809);
not I_17136 (I294062,I2709);
not I_17137 (I294079,I645760);
nor I_17138 (I294096,I645778,I645769);
nand I_17139 (I294113,I294096,I645775);
nor I_17140 (I294130,I294079,I645778);
nand I_17141 (I294147,I294130,I645781);
not I_17142 (I294164,I294147);
not I_17143 (I294181,I645778);
nor I_17144 (I294051,I294147,I294181);
not I_17145 (I294212,I294181);
nand I_17146 (I294036,I294147,I294212);
not I_17147 (I294243,I645757);
nor I_17148 (I294260,I294243,I645772);
and I_17149 (I294277,I294260,I645754);
or I_17150 (I294294,I294277,I645763);
DFFARX1 I_17151  ( .D(I294294), .CLK(I2702), .RSTB(I294062), .Q(I294311) );
nor I_17152 (I294328,I294311,I294164);
DFFARX1 I_17153  ( .D(I294311), .CLK(I2702), .RSTB(I294062), .Q(I294345) );
not I_17154 (I294033,I294345);
nand I_17155 (I294376,I294079,I645757);
and I_17156 (I294393,I294376,I294328);
DFFARX1 I_17157  ( .D(I294376), .CLK(I2702), .RSTB(I294062), .Q(I294030) );
DFFARX1 I_17158  ( .D(I645766), .CLK(I2702), .RSTB(I294062), .Q(I294424) );
nor I_17159 (I294441,I294424,I294147);
nand I_17160 (I294048,I294311,I294441);
nor I_17161 (I294472,I294424,I294212);
not I_17162 (I294045,I294424);
nand I_17163 (I294503,I294424,I294113);
and I_17164 (I294520,I294181,I294503);
DFFARX1 I_17165  ( .D(I294520), .CLK(I2702), .RSTB(I294062), .Q(I294024) );
DFFARX1 I_17166  ( .D(I294424), .CLK(I2702), .RSTB(I294062), .Q(I294027) );
DFFARX1 I_17167  ( .D(I645784), .CLK(I2702), .RSTB(I294062), .Q(I294565) );
not I_17168 (I294582,I294565);
nand I_17169 (I294599,I294582,I294147);
and I_17170 (I294616,I294376,I294599);
DFFARX1 I_17171  ( .D(I294616), .CLK(I2702), .RSTB(I294062), .Q(I294054) );
or I_17172 (I294647,I294582,I294393);
DFFARX1 I_17173  ( .D(I294647), .CLK(I2702), .RSTB(I294062), .Q(I294039) );
nand I_17174 (I294042,I294582,I294472);
not I_17175 (I294725,I2709);
not I_17176 (I294742,I642615);
nor I_17177 (I294759,I642633,I642624);
nand I_17178 (I294776,I294759,I642630);
nor I_17179 (I294793,I294742,I642633);
nand I_17180 (I294810,I294793,I642636);
not I_17181 (I294827,I294810);
not I_17182 (I294844,I642633);
nor I_17183 (I294714,I294810,I294844);
not I_17184 (I294875,I294844);
nand I_17185 (I294699,I294810,I294875);
not I_17186 (I294906,I642612);
nor I_17187 (I294923,I294906,I642627);
and I_17188 (I294940,I294923,I642609);
or I_17189 (I294957,I294940,I642618);
DFFARX1 I_17190  ( .D(I294957), .CLK(I2702), .RSTB(I294725), .Q(I294974) );
nor I_17191 (I294991,I294974,I294827);
DFFARX1 I_17192  ( .D(I294974), .CLK(I2702), .RSTB(I294725), .Q(I295008) );
not I_17193 (I294696,I295008);
nand I_17194 (I295039,I294742,I642612);
and I_17195 (I295056,I295039,I294991);
DFFARX1 I_17196  ( .D(I295039), .CLK(I2702), .RSTB(I294725), .Q(I294693) );
DFFARX1 I_17197  ( .D(I642621), .CLK(I2702), .RSTB(I294725), .Q(I295087) );
nor I_17198 (I295104,I295087,I294810);
nand I_17199 (I294711,I294974,I295104);
nor I_17200 (I295135,I295087,I294875);
not I_17201 (I294708,I295087);
nand I_17202 (I295166,I295087,I294776);
and I_17203 (I295183,I294844,I295166);
DFFARX1 I_17204  ( .D(I295183), .CLK(I2702), .RSTB(I294725), .Q(I294687) );
DFFARX1 I_17205  ( .D(I295087), .CLK(I2702), .RSTB(I294725), .Q(I294690) );
DFFARX1 I_17206  ( .D(I642639), .CLK(I2702), .RSTB(I294725), .Q(I295228) );
not I_17207 (I295245,I295228);
nand I_17208 (I295262,I295245,I294810);
and I_17209 (I295279,I295039,I295262);
DFFARX1 I_17210  ( .D(I295279), .CLK(I2702), .RSTB(I294725), .Q(I294717) );
or I_17211 (I295310,I295245,I295056);
DFFARX1 I_17212  ( .D(I295310), .CLK(I2702), .RSTB(I294725), .Q(I294702) );
nand I_17213 (I294705,I295245,I295135);
not I_17214 (I295388,I2709);
not I_17215 (I295405,I125985);
nor I_17216 (I295422,I125982,I126006);
nand I_17217 (I295439,I295422,I126003);
nor I_17218 (I295456,I295405,I125982);
nand I_17219 (I295473,I295456,I126009);
not I_17220 (I295490,I295473);
not I_17221 (I295507,I125982);
nor I_17222 (I295377,I295473,I295507);
not I_17223 (I295538,I295507);
nand I_17224 (I295362,I295473,I295538);
not I_17225 (I295569,I126000);
nor I_17226 (I295586,I295569,I125991);
and I_17227 (I295603,I295586,I125988);
or I_17228 (I295620,I295603,I125997);
DFFARX1 I_17229  ( .D(I295620), .CLK(I2702), .RSTB(I295388), .Q(I295637) );
nor I_17230 (I295654,I295637,I295490);
DFFARX1 I_17231  ( .D(I295637), .CLK(I2702), .RSTB(I295388), .Q(I295671) );
not I_17232 (I295359,I295671);
nand I_17233 (I295702,I295405,I126000);
and I_17234 (I295719,I295702,I295654);
DFFARX1 I_17235  ( .D(I295702), .CLK(I2702), .RSTB(I295388), .Q(I295356) );
DFFARX1 I_17236  ( .D(I125979), .CLK(I2702), .RSTB(I295388), .Q(I295750) );
nor I_17237 (I295767,I295750,I295473);
nand I_17238 (I295374,I295637,I295767);
nor I_17239 (I295798,I295750,I295538);
not I_17240 (I295371,I295750);
nand I_17241 (I295829,I295750,I295439);
and I_17242 (I295846,I295507,I295829);
DFFARX1 I_17243  ( .D(I295846), .CLK(I2702), .RSTB(I295388), .Q(I295350) );
DFFARX1 I_17244  ( .D(I295750), .CLK(I2702), .RSTB(I295388), .Q(I295353) );
DFFARX1 I_17245  ( .D(I125994), .CLK(I2702), .RSTB(I295388), .Q(I295891) );
not I_17246 (I295908,I295891);
nand I_17247 (I295925,I295908,I295473);
and I_17248 (I295942,I295702,I295925);
DFFARX1 I_17249  ( .D(I295942), .CLK(I2702), .RSTB(I295388), .Q(I295380) );
or I_17250 (I295973,I295908,I295719);
DFFARX1 I_17251  ( .D(I295973), .CLK(I2702), .RSTB(I295388), .Q(I295365) );
nand I_17252 (I295368,I295908,I295798);
not I_17253 (I296051,I2709);
not I_17254 (I296068,I357055);
nor I_17255 (I296085,I357052,I357070);
nand I_17256 (I296102,I296085,I357073);
nor I_17257 (I296119,I296068,I357052);
nand I_17258 (I296136,I296119,I357058);
not I_17259 (I296153,I296136);
not I_17260 (I296170,I357052);
nor I_17261 (I296040,I296136,I296170);
not I_17262 (I296201,I296170);
nand I_17263 (I296025,I296136,I296201);
not I_17264 (I296232,I357067);
nor I_17265 (I296249,I296232,I357049);
and I_17266 (I296266,I296249,I357043);
or I_17267 (I296283,I296266,I357061);
DFFARX1 I_17268  ( .D(I296283), .CLK(I2702), .RSTB(I296051), .Q(I296300) );
nor I_17269 (I296317,I296300,I296153);
DFFARX1 I_17270  ( .D(I296300), .CLK(I2702), .RSTB(I296051), .Q(I296334) );
not I_17271 (I296022,I296334);
nand I_17272 (I296365,I296068,I357067);
and I_17273 (I296382,I296365,I296317);
DFFARX1 I_17274  ( .D(I296365), .CLK(I2702), .RSTB(I296051), .Q(I296019) );
DFFARX1 I_17275  ( .D(I357046), .CLK(I2702), .RSTB(I296051), .Q(I296413) );
nor I_17276 (I296430,I296413,I296136);
nand I_17277 (I296037,I296300,I296430);
nor I_17278 (I296461,I296413,I296201);
not I_17279 (I296034,I296413);
nand I_17280 (I296492,I296413,I296102);
and I_17281 (I296509,I296170,I296492);
DFFARX1 I_17282  ( .D(I296509), .CLK(I2702), .RSTB(I296051), .Q(I296013) );
DFFARX1 I_17283  ( .D(I296413), .CLK(I2702), .RSTB(I296051), .Q(I296016) );
DFFARX1 I_17284  ( .D(I357064), .CLK(I2702), .RSTB(I296051), .Q(I296554) );
not I_17285 (I296571,I296554);
nand I_17286 (I296588,I296571,I296136);
and I_17287 (I296605,I296365,I296588);
DFFARX1 I_17288  ( .D(I296605), .CLK(I2702), .RSTB(I296051), .Q(I296043) );
or I_17289 (I296636,I296571,I296382);
DFFARX1 I_17290  ( .D(I296636), .CLK(I2702), .RSTB(I296051), .Q(I296028) );
nand I_17291 (I296031,I296571,I296461);
not I_17292 (I296714,I2709);
not I_17293 (I296731,I591117);
nor I_17294 (I296748,I591114,I591105);
nand I_17295 (I296765,I296748,I591108);
nor I_17296 (I296782,I296731,I591114);
nand I_17297 (I296799,I296782,I591102);
not I_17298 (I296816,I296799);
not I_17299 (I296833,I591114);
nor I_17300 (I296703,I296799,I296833);
not I_17301 (I296864,I296833);
nand I_17302 (I296688,I296799,I296864);
not I_17303 (I296895,I591123);
nor I_17304 (I296912,I296895,I591126);
and I_17305 (I296929,I296912,I591111);
or I_17306 (I296946,I296929,I591099);
DFFARX1 I_17307  ( .D(I296946), .CLK(I2702), .RSTB(I296714), .Q(I296963) );
nor I_17308 (I296980,I296963,I296816);
DFFARX1 I_17309  ( .D(I296963), .CLK(I2702), .RSTB(I296714), .Q(I296997) );
not I_17310 (I296685,I296997);
nand I_17311 (I297028,I296731,I591123);
and I_17312 (I297045,I297028,I296980);
DFFARX1 I_17313  ( .D(I297028), .CLK(I2702), .RSTB(I296714), .Q(I296682) );
DFFARX1 I_17314  ( .D(I591120), .CLK(I2702), .RSTB(I296714), .Q(I297076) );
nor I_17315 (I297093,I297076,I296799);
nand I_17316 (I296700,I296963,I297093);
nor I_17317 (I297124,I297076,I296864);
not I_17318 (I296697,I297076);
nand I_17319 (I297155,I297076,I296765);
and I_17320 (I297172,I296833,I297155);
DFFARX1 I_17321  ( .D(I297172), .CLK(I2702), .RSTB(I296714), .Q(I296676) );
DFFARX1 I_17322  ( .D(I297076), .CLK(I2702), .RSTB(I296714), .Q(I296679) );
DFFARX1 I_17323  ( .D(I591129), .CLK(I2702), .RSTB(I296714), .Q(I297217) );
not I_17324 (I297234,I297217);
nand I_17325 (I297251,I297234,I296799);
and I_17326 (I297268,I297028,I297251);
DFFARX1 I_17327  ( .D(I297268), .CLK(I2702), .RSTB(I296714), .Q(I296706) );
or I_17328 (I297299,I297234,I297045);
DFFARX1 I_17329  ( .D(I297299), .CLK(I2702), .RSTB(I296714), .Q(I296691) );
nand I_17330 (I296694,I297234,I297124);
not I_17331 (I297377,I2709);
not I_17332 (I297394,I245720);
nor I_17333 (I297411,I245693,I245696);
nand I_17334 (I297428,I297411,I245708);
nor I_17335 (I297445,I297394,I245693);
nand I_17336 (I297462,I297445,I245714);
not I_17337 (I297479,I297462);
not I_17338 (I297496,I245693);
nor I_17339 (I297366,I297462,I297496);
not I_17340 (I297527,I297496);
nand I_17341 (I297351,I297462,I297527);
not I_17342 (I297558,I245717);
nor I_17343 (I297575,I297558,I245699);
and I_17344 (I297592,I297575,I245702);
or I_17345 (I297609,I297592,I245723);
DFFARX1 I_17346  ( .D(I297609), .CLK(I2702), .RSTB(I297377), .Q(I297626) );
nor I_17347 (I297643,I297626,I297479);
DFFARX1 I_17348  ( .D(I297626), .CLK(I2702), .RSTB(I297377), .Q(I297660) );
not I_17349 (I297348,I297660);
nand I_17350 (I297691,I297394,I245717);
and I_17351 (I297708,I297691,I297643);
DFFARX1 I_17352  ( .D(I297691), .CLK(I2702), .RSTB(I297377), .Q(I297345) );
DFFARX1 I_17353  ( .D(I245705), .CLK(I2702), .RSTB(I297377), .Q(I297739) );
nor I_17354 (I297756,I297739,I297462);
nand I_17355 (I297363,I297626,I297756);
nor I_17356 (I297787,I297739,I297527);
not I_17357 (I297360,I297739);
nand I_17358 (I297818,I297739,I297428);
and I_17359 (I297835,I297496,I297818);
DFFARX1 I_17360  ( .D(I297835), .CLK(I2702), .RSTB(I297377), .Q(I297339) );
DFFARX1 I_17361  ( .D(I297739), .CLK(I2702), .RSTB(I297377), .Q(I297342) );
DFFARX1 I_17362  ( .D(I245711), .CLK(I2702), .RSTB(I297377), .Q(I297880) );
not I_17363 (I297897,I297880);
nand I_17364 (I297914,I297897,I297462);
and I_17365 (I297931,I297691,I297914);
DFFARX1 I_17366  ( .D(I297931), .CLK(I2702), .RSTB(I297377), .Q(I297369) );
or I_17367 (I297962,I297897,I297708);
DFFARX1 I_17368  ( .D(I297962), .CLK(I2702), .RSTB(I297377), .Q(I297354) );
nand I_17369 (I297357,I297897,I297787);
not I_17370 (I298040,I2709);
not I_17371 (I298057,I647018);
nor I_17372 (I298074,I647036,I647027);
nand I_17373 (I298091,I298074,I647033);
nor I_17374 (I298108,I298057,I647036);
nand I_17375 (I298125,I298108,I647039);
not I_17376 (I298142,I298125);
not I_17377 (I298159,I647036);
nor I_17378 (I298029,I298125,I298159);
not I_17379 (I298190,I298159);
nand I_17380 (I298014,I298125,I298190);
not I_17381 (I298221,I647015);
nor I_17382 (I298238,I298221,I647030);
and I_17383 (I298255,I298238,I647012);
or I_17384 (I298272,I298255,I647021);
DFFARX1 I_17385  ( .D(I298272), .CLK(I2702), .RSTB(I298040), .Q(I298289) );
nor I_17386 (I298306,I298289,I298142);
DFFARX1 I_17387  ( .D(I298289), .CLK(I2702), .RSTB(I298040), .Q(I298323) );
not I_17388 (I298011,I298323);
nand I_17389 (I298354,I298057,I647015);
and I_17390 (I298371,I298354,I298306);
DFFARX1 I_17391  ( .D(I298354), .CLK(I2702), .RSTB(I298040), .Q(I298008) );
DFFARX1 I_17392  ( .D(I647024), .CLK(I2702), .RSTB(I298040), .Q(I298402) );
nor I_17393 (I298419,I298402,I298125);
nand I_17394 (I298026,I298289,I298419);
nor I_17395 (I298450,I298402,I298190);
not I_17396 (I298023,I298402);
nand I_17397 (I298481,I298402,I298091);
and I_17398 (I298498,I298159,I298481);
DFFARX1 I_17399  ( .D(I298498), .CLK(I2702), .RSTB(I298040), .Q(I298002) );
DFFARX1 I_17400  ( .D(I298402), .CLK(I2702), .RSTB(I298040), .Q(I298005) );
DFFARX1 I_17401  ( .D(I647042), .CLK(I2702), .RSTB(I298040), .Q(I298543) );
not I_17402 (I298560,I298543);
nand I_17403 (I298577,I298560,I298125);
and I_17404 (I298594,I298354,I298577);
DFFARX1 I_17405  ( .D(I298594), .CLK(I2702), .RSTB(I298040), .Q(I298032) );
or I_17406 (I298625,I298560,I298371);
DFFARX1 I_17407  ( .D(I298625), .CLK(I2702), .RSTB(I298040), .Q(I298017) );
nand I_17408 (I298020,I298560,I298450);
not I_17409 (I298703,I2709);
not I_17410 (I298720,I491327);
nor I_17411 (I298737,I491324,I491321);
nand I_17412 (I298754,I298737,I491309);
nor I_17413 (I298771,I298720,I491324);
nand I_17414 (I298788,I298771,I491330);
not I_17415 (I298805,I298788);
not I_17416 (I298822,I491324);
nor I_17417 (I298692,I298788,I298822);
not I_17418 (I298853,I298822);
nand I_17419 (I298677,I298788,I298853);
not I_17420 (I298884,I491312);
nor I_17421 (I298901,I298884,I491318);
and I_17422 (I298918,I298901,I491315);
or I_17423 (I298935,I298918,I491339);
DFFARX1 I_17424  ( .D(I298935), .CLK(I2702), .RSTB(I298703), .Q(I298952) );
nor I_17425 (I298969,I298952,I298805);
DFFARX1 I_17426  ( .D(I298952), .CLK(I2702), .RSTB(I298703), .Q(I298986) );
not I_17427 (I298674,I298986);
nand I_17428 (I299017,I298720,I491312);
and I_17429 (I299034,I299017,I298969);
DFFARX1 I_17430  ( .D(I299017), .CLK(I2702), .RSTB(I298703), .Q(I298671) );
DFFARX1 I_17431  ( .D(I491336), .CLK(I2702), .RSTB(I298703), .Q(I299065) );
nor I_17432 (I299082,I299065,I298788);
nand I_17433 (I298689,I298952,I299082);
nor I_17434 (I299113,I299065,I298853);
not I_17435 (I298686,I299065);
nand I_17436 (I299144,I299065,I298754);
and I_17437 (I299161,I298822,I299144);
DFFARX1 I_17438  ( .D(I299161), .CLK(I2702), .RSTB(I298703), .Q(I298665) );
DFFARX1 I_17439  ( .D(I299065), .CLK(I2702), .RSTB(I298703), .Q(I298668) );
DFFARX1 I_17440  ( .D(I491333), .CLK(I2702), .RSTB(I298703), .Q(I299206) );
not I_17441 (I299223,I299206);
nand I_17442 (I299240,I299223,I298788);
and I_17443 (I299257,I299017,I299240);
DFFARX1 I_17444  ( .D(I299257), .CLK(I2702), .RSTB(I298703), .Q(I298695) );
or I_17445 (I299288,I299223,I299034);
DFFARX1 I_17446  ( .D(I299288), .CLK(I2702), .RSTB(I298703), .Q(I298680) );
nand I_17447 (I298683,I299223,I299113);
not I_17448 (I299366,I2709);
not I_17449 (I299383,I60739);
nor I_17450 (I299400,I60736,I60760);
nand I_17451 (I299417,I299400,I60757);
nor I_17452 (I299434,I299383,I60736);
nand I_17453 (I299451,I299434,I60763);
not I_17454 (I299468,I299451);
not I_17455 (I299485,I60736);
nor I_17456 (I299355,I299451,I299485);
not I_17457 (I299516,I299485);
nand I_17458 (I299340,I299451,I299516);
not I_17459 (I299547,I60754);
nor I_17460 (I299564,I299547,I60745);
and I_17461 (I299581,I299564,I60742);
or I_17462 (I299598,I299581,I60751);
DFFARX1 I_17463  ( .D(I299598), .CLK(I2702), .RSTB(I299366), .Q(I299615) );
nor I_17464 (I299632,I299615,I299468);
DFFARX1 I_17465  ( .D(I299615), .CLK(I2702), .RSTB(I299366), .Q(I299649) );
not I_17466 (I299337,I299649);
nand I_17467 (I299680,I299383,I60754);
and I_17468 (I299697,I299680,I299632);
DFFARX1 I_17469  ( .D(I299680), .CLK(I2702), .RSTB(I299366), .Q(I299334) );
DFFARX1 I_17470  ( .D(I60733), .CLK(I2702), .RSTB(I299366), .Q(I299728) );
nor I_17471 (I299745,I299728,I299451);
nand I_17472 (I299352,I299615,I299745);
nor I_17473 (I299776,I299728,I299516);
not I_17474 (I299349,I299728);
nand I_17475 (I299807,I299728,I299417);
and I_17476 (I299824,I299485,I299807);
DFFARX1 I_17477  ( .D(I299824), .CLK(I2702), .RSTB(I299366), .Q(I299328) );
DFFARX1 I_17478  ( .D(I299728), .CLK(I2702), .RSTB(I299366), .Q(I299331) );
DFFARX1 I_17479  ( .D(I60748), .CLK(I2702), .RSTB(I299366), .Q(I299869) );
not I_17480 (I299886,I299869);
nand I_17481 (I299903,I299886,I299451);
and I_17482 (I299920,I299680,I299903);
DFFARX1 I_17483  ( .D(I299920), .CLK(I2702), .RSTB(I299366), .Q(I299358) );
or I_17484 (I299951,I299886,I299697);
DFFARX1 I_17485  ( .D(I299951), .CLK(I2702), .RSTB(I299366), .Q(I299343) );
nand I_17486 (I299346,I299886,I299776);
not I_17487 (I300029,I2709);
not I_17488 (I300046,I406797);
nor I_17489 (I300063,I406794,I406812);
nand I_17490 (I300080,I300063,I406815);
nor I_17491 (I300097,I300046,I406794);
nand I_17492 (I300114,I300097,I406800);
not I_17493 (I300131,I300114);
not I_17494 (I300148,I406794);
nor I_17495 (I300018,I300114,I300148);
not I_17496 (I300179,I300148);
nand I_17497 (I300003,I300114,I300179);
not I_17498 (I300210,I406809);
nor I_17499 (I300227,I300210,I406791);
and I_17500 (I300244,I300227,I406785);
or I_17501 (I300261,I300244,I406803);
DFFARX1 I_17502  ( .D(I300261), .CLK(I2702), .RSTB(I300029), .Q(I300278) );
nor I_17503 (I300295,I300278,I300131);
DFFARX1 I_17504  ( .D(I300278), .CLK(I2702), .RSTB(I300029), .Q(I300312) );
not I_17505 (I300000,I300312);
nand I_17506 (I300343,I300046,I406809);
and I_17507 (I300360,I300343,I300295);
DFFARX1 I_17508  ( .D(I300343), .CLK(I2702), .RSTB(I300029), .Q(I299997) );
DFFARX1 I_17509  ( .D(I406788), .CLK(I2702), .RSTB(I300029), .Q(I300391) );
nor I_17510 (I300408,I300391,I300114);
nand I_17511 (I300015,I300278,I300408);
nor I_17512 (I300439,I300391,I300179);
not I_17513 (I300012,I300391);
nand I_17514 (I300470,I300391,I300080);
and I_17515 (I300487,I300148,I300470);
DFFARX1 I_17516  ( .D(I300487), .CLK(I2702), .RSTB(I300029), .Q(I299991) );
DFFARX1 I_17517  ( .D(I300391), .CLK(I2702), .RSTB(I300029), .Q(I299994) );
DFFARX1 I_17518  ( .D(I406806), .CLK(I2702), .RSTB(I300029), .Q(I300532) );
not I_17519 (I300549,I300532);
nand I_17520 (I300566,I300549,I300114);
and I_17521 (I300583,I300343,I300566);
DFFARX1 I_17522  ( .D(I300583), .CLK(I2702), .RSTB(I300029), .Q(I300021) );
or I_17523 (I300614,I300549,I300360);
DFFARX1 I_17524  ( .D(I300614), .CLK(I2702), .RSTB(I300029), .Q(I300006) );
nand I_17525 (I300009,I300549,I300439);
not I_17526 (I300692,I2709);
not I_17527 (I300709,I524477);
nor I_17528 (I300726,I524486,I524468);
nand I_17529 (I300743,I300726,I524489);
nor I_17530 (I300760,I300709,I524486);
nand I_17531 (I300777,I300760,I524480);
not I_17532 (I300794,I300777);
not I_17533 (I300811,I524486);
nor I_17534 (I300681,I300777,I300811);
not I_17535 (I300842,I300811);
nand I_17536 (I300666,I300777,I300842);
not I_17537 (I300873,I524474);
nor I_17538 (I300890,I300873,I524465);
and I_17539 (I300907,I300890,I524462);
or I_17540 (I300924,I300907,I524459);
DFFARX1 I_17541  ( .D(I300924), .CLK(I2702), .RSTB(I300692), .Q(I300941) );
nor I_17542 (I300958,I300941,I300794);
DFFARX1 I_17543  ( .D(I300941), .CLK(I2702), .RSTB(I300692), .Q(I300975) );
not I_17544 (I300663,I300975);
nand I_17545 (I301006,I300709,I524474);
and I_17546 (I301023,I301006,I300958);
DFFARX1 I_17547  ( .D(I301006), .CLK(I2702), .RSTB(I300692), .Q(I300660) );
DFFARX1 I_17548  ( .D(I524483), .CLK(I2702), .RSTB(I300692), .Q(I301054) );
nor I_17549 (I301071,I301054,I300777);
nand I_17550 (I300678,I300941,I301071);
nor I_17551 (I301102,I301054,I300842);
not I_17552 (I300675,I301054);
nand I_17553 (I301133,I301054,I300743);
and I_17554 (I301150,I300811,I301133);
DFFARX1 I_17555  ( .D(I301150), .CLK(I2702), .RSTB(I300692), .Q(I300654) );
DFFARX1 I_17556  ( .D(I301054), .CLK(I2702), .RSTB(I300692), .Q(I300657) );
DFFARX1 I_17557  ( .D(I524471), .CLK(I2702), .RSTB(I300692), .Q(I301195) );
not I_17558 (I301212,I301195);
nand I_17559 (I301229,I301212,I300777);
and I_17560 (I301246,I301006,I301229);
DFFARX1 I_17561  ( .D(I301246), .CLK(I2702), .RSTB(I300692), .Q(I300684) );
or I_17562 (I301277,I301212,I301023);
DFFARX1 I_17563  ( .D(I301277), .CLK(I2702), .RSTB(I300692), .Q(I300669) );
nand I_17564 (I300672,I301212,I301102);
not I_17565 (I301355,I2709);
not I_17566 (I301372,I354471);
nor I_17567 (I301389,I354468,I354486);
nand I_17568 (I301406,I301389,I354489);
nor I_17569 (I301423,I301372,I354468);
nand I_17570 (I301440,I301423,I354474);
not I_17571 (I301457,I301440);
not I_17572 (I301474,I354468);
nor I_17573 (I301344,I301440,I301474);
not I_17574 (I301505,I301474);
nand I_17575 (I301329,I301440,I301505);
not I_17576 (I301536,I354483);
nor I_17577 (I301553,I301536,I354465);
and I_17578 (I301570,I301553,I354459);
or I_17579 (I301587,I301570,I354477);
DFFARX1 I_17580  ( .D(I301587), .CLK(I2702), .RSTB(I301355), .Q(I301604) );
nor I_17581 (I301621,I301604,I301457);
DFFARX1 I_17582  ( .D(I301604), .CLK(I2702), .RSTB(I301355), .Q(I301638) );
not I_17583 (I301326,I301638);
nand I_17584 (I301669,I301372,I354483);
and I_17585 (I301686,I301669,I301621);
DFFARX1 I_17586  ( .D(I301669), .CLK(I2702), .RSTB(I301355), .Q(I301323) );
DFFARX1 I_17587  ( .D(I354462), .CLK(I2702), .RSTB(I301355), .Q(I301717) );
nor I_17588 (I301734,I301717,I301440);
nand I_17589 (I301341,I301604,I301734);
nor I_17590 (I301765,I301717,I301505);
not I_17591 (I301338,I301717);
nand I_17592 (I301796,I301717,I301406);
and I_17593 (I301813,I301474,I301796);
DFFARX1 I_17594  ( .D(I301813), .CLK(I2702), .RSTB(I301355), .Q(I301317) );
DFFARX1 I_17595  ( .D(I301717), .CLK(I2702), .RSTB(I301355), .Q(I301320) );
DFFARX1 I_17596  ( .D(I354480), .CLK(I2702), .RSTB(I301355), .Q(I301858) );
not I_17597 (I301875,I301858);
nand I_17598 (I301892,I301875,I301440);
and I_17599 (I301909,I301669,I301892);
DFFARX1 I_17600  ( .D(I301909), .CLK(I2702), .RSTB(I301355), .Q(I301347) );
or I_17601 (I301940,I301875,I301686);
DFFARX1 I_17602  ( .D(I301940), .CLK(I2702), .RSTB(I301355), .Q(I301332) );
nand I_17603 (I301335,I301875,I301765);
not I_17604 (I302018,I2709);
not I_17605 (I302035,I690374);
nor I_17606 (I302052,I690365,I690371);
nand I_17607 (I302069,I302052,I690383);
nor I_17608 (I302086,I302035,I690365);
nand I_17609 (I302103,I302086,I690368);
not I_17610 (I302120,I302103);
not I_17611 (I302137,I690365);
nor I_17612 (I302007,I302103,I302137);
not I_17613 (I302168,I302137);
nand I_17614 (I301992,I302103,I302168);
not I_17615 (I302199,I690392);
nor I_17616 (I302216,I302199,I690386);
and I_17617 (I302233,I302216,I690377);
or I_17618 (I302250,I302233,I690362);
DFFARX1 I_17619  ( .D(I302250), .CLK(I2702), .RSTB(I302018), .Q(I302267) );
nor I_17620 (I302284,I302267,I302120);
DFFARX1 I_17621  ( .D(I302267), .CLK(I2702), .RSTB(I302018), .Q(I302301) );
not I_17622 (I301989,I302301);
nand I_17623 (I302332,I302035,I690392);
and I_17624 (I302349,I302332,I302284);
DFFARX1 I_17625  ( .D(I302332), .CLK(I2702), .RSTB(I302018), .Q(I301986) );
DFFARX1 I_17626  ( .D(I690380), .CLK(I2702), .RSTB(I302018), .Q(I302380) );
nor I_17627 (I302397,I302380,I302103);
nand I_17628 (I302004,I302267,I302397);
nor I_17629 (I302428,I302380,I302168);
not I_17630 (I302001,I302380);
nand I_17631 (I302459,I302380,I302069);
and I_17632 (I302476,I302137,I302459);
DFFARX1 I_17633  ( .D(I302476), .CLK(I2702), .RSTB(I302018), .Q(I301980) );
DFFARX1 I_17634  ( .D(I302380), .CLK(I2702), .RSTB(I302018), .Q(I301983) );
DFFARX1 I_17635  ( .D(I690389), .CLK(I2702), .RSTB(I302018), .Q(I302521) );
not I_17636 (I302538,I302521);
nand I_17637 (I302555,I302538,I302103);
and I_17638 (I302572,I302332,I302555);
DFFARX1 I_17639  ( .D(I302572), .CLK(I2702), .RSTB(I302018), .Q(I302010) );
or I_17640 (I302603,I302538,I302349);
DFFARX1 I_17641  ( .D(I302603), .CLK(I2702), .RSTB(I302018), .Q(I301995) );
nand I_17642 (I301998,I302538,I302428);
not I_17643 (I302681,I2709);
not I_17644 (I302698,I700778);
nor I_17645 (I302715,I700769,I700775);
nand I_17646 (I302732,I302715,I700787);
nor I_17647 (I302749,I302698,I700769);
nand I_17648 (I302766,I302749,I700772);
not I_17649 (I302783,I302766);
not I_17650 (I302800,I700769);
nor I_17651 (I302670,I302766,I302800);
not I_17652 (I302831,I302800);
nand I_17653 (I302655,I302766,I302831);
not I_17654 (I302862,I700796);
nor I_17655 (I302879,I302862,I700790);
and I_17656 (I302896,I302879,I700781);
or I_17657 (I302913,I302896,I700766);
DFFARX1 I_17658  ( .D(I302913), .CLK(I2702), .RSTB(I302681), .Q(I302930) );
nor I_17659 (I302947,I302930,I302783);
DFFARX1 I_17660  ( .D(I302930), .CLK(I2702), .RSTB(I302681), .Q(I302964) );
not I_17661 (I302652,I302964);
nand I_17662 (I302995,I302698,I700796);
and I_17663 (I303012,I302995,I302947);
DFFARX1 I_17664  ( .D(I302995), .CLK(I2702), .RSTB(I302681), .Q(I302649) );
DFFARX1 I_17665  ( .D(I700784), .CLK(I2702), .RSTB(I302681), .Q(I303043) );
nor I_17666 (I303060,I303043,I302766);
nand I_17667 (I302667,I302930,I303060);
nor I_17668 (I303091,I303043,I302831);
not I_17669 (I302664,I303043);
nand I_17670 (I303122,I303043,I302732);
and I_17671 (I303139,I302800,I303122);
DFFARX1 I_17672  ( .D(I303139), .CLK(I2702), .RSTB(I302681), .Q(I302643) );
DFFARX1 I_17673  ( .D(I303043), .CLK(I2702), .RSTB(I302681), .Q(I302646) );
DFFARX1 I_17674  ( .D(I700793), .CLK(I2702), .RSTB(I302681), .Q(I303184) );
not I_17675 (I303201,I303184);
nand I_17676 (I303218,I303201,I302766);
and I_17677 (I303235,I302995,I303218);
DFFARX1 I_17678  ( .D(I303235), .CLK(I2702), .RSTB(I302681), .Q(I302673) );
or I_17679 (I303266,I303201,I303012);
DFFARX1 I_17680  ( .D(I303266), .CLK(I2702), .RSTB(I302681), .Q(I302658) );
nand I_17681 (I302661,I303201,I303091);
not I_17682 (I303344,I2709);
not I_17683 (I303361,I155460);
nor I_17684 (I303378,I155466,I155472);
nand I_17685 (I303395,I303378,I155475);
nor I_17686 (I303412,I303361,I155466);
nand I_17687 (I303429,I303412,I155457);
not I_17688 (I303446,I303429);
not I_17689 (I303463,I155466);
nor I_17690 (I303333,I303429,I303463);
not I_17691 (I303494,I303463);
nand I_17692 (I303318,I303429,I303494);
not I_17693 (I303525,I155469);
nor I_17694 (I303542,I303525,I155463);
and I_17695 (I303559,I303542,I155478);
or I_17696 (I303576,I303559,I155484);
DFFARX1 I_17697  ( .D(I303576), .CLK(I2702), .RSTB(I303344), .Q(I303593) );
nor I_17698 (I303610,I303593,I303446);
DFFARX1 I_17699  ( .D(I303593), .CLK(I2702), .RSTB(I303344), .Q(I303627) );
not I_17700 (I303315,I303627);
nand I_17701 (I303658,I303361,I155469);
and I_17702 (I303675,I303658,I303610);
DFFARX1 I_17703  ( .D(I303658), .CLK(I2702), .RSTB(I303344), .Q(I303312) );
DFFARX1 I_17704  ( .D(I155481), .CLK(I2702), .RSTB(I303344), .Q(I303706) );
nor I_17705 (I303723,I303706,I303429);
nand I_17706 (I303330,I303593,I303723);
nor I_17707 (I303754,I303706,I303494);
not I_17708 (I303327,I303706);
nand I_17709 (I303785,I303706,I303395);
and I_17710 (I303802,I303463,I303785);
DFFARX1 I_17711  ( .D(I303802), .CLK(I2702), .RSTB(I303344), .Q(I303306) );
DFFARX1 I_17712  ( .D(I303706), .CLK(I2702), .RSTB(I303344), .Q(I303309) );
DFFARX1 I_17713  ( .D(I155487), .CLK(I2702), .RSTB(I303344), .Q(I303847) );
not I_17714 (I303864,I303847);
nand I_17715 (I303881,I303864,I303429);
and I_17716 (I303898,I303658,I303881);
DFFARX1 I_17717  ( .D(I303898), .CLK(I2702), .RSTB(I303344), .Q(I303336) );
or I_17718 (I303929,I303864,I303675);
DFFARX1 I_17719  ( .D(I303929), .CLK(I2702), .RSTB(I303344), .Q(I303321) );
nand I_17720 (I303324,I303864,I303754);
not I_17721 (I304007,I2709);
not I_17722 (I304024,I577432);
nor I_17723 (I304041,I577429,I577420);
nand I_17724 (I304058,I304041,I577423);
nor I_17725 (I304075,I304024,I577429);
nand I_17726 (I304092,I304075,I577417);
not I_17727 (I304109,I304092);
not I_17728 (I304126,I577429);
nor I_17729 (I303996,I304092,I304126);
not I_17730 (I304157,I304126);
nand I_17731 (I303981,I304092,I304157);
not I_17732 (I304188,I577438);
nor I_17733 (I304205,I304188,I577441);
and I_17734 (I304222,I304205,I577426);
or I_17735 (I304239,I304222,I577414);
DFFARX1 I_17736  ( .D(I304239), .CLK(I2702), .RSTB(I304007), .Q(I304256) );
nor I_17737 (I304273,I304256,I304109);
DFFARX1 I_17738  ( .D(I304256), .CLK(I2702), .RSTB(I304007), .Q(I304290) );
not I_17739 (I303978,I304290);
nand I_17740 (I304321,I304024,I577438);
and I_17741 (I304338,I304321,I304273);
DFFARX1 I_17742  ( .D(I304321), .CLK(I2702), .RSTB(I304007), .Q(I303975) );
DFFARX1 I_17743  ( .D(I577435), .CLK(I2702), .RSTB(I304007), .Q(I304369) );
nor I_17744 (I304386,I304369,I304092);
nand I_17745 (I303993,I304256,I304386);
nor I_17746 (I304417,I304369,I304157);
not I_17747 (I303990,I304369);
nand I_17748 (I304448,I304369,I304058);
and I_17749 (I304465,I304126,I304448);
DFFARX1 I_17750  ( .D(I304465), .CLK(I2702), .RSTB(I304007), .Q(I303969) );
DFFARX1 I_17751  ( .D(I304369), .CLK(I2702), .RSTB(I304007), .Q(I303972) );
DFFARX1 I_17752  ( .D(I577444), .CLK(I2702), .RSTB(I304007), .Q(I304510) );
not I_17753 (I304527,I304510);
nand I_17754 (I304544,I304527,I304092);
and I_17755 (I304561,I304321,I304544);
DFFARX1 I_17756  ( .D(I304561), .CLK(I2702), .RSTB(I304007), .Q(I303999) );
or I_17757 (I304592,I304527,I304338);
DFFARX1 I_17758  ( .D(I304592), .CLK(I2702), .RSTB(I304007), .Q(I303984) );
nand I_17759 (I303987,I304527,I304417);
not I_17760 (I304670,I2709);
not I_17761 (I304687,I514957);
nor I_17762 (I304704,I514966,I514948);
nand I_17763 (I304721,I304704,I514969);
nor I_17764 (I304738,I304687,I514966);
nand I_17765 (I304755,I304738,I514960);
not I_17766 (I304772,I304755);
not I_17767 (I304789,I514966);
nor I_17768 (I304659,I304755,I304789);
not I_17769 (I304820,I304789);
nand I_17770 (I304644,I304755,I304820);
not I_17771 (I304851,I514954);
nor I_17772 (I304868,I304851,I514945);
and I_17773 (I304885,I304868,I514942);
or I_17774 (I304902,I304885,I514939);
DFFARX1 I_17775  ( .D(I304902), .CLK(I2702), .RSTB(I304670), .Q(I304919) );
nor I_17776 (I304936,I304919,I304772);
DFFARX1 I_17777  ( .D(I304919), .CLK(I2702), .RSTB(I304670), .Q(I304953) );
not I_17778 (I304641,I304953);
nand I_17779 (I304984,I304687,I514954);
and I_17780 (I305001,I304984,I304936);
DFFARX1 I_17781  ( .D(I304984), .CLK(I2702), .RSTB(I304670), .Q(I304638) );
DFFARX1 I_17782  ( .D(I514963), .CLK(I2702), .RSTB(I304670), .Q(I305032) );
nor I_17783 (I305049,I305032,I304755);
nand I_17784 (I304656,I304919,I305049);
nor I_17785 (I305080,I305032,I304820);
not I_17786 (I304653,I305032);
nand I_17787 (I305111,I305032,I304721);
and I_17788 (I305128,I304789,I305111);
DFFARX1 I_17789  ( .D(I305128), .CLK(I2702), .RSTB(I304670), .Q(I304632) );
DFFARX1 I_17790  ( .D(I305032), .CLK(I2702), .RSTB(I304670), .Q(I304635) );
DFFARX1 I_17791  ( .D(I514951), .CLK(I2702), .RSTB(I304670), .Q(I305173) );
not I_17792 (I305190,I305173);
nand I_17793 (I305207,I305190,I304755);
and I_17794 (I305224,I304984,I305207);
DFFARX1 I_17795  ( .D(I305224), .CLK(I2702), .RSTB(I304670), .Q(I304662) );
or I_17796 (I305255,I305190,I305001);
DFFARX1 I_17797  ( .D(I305255), .CLK(I2702), .RSTB(I304670), .Q(I304647) );
nand I_17798 (I304650,I305190,I305080);
not I_17799 (I305333,I2709);
not I_17800 (I305350,I710604);
nor I_17801 (I305367,I710595,I710601);
nand I_17802 (I305384,I305367,I710613);
nor I_17803 (I305401,I305350,I710595);
nand I_17804 (I305418,I305401,I710598);
not I_17805 (I305435,I305418);
not I_17806 (I305452,I710595);
nor I_17807 (I305322,I305418,I305452);
not I_17808 (I305483,I305452);
nand I_17809 (I305307,I305418,I305483);
not I_17810 (I305514,I710622);
nor I_17811 (I305531,I305514,I710616);
and I_17812 (I305548,I305531,I710607);
or I_17813 (I305565,I305548,I710592);
DFFARX1 I_17814  ( .D(I305565), .CLK(I2702), .RSTB(I305333), .Q(I305582) );
nor I_17815 (I305599,I305582,I305435);
DFFARX1 I_17816  ( .D(I305582), .CLK(I2702), .RSTB(I305333), .Q(I305616) );
not I_17817 (I305304,I305616);
nand I_17818 (I305647,I305350,I710622);
and I_17819 (I305664,I305647,I305599);
DFFARX1 I_17820  ( .D(I305647), .CLK(I2702), .RSTB(I305333), .Q(I305301) );
DFFARX1 I_17821  ( .D(I710610), .CLK(I2702), .RSTB(I305333), .Q(I305695) );
nor I_17822 (I305712,I305695,I305418);
nand I_17823 (I305319,I305582,I305712);
nor I_17824 (I305743,I305695,I305483);
not I_17825 (I305316,I305695);
nand I_17826 (I305774,I305695,I305384);
and I_17827 (I305791,I305452,I305774);
DFFARX1 I_17828  ( .D(I305791), .CLK(I2702), .RSTB(I305333), .Q(I305295) );
DFFARX1 I_17829  ( .D(I305695), .CLK(I2702), .RSTB(I305333), .Q(I305298) );
DFFARX1 I_17830  ( .D(I710619), .CLK(I2702), .RSTB(I305333), .Q(I305836) );
not I_17831 (I305853,I305836);
nand I_17832 (I305870,I305853,I305418);
and I_17833 (I305887,I305647,I305870);
DFFARX1 I_17834  ( .D(I305887), .CLK(I2702), .RSTB(I305333), .Q(I305325) );
or I_17835 (I305918,I305853,I305664);
DFFARX1 I_17836  ( .D(I305918), .CLK(I2702), .RSTB(I305333), .Q(I305310) );
nand I_17837 (I305313,I305853,I305743);
not I_17838 (I305996,I2709);
not I_17839 (I306013,I211201);
nor I_17840 (I306030,I211195,I211186);
nand I_17841 (I306047,I306030,I211198);
nor I_17842 (I306064,I306013,I211195);
nand I_17843 (I306081,I306064,I211213);
not I_17844 (I306098,I306081);
not I_17845 (I306115,I211195);
nor I_17846 (I305985,I306081,I306115);
not I_17847 (I306146,I306115);
nand I_17848 (I305970,I306081,I306146);
not I_17849 (I306177,I211189);
nor I_17850 (I306194,I306177,I211183);
and I_17851 (I306211,I306194,I211210);
or I_17852 (I306228,I306211,I211207);
DFFARX1 I_17853  ( .D(I306228), .CLK(I2702), .RSTB(I305996), .Q(I306245) );
nor I_17854 (I306262,I306245,I306098);
DFFARX1 I_17855  ( .D(I306245), .CLK(I2702), .RSTB(I305996), .Q(I306279) );
not I_17856 (I305967,I306279);
nand I_17857 (I306310,I306013,I211189);
and I_17858 (I306327,I306310,I306262);
DFFARX1 I_17859  ( .D(I306310), .CLK(I2702), .RSTB(I305996), .Q(I305964) );
DFFARX1 I_17860  ( .D(I211204), .CLK(I2702), .RSTB(I305996), .Q(I306358) );
nor I_17861 (I306375,I306358,I306081);
nand I_17862 (I305982,I306245,I306375);
nor I_17863 (I306406,I306358,I306146);
not I_17864 (I305979,I306358);
nand I_17865 (I306437,I306358,I306047);
and I_17866 (I306454,I306115,I306437);
DFFARX1 I_17867  ( .D(I306454), .CLK(I2702), .RSTB(I305996), .Q(I305958) );
DFFARX1 I_17868  ( .D(I306358), .CLK(I2702), .RSTB(I305996), .Q(I305961) );
DFFARX1 I_17869  ( .D(I211192), .CLK(I2702), .RSTB(I305996), .Q(I306499) );
not I_17870 (I306516,I306499);
nand I_17871 (I306533,I306516,I306081);
and I_17872 (I306550,I306310,I306533);
DFFARX1 I_17873  ( .D(I306550), .CLK(I2702), .RSTB(I305996), .Q(I305988) );
or I_17874 (I306581,I306516,I306327);
DFFARX1 I_17875  ( .D(I306581), .CLK(I2702), .RSTB(I305996), .Q(I305973) );
nand I_17876 (I305976,I306516,I306406);
not I_17877 (I306659,I2709);
not I_17878 (I306676,I420527);
nor I_17879 (I306693,I420530,I420536);
nand I_17880 (I306710,I306693,I420542);
nor I_17881 (I306727,I306676,I420530);
nand I_17882 (I306744,I306727,I420521);
not I_17883 (I306761,I306744);
not I_17884 (I306778,I420530);
nor I_17885 (I306648,I306744,I306778);
not I_17886 (I306809,I306778);
nand I_17887 (I306633,I306744,I306809);
not I_17888 (I306840,I420533);
nor I_17889 (I306857,I306840,I420548);
and I_17890 (I306874,I306857,I420551);
or I_17891 (I306891,I306874,I420524);
DFFARX1 I_17892  ( .D(I306891), .CLK(I2702), .RSTB(I306659), .Q(I306908) );
nor I_17893 (I306925,I306908,I306761);
DFFARX1 I_17894  ( .D(I306908), .CLK(I2702), .RSTB(I306659), .Q(I306942) );
not I_17895 (I306630,I306942);
nand I_17896 (I306973,I306676,I420533);
and I_17897 (I306990,I306973,I306925);
DFFARX1 I_17898  ( .D(I306973), .CLK(I2702), .RSTB(I306659), .Q(I306627) );
DFFARX1 I_17899  ( .D(I420545), .CLK(I2702), .RSTB(I306659), .Q(I307021) );
nor I_17900 (I307038,I307021,I306744);
nand I_17901 (I306645,I306908,I307038);
nor I_17902 (I307069,I307021,I306809);
not I_17903 (I306642,I307021);
nand I_17904 (I307100,I307021,I306710);
and I_17905 (I307117,I306778,I307100);
DFFARX1 I_17906  ( .D(I307117), .CLK(I2702), .RSTB(I306659), .Q(I306621) );
DFFARX1 I_17907  ( .D(I307021), .CLK(I2702), .RSTB(I306659), .Q(I306624) );
DFFARX1 I_17908  ( .D(I420539), .CLK(I2702), .RSTB(I306659), .Q(I307162) );
not I_17909 (I307179,I307162);
nand I_17910 (I307196,I307179,I306744);
and I_17911 (I307213,I306973,I307196);
DFFARX1 I_17912  ( .D(I307213), .CLK(I2702), .RSTB(I306659), .Q(I306651) );
or I_17913 (I307244,I307179,I306990);
DFFARX1 I_17914  ( .D(I307244), .CLK(I2702), .RSTB(I306659), .Q(I306636) );
nand I_17915 (I306639,I307179,I307069);
not I_17916 (I307322,I2709);
not I_17917 (I307339,I567317);
nor I_17918 (I307356,I567326,I567308);
nand I_17919 (I307373,I307356,I567329);
nor I_17920 (I307390,I307339,I567326);
nand I_17921 (I307407,I307390,I567320);
not I_17922 (I307424,I307407);
not I_17923 (I307441,I567326);
nor I_17924 (I307311,I307407,I307441);
not I_17925 (I307472,I307441);
nand I_17926 (I307296,I307407,I307472);
not I_17927 (I307503,I567314);
nor I_17928 (I307520,I307503,I567305);
and I_17929 (I307537,I307520,I567302);
or I_17930 (I307554,I307537,I567299);
DFFARX1 I_17931  ( .D(I307554), .CLK(I2702), .RSTB(I307322), .Q(I307571) );
nor I_17932 (I307588,I307571,I307424);
DFFARX1 I_17933  ( .D(I307571), .CLK(I2702), .RSTB(I307322), .Q(I307605) );
not I_17934 (I307293,I307605);
nand I_17935 (I307636,I307339,I567314);
and I_17936 (I307653,I307636,I307588);
DFFARX1 I_17937  ( .D(I307636), .CLK(I2702), .RSTB(I307322), .Q(I307290) );
DFFARX1 I_17938  ( .D(I567323), .CLK(I2702), .RSTB(I307322), .Q(I307684) );
nor I_17939 (I307701,I307684,I307407);
nand I_17940 (I307308,I307571,I307701);
nor I_17941 (I307732,I307684,I307472);
not I_17942 (I307305,I307684);
nand I_17943 (I307763,I307684,I307373);
and I_17944 (I307780,I307441,I307763);
DFFARX1 I_17945  ( .D(I307780), .CLK(I2702), .RSTB(I307322), .Q(I307284) );
DFFARX1 I_17946  ( .D(I307684), .CLK(I2702), .RSTB(I307322), .Q(I307287) );
DFFARX1 I_17947  ( .D(I567311), .CLK(I2702), .RSTB(I307322), .Q(I307825) );
not I_17948 (I307842,I307825);
nand I_17949 (I307859,I307842,I307407);
and I_17950 (I307876,I307636,I307859);
DFFARX1 I_17951  ( .D(I307876), .CLK(I2702), .RSTB(I307322), .Q(I307314) );
or I_17952 (I307907,I307842,I307653);
DFFARX1 I_17953  ( .D(I307907), .CLK(I2702), .RSTB(I307322), .Q(I307299) );
nand I_17954 (I307302,I307842,I307732);
not I_17955 (I307985,I2709);
not I_17956 (I308002,I172035);
nor I_17957 (I308019,I172041,I172047);
nand I_17958 (I308036,I308019,I172050);
nor I_17959 (I308053,I308002,I172041);
nand I_17960 (I308070,I308053,I172032);
not I_17961 (I308087,I308070);
not I_17962 (I308104,I172041);
nor I_17963 (I307974,I308070,I308104);
not I_17964 (I308135,I308104);
nand I_17965 (I307959,I308070,I308135);
not I_17966 (I308166,I172044);
nor I_17967 (I308183,I308166,I172038);
and I_17968 (I308200,I308183,I172053);
or I_17969 (I308217,I308200,I172059);
DFFARX1 I_17970  ( .D(I308217), .CLK(I2702), .RSTB(I307985), .Q(I308234) );
nor I_17971 (I308251,I308234,I308087);
DFFARX1 I_17972  ( .D(I308234), .CLK(I2702), .RSTB(I307985), .Q(I308268) );
not I_17973 (I307956,I308268);
nand I_17974 (I308299,I308002,I172044);
and I_17975 (I308316,I308299,I308251);
DFFARX1 I_17976  ( .D(I308299), .CLK(I2702), .RSTB(I307985), .Q(I307953) );
DFFARX1 I_17977  ( .D(I172056), .CLK(I2702), .RSTB(I307985), .Q(I308347) );
nor I_17978 (I308364,I308347,I308070);
nand I_17979 (I307971,I308234,I308364);
nor I_17980 (I308395,I308347,I308135);
not I_17981 (I307968,I308347);
nand I_17982 (I308426,I308347,I308036);
and I_17983 (I308443,I308104,I308426);
DFFARX1 I_17984  ( .D(I308443), .CLK(I2702), .RSTB(I307985), .Q(I307947) );
DFFARX1 I_17985  ( .D(I308347), .CLK(I2702), .RSTB(I307985), .Q(I307950) );
DFFARX1 I_17986  ( .D(I172062), .CLK(I2702), .RSTB(I307985), .Q(I308488) );
not I_17987 (I308505,I308488);
nand I_17988 (I308522,I308505,I308070);
and I_17989 (I308539,I308299,I308522);
DFFARX1 I_17990  ( .D(I308539), .CLK(I2702), .RSTB(I307985), .Q(I307977) );
or I_17991 (I308570,I308505,I308316);
DFFARX1 I_17992  ( .D(I308570), .CLK(I2702), .RSTB(I307985), .Q(I307962) );
nand I_17993 (I307965,I308505,I308395);
not I_17994 (I308648,I2709);
not I_17995 (I308665,I373205);
nor I_17996 (I308682,I373202,I373220);
nand I_17997 (I308699,I308682,I373223);
nor I_17998 (I308716,I308665,I373202);
nand I_17999 (I308733,I308716,I373208);
not I_18000 (I308750,I308733);
not I_18001 (I308767,I373202);
nor I_18002 (I308637,I308733,I308767);
not I_18003 (I308798,I308767);
nand I_18004 (I308622,I308733,I308798);
not I_18005 (I308829,I373217);
nor I_18006 (I308846,I308829,I373199);
and I_18007 (I308863,I308846,I373193);
or I_18008 (I308880,I308863,I373211);
DFFARX1 I_18009  ( .D(I308880), .CLK(I2702), .RSTB(I308648), .Q(I308897) );
nor I_18010 (I308914,I308897,I308750);
DFFARX1 I_18011  ( .D(I308897), .CLK(I2702), .RSTB(I308648), .Q(I308931) );
not I_18012 (I308619,I308931);
nand I_18013 (I308962,I308665,I373217);
and I_18014 (I308979,I308962,I308914);
DFFARX1 I_18015  ( .D(I308962), .CLK(I2702), .RSTB(I308648), .Q(I308616) );
DFFARX1 I_18016  ( .D(I373196), .CLK(I2702), .RSTB(I308648), .Q(I309010) );
nor I_18017 (I309027,I309010,I308733);
nand I_18018 (I308634,I308897,I309027);
nor I_18019 (I309058,I309010,I308798);
not I_18020 (I308631,I309010);
nand I_18021 (I309089,I309010,I308699);
and I_18022 (I309106,I308767,I309089);
DFFARX1 I_18023  ( .D(I309106), .CLK(I2702), .RSTB(I308648), .Q(I308610) );
DFFARX1 I_18024  ( .D(I309010), .CLK(I2702), .RSTB(I308648), .Q(I308613) );
DFFARX1 I_18025  ( .D(I373214), .CLK(I2702), .RSTB(I308648), .Q(I309151) );
not I_18026 (I309168,I309151);
nand I_18027 (I309185,I309168,I308733);
and I_18028 (I309202,I308962,I309185);
DFFARX1 I_18029  ( .D(I309202), .CLK(I2702), .RSTB(I308648), .Q(I308640) );
or I_18030 (I309233,I309168,I308979);
DFFARX1 I_18031  ( .D(I309233), .CLK(I2702), .RSTB(I308648), .Q(I308625) );
nand I_18032 (I308628,I309168,I309058);
not I_18033 (I309311,I2709);
not I_18034 (I309328,I569697);
nor I_18035 (I309345,I569706,I569688);
nand I_18036 (I309362,I309345,I569709);
nor I_18037 (I309379,I309328,I569706);
nand I_18038 (I309396,I309379,I569700);
not I_18039 (I309413,I309396);
not I_18040 (I309430,I569706);
nor I_18041 (I309300,I309396,I309430);
not I_18042 (I309461,I309430);
nand I_18043 (I309285,I309396,I309461);
not I_18044 (I309492,I569694);
nor I_18045 (I309509,I309492,I569685);
and I_18046 (I309526,I309509,I569682);
or I_18047 (I309543,I309526,I569679);
DFFARX1 I_18048  ( .D(I309543), .CLK(I2702), .RSTB(I309311), .Q(I309560) );
nor I_18049 (I309577,I309560,I309413);
DFFARX1 I_18050  ( .D(I309560), .CLK(I2702), .RSTB(I309311), .Q(I309594) );
not I_18051 (I309282,I309594);
nand I_18052 (I309625,I309328,I569694);
and I_18053 (I309642,I309625,I309577);
DFFARX1 I_18054  ( .D(I309625), .CLK(I2702), .RSTB(I309311), .Q(I309279) );
DFFARX1 I_18055  ( .D(I569703), .CLK(I2702), .RSTB(I309311), .Q(I309673) );
nor I_18056 (I309690,I309673,I309396);
nand I_18057 (I309297,I309560,I309690);
nor I_18058 (I309721,I309673,I309461);
not I_18059 (I309294,I309673);
nand I_18060 (I309752,I309673,I309362);
and I_18061 (I309769,I309430,I309752);
DFFARX1 I_18062  ( .D(I309769), .CLK(I2702), .RSTB(I309311), .Q(I309273) );
DFFARX1 I_18063  ( .D(I309673), .CLK(I2702), .RSTB(I309311), .Q(I309276) );
DFFARX1 I_18064  ( .D(I569691), .CLK(I2702), .RSTB(I309311), .Q(I309814) );
not I_18065 (I309831,I309814);
nand I_18066 (I309848,I309831,I309396);
and I_18067 (I309865,I309625,I309848);
DFFARX1 I_18068  ( .D(I309865), .CLK(I2702), .RSTB(I309311), .Q(I309303) );
or I_18069 (I309896,I309831,I309642);
DFFARX1 I_18070  ( .D(I309896), .CLK(I2702), .RSTB(I309311), .Q(I309288) );
nand I_18071 (I309291,I309831,I309721);
not I_18072 (I309974,I2709);
not I_18073 (I309991,I162753);
nor I_18074 (I310008,I162759,I162765);
nand I_18075 (I310025,I310008,I162768);
nor I_18076 (I310042,I309991,I162759);
nand I_18077 (I310059,I310042,I162750);
not I_18078 (I310076,I310059);
not I_18079 (I310093,I162759);
nor I_18080 (I309963,I310059,I310093);
not I_18081 (I310124,I310093);
nand I_18082 (I309948,I310059,I310124);
not I_18083 (I310155,I162762);
nor I_18084 (I310172,I310155,I162756);
and I_18085 (I310189,I310172,I162771);
or I_18086 (I310206,I310189,I162777);
DFFARX1 I_18087  ( .D(I310206), .CLK(I2702), .RSTB(I309974), .Q(I310223) );
nor I_18088 (I310240,I310223,I310076);
DFFARX1 I_18089  ( .D(I310223), .CLK(I2702), .RSTB(I309974), .Q(I310257) );
not I_18090 (I309945,I310257);
nand I_18091 (I310288,I309991,I162762);
and I_18092 (I310305,I310288,I310240);
DFFARX1 I_18093  ( .D(I310288), .CLK(I2702), .RSTB(I309974), .Q(I309942) );
DFFARX1 I_18094  ( .D(I162774), .CLK(I2702), .RSTB(I309974), .Q(I310336) );
nor I_18095 (I310353,I310336,I310059);
nand I_18096 (I309960,I310223,I310353);
nor I_18097 (I310384,I310336,I310124);
not I_18098 (I309957,I310336);
nand I_18099 (I310415,I310336,I310025);
and I_18100 (I310432,I310093,I310415);
DFFARX1 I_18101  ( .D(I310432), .CLK(I2702), .RSTB(I309974), .Q(I309936) );
DFFARX1 I_18102  ( .D(I310336), .CLK(I2702), .RSTB(I309974), .Q(I309939) );
DFFARX1 I_18103  ( .D(I162780), .CLK(I2702), .RSTB(I309974), .Q(I310477) );
not I_18104 (I310494,I310477);
nand I_18105 (I310511,I310494,I310059);
and I_18106 (I310528,I310288,I310511);
DFFARX1 I_18107  ( .D(I310528), .CLK(I2702), .RSTB(I309974), .Q(I309966) );
or I_18108 (I310559,I310494,I310305);
DFFARX1 I_18109  ( .D(I310559), .CLK(I2702), .RSTB(I309974), .Q(I309951) );
nand I_18110 (I309954,I310494,I310384);
not I_18111 (I310637,I2709);
not I_18112 (I310654,I447158);
nor I_18113 (I310671,I447170,I447152);
nand I_18114 (I310688,I310671,I447173);
nor I_18115 (I310705,I310654,I447170);
nand I_18116 (I310722,I310705,I447164);
not I_18117 (I310739,I310722);
not I_18118 (I310756,I447170);
nor I_18119 (I310626,I310722,I310756);
not I_18120 (I310787,I310756);
nand I_18121 (I310611,I310722,I310787);
not I_18122 (I310818,I447155);
nor I_18123 (I310835,I310818,I447149);
and I_18124 (I310852,I310835,I447161);
or I_18125 (I310869,I310852,I447146);
DFFARX1 I_18126  ( .D(I310869), .CLK(I2702), .RSTB(I310637), .Q(I310886) );
nor I_18127 (I310903,I310886,I310739);
DFFARX1 I_18128  ( .D(I310886), .CLK(I2702), .RSTB(I310637), .Q(I310920) );
not I_18129 (I310608,I310920);
nand I_18130 (I310951,I310654,I447155);
and I_18131 (I310968,I310951,I310903);
DFFARX1 I_18132  ( .D(I310951), .CLK(I2702), .RSTB(I310637), .Q(I310605) );
DFFARX1 I_18133  ( .D(I447143), .CLK(I2702), .RSTB(I310637), .Q(I310999) );
nor I_18134 (I311016,I310999,I310722);
nand I_18135 (I310623,I310886,I311016);
nor I_18136 (I311047,I310999,I310787);
not I_18137 (I310620,I310999);
nand I_18138 (I311078,I310999,I310688);
and I_18139 (I311095,I310756,I311078);
DFFARX1 I_18140  ( .D(I311095), .CLK(I2702), .RSTB(I310637), .Q(I310599) );
DFFARX1 I_18141  ( .D(I310999), .CLK(I2702), .RSTB(I310637), .Q(I310602) );
DFFARX1 I_18142  ( .D(I447167), .CLK(I2702), .RSTB(I310637), .Q(I311140) );
not I_18143 (I311157,I311140);
nand I_18144 (I311174,I311157,I310722);
and I_18145 (I311191,I310951,I311174);
DFFARX1 I_18146  ( .D(I311191), .CLK(I2702), .RSTB(I310637), .Q(I310629) );
or I_18147 (I311222,I311157,I310968);
DFFARX1 I_18148  ( .D(I311222), .CLK(I2702), .RSTB(I310637), .Q(I310614) );
nand I_18149 (I310617,I311157,I311047);
not I_18150 (I311300,I2709);
not I_18151 (I311317,I675952);
nor I_18152 (I311334,I675970,I675961);
nand I_18153 (I311351,I311334,I675967);
nor I_18154 (I311368,I311317,I675970);
nand I_18155 (I311385,I311368,I675973);
not I_18156 (I311402,I311385);
not I_18157 (I311419,I675970);
nor I_18158 (I311289,I311385,I311419);
not I_18159 (I311450,I311419);
nand I_18160 (I311274,I311385,I311450);
not I_18161 (I311481,I675949);
nor I_18162 (I311498,I311481,I675964);
and I_18163 (I311515,I311498,I675946);
or I_18164 (I311532,I311515,I675955);
DFFARX1 I_18165  ( .D(I311532), .CLK(I2702), .RSTB(I311300), .Q(I311549) );
nor I_18166 (I311566,I311549,I311402);
DFFARX1 I_18167  ( .D(I311549), .CLK(I2702), .RSTB(I311300), .Q(I311583) );
not I_18168 (I311271,I311583);
nand I_18169 (I311614,I311317,I675949);
and I_18170 (I311631,I311614,I311566);
DFFARX1 I_18171  ( .D(I311614), .CLK(I2702), .RSTB(I311300), .Q(I311268) );
DFFARX1 I_18172  ( .D(I675958), .CLK(I2702), .RSTB(I311300), .Q(I311662) );
nor I_18173 (I311679,I311662,I311385);
nand I_18174 (I311286,I311549,I311679);
nor I_18175 (I311710,I311662,I311450);
not I_18176 (I311283,I311662);
nand I_18177 (I311741,I311662,I311351);
and I_18178 (I311758,I311419,I311741);
DFFARX1 I_18179  ( .D(I311758), .CLK(I2702), .RSTB(I311300), .Q(I311262) );
DFFARX1 I_18180  ( .D(I311662), .CLK(I2702), .RSTB(I311300), .Q(I311265) );
DFFARX1 I_18181  ( .D(I675976), .CLK(I2702), .RSTB(I311300), .Q(I311803) );
not I_18182 (I311820,I311803);
nand I_18183 (I311837,I311820,I311385);
and I_18184 (I311854,I311614,I311837);
DFFARX1 I_18185  ( .D(I311854), .CLK(I2702), .RSTB(I311300), .Q(I311292) );
or I_18186 (I311885,I311820,I311631);
DFFARX1 I_18187  ( .D(I311885), .CLK(I2702), .RSTB(I311300), .Q(I311277) );
nand I_18188 (I311280,I311820,I311710);
not I_18189 (I311963,I2709);
not I_18190 (I311980,I224291);
nor I_18191 (I311997,I224285,I224276);
nand I_18192 (I312014,I311997,I224288);
nor I_18193 (I312031,I311980,I224285);
nand I_18194 (I312048,I312031,I224303);
not I_18195 (I312065,I312048);
not I_18196 (I312082,I224285);
nor I_18197 (I311952,I312048,I312082);
not I_18198 (I312113,I312082);
nand I_18199 (I311937,I312048,I312113);
not I_18200 (I312144,I224279);
nor I_18201 (I312161,I312144,I224273);
and I_18202 (I312178,I312161,I224300);
or I_18203 (I312195,I312178,I224297);
DFFARX1 I_18204  ( .D(I312195), .CLK(I2702), .RSTB(I311963), .Q(I312212) );
nor I_18205 (I312229,I312212,I312065);
DFFARX1 I_18206  ( .D(I312212), .CLK(I2702), .RSTB(I311963), .Q(I312246) );
not I_18207 (I311934,I312246);
nand I_18208 (I312277,I311980,I224279);
and I_18209 (I312294,I312277,I312229);
DFFARX1 I_18210  ( .D(I312277), .CLK(I2702), .RSTB(I311963), .Q(I311931) );
DFFARX1 I_18211  ( .D(I224294), .CLK(I2702), .RSTB(I311963), .Q(I312325) );
nor I_18212 (I312342,I312325,I312048);
nand I_18213 (I311949,I312212,I312342);
nor I_18214 (I312373,I312325,I312113);
not I_18215 (I311946,I312325);
nand I_18216 (I312404,I312325,I312014);
and I_18217 (I312421,I312082,I312404);
DFFARX1 I_18218  ( .D(I312421), .CLK(I2702), .RSTB(I311963), .Q(I311925) );
DFFARX1 I_18219  ( .D(I312325), .CLK(I2702), .RSTB(I311963), .Q(I311928) );
DFFARX1 I_18220  ( .D(I224282), .CLK(I2702), .RSTB(I311963), .Q(I312466) );
not I_18221 (I312483,I312466);
nand I_18222 (I312500,I312483,I312048);
and I_18223 (I312517,I312277,I312500);
DFFARX1 I_18224  ( .D(I312517), .CLK(I2702), .RSTB(I311963), .Q(I311955) );
or I_18225 (I312548,I312483,I312294);
DFFARX1 I_18226  ( .D(I312548), .CLK(I2702), .RSTB(I311963), .Q(I311940) );
nand I_18227 (I311943,I312483,I312373);
not I_18228 (I312626,I2709);
not I_18229 (I312643,I670291);
nor I_18230 (I312660,I670309,I670300);
nand I_18231 (I312677,I312660,I670306);
nor I_18232 (I312694,I312643,I670309);
nand I_18233 (I312711,I312694,I670312);
not I_18234 (I312728,I312711);
not I_18235 (I312745,I670309);
nor I_18236 (I312615,I312711,I312745);
not I_18237 (I312776,I312745);
nand I_18238 (I312600,I312711,I312776);
not I_18239 (I312807,I670288);
nor I_18240 (I312824,I312807,I670303);
and I_18241 (I312841,I312824,I670285);
or I_18242 (I312858,I312841,I670294);
DFFARX1 I_18243  ( .D(I312858), .CLK(I2702), .RSTB(I312626), .Q(I312875) );
nor I_18244 (I312892,I312875,I312728);
DFFARX1 I_18245  ( .D(I312875), .CLK(I2702), .RSTB(I312626), .Q(I312909) );
not I_18246 (I312597,I312909);
nand I_18247 (I312940,I312643,I670288);
and I_18248 (I312957,I312940,I312892);
DFFARX1 I_18249  ( .D(I312940), .CLK(I2702), .RSTB(I312626), .Q(I312594) );
DFFARX1 I_18250  ( .D(I670297), .CLK(I2702), .RSTB(I312626), .Q(I312988) );
nor I_18251 (I313005,I312988,I312711);
nand I_18252 (I312612,I312875,I313005);
nor I_18253 (I313036,I312988,I312776);
not I_18254 (I312609,I312988);
nand I_18255 (I313067,I312988,I312677);
and I_18256 (I313084,I312745,I313067);
DFFARX1 I_18257  ( .D(I313084), .CLK(I2702), .RSTB(I312626), .Q(I312588) );
DFFARX1 I_18258  ( .D(I312988), .CLK(I2702), .RSTB(I312626), .Q(I312591) );
DFFARX1 I_18259  ( .D(I670315), .CLK(I2702), .RSTB(I312626), .Q(I313129) );
not I_18260 (I313146,I313129);
nand I_18261 (I313163,I313146,I312711);
and I_18262 (I313180,I312940,I313163);
DFFARX1 I_18263  ( .D(I313180), .CLK(I2702), .RSTB(I312626), .Q(I312618) );
or I_18264 (I313211,I313146,I312957);
DFFARX1 I_18265  ( .D(I313211), .CLK(I2702), .RSTB(I312626), .Q(I312603) );
nand I_18266 (I312606,I313146,I313036);
not I_18267 (I313289,I2709);
not I_18268 (I313306,I519717);
nor I_18269 (I313323,I519726,I519708);
nand I_18270 (I313340,I313323,I519729);
nor I_18271 (I313357,I313306,I519726);
nand I_18272 (I313374,I313357,I519720);
not I_18273 (I313391,I313374);
not I_18274 (I313408,I519726);
nor I_18275 (I313278,I313374,I313408);
not I_18276 (I313439,I313408);
nand I_18277 (I313263,I313374,I313439);
not I_18278 (I313470,I519714);
nor I_18279 (I313487,I313470,I519705);
and I_18280 (I313504,I313487,I519702);
or I_18281 (I313521,I313504,I519699);
DFFARX1 I_18282  ( .D(I313521), .CLK(I2702), .RSTB(I313289), .Q(I313538) );
nor I_18283 (I313555,I313538,I313391);
DFFARX1 I_18284  ( .D(I313538), .CLK(I2702), .RSTB(I313289), .Q(I313572) );
not I_18285 (I313260,I313572);
nand I_18286 (I313603,I313306,I519714);
and I_18287 (I313620,I313603,I313555);
DFFARX1 I_18288  ( .D(I313603), .CLK(I2702), .RSTB(I313289), .Q(I313257) );
DFFARX1 I_18289  ( .D(I519723), .CLK(I2702), .RSTB(I313289), .Q(I313651) );
nor I_18290 (I313668,I313651,I313374);
nand I_18291 (I313275,I313538,I313668);
nor I_18292 (I313699,I313651,I313439);
not I_18293 (I313272,I313651);
nand I_18294 (I313730,I313651,I313340);
and I_18295 (I313747,I313408,I313730);
DFFARX1 I_18296  ( .D(I313747), .CLK(I2702), .RSTB(I313289), .Q(I313251) );
DFFARX1 I_18297  ( .D(I313651), .CLK(I2702), .RSTB(I313289), .Q(I313254) );
DFFARX1 I_18298  ( .D(I519711), .CLK(I2702), .RSTB(I313289), .Q(I313792) );
not I_18299 (I313809,I313792);
nand I_18300 (I313826,I313809,I313374);
and I_18301 (I313843,I313603,I313826);
DFFARX1 I_18302  ( .D(I313843), .CLK(I2702), .RSTB(I313289), .Q(I313281) );
or I_18303 (I313874,I313809,I313620);
DFFARX1 I_18304  ( .D(I313874), .CLK(I2702), .RSTB(I313289), .Q(I313266) );
nand I_18305 (I313269,I313809,I313699);
not I_18306 (I313952,I2709);
not I_18307 (I313969,I699044);
nor I_18308 (I313986,I699035,I699041);
nand I_18309 (I314003,I313986,I699053);
nor I_18310 (I314020,I313969,I699035);
nand I_18311 (I314037,I314020,I699038);
not I_18312 (I314054,I314037);
not I_18313 (I314071,I699035);
nor I_18314 (I313941,I314037,I314071);
not I_18315 (I314102,I314071);
nand I_18316 (I313926,I314037,I314102);
not I_18317 (I314133,I699062);
nor I_18318 (I314150,I314133,I699056);
and I_18319 (I314167,I314150,I699047);
or I_18320 (I314184,I314167,I699032);
DFFARX1 I_18321  ( .D(I314184), .CLK(I2702), .RSTB(I313952), .Q(I314201) );
nor I_18322 (I314218,I314201,I314054);
DFFARX1 I_18323  ( .D(I314201), .CLK(I2702), .RSTB(I313952), .Q(I314235) );
not I_18324 (I313923,I314235);
nand I_18325 (I314266,I313969,I699062);
and I_18326 (I314283,I314266,I314218);
DFFARX1 I_18327  ( .D(I314266), .CLK(I2702), .RSTB(I313952), .Q(I313920) );
DFFARX1 I_18328  ( .D(I699050), .CLK(I2702), .RSTB(I313952), .Q(I314314) );
nor I_18329 (I314331,I314314,I314037);
nand I_18330 (I313938,I314201,I314331);
nor I_18331 (I314362,I314314,I314102);
not I_18332 (I313935,I314314);
nand I_18333 (I314393,I314314,I314003);
and I_18334 (I314410,I314071,I314393);
DFFARX1 I_18335  ( .D(I314410), .CLK(I2702), .RSTB(I313952), .Q(I313914) );
DFFARX1 I_18336  ( .D(I314314), .CLK(I2702), .RSTB(I313952), .Q(I313917) );
DFFARX1 I_18337  ( .D(I699059), .CLK(I2702), .RSTB(I313952), .Q(I314455) );
not I_18338 (I314472,I314455);
nand I_18339 (I314489,I314472,I314037);
and I_18340 (I314506,I314266,I314489);
DFFARX1 I_18341  ( .D(I314506), .CLK(I2702), .RSTB(I313952), .Q(I313944) );
or I_18342 (I314537,I314472,I314283);
DFFARX1 I_18343  ( .D(I314537), .CLK(I2702), .RSTB(I313952), .Q(I313929) );
nand I_18344 (I313932,I314472,I314362);
not I_18345 (I314615,I2709);
not I_18346 (I314632,I149493);
nor I_18347 (I314649,I149499,I149505);
nand I_18348 (I314666,I314649,I149508);
nor I_18349 (I314683,I314632,I149499);
nand I_18350 (I314700,I314683,I149490);
not I_18351 (I314717,I314700);
not I_18352 (I314734,I149499);
nor I_18353 (I314604,I314700,I314734);
not I_18354 (I314765,I314734);
nand I_18355 (I314589,I314700,I314765);
not I_18356 (I314796,I149502);
nor I_18357 (I314813,I314796,I149496);
and I_18358 (I314830,I314813,I149511);
or I_18359 (I314847,I314830,I149517);
DFFARX1 I_18360  ( .D(I314847), .CLK(I2702), .RSTB(I314615), .Q(I314864) );
nor I_18361 (I314881,I314864,I314717);
DFFARX1 I_18362  ( .D(I314864), .CLK(I2702), .RSTB(I314615), .Q(I314898) );
not I_18363 (I314586,I314898);
nand I_18364 (I314929,I314632,I149502);
and I_18365 (I314946,I314929,I314881);
DFFARX1 I_18366  ( .D(I314929), .CLK(I2702), .RSTB(I314615), .Q(I314583) );
DFFARX1 I_18367  ( .D(I149514), .CLK(I2702), .RSTB(I314615), .Q(I314977) );
nor I_18368 (I314994,I314977,I314700);
nand I_18369 (I314601,I314864,I314994);
nor I_18370 (I315025,I314977,I314765);
not I_18371 (I314598,I314977);
nand I_18372 (I315056,I314977,I314666);
and I_18373 (I315073,I314734,I315056);
DFFARX1 I_18374  ( .D(I315073), .CLK(I2702), .RSTB(I314615), .Q(I314577) );
DFFARX1 I_18375  ( .D(I314977), .CLK(I2702), .RSTB(I314615), .Q(I314580) );
DFFARX1 I_18376  ( .D(I149520), .CLK(I2702), .RSTB(I314615), .Q(I315118) );
not I_18377 (I315135,I315118);
nand I_18378 (I315152,I315135,I314700);
and I_18379 (I315169,I314929,I315152);
DFFARX1 I_18380  ( .D(I315169), .CLK(I2702), .RSTB(I314615), .Q(I314607) );
or I_18381 (I315200,I315135,I314946);
DFFARX1 I_18382  ( .D(I315200), .CLK(I2702), .RSTB(I314615), .Q(I314592) );
nand I_18383 (I314595,I315135,I315025);
not I_18384 (I315278,I2709);
not I_18385 (I315295,I2111);
nor I_18386 (I315312,I1823,I1311);
nand I_18387 (I315329,I315312,I2087);
nor I_18388 (I315346,I315295,I1823);
nand I_18389 (I315363,I315346,I1663);
not I_18390 (I315380,I315363);
not I_18391 (I315397,I1823);
nor I_18392 (I315267,I315363,I315397);
not I_18393 (I315428,I315397);
nand I_18394 (I315252,I315363,I315428);
not I_18395 (I315459,I2175);
nor I_18396 (I315476,I315459,I2463);
and I_18397 (I315493,I315476,I2247);
or I_18398 (I315510,I315493,I2399);
DFFARX1 I_18399  ( .D(I315510), .CLK(I2702), .RSTB(I315278), .Q(I315527) );
nor I_18400 (I315544,I315527,I315380);
DFFARX1 I_18401  ( .D(I315527), .CLK(I2702), .RSTB(I315278), .Q(I315561) );
not I_18402 (I315249,I315561);
nand I_18403 (I315592,I315295,I2175);
and I_18404 (I315609,I315592,I315544);
DFFARX1 I_18405  ( .D(I315592), .CLK(I2702), .RSTB(I315278), .Q(I315246) );
DFFARX1 I_18406  ( .D(I2583), .CLK(I2702), .RSTB(I315278), .Q(I315640) );
nor I_18407 (I315657,I315640,I315363);
nand I_18408 (I315264,I315527,I315657);
nor I_18409 (I315688,I315640,I315428);
not I_18410 (I315261,I315640);
nand I_18411 (I315719,I315640,I315329);
and I_18412 (I315736,I315397,I315719);
DFFARX1 I_18413  ( .D(I315736), .CLK(I2702), .RSTB(I315278), .Q(I315240) );
DFFARX1 I_18414  ( .D(I315640), .CLK(I2702), .RSTB(I315278), .Q(I315243) );
DFFARX1 I_18415  ( .D(I2015), .CLK(I2702), .RSTB(I315278), .Q(I315781) );
not I_18416 (I315798,I315781);
nand I_18417 (I315815,I315798,I315363);
and I_18418 (I315832,I315592,I315815);
DFFARX1 I_18419  ( .D(I315832), .CLK(I2702), .RSTB(I315278), .Q(I315270) );
or I_18420 (I315863,I315798,I315609);
DFFARX1 I_18421  ( .D(I315863), .CLK(I2702), .RSTB(I315278), .Q(I315255) );
nand I_18422 (I315258,I315798,I315688);
not I_18423 (I315941,I2709);
not I_18424 (I315958,I355763);
nor I_18425 (I315975,I355760,I355778);
nand I_18426 (I315992,I315975,I355781);
nor I_18427 (I316009,I315958,I355760);
nand I_18428 (I316026,I316009,I355766);
not I_18429 (I316043,I316026);
not I_18430 (I316060,I355760);
nor I_18431 (I315930,I316026,I316060);
not I_18432 (I316091,I316060);
nand I_18433 (I315915,I316026,I316091);
not I_18434 (I316122,I355775);
nor I_18435 (I316139,I316122,I355757);
and I_18436 (I316156,I316139,I355751);
or I_18437 (I316173,I316156,I355769);
DFFARX1 I_18438  ( .D(I316173), .CLK(I2702), .RSTB(I315941), .Q(I316190) );
nor I_18439 (I316207,I316190,I316043);
DFFARX1 I_18440  ( .D(I316190), .CLK(I2702), .RSTB(I315941), .Q(I316224) );
not I_18441 (I315912,I316224);
nand I_18442 (I316255,I315958,I355775);
and I_18443 (I316272,I316255,I316207);
DFFARX1 I_18444  ( .D(I316255), .CLK(I2702), .RSTB(I315941), .Q(I315909) );
DFFARX1 I_18445  ( .D(I355754), .CLK(I2702), .RSTB(I315941), .Q(I316303) );
nor I_18446 (I316320,I316303,I316026);
nand I_18447 (I315927,I316190,I316320);
nor I_18448 (I316351,I316303,I316091);
not I_18449 (I315924,I316303);
nand I_18450 (I316382,I316303,I315992);
and I_18451 (I316399,I316060,I316382);
DFFARX1 I_18452  ( .D(I316399), .CLK(I2702), .RSTB(I315941), .Q(I315903) );
DFFARX1 I_18453  ( .D(I316303), .CLK(I2702), .RSTB(I315941), .Q(I315906) );
DFFARX1 I_18454  ( .D(I355772), .CLK(I2702), .RSTB(I315941), .Q(I316444) );
not I_18455 (I316461,I316444);
nand I_18456 (I316478,I316461,I316026);
and I_18457 (I316495,I316255,I316478);
DFFARX1 I_18458  ( .D(I316495), .CLK(I2702), .RSTB(I315941), .Q(I315933) );
or I_18459 (I316526,I316461,I316272);
DFFARX1 I_18460  ( .D(I316526), .CLK(I2702), .RSTB(I315941), .Q(I315918) );
nand I_18461 (I315921,I316461,I316351);
not I_18462 (I316604,I2709);
not I_18463 (I316621,I217151);
nor I_18464 (I316638,I217145,I217136);
nand I_18465 (I316655,I316638,I217148);
nor I_18466 (I316672,I316621,I217145);
nand I_18467 (I316689,I316672,I217163);
not I_18468 (I316706,I316689);
not I_18469 (I316723,I217145);
nor I_18470 (I316593,I316689,I316723);
not I_18471 (I316754,I316723);
nand I_18472 (I316578,I316689,I316754);
not I_18473 (I316785,I217139);
nor I_18474 (I316802,I316785,I217133);
and I_18475 (I316819,I316802,I217160);
or I_18476 (I316836,I316819,I217157);
DFFARX1 I_18477  ( .D(I316836), .CLK(I2702), .RSTB(I316604), .Q(I316853) );
nor I_18478 (I316870,I316853,I316706);
DFFARX1 I_18479  ( .D(I316853), .CLK(I2702), .RSTB(I316604), .Q(I316887) );
not I_18480 (I316575,I316887);
nand I_18481 (I316918,I316621,I217139);
and I_18482 (I316935,I316918,I316870);
DFFARX1 I_18483  ( .D(I316918), .CLK(I2702), .RSTB(I316604), .Q(I316572) );
DFFARX1 I_18484  ( .D(I217154), .CLK(I2702), .RSTB(I316604), .Q(I316966) );
nor I_18485 (I316983,I316966,I316689);
nand I_18486 (I316590,I316853,I316983);
nor I_18487 (I317014,I316966,I316754);
not I_18488 (I316587,I316966);
nand I_18489 (I317045,I316966,I316655);
and I_18490 (I317062,I316723,I317045);
DFFARX1 I_18491  ( .D(I317062), .CLK(I2702), .RSTB(I316604), .Q(I316566) );
DFFARX1 I_18492  ( .D(I316966), .CLK(I2702), .RSTB(I316604), .Q(I316569) );
DFFARX1 I_18493  ( .D(I217142), .CLK(I2702), .RSTB(I316604), .Q(I317107) );
not I_18494 (I317124,I317107);
nand I_18495 (I317141,I317124,I316689);
and I_18496 (I317158,I316918,I317141);
DFFARX1 I_18497  ( .D(I317158), .CLK(I2702), .RSTB(I316604), .Q(I316596) );
or I_18498 (I317189,I317124,I316935);
DFFARX1 I_18499  ( .D(I317189), .CLK(I2702), .RSTB(I316604), .Q(I316581) );
nand I_18500 (I316584,I317124,I317014);
not I_18501 (I317267,I2709);
not I_18502 (I317284,I727366);
nor I_18503 (I317301,I727357,I727363);
nand I_18504 (I317318,I317301,I727375);
nor I_18505 (I317335,I317284,I727357);
nand I_18506 (I317352,I317335,I727360);
not I_18507 (I317369,I317352);
not I_18508 (I317386,I727357);
nor I_18509 (I317256,I317352,I317386);
not I_18510 (I317417,I317386);
nand I_18511 (I317241,I317352,I317417);
not I_18512 (I317448,I727384);
nor I_18513 (I317465,I317448,I727378);
and I_18514 (I317482,I317465,I727369);
or I_18515 (I317499,I317482,I727354);
DFFARX1 I_18516  ( .D(I317499), .CLK(I2702), .RSTB(I317267), .Q(I317516) );
nor I_18517 (I317533,I317516,I317369);
DFFARX1 I_18518  ( .D(I317516), .CLK(I2702), .RSTB(I317267), .Q(I317550) );
not I_18519 (I317238,I317550);
nand I_18520 (I317581,I317284,I727384);
and I_18521 (I317598,I317581,I317533);
DFFARX1 I_18522  ( .D(I317581), .CLK(I2702), .RSTB(I317267), .Q(I317235) );
DFFARX1 I_18523  ( .D(I727372), .CLK(I2702), .RSTB(I317267), .Q(I317629) );
nor I_18524 (I317646,I317629,I317352);
nand I_18525 (I317253,I317516,I317646);
nor I_18526 (I317677,I317629,I317417);
not I_18527 (I317250,I317629);
nand I_18528 (I317708,I317629,I317318);
and I_18529 (I317725,I317386,I317708);
DFFARX1 I_18530  ( .D(I317725), .CLK(I2702), .RSTB(I317267), .Q(I317229) );
DFFARX1 I_18531  ( .D(I317629), .CLK(I2702), .RSTB(I317267), .Q(I317232) );
DFFARX1 I_18532  ( .D(I727381), .CLK(I2702), .RSTB(I317267), .Q(I317770) );
not I_18533 (I317787,I317770);
nand I_18534 (I317804,I317787,I317352);
and I_18535 (I317821,I317581,I317804);
DFFARX1 I_18536  ( .D(I317821), .CLK(I2702), .RSTB(I317267), .Q(I317259) );
or I_18537 (I317852,I317787,I317598);
DFFARX1 I_18538  ( .D(I317852), .CLK(I2702), .RSTB(I317267), .Q(I317244) );
nand I_18539 (I317247,I317787,I317677);
not I_18540 (I317930,I2709);
not I_18541 (I317947,I168057);
nor I_18542 (I317964,I168063,I168069);
nand I_18543 (I317981,I317964,I168072);
nor I_18544 (I317998,I317947,I168063);
nand I_18545 (I318015,I317998,I168054);
not I_18546 (I318032,I318015);
not I_18547 (I318049,I168063);
nor I_18548 (I317919,I318015,I318049);
not I_18549 (I318080,I318049);
nand I_18550 (I317904,I318015,I318080);
not I_18551 (I318111,I168066);
nor I_18552 (I318128,I318111,I168060);
and I_18553 (I318145,I318128,I168075);
or I_18554 (I318162,I318145,I168081);
DFFARX1 I_18555  ( .D(I318162), .CLK(I2702), .RSTB(I317930), .Q(I318179) );
nor I_18556 (I318196,I318179,I318032);
DFFARX1 I_18557  ( .D(I318179), .CLK(I2702), .RSTB(I317930), .Q(I318213) );
not I_18558 (I317901,I318213);
nand I_18559 (I318244,I317947,I168066);
and I_18560 (I318261,I318244,I318196);
DFFARX1 I_18561  ( .D(I318244), .CLK(I2702), .RSTB(I317930), .Q(I317898) );
DFFARX1 I_18562  ( .D(I168078), .CLK(I2702), .RSTB(I317930), .Q(I318292) );
nor I_18563 (I318309,I318292,I318015);
nand I_18564 (I317916,I318179,I318309);
nor I_18565 (I318340,I318292,I318080);
not I_18566 (I317913,I318292);
nand I_18567 (I318371,I318292,I317981);
and I_18568 (I318388,I318049,I318371);
DFFARX1 I_18569  ( .D(I318388), .CLK(I2702), .RSTB(I317930), .Q(I317892) );
DFFARX1 I_18570  ( .D(I318292), .CLK(I2702), .RSTB(I317930), .Q(I317895) );
DFFARX1 I_18571  ( .D(I168084), .CLK(I2702), .RSTB(I317930), .Q(I318433) );
not I_18572 (I318450,I318433);
nand I_18573 (I318467,I318450,I318015);
and I_18574 (I318484,I318244,I318467);
DFFARX1 I_18575  ( .D(I318484), .CLK(I2702), .RSTB(I317930), .Q(I317922) );
or I_18576 (I318515,I318450,I318261);
DFFARX1 I_18577  ( .D(I318515), .CLK(I2702), .RSTB(I317930), .Q(I317907) );
nand I_18578 (I317910,I318450,I318340);
not I_18579 (I318593,I2709);
not I_18580 (I318610,I624374);
nor I_18581 (I318627,I624392,I624383);
nand I_18582 (I318644,I318627,I624389);
nor I_18583 (I318661,I318610,I624392);
nand I_18584 (I318678,I318661,I624395);
not I_18585 (I318695,I318678);
not I_18586 (I318712,I624392);
nor I_18587 (I318582,I318678,I318712);
not I_18588 (I318743,I318712);
nand I_18589 (I318567,I318678,I318743);
not I_18590 (I318774,I624371);
nor I_18591 (I318791,I318774,I624386);
and I_18592 (I318808,I318791,I624368);
or I_18593 (I318825,I318808,I624377);
DFFARX1 I_18594  ( .D(I318825), .CLK(I2702), .RSTB(I318593), .Q(I318842) );
nor I_18595 (I318859,I318842,I318695);
DFFARX1 I_18596  ( .D(I318842), .CLK(I2702), .RSTB(I318593), .Q(I318876) );
not I_18597 (I318564,I318876);
nand I_18598 (I318907,I318610,I624371);
and I_18599 (I318924,I318907,I318859);
DFFARX1 I_18600  ( .D(I318907), .CLK(I2702), .RSTB(I318593), .Q(I318561) );
DFFARX1 I_18601  ( .D(I624380), .CLK(I2702), .RSTB(I318593), .Q(I318955) );
nor I_18602 (I318972,I318955,I318678);
nand I_18603 (I318579,I318842,I318972);
nor I_18604 (I319003,I318955,I318743);
not I_18605 (I318576,I318955);
nand I_18606 (I319034,I318955,I318644);
and I_18607 (I319051,I318712,I319034);
DFFARX1 I_18608  ( .D(I319051), .CLK(I2702), .RSTB(I318593), .Q(I318555) );
DFFARX1 I_18609  ( .D(I318955), .CLK(I2702), .RSTB(I318593), .Q(I318558) );
DFFARX1 I_18610  ( .D(I624398), .CLK(I2702), .RSTB(I318593), .Q(I319096) );
not I_18611 (I319113,I319096);
nand I_18612 (I319130,I319113,I318678);
and I_18613 (I319147,I318907,I319130);
DFFARX1 I_18614  ( .D(I319147), .CLK(I2702), .RSTB(I318593), .Q(I318585) );
or I_18615 (I319178,I319113,I318924);
DFFARX1 I_18616  ( .D(I319178), .CLK(I2702), .RSTB(I318593), .Q(I318570) );
nand I_18617 (I318573,I319113,I319003);
not I_18618 (I319256,I2709);
not I_18619 (I319273,I231440);
nor I_18620 (I319290,I231413,I231416);
nand I_18621 (I319307,I319290,I231428);
nor I_18622 (I319324,I319273,I231413);
nand I_18623 (I319341,I319324,I231434);
not I_18624 (I319358,I319341);
not I_18625 (I319375,I231413);
nor I_18626 (I319245,I319341,I319375);
not I_18627 (I319406,I319375);
nand I_18628 (I319230,I319341,I319406);
not I_18629 (I319437,I231437);
nor I_18630 (I319454,I319437,I231419);
and I_18631 (I319471,I319454,I231422);
or I_18632 (I319488,I319471,I231443);
DFFARX1 I_18633  ( .D(I319488), .CLK(I2702), .RSTB(I319256), .Q(I319505) );
nor I_18634 (I319522,I319505,I319358);
DFFARX1 I_18635  ( .D(I319505), .CLK(I2702), .RSTB(I319256), .Q(I319539) );
not I_18636 (I319227,I319539);
nand I_18637 (I319570,I319273,I231437);
and I_18638 (I319587,I319570,I319522);
DFFARX1 I_18639  ( .D(I319570), .CLK(I2702), .RSTB(I319256), .Q(I319224) );
DFFARX1 I_18640  ( .D(I231425), .CLK(I2702), .RSTB(I319256), .Q(I319618) );
nor I_18641 (I319635,I319618,I319341);
nand I_18642 (I319242,I319505,I319635);
nor I_18643 (I319666,I319618,I319406);
not I_18644 (I319239,I319618);
nand I_18645 (I319697,I319618,I319307);
and I_18646 (I319714,I319375,I319697);
DFFARX1 I_18647  ( .D(I319714), .CLK(I2702), .RSTB(I319256), .Q(I319218) );
DFFARX1 I_18648  ( .D(I319618), .CLK(I2702), .RSTB(I319256), .Q(I319221) );
DFFARX1 I_18649  ( .D(I231431), .CLK(I2702), .RSTB(I319256), .Q(I319759) );
not I_18650 (I319776,I319759);
nand I_18651 (I319793,I319776,I319341);
and I_18652 (I319810,I319570,I319793);
DFFARX1 I_18653  ( .D(I319810), .CLK(I2702), .RSTB(I319256), .Q(I319248) );
or I_18654 (I319841,I319776,I319587);
DFFARX1 I_18655  ( .D(I319841), .CLK(I2702), .RSTB(I319256), .Q(I319233) );
nand I_18656 (I319236,I319776,I319666);
not I_18657 (I319919,I2709);
not I_18658 (I319936,I219531);
nor I_18659 (I319953,I219525,I219516);
nand I_18660 (I319970,I319953,I219528);
nor I_18661 (I319987,I319936,I219525);
nand I_18662 (I320004,I319987,I219543);
not I_18663 (I320021,I320004);
not I_18664 (I320038,I219525);
nor I_18665 (I319908,I320004,I320038);
not I_18666 (I320069,I320038);
nand I_18667 (I319893,I320004,I320069);
not I_18668 (I320100,I219519);
nor I_18669 (I320117,I320100,I219513);
and I_18670 (I320134,I320117,I219540);
or I_18671 (I320151,I320134,I219537);
DFFARX1 I_18672  ( .D(I320151), .CLK(I2702), .RSTB(I319919), .Q(I320168) );
nor I_18673 (I320185,I320168,I320021);
DFFARX1 I_18674  ( .D(I320168), .CLK(I2702), .RSTB(I319919), .Q(I320202) );
not I_18675 (I319890,I320202);
nand I_18676 (I320233,I319936,I219519);
and I_18677 (I320250,I320233,I320185);
DFFARX1 I_18678  ( .D(I320233), .CLK(I2702), .RSTB(I319919), .Q(I319887) );
DFFARX1 I_18679  ( .D(I219534), .CLK(I2702), .RSTB(I319919), .Q(I320281) );
nor I_18680 (I320298,I320281,I320004);
nand I_18681 (I319905,I320168,I320298);
nor I_18682 (I320329,I320281,I320069);
not I_18683 (I319902,I320281);
nand I_18684 (I320360,I320281,I319970);
and I_18685 (I320377,I320038,I320360);
DFFARX1 I_18686  ( .D(I320377), .CLK(I2702), .RSTB(I319919), .Q(I319881) );
DFFARX1 I_18687  ( .D(I320281), .CLK(I2702), .RSTB(I319919), .Q(I319884) );
DFFARX1 I_18688  ( .D(I219522), .CLK(I2702), .RSTB(I319919), .Q(I320422) );
not I_18689 (I320439,I320422);
nand I_18690 (I320456,I320439,I320004);
and I_18691 (I320473,I320233,I320456);
DFFARX1 I_18692  ( .D(I320473), .CLK(I2702), .RSTB(I319919), .Q(I319911) );
or I_18693 (I320504,I320439,I320250);
DFFARX1 I_18694  ( .D(I320504), .CLK(I2702), .RSTB(I319919), .Q(I319896) );
nand I_18695 (I319899,I320439,I320329);
not I_18696 (I320582,I2709);
not I_18697 (I320599,I109835);
nor I_18698 (I320616,I109832,I109856);
nand I_18699 (I320633,I320616,I109853);
nor I_18700 (I320650,I320599,I109832);
nand I_18701 (I320667,I320650,I109859);
not I_18702 (I320684,I320667);
not I_18703 (I320701,I109832);
nor I_18704 (I320571,I320667,I320701);
not I_18705 (I320732,I320701);
nand I_18706 (I320556,I320667,I320732);
not I_18707 (I320763,I109850);
nor I_18708 (I320780,I320763,I109841);
and I_18709 (I320797,I320780,I109838);
or I_18710 (I320814,I320797,I109847);
DFFARX1 I_18711  ( .D(I320814), .CLK(I2702), .RSTB(I320582), .Q(I320831) );
nor I_18712 (I320848,I320831,I320684);
DFFARX1 I_18713  ( .D(I320831), .CLK(I2702), .RSTB(I320582), .Q(I320865) );
not I_18714 (I320553,I320865);
nand I_18715 (I320896,I320599,I109850);
and I_18716 (I320913,I320896,I320848);
DFFARX1 I_18717  ( .D(I320896), .CLK(I2702), .RSTB(I320582), .Q(I320550) );
DFFARX1 I_18718  ( .D(I109829), .CLK(I2702), .RSTB(I320582), .Q(I320944) );
nor I_18719 (I320961,I320944,I320667);
nand I_18720 (I320568,I320831,I320961);
nor I_18721 (I320992,I320944,I320732);
not I_18722 (I320565,I320944);
nand I_18723 (I321023,I320944,I320633);
and I_18724 (I321040,I320701,I321023);
DFFARX1 I_18725  ( .D(I321040), .CLK(I2702), .RSTB(I320582), .Q(I320544) );
DFFARX1 I_18726  ( .D(I320944), .CLK(I2702), .RSTB(I320582), .Q(I320547) );
DFFARX1 I_18727  ( .D(I109844), .CLK(I2702), .RSTB(I320582), .Q(I321085) );
not I_18728 (I321102,I321085);
nand I_18729 (I321119,I321102,I320667);
and I_18730 (I321136,I320896,I321119);
DFFARX1 I_18731  ( .D(I321136), .CLK(I2702), .RSTB(I320582), .Q(I320574) );
or I_18732 (I321167,I321102,I320913);
DFFARX1 I_18733  ( .D(I321167), .CLK(I2702), .RSTB(I320582), .Q(I320559) );
nand I_18734 (I320562,I321102,I320992);
not I_18735 (I321245,I2709);
not I_18736 (I321262,I30219);
nor I_18737 (I321279,I30225,I30228);
nand I_18738 (I321296,I321279,I30204);
nor I_18739 (I321313,I321262,I30225);
nand I_18740 (I321330,I321313,I30213);
not I_18741 (I321347,I321330);
not I_18742 (I321364,I30225);
nor I_18743 (I321234,I321330,I321364);
not I_18744 (I321395,I321364);
nand I_18745 (I321219,I321330,I321395);
not I_18746 (I321426,I30207);
nor I_18747 (I321443,I321426,I30231);
and I_18748 (I321460,I321443,I30201);
or I_18749 (I321477,I321460,I30210);
DFFARX1 I_18750  ( .D(I321477), .CLK(I2702), .RSTB(I321245), .Q(I321494) );
nor I_18751 (I321511,I321494,I321347);
DFFARX1 I_18752  ( .D(I321494), .CLK(I2702), .RSTB(I321245), .Q(I321528) );
not I_18753 (I321216,I321528);
nand I_18754 (I321559,I321262,I30207);
and I_18755 (I321576,I321559,I321511);
DFFARX1 I_18756  ( .D(I321559), .CLK(I2702), .RSTB(I321245), .Q(I321213) );
DFFARX1 I_18757  ( .D(I30216), .CLK(I2702), .RSTB(I321245), .Q(I321607) );
nor I_18758 (I321624,I321607,I321330);
nand I_18759 (I321231,I321494,I321624);
nor I_18760 (I321655,I321607,I321395);
not I_18761 (I321228,I321607);
nand I_18762 (I321686,I321607,I321296);
and I_18763 (I321703,I321364,I321686);
DFFARX1 I_18764  ( .D(I321703), .CLK(I2702), .RSTB(I321245), .Q(I321207) );
DFFARX1 I_18765  ( .D(I321607), .CLK(I2702), .RSTB(I321245), .Q(I321210) );
DFFARX1 I_18766  ( .D(I30222), .CLK(I2702), .RSTB(I321245), .Q(I321748) );
not I_18767 (I321765,I321748);
nand I_18768 (I321782,I321765,I321330);
and I_18769 (I321799,I321559,I321782);
DFFARX1 I_18770  ( .D(I321799), .CLK(I2702), .RSTB(I321245), .Q(I321237) );
or I_18771 (I321830,I321765,I321576);
DFFARX1 I_18772  ( .D(I321830), .CLK(I2702), .RSTB(I321245), .Q(I321222) );
nand I_18773 (I321225,I321765,I321655);
not I_18774 (I321908,I2709);
not I_18775 (I321925,I398399);
nor I_18776 (I321942,I398396,I398414);
nand I_18777 (I321959,I321942,I398417);
nor I_18778 (I321976,I321925,I398396);
nand I_18779 (I321993,I321976,I398402);
not I_18780 (I322010,I321993);
not I_18781 (I322027,I398396);
nor I_18782 (I321897,I321993,I322027);
not I_18783 (I322058,I322027);
nand I_18784 (I321882,I321993,I322058);
not I_18785 (I322089,I398411);
nor I_18786 (I322106,I322089,I398393);
and I_18787 (I322123,I322106,I398387);
or I_18788 (I322140,I322123,I398405);
DFFARX1 I_18789  ( .D(I322140), .CLK(I2702), .RSTB(I321908), .Q(I322157) );
nor I_18790 (I322174,I322157,I322010);
DFFARX1 I_18791  ( .D(I322157), .CLK(I2702), .RSTB(I321908), .Q(I322191) );
not I_18792 (I321879,I322191);
nand I_18793 (I322222,I321925,I398411);
and I_18794 (I322239,I322222,I322174);
DFFARX1 I_18795  ( .D(I322222), .CLK(I2702), .RSTB(I321908), .Q(I321876) );
DFFARX1 I_18796  ( .D(I398390), .CLK(I2702), .RSTB(I321908), .Q(I322270) );
nor I_18797 (I322287,I322270,I321993);
nand I_18798 (I321894,I322157,I322287);
nor I_18799 (I322318,I322270,I322058);
not I_18800 (I321891,I322270);
nand I_18801 (I322349,I322270,I321959);
and I_18802 (I322366,I322027,I322349);
DFFARX1 I_18803  ( .D(I322366), .CLK(I2702), .RSTB(I321908), .Q(I321870) );
DFFARX1 I_18804  ( .D(I322270), .CLK(I2702), .RSTB(I321908), .Q(I321873) );
DFFARX1 I_18805  ( .D(I398408), .CLK(I2702), .RSTB(I321908), .Q(I322411) );
not I_18806 (I322428,I322411);
nand I_18807 (I322445,I322428,I321993);
and I_18808 (I322462,I322222,I322445);
DFFARX1 I_18809  ( .D(I322462), .CLK(I2702), .RSTB(I321908), .Q(I321900) );
or I_18810 (I322493,I322428,I322239);
DFFARX1 I_18811  ( .D(I322493), .CLK(I2702), .RSTB(I321908), .Q(I321885) );
nand I_18812 (I321888,I322428,I322318);
not I_18813 (I322571,I2709);
not I_18814 (I322588,I229060);
nor I_18815 (I322605,I229033,I229036);
nand I_18816 (I322622,I322605,I229048);
nor I_18817 (I322639,I322588,I229033);
nand I_18818 (I322656,I322639,I229054);
not I_18819 (I322673,I322656);
not I_18820 (I322690,I229033);
nor I_18821 (I322560,I322656,I322690);
not I_18822 (I322721,I322690);
nand I_18823 (I322545,I322656,I322721);
not I_18824 (I322752,I229057);
nor I_18825 (I322769,I322752,I229039);
and I_18826 (I322786,I322769,I229042);
or I_18827 (I322803,I322786,I229063);
DFFARX1 I_18828  ( .D(I322803), .CLK(I2702), .RSTB(I322571), .Q(I322820) );
nor I_18829 (I322837,I322820,I322673);
DFFARX1 I_18830  ( .D(I322820), .CLK(I2702), .RSTB(I322571), .Q(I322854) );
not I_18831 (I322542,I322854);
nand I_18832 (I322885,I322588,I229057);
and I_18833 (I322902,I322885,I322837);
DFFARX1 I_18834  ( .D(I322885), .CLK(I2702), .RSTB(I322571), .Q(I322539) );
DFFARX1 I_18835  ( .D(I229045), .CLK(I2702), .RSTB(I322571), .Q(I322933) );
nor I_18836 (I322950,I322933,I322656);
nand I_18837 (I322557,I322820,I322950);
nor I_18838 (I322981,I322933,I322721);
not I_18839 (I322554,I322933);
nand I_18840 (I323012,I322933,I322622);
and I_18841 (I323029,I322690,I323012);
DFFARX1 I_18842  ( .D(I323029), .CLK(I2702), .RSTB(I322571), .Q(I322533) );
DFFARX1 I_18843  ( .D(I322933), .CLK(I2702), .RSTB(I322571), .Q(I322536) );
DFFARX1 I_18844  ( .D(I229051), .CLK(I2702), .RSTB(I322571), .Q(I323074) );
not I_18845 (I323091,I323074);
nand I_18846 (I323108,I323091,I322656);
and I_18847 (I323125,I322885,I323108);
DFFARX1 I_18848  ( .D(I323125), .CLK(I2702), .RSTB(I322571), .Q(I322563) );
or I_18849 (I323156,I323091,I322902);
DFFARX1 I_18850  ( .D(I323156), .CLK(I2702), .RSTB(I322571), .Q(I322548) );
nand I_18851 (I322551,I323091,I322981);
not I_18852 (I323234,I2709);
not I_18853 (I323251,I582787);
nor I_18854 (I323268,I582784,I582775);
nand I_18855 (I323285,I323268,I582778);
nor I_18856 (I323302,I323251,I582784);
nand I_18857 (I323319,I323302,I582772);
not I_18858 (I323336,I323319);
not I_18859 (I323353,I582784);
nor I_18860 (I323223,I323319,I323353);
not I_18861 (I323384,I323353);
nand I_18862 (I323208,I323319,I323384);
not I_18863 (I323415,I582793);
nor I_18864 (I323432,I323415,I582796);
and I_18865 (I323449,I323432,I582781);
or I_18866 (I323466,I323449,I582769);
DFFARX1 I_18867  ( .D(I323466), .CLK(I2702), .RSTB(I323234), .Q(I323483) );
nor I_18868 (I323500,I323483,I323336);
DFFARX1 I_18869  ( .D(I323483), .CLK(I2702), .RSTB(I323234), .Q(I323517) );
not I_18870 (I323205,I323517);
nand I_18871 (I323548,I323251,I582793);
and I_18872 (I323565,I323548,I323500);
DFFARX1 I_18873  ( .D(I323548), .CLK(I2702), .RSTB(I323234), .Q(I323202) );
DFFARX1 I_18874  ( .D(I582790), .CLK(I2702), .RSTB(I323234), .Q(I323596) );
nor I_18875 (I323613,I323596,I323319);
nand I_18876 (I323220,I323483,I323613);
nor I_18877 (I323644,I323596,I323384);
not I_18878 (I323217,I323596);
nand I_18879 (I323675,I323596,I323285);
and I_18880 (I323692,I323353,I323675);
DFFARX1 I_18881  ( .D(I323692), .CLK(I2702), .RSTB(I323234), .Q(I323196) );
DFFARX1 I_18882  ( .D(I323596), .CLK(I2702), .RSTB(I323234), .Q(I323199) );
DFFARX1 I_18883  ( .D(I582799), .CLK(I2702), .RSTB(I323234), .Q(I323737) );
not I_18884 (I323754,I323737);
nand I_18885 (I323771,I323754,I323319);
and I_18886 (I323788,I323548,I323771);
DFFARX1 I_18887  ( .D(I323788), .CLK(I2702), .RSTB(I323234), .Q(I323226) );
or I_18888 (I323819,I323754,I323565);
DFFARX1 I_18889  ( .D(I323819), .CLK(I2702), .RSTB(I323234), .Q(I323211) );
nand I_18890 (I323214,I323754,I323644);
not I_18891 (I323897,I2709);
not I_18892 (I323914,I208821);
nor I_18893 (I323931,I208815,I208806);
nand I_18894 (I323948,I323931,I208818);
nor I_18895 (I323965,I323914,I208815);
nand I_18896 (I323982,I323965,I208833);
not I_18897 (I323999,I323982);
not I_18898 (I324016,I208815);
nor I_18899 (I323886,I323982,I324016);
not I_18900 (I324047,I324016);
nand I_18901 (I323871,I323982,I324047);
not I_18902 (I324078,I208809);
nor I_18903 (I324095,I324078,I208803);
and I_18904 (I324112,I324095,I208830);
or I_18905 (I324129,I324112,I208827);
DFFARX1 I_18906  ( .D(I324129), .CLK(I2702), .RSTB(I323897), .Q(I324146) );
nor I_18907 (I324163,I324146,I323999);
DFFARX1 I_18908  ( .D(I324146), .CLK(I2702), .RSTB(I323897), .Q(I324180) );
not I_18909 (I323868,I324180);
nand I_18910 (I324211,I323914,I208809);
and I_18911 (I324228,I324211,I324163);
DFFARX1 I_18912  ( .D(I324211), .CLK(I2702), .RSTB(I323897), .Q(I323865) );
DFFARX1 I_18913  ( .D(I208824), .CLK(I2702), .RSTB(I323897), .Q(I324259) );
nor I_18914 (I324276,I324259,I323982);
nand I_18915 (I323883,I324146,I324276);
nor I_18916 (I324307,I324259,I324047);
not I_18917 (I323880,I324259);
nand I_18918 (I324338,I324259,I323948);
and I_18919 (I324355,I324016,I324338);
DFFARX1 I_18920  ( .D(I324355), .CLK(I2702), .RSTB(I323897), .Q(I323859) );
DFFARX1 I_18921  ( .D(I324259), .CLK(I2702), .RSTB(I323897), .Q(I323862) );
DFFARX1 I_18922  ( .D(I208812), .CLK(I2702), .RSTB(I323897), .Q(I324400) );
not I_18923 (I324417,I324400);
nand I_18924 (I324434,I324417,I323982);
and I_18925 (I324451,I324211,I324434);
DFFARX1 I_18926  ( .D(I324451), .CLK(I2702), .RSTB(I323897), .Q(I323889) );
or I_18927 (I324482,I324417,I324228);
DFFARX1 I_18928  ( .D(I324482), .CLK(I2702), .RSTB(I323897), .Q(I323874) );
nand I_18929 (I323877,I324417,I324307);
not I_18930 (I324560,I2709);
not I_18931 (I324577,I54925);
nor I_18932 (I324594,I54922,I54946);
nand I_18933 (I324611,I324594,I54943);
nor I_18934 (I324628,I324577,I54922);
nand I_18935 (I324645,I324628,I54949);
not I_18936 (I324662,I324645);
not I_18937 (I324679,I54922);
nor I_18938 (I324549,I324645,I324679);
not I_18939 (I324710,I324679);
nand I_18940 (I324534,I324645,I324710);
not I_18941 (I324741,I54940);
nor I_18942 (I324758,I324741,I54931);
and I_18943 (I324775,I324758,I54928);
or I_18944 (I324792,I324775,I54937);
DFFARX1 I_18945  ( .D(I324792), .CLK(I2702), .RSTB(I324560), .Q(I324809) );
nor I_18946 (I324826,I324809,I324662);
DFFARX1 I_18947  ( .D(I324809), .CLK(I2702), .RSTB(I324560), .Q(I324843) );
not I_18948 (I324531,I324843);
nand I_18949 (I324874,I324577,I54940);
and I_18950 (I324891,I324874,I324826);
DFFARX1 I_18951  ( .D(I324874), .CLK(I2702), .RSTB(I324560), .Q(I324528) );
DFFARX1 I_18952  ( .D(I54919), .CLK(I2702), .RSTB(I324560), .Q(I324922) );
nor I_18953 (I324939,I324922,I324645);
nand I_18954 (I324546,I324809,I324939);
nor I_18955 (I324970,I324922,I324710);
not I_18956 (I324543,I324922);
nand I_18957 (I325001,I324922,I324611);
and I_18958 (I325018,I324679,I325001);
DFFARX1 I_18959  ( .D(I325018), .CLK(I2702), .RSTB(I324560), .Q(I324522) );
DFFARX1 I_18960  ( .D(I324922), .CLK(I2702), .RSTB(I324560), .Q(I324525) );
DFFARX1 I_18961  ( .D(I54934), .CLK(I2702), .RSTB(I324560), .Q(I325063) );
not I_18962 (I325080,I325063);
nand I_18963 (I325097,I325080,I324645);
and I_18964 (I325114,I324874,I325097);
DFFARX1 I_18965  ( .D(I325114), .CLK(I2702), .RSTB(I324560), .Q(I324552) );
or I_18966 (I325145,I325080,I324891);
DFFARX1 I_18967  ( .D(I325145), .CLK(I2702), .RSTB(I324560), .Q(I324537) );
nand I_18968 (I324540,I325080,I324970);
not I_18969 (I325223,I2709);
not I_18970 (I325240,I133091);
nor I_18971 (I325257,I133088,I133112);
nand I_18972 (I325274,I325257,I133109);
nor I_18973 (I325291,I325240,I133088);
nand I_18974 (I325308,I325291,I133115);
not I_18975 (I325325,I325308);
not I_18976 (I325342,I133088);
nor I_18977 (I325212,I325308,I325342);
not I_18978 (I325373,I325342);
nand I_18979 (I325197,I325308,I325373);
not I_18980 (I325404,I133106);
nor I_18981 (I325421,I325404,I133097);
and I_18982 (I325438,I325421,I133094);
or I_18983 (I325455,I325438,I133103);
DFFARX1 I_18984  ( .D(I325455), .CLK(I2702), .RSTB(I325223), .Q(I325472) );
nor I_18985 (I325489,I325472,I325325);
DFFARX1 I_18986  ( .D(I325472), .CLK(I2702), .RSTB(I325223), .Q(I325506) );
not I_18987 (I325194,I325506);
nand I_18988 (I325537,I325240,I133106);
and I_18989 (I325554,I325537,I325489);
DFFARX1 I_18990  ( .D(I325537), .CLK(I2702), .RSTB(I325223), .Q(I325191) );
DFFARX1 I_18991  ( .D(I133085), .CLK(I2702), .RSTB(I325223), .Q(I325585) );
nor I_18992 (I325602,I325585,I325308);
nand I_18993 (I325209,I325472,I325602);
nor I_18994 (I325633,I325585,I325373);
not I_18995 (I325206,I325585);
nand I_18996 (I325664,I325585,I325274);
and I_18997 (I325681,I325342,I325664);
DFFARX1 I_18998  ( .D(I325681), .CLK(I2702), .RSTB(I325223), .Q(I325185) );
DFFARX1 I_18999  ( .D(I325585), .CLK(I2702), .RSTB(I325223), .Q(I325188) );
DFFARX1 I_19000  ( .D(I133100), .CLK(I2702), .RSTB(I325223), .Q(I325726) );
not I_19001 (I325743,I325726);
nand I_19002 (I325760,I325743,I325308);
and I_19003 (I325777,I325537,I325760);
DFFARX1 I_19004  ( .D(I325777), .CLK(I2702), .RSTB(I325223), .Q(I325215) );
or I_19005 (I325808,I325743,I325554);
DFFARX1 I_19006  ( .D(I325808), .CLK(I2702), .RSTB(I325223), .Q(I325200) );
nand I_19007 (I325203,I325743,I325633);
not I_19008 (I325886,I2709);
not I_19009 (I325903,I220126);
nor I_19010 (I325920,I220120,I220111);
nand I_19011 (I325937,I325920,I220123);
nor I_19012 (I325954,I325903,I220120);
nand I_19013 (I325971,I325954,I220138);
not I_19014 (I325988,I325971);
not I_19015 (I326005,I220120);
nor I_19016 (I325875,I325971,I326005);
not I_19017 (I326036,I326005);
nand I_19018 (I325860,I325971,I326036);
not I_19019 (I326067,I220114);
nor I_19020 (I326084,I326067,I220108);
and I_19021 (I326101,I326084,I220135);
or I_19022 (I326118,I326101,I220132);
DFFARX1 I_19023  ( .D(I326118), .CLK(I2702), .RSTB(I325886), .Q(I326135) );
nor I_19024 (I326152,I326135,I325988);
DFFARX1 I_19025  ( .D(I326135), .CLK(I2702), .RSTB(I325886), .Q(I326169) );
not I_19026 (I325857,I326169);
nand I_19027 (I326200,I325903,I220114);
and I_19028 (I326217,I326200,I326152);
DFFARX1 I_19029  ( .D(I326200), .CLK(I2702), .RSTB(I325886), .Q(I325854) );
DFFARX1 I_19030  ( .D(I220129), .CLK(I2702), .RSTB(I325886), .Q(I326248) );
nor I_19031 (I326265,I326248,I325971);
nand I_19032 (I325872,I326135,I326265);
nor I_19033 (I326296,I326248,I326036);
not I_19034 (I325869,I326248);
nand I_19035 (I326327,I326248,I325937);
and I_19036 (I326344,I326005,I326327);
DFFARX1 I_19037  ( .D(I326344), .CLK(I2702), .RSTB(I325886), .Q(I325848) );
DFFARX1 I_19038  ( .D(I326248), .CLK(I2702), .RSTB(I325886), .Q(I325851) );
DFFARX1 I_19039  ( .D(I220117), .CLK(I2702), .RSTB(I325886), .Q(I326389) );
not I_19040 (I326406,I326389);
nand I_19041 (I326423,I326406,I325971);
and I_19042 (I326440,I326200,I326423);
DFFARX1 I_19043  ( .D(I326440), .CLK(I2702), .RSTB(I325886), .Q(I325878) );
or I_19044 (I326471,I326406,I326217);
DFFARX1 I_19045  ( .D(I326471), .CLK(I2702), .RSTB(I325886), .Q(I325863) );
nand I_19046 (I325866,I326406,I326296);
not I_19047 (I326549,I2709);
not I_19048 (I326566,I2527);
nor I_19049 (I326583,I1743,I2671);
nand I_19050 (I326600,I326583,I1759);
nor I_19051 (I326617,I326566,I1743);
nand I_19052 (I326634,I326617,I2343);
not I_19053 (I326651,I326634);
not I_19054 (I326668,I1743);
nor I_19055 (I326538,I326634,I326668);
not I_19056 (I326699,I326668);
nand I_19057 (I326523,I326634,I326699);
not I_19058 (I326730,I2519);
nor I_19059 (I326747,I326730,I2367);
and I_19060 (I326764,I326747,I1943);
or I_19061 (I326781,I326764,I2023);
DFFARX1 I_19062  ( .D(I326781), .CLK(I2702), .RSTB(I326549), .Q(I326798) );
nor I_19063 (I326815,I326798,I326651);
DFFARX1 I_19064  ( .D(I326798), .CLK(I2702), .RSTB(I326549), .Q(I326832) );
not I_19065 (I326520,I326832);
nand I_19066 (I326863,I326566,I2519);
and I_19067 (I326880,I326863,I326815);
DFFARX1 I_19068  ( .D(I326863), .CLK(I2702), .RSTB(I326549), .Q(I326517) );
DFFARX1 I_19069  ( .D(I2647), .CLK(I2702), .RSTB(I326549), .Q(I326911) );
nor I_19070 (I326928,I326911,I326634);
nand I_19071 (I326535,I326798,I326928);
nor I_19072 (I326959,I326911,I326699);
not I_19073 (I326532,I326911);
nand I_19074 (I326990,I326911,I326600);
and I_19075 (I327007,I326668,I326990);
DFFARX1 I_19076  ( .D(I327007), .CLK(I2702), .RSTB(I326549), .Q(I326511) );
DFFARX1 I_19077  ( .D(I326911), .CLK(I2702), .RSTB(I326549), .Q(I326514) );
DFFARX1 I_19078  ( .D(I2479), .CLK(I2702), .RSTB(I326549), .Q(I327052) );
not I_19079 (I327069,I327052);
nand I_19080 (I327086,I327069,I326634);
and I_19081 (I327103,I326863,I327086);
DFFARX1 I_19082  ( .D(I327103), .CLK(I2702), .RSTB(I326549), .Q(I326541) );
or I_19083 (I327134,I327069,I326880);
DFFARX1 I_19084  ( .D(I327134), .CLK(I2702), .RSTB(I326549), .Q(I326526) );
nand I_19085 (I326529,I327069,I326959);
not I_19086 (I327212,I2709);
not I_19087 (I327229,I633809);
nor I_19088 (I327246,I633827,I633818);
nand I_19089 (I327263,I327246,I633824);
nor I_19090 (I327280,I327229,I633827);
nand I_19091 (I327297,I327280,I633830);
not I_19092 (I327314,I327297);
not I_19093 (I327331,I633827);
nor I_19094 (I327201,I327297,I327331);
not I_19095 (I327362,I327331);
nand I_19096 (I327186,I327297,I327362);
not I_19097 (I327393,I633806);
nor I_19098 (I327410,I327393,I633821);
and I_19099 (I327427,I327410,I633803);
or I_19100 (I327444,I327427,I633812);
DFFARX1 I_19101  ( .D(I327444), .CLK(I2702), .RSTB(I327212), .Q(I327461) );
nor I_19102 (I327478,I327461,I327314);
DFFARX1 I_19103  ( .D(I327461), .CLK(I2702), .RSTB(I327212), .Q(I327495) );
not I_19104 (I327183,I327495);
nand I_19105 (I327526,I327229,I633806);
and I_19106 (I327543,I327526,I327478);
DFFARX1 I_19107  ( .D(I327526), .CLK(I2702), .RSTB(I327212), .Q(I327180) );
DFFARX1 I_19108  ( .D(I633815), .CLK(I2702), .RSTB(I327212), .Q(I327574) );
nor I_19109 (I327591,I327574,I327297);
nand I_19110 (I327198,I327461,I327591);
nor I_19111 (I327622,I327574,I327362);
not I_19112 (I327195,I327574);
nand I_19113 (I327653,I327574,I327263);
and I_19114 (I327670,I327331,I327653);
DFFARX1 I_19115  ( .D(I327670), .CLK(I2702), .RSTB(I327212), .Q(I327174) );
DFFARX1 I_19116  ( .D(I327574), .CLK(I2702), .RSTB(I327212), .Q(I327177) );
DFFARX1 I_19117  ( .D(I633833), .CLK(I2702), .RSTB(I327212), .Q(I327715) );
not I_19118 (I327732,I327715);
nand I_19119 (I327749,I327732,I327297);
and I_19120 (I327766,I327526,I327749);
DFFARX1 I_19121  ( .D(I327766), .CLK(I2702), .RSTB(I327212), .Q(I327204) );
or I_19122 (I327797,I327732,I327543);
DFFARX1 I_19123  ( .D(I327797), .CLK(I2702), .RSTB(I327212), .Q(I327189) );
nand I_19124 (I327192,I327732,I327622);
not I_19125 (I327875,I2709);
not I_19126 (I327892,I626261);
nor I_19127 (I327909,I626279,I626270);
nand I_19128 (I327926,I327909,I626276);
nor I_19129 (I327943,I327892,I626279);
nand I_19130 (I327960,I327943,I626282);
not I_19131 (I327977,I327960);
not I_19132 (I327994,I626279);
nor I_19133 (I327864,I327960,I327994);
not I_19134 (I328025,I327994);
nand I_19135 (I327849,I327960,I328025);
not I_19136 (I328056,I626258);
nor I_19137 (I328073,I328056,I626273);
and I_19138 (I328090,I328073,I626255);
or I_19139 (I328107,I328090,I626264);
DFFARX1 I_19140  ( .D(I328107), .CLK(I2702), .RSTB(I327875), .Q(I328124) );
nor I_19141 (I328141,I328124,I327977);
DFFARX1 I_19142  ( .D(I328124), .CLK(I2702), .RSTB(I327875), .Q(I328158) );
not I_19143 (I327846,I328158);
nand I_19144 (I328189,I327892,I626258);
and I_19145 (I328206,I328189,I328141);
DFFARX1 I_19146  ( .D(I328189), .CLK(I2702), .RSTB(I327875), .Q(I327843) );
DFFARX1 I_19147  ( .D(I626267), .CLK(I2702), .RSTB(I327875), .Q(I328237) );
nor I_19148 (I328254,I328237,I327960);
nand I_19149 (I327861,I328124,I328254);
nor I_19150 (I328285,I328237,I328025);
not I_19151 (I327858,I328237);
nand I_19152 (I328316,I328237,I327926);
and I_19153 (I328333,I327994,I328316);
DFFARX1 I_19154  ( .D(I328333), .CLK(I2702), .RSTB(I327875), .Q(I327837) );
DFFARX1 I_19155  ( .D(I328237), .CLK(I2702), .RSTB(I327875), .Q(I327840) );
DFFARX1 I_19156  ( .D(I626285), .CLK(I2702), .RSTB(I327875), .Q(I328378) );
not I_19157 (I328395,I328378);
nand I_19158 (I328412,I328395,I327960);
and I_19159 (I328429,I328189,I328412);
DFFARX1 I_19160  ( .D(I328429), .CLK(I2702), .RSTB(I327875), .Q(I327867) );
or I_19161 (I328460,I328395,I328206);
DFFARX1 I_19162  ( .D(I328460), .CLK(I2702), .RSTB(I327875), .Q(I327852) );
nand I_19163 (I327855,I328395,I328285);
not I_19164 (I328538,I2709);
not I_19165 (I328555,I482994);
nor I_19166 (I328572,I483006,I482988);
nand I_19167 (I328589,I328572,I483009);
nor I_19168 (I328606,I328555,I483006);
nand I_19169 (I328623,I328606,I483000);
not I_19170 (I328640,I328623);
not I_19171 (I328657,I483006);
nor I_19172 (I328527,I328623,I328657);
not I_19173 (I328688,I328657);
nand I_19174 (I328512,I328623,I328688);
not I_19175 (I328719,I482991);
nor I_19176 (I328736,I328719,I482985);
and I_19177 (I328753,I328736,I482997);
or I_19178 (I328770,I328753,I482982);
DFFARX1 I_19179  ( .D(I328770), .CLK(I2702), .RSTB(I328538), .Q(I328787) );
nor I_19180 (I328804,I328787,I328640);
DFFARX1 I_19181  ( .D(I328787), .CLK(I2702), .RSTB(I328538), .Q(I328821) );
not I_19182 (I328509,I328821);
nand I_19183 (I328852,I328555,I482991);
and I_19184 (I328869,I328852,I328804);
DFFARX1 I_19185  ( .D(I328852), .CLK(I2702), .RSTB(I328538), .Q(I328506) );
DFFARX1 I_19186  ( .D(I482979), .CLK(I2702), .RSTB(I328538), .Q(I328900) );
nor I_19187 (I328917,I328900,I328623);
nand I_19188 (I328524,I328787,I328917);
nor I_19189 (I328948,I328900,I328688);
not I_19190 (I328521,I328900);
nand I_19191 (I328979,I328900,I328589);
and I_19192 (I328996,I328657,I328979);
DFFARX1 I_19193  ( .D(I328996), .CLK(I2702), .RSTB(I328538), .Q(I328500) );
DFFARX1 I_19194  ( .D(I328900), .CLK(I2702), .RSTB(I328538), .Q(I328503) );
DFFARX1 I_19195  ( .D(I483003), .CLK(I2702), .RSTB(I328538), .Q(I329041) );
not I_19196 (I329058,I329041);
nand I_19197 (I329075,I329058,I328623);
and I_19198 (I329092,I328852,I329075);
DFFARX1 I_19199  ( .D(I329092), .CLK(I2702), .RSTB(I328538), .Q(I328530) );
or I_19200 (I329123,I329058,I328869);
DFFARX1 I_19201  ( .D(I329123), .CLK(I2702), .RSTB(I328538), .Q(I328515) );
nand I_19202 (I328518,I329058,I328948);
not I_19203 (I329201,I2709);
not I_19204 (I329218,I479526);
nor I_19205 (I329235,I479538,I479520);
nand I_19206 (I329252,I329235,I479541);
nor I_19207 (I329269,I329218,I479538);
nand I_19208 (I329286,I329269,I479532);
not I_19209 (I329303,I329286);
not I_19210 (I329320,I479538);
nor I_19211 (I329190,I329286,I329320);
not I_19212 (I329351,I329320);
nand I_19213 (I329175,I329286,I329351);
not I_19214 (I329382,I479523);
nor I_19215 (I329399,I329382,I479517);
and I_19216 (I329416,I329399,I479529);
or I_19217 (I329433,I329416,I479514);
DFFARX1 I_19218  ( .D(I329433), .CLK(I2702), .RSTB(I329201), .Q(I329450) );
nor I_19219 (I329467,I329450,I329303);
DFFARX1 I_19220  ( .D(I329450), .CLK(I2702), .RSTB(I329201), .Q(I329484) );
not I_19221 (I329172,I329484);
nand I_19222 (I329515,I329218,I479523);
and I_19223 (I329532,I329515,I329467);
DFFARX1 I_19224  ( .D(I329515), .CLK(I2702), .RSTB(I329201), .Q(I329169) );
DFFARX1 I_19225  ( .D(I479511), .CLK(I2702), .RSTB(I329201), .Q(I329563) );
nor I_19226 (I329580,I329563,I329286);
nand I_19227 (I329187,I329450,I329580);
nor I_19228 (I329611,I329563,I329351);
not I_19229 (I329184,I329563);
nand I_19230 (I329642,I329563,I329252);
and I_19231 (I329659,I329320,I329642);
DFFARX1 I_19232  ( .D(I329659), .CLK(I2702), .RSTB(I329201), .Q(I329163) );
DFFARX1 I_19233  ( .D(I329563), .CLK(I2702), .RSTB(I329201), .Q(I329166) );
DFFARX1 I_19234  ( .D(I479535), .CLK(I2702), .RSTB(I329201), .Q(I329704) );
not I_19235 (I329721,I329704);
nand I_19236 (I329738,I329721,I329286);
and I_19237 (I329755,I329515,I329738);
DFFARX1 I_19238  ( .D(I329755), .CLK(I2702), .RSTB(I329201), .Q(I329193) );
or I_19239 (I329786,I329721,I329532);
DFFARX1 I_19240  ( .D(I329786), .CLK(I2702), .RSTB(I329201), .Q(I329178) );
nand I_19241 (I329181,I329721,I329611);
not I_19242 (I329864,I2709);
not I_19243 (I329881,I375789);
nor I_19244 (I329898,I375786,I375804);
nand I_19245 (I329915,I329898,I375807);
nor I_19246 (I329932,I329881,I375786);
nand I_19247 (I329949,I329932,I375792);
not I_19248 (I329966,I329949);
not I_19249 (I329983,I375786);
nor I_19250 (I329853,I329949,I329983);
not I_19251 (I330014,I329983);
nand I_19252 (I329838,I329949,I330014);
not I_19253 (I330045,I375801);
nor I_19254 (I330062,I330045,I375783);
and I_19255 (I330079,I330062,I375777);
or I_19256 (I330096,I330079,I375795);
DFFARX1 I_19257  ( .D(I330096), .CLK(I2702), .RSTB(I329864), .Q(I330113) );
nor I_19258 (I330130,I330113,I329966);
DFFARX1 I_19259  ( .D(I330113), .CLK(I2702), .RSTB(I329864), .Q(I330147) );
not I_19260 (I329835,I330147);
nand I_19261 (I330178,I329881,I375801);
and I_19262 (I330195,I330178,I330130);
DFFARX1 I_19263  ( .D(I330178), .CLK(I2702), .RSTB(I329864), .Q(I329832) );
DFFARX1 I_19264  ( .D(I375780), .CLK(I2702), .RSTB(I329864), .Q(I330226) );
nor I_19265 (I330243,I330226,I329949);
nand I_19266 (I329850,I330113,I330243);
nor I_19267 (I330274,I330226,I330014);
not I_19268 (I329847,I330226);
nand I_19269 (I330305,I330226,I329915);
and I_19270 (I330322,I329983,I330305);
DFFARX1 I_19271  ( .D(I330322), .CLK(I2702), .RSTB(I329864), .Q(I329826) );
DFFARX1 I_19272  ( .D(I330226), .CLK(I2702), .RSTB(I329864), .Q(I329829) );
DFFARX1 I_19273  ( .D(I375798), .CLK(I2702), .RSTB(I329864), .Q(I330367) );
not I_19274 (I330384,I330367);
nand I_19275 (I330401,I330384,I329949);
and I_19276 (I330418,I330178,I330401);
DFFARX1 I_19277  ( .D(I330418), .CLK(I2702), .RSTB(I329864), .Q(I329856) );
or I_19278 (I330449,I330384,I330195);
DFFARX1 I_19279  ( .D(I330449), .CLK(I2702), .RSTB(I329864), .Q(I329841) );
nand I_19280 (I329844,I330384,I330274);
not I_19281 (I330527,I2709);
not I_19282 (I330544,I178665);
nor I_19283 (I330561,I178671,I178677);
nand I_19284 (I330578,I330561,I178680);
nor I_19285 (I330595,I330544,I178671);
nand I_19286 (I330612,I330595,I178662);
not I_19287 (I330629,I330612);
not I_19288 (I330646,I178671);
nor I_19289 (I330516,I330612,I330646);
not I_19290 (I330677,I330646);
nand I_19291 (I330501,I330612,I330677);
not I_19292 (I330708,I178674);
nor I_19293 (I330725,I330708,I178668);
and I_19294 (I330742,I330725,I178683);
or I_19295 (I330759,I330742,I178689);
DFFARX1 I_19296  ( .D(I330759), .CLK(I2702), .RSTB(I330527), .Q(I330776) );
nor I_19297 (I330793,I330776,I330629);
DFFARX1 I_19298  ( .D(I330776), .CLK(I2702), .RSTB(I330527), .Q(I330810) );
not I_19299 (I330498,I330810);
nand I_19300 (I330841,I330544,I178674);
and I_19301 (I330858,I330841,I330793);
DFFARX1 I_19302  ( .D(I330841), .CLK(I2702), .RSTB(I330527), .Q(I330495) );
DFFARX1 I_19303  ( .D(I178686), .CLK(I2702), .RSTB(I330527), .Q(I330889) );
nor I_19304 (I330906,I330889,I330612);
nand I_19305 (I330513,I330776,I330906);
nor I_19306 (I330937,I330889,I330677);
not I_19307 (I330510,I330889);
nand I_19308 (I330968,I330889,I330578);
and I_19309 (I330985,I330646,I330968);
DFFARX1 I_19310  ( .D(I330985), .CLK(I2702), .RSTB(I330527), .Q(I330489) );
DFFARX1 I_19311  ( .D(I330889), .CLK(I2702), .RSTB(I330527), .Q(I330492) );
DFFARX1 I_19312  ( .D(I178692), .CLK(I2702), .RSTB(I330527), .Q(I331030) );
not I_19313 (I331047,I331030);
nand I_19314 (I331064,I331047,I330612);
and I_19315 (I331081,I330841,I331064);
DFFARX1 I_19316  ( .D(I331081), .CLK(I2702), .RSTB(I330527), .Q(I330519) );
or I_19317 (I331112,I331047,I330858);
DFFARX1 I_19318  ( .D(I331112), .CLK(I2702), .RSTB(I330527), .Q(I330504) );
nand I_19319 (I330507,I331047,I330937);
not I_19320 (I331190,I2709);
not I_19321 (I331207,I477792);
nor I_19322 (I331224,I477804,I477786);
nand I_19323 (I331241,I331224,I477807);
nor I_19324 (I331258,I331207,I477804);
nand I_19325 (I331275,I331258,I477798);
not I_19326 (I331292,I331275);
not I_19327 (I331309,I477804);
nor I_19328 (I331179,I331275,I331309);
not I_19329 (I331340,I331309);
nand I_19330 (I331164,I331275,I331340);
not I_19331 (I331371,I477789);
nor I_19332 (I331388,I331371,I477783);
and I_19333 (I331405,I331388,I477795);
or I_19334 (I331422,I331405,I477780);
DFFARX1 I_19335  ( .D(I331422), .CLK(I2702), .RSTB(I331190), .Q(I331439) );
nor I_19336 (I331456,I331439,I331292);
DFFARX1 I_19337  ( .D(I331439), .CLK(I2702), .RSTB(I331190), .Q(I331473) );
not I_19338 (I331161,I331473);
nand I_19339 (I331504,I331207,I477789);
and I_19340 (I331521,I331504,I331456);
DFFARX1 I_19341  ( .D(I331504), .CLK(I2702), .RSTB(I331190), .Q(I331158) );
DFFARX1 I_19342  ( .D(I477777), .CLK(I2702), .RSTB(I331190), .Q(I331552) );
nor I_19343 (I331569,I331552,I331275);
nand I_19344 (I331176,I331439,I331569);
nor I_19345 (I331600,I331552,I331340);
not I_19346 (I331173,I331552);
nand I_19347 (I331631,I331552,I331241);
and I_19348 (I331648,I331309,I331631);
DFFARX1 I_19349  ( .D(I331648), .CLK(I2702), .RSTB(I331190), .Q(I331152) );
DFFARX1 I_19350  ( .D(I331552), .CLK(I2702), .RSTB(I331190), .Q(I331155) );
DFFARX1 I_19351  ( .D(I477801), .CLK(I2702), .RSTB(I331190), .Q(I331693) );
not I_19352 (I331710,I331693);
nand I_19353 (I331727,I331710,I331275);
and I_19354 (I331744,I331504,I331727);
DFFARX1 I_19355  ( .D(I331744), .CLK(I2702), .RSTB(I331190), .Q(I331182) );
or I_19356 (I331775,I331710,I331521);
DFFARX1 I_19357  ( .D(I331775), .CLK(I2702), .RSTB(I331190), .Q(I331167) );
nand I_19358 (I331170,I331710,I331600);
not I_19359 (I331853,I2709);
not I_19360 (I331870,I488267);
nor I_19361 (I331887,I488264,I488261);
nand I_19362 (I331904,I331887,I488249);
nor I_19363 (I331921,I331870,I488264);
nand I_19364 (I331938,I331921,I488270);
not I_19365 (I331955,I331938);
not I_19366 (I331972,I488264);
nor I_19367 (I331842,I331938,I331972);
not I_19368 (I332003,I331972);
nand I_19369 (I331827,I331938,I332003);
not I_19370 (I332034,I488252);
nor I_19371 (I332051,I332034,I488258);
and I_19372 (I332068,I332051,I488255);
or I_19373 (I332085,I332068,I488279);
DFFARX1 I_19374  ( .D(I332085), .CLK(I2702), .RSTB(I331853), .Q(I332102) );
nor I_19375 (I332119,I332102,I331955);
DFFARX1 I_19376  ( .D(I332102), .CLK(I2702), .RSTB(I331853), .Q(I332136) );
not I_19377 (I331824,I332136);
nand I_19378 (I332167,I331870,I488252);
and I_19379 (I332184,I332167,I332119);
DFFARX1 I_19380  ( .D(I332167), .CLK(I2702), .RSTB(I331853), .Q(I331821) );
DFFARX1 I_19381  ( .D(I488276), .CLK(I2702), .RSTB(I331853), .Q(I332215) );
nor I_19382 (I332232,I332215,I331938);
nand I_19383 (I331839,I332102,I332232);
nor I_19384 (I332263,I332215,I332003);
not I_19385 (I331836,I332215);
nand I_19386 (I332294,I332215,I331904);
and I_19387 (I332311,I331972,I332294);
DFFARX1 I_19388  ( .D(I332311), .CLK(I2702), .RSTB(I331853), .Q(I331815) );
DFFARX1 I_19389  ( .D(I332215), .CLK(I2702), .RSTB(I331853), .Q(I331818) );
DFFARX1 I_19390  ( .D(I488273), .CLK(I2702), .RSTB(I331853), .Q(I332356) );
not I_19391 (I332373,I332356);
nand I_19392 (I332390,I332373,I331938);
and I_19393 (I332407,I332167,I332390);
DFFARX1 I_19394  ( .D(I332407), .CLK(I2702), .RSTB(I331853), .Q(I331845) );
or I_19395 (I332438,I332373,I332184);
DFFARX1 I_19396  ( .D(I332438), .CLK(I2702), .RSTB(I331853), .Q(I331830) );
nand I_19397 (I331833,I332373,I332263);
not I_19398 (I332516,I2709);
not I_19399 (I332533,I207036);
nor I_19400 (I332550,I207030,I207021);
nand I_19401 (I332567,I332550,I207033);
nor I_19402 (I332584,I332533,I207030);
nand I_19403 (I332601,I332584,I207048);
not I_19404 (I332618,I332601);
not I_19405 (I332635,I207030);
nor I_19406 (I332505,I332601,I332635);
not I_19407 (I332666,I332635);
nand I_19408 (I332490,I332601,I332666);
not I_19409 (I332697,I207024);
nor I_19410 (I332714,I332697,I207018);
and I_19411 (I332731,I332714,I207045);
or I_19412 (I332748,I332731,I207042);
DFFARX1 I_19413  ( .D(I332748), .CLK(I2702), .RSTB(I332516), .Q(I332765) );
nor I_19414 (I332782,I332765,I332618);
DFFARX1 I_19415  ( .D(I332765), .CLK(I2702), .RSTB(I332516), .Q(I332799) );
not I_19416 (I332487,I332799);
nand I_19417 (I332830,I332533,I207024);
and I_19418 (I332847,I332830,I332782);
DFFARX1 I_19419  ( .D(I332830), .CLK(I2702), .RSTB(I332516), .Q(I332484) );
DFFARX1 I_19420  ( .D(I207039), .CLK(I2702), .RSTB(I332516), .Q(I332878) );
nor I_19421 (I332895,I332878,I332601);
nand I_19422 (I332502,I332765,I332895);
nor I_19423 (I332926,I332878,I332666);
not I_19424 (I332499,I332878);
nand I_19425 (I332957,I332878,I332567);
and I_19426 (I332974,I332635,I332957);
DFFARX1 I_19427  ( .D(I332974), .CLK(I2702), .RSTB(I332516), .Q(I332478) );
DFFARX1 I_19428  ( .D(I332878), .CLK(I2702), .RSTB(I332516), .Q(I332481) );
DFFARX1 I_19429  ( .D(I207027), .CLK(I2702), .RSTB(I332516), .Q(I333019) );
not I_19430 (I333036,I333019);
nand I_19431 (I333053,I333036,I332601);
and I_19432 (I333070,I332830,I333053);
DFFARX1 I_19433  ( .D(I333070), .CLK(I2702), .RSTB(I332516), .Q(I332508) );
or I_19434 (I333101,I333036,I332847);
DFFARX1 I_19435  ( .D(I333101), .CLK(I2702), .RSTB(I332516), .Q(I332493) );
nand I_19436 (I332496,I333036,I332926);
not I_19437 (I333179,I2709);
not I_19438 (I333196,I89178);
nor I_19439 (I333213,I89169,I89160);
nand I_19440 (I333230,I333213,I89175);
nor I_19441 (I333247,I333196,I89169);
nand I_19442 (I333264,I333247,I89172);
DFFARX1 I_19443  ( .D(I333264), .CLK(I2702), .RSTB(I333179), .Q(I333281) );
not I_19444 (I333150,I333281);
not I_19445 (I333312,I89169);
not I_19446 (I333329,I333312);
not I_19447 (I333346,I89181);
nor I_19448 (I333363,I333346,I89166);
and I_19449 (I333380,I333363,I89184);
or I_19450 (I333397,I333380,I89157);
DFFARX1 I_19451  ( .D(I333397), .CLK(I2702), .RSTB(I333179), .Q(I333414) );
DFFARX1 I_19452  ( .D(I333414), .CLK(I2702), .RSTB(I333179), .Q(I333147) );
DFFARX1 I_19453  ( .D(I333414), .CLK(I2702), .RSTB(I333179), .Q(I333445) );
DFFARX1 I_19454  ( .D(I333414), .CLK(I2702), .RSTB(I333179), .Q(I333141) );
nand I_19455 (I333476,I333196,I89181);
nand I_19456 (I333493,I333476,I333230);
and I_19457 (I333510,I333312,I333493);
DFFARX1 I_19458  ( .D(I333510), .CLK(I2702), .RSTB(I333179), .Q(I333171) );
and I_19459 (I333144,I333476,I333445);
DFFARX1 I_19460  ( .D(I89187), .CLK(I2702), .RSTB(I333179), .Q(I333555) );
nor I_19461 (I333168,I333555,I333476);
nor I_19462 (I333586,I333555,I333230);
nand I_19463 (I333165,I333264,I333586);
not I_19464 (I333162,I333555);
DFFARX1 I_19465  ( .D(I89163), .CLK(I2702), .RSTB(I333179), .Q(I333631) );
not I_19466 (I333648,I333631);
nor I_19467 (I333665,I333648,I333329);
and I_19468 (I333682,I333555,I333665);
or I_19469 (I333699,I333476,I333682);
DFFARX1 I_19470  ( .D(I333699), .CLK(I2702), .RSTB(I333179), .Q(I333156) );
not I_19471 (I333730,I333648);
nor I_19472 (I333747,I333555,I333730);
nand I_19473 (I333159,I333648,I333747);
nand I_19474 (I333153,I333312,I333730);
not I_19475 (I333825,I2709);
not I_19476 (I333842,I160764);
nor I_19477 (I333859,I160785,I160767);
nand I_19478 (I333876,I333859,I160791);
nor I_19479 (I333893,I333842,I160785);
nand I_19480 (I333910,I333893,I160788);
DFFARX1 I_19481  ( .D(I333910), .CLK(I2702), .RSTB(I333825), .Q(I333927) );
not I_19482 (I333796,I333927);
not I_19483 (I333958,I160785);
not I_19484 (I333975,I333958);
not I_19485 (I333992,I160782);
nor I_19486 (I334009,I333992,I160761);
and I_19487 (I334026,I334009,I160773);
or I_19488 (I334043,I334026,I160770);
DFFARX1 I_19489  ( .D(I334043), .CLK(I2702), .RSTB(I333825), .Q(I334060) );
DFFARX1 I_19490  ( .D(I334060), .CLK(I2702), .RSTB(I333825), .Q(I333793) );
DFFARX1 I_19491  ( .D(I334060), .CLK(I2702), .RSTB(I333825), .Q(I334091) );
DFFARX1 I_19492  ( .D(I334060), .CLK(I2702), .RSTB(I333825), .Q(I333787) );
nand I_19493 (I334122,I333842,I160782);
nand I_19494 (I334139,I334122,I333876);
and I_19495 (I334156,I333958,I334139);
DFFARX1 I_19496  ( .D(I334156), .CLK(I2702), .RSTB(I333825), .Q(I333817) );
and I_19497 (I333790,I334122,I334091);
DFFARX1 I_19498  ( .D(I160776), .CLK(I2702), .RSTB(I333825), .Q(I334201) );
nor I_19499 (I333814,I334201,I334122);
nor I_19500 (I334232,I334201,I333876);
nand I_19501 (I333811,I333910,I334232);
not I_19502 (I333808,I334201);
DFFARX1 I_19503  ( .D(I160779), .CLK(I2702), .RSTB(I333825), .Q(I334277) );
not I_19504 (I334294,I334277);
nor I_19505 (I334311,I334294,I333975);
and I_19506 (I334328,I334201,I334311);
or I_19507 (I334345,I334122,I334328);
DFFARX1 I_19508  ( .D(I334345), .CLK(I2702), .RSTB(I333825), .Q(I333802) );
not I_19509 (I334376,I334294);
nor I_19510 (I334393,I334201,I334376);
nand I_19511 (I333805,I334294,I334393);
nand I_19512 (I333799,I333958,I334376);
not I_19513 (I334471,I2709);
not I_19514 (I334488,I313275);
nor I_19515 (I334505,I313254,I313266);
nand I_19516 (I334522,I334505,I313269);
nor I_19517 (I334539,I334488,I313254);
nand I_19518 (I334556,I334539,I313251);
DFFARX1 I_19519  ( .D(I334556), .CLK(I2702), .RSTB(I334471), .Q(I334573) );
not I_19520 (I334442,I334573);
not I_19521 (I334604,I313254);
not I_19522 (I334621,I334604);
not I_19523 (I334638,I313272);
nor I_19524 (I334655,I334638,I313263);
and I_19525 (I334672,I334655,I313257);
or I_19526 (I334689,I334672,I313281);
DFFARX1 I_19527  ( .D(I334689), .CLK(I2702), .RSTB(I334471), .Q(I334706) );
DFFARX1 I_19528  ( .D(I334706), .CLK(I2702), .RSTB(I334471), .Q(I334439) );
DFFARX1 I_19529  ( .D(I334706), .CLK(I2702), .RSTB(I334471), .Q(I334737) );
DFFARX1 I_19530  ( .D(I334706), .CLK(I2702), .RSTB(I334471), .Q(I334433) );
nand I_19531 (I334768,I334488,I313272);
nand I_19532 (I334785,I334768,I334522);
and I_19533 (I334802,I334604,I334785);
DFFARX1 I_19534  ( .D(I334802), .CLK(I2702), .RSTB(I334471), .Q(I334463) );
and I_19535 (I334436,I334768,I334737);
DFFARX1 I_19536  ( .D(I313278), .CLK(I2702), .RSTB(I334471), .Q(I334847) );
nor I_19537 (I334460,I334847,I334768);
nor I_19538 (I334878,I334847,I334522);
nand I_19539 (I334457,I334556,I334878);
not I_19540 (I334454,I334847);
DFFARX1 I_19541  ( .D(I313260), .CLK(I2702), .RSTB(I334471), .Q(I334923) );
not I_19542 (I334940,I334923);
nor I_19543 (I334957,I334940,I334621);
and I_19544 (I334974,I334847,I334957);
or I_19545 (I334991,I334768,I334974);
DFFARX1 I_19546  ( .D(I334991), .CLK(I2702), .RSTB(I334471), .Q(I334448) );
not I_19547 (I335022,I334940);
nor I_19548 (I335039,I334847,I335022);
nand I_19549 (I334451,I334940,I335039);
nand I_19550 (I334445,I334604,I335022);
not I_19551 (I335117,I2709);
not I_19552 (I335134,I272832);
nor I_19553 (I335151,I272811,I272823);
nand I_19554 (I335168,I335151,I272826);
nor I_19555 (I335185,I335134,I272811);
nand I_19556 (I335202,I335185,I272808);
DFFARX1 I_19557  ( .D(I335202), .CLK(I2702), .RSTB(I335117), .Q(I335219) );
not I_19558 (I335088,I335219);
not I_19559 (I335250,I272811);
not I_19560 (I335267,I335250);
not I_19561 (I335284,I272829);
nor I_19562 (I335301,I335284,I272820);
and I_19563 (I335318,I335301,I272814);
or I_19564 (I335335,I335318,I272838);
DFFARX1 I_19565  ( .D(I335335), .CLK(I2702), .RSTB(I335117), .Q(I335352) );
DFFARX1 I_19566  ( .D(I335352), .CLK(I2702), .RSTB(I335117), .Q(I335085) );
DFFARX1 I_19567  ( .D(I335352), .CLK(I2702), .RSTB(I335117), .Q(I335383) );
DFFARX1 I_19568  ( .D(I335352), .CLK(I2702), .RSTB(I335117), .Q(I335079) );
nand I_19569 (I335414,I335134,I272829);
nand I_19570 (I335431,I335414,I335168);
and I_19571 (I335448,I335250,I335431);
DFFARX1 I_19572  ( .D(I335448), .CLK(I2702), .RSTB(I335117), .Q(I335109) );
and I_19573 (I335082,I335414,I335383);
DFFARX1 I_19574  ( .D(I272835), .CLK(I2702), .RSTB(I335117), .Q(I335493) );
nor I_19575 (I335106,I335493,I335414);
nor I_19576 (I335524,I335493,I335168);
nand I_19577 (I335103,I335202,I335524);
not I_19578 (I335100,I335493);
DFFARX1 I_19579  ( .D(I272817), .CLK(I2702), .RSTB(I335117), .Q(I335569) );
not I_19580 (I335586,I335569);
nor I_19581 (I335603,I335586,I335267);
and I_19582 (I335620,I335493,I335603);
or I_19583 (I335637,I335414,I335620);
DFFARX1 I_19584  ( .D(I335637), .CLK(I2702), .RSTB(I335117), .Q(I335094) );
not I_19585 (I335668,I335586);
nor I_19586 (I335685,I335493,I335668);
nand I_19587 (I335097,I335586,I335685);
nand I_19588 (I335091,I335250,I335668);
not I_19589 (I335763,I2709);
not I_19590 (I335780,I636340);
nor I_19591 (I335797,I636337,I636322);
nand I_19592 (I335814,I335797,I636331);
nor I_19593 (I335831,I335780,I636337);
nand I_19594 (I335848,I335831,I636346);
DFFARX1 I_19595  ( .D(I335848), .CLK(I2702), .RSTB(I335763), .Q(I335865) );
not I_19596 (I335734,I335865);
not I_19597 (I335896,I636337);
not I_19598 (I335913,I335896);
not I_19599 (I335930,I636319);
nor I_19600 (I335947,I335930,I636325);
and I_19601 (I335964,I335947,I636349);
or I_19602 (I335981,I335964,I636343);
DFFARX1 I_19603  ( .D(I335981), .CLK(I2702), .RSTB(I335763), .Q(I335998) );
DFFARX1 I_19604  ( .D(I335998), .CLK(I2702), .RSTB(I335763), .Q(I335731) );
DFFARX1 I_19605  ( .D(I335998), .CLK(I2702), .RSTB(I335763), .Q(I336029) );
DFFARX1 I_19606  ( .D(I335998), .CLK(I2702), .RSTB(I335763), .Q(I335725) );
nand I_19607 (I336060,I335780,I636319);
nand I_19608 (I336077,I336060,I335814);
and I_19609 (I336094,I335896,I336077);
DFFARX1 I_19610  ( .D(I336094), .CLK(I2702), .RSTB(I335763), .Q(I335755) );
and I_19611 (I335728,I336060,I336029);
DFFARX1 I_19612  ( .D(I636328), .CLK(I2702), .RSTB(I335763), .Q(I336139) );
nor I_19613 (I335752,I336139,I336060);
nor I_19614 (I336170,I336139,I335814);
nand I_19615 (I335749,I335848,I336170);
not I_19616 (I335746,I336139);
DFFARX1 I_19617  ( .D(I636334), .CLK(I2702), .RSTB(I335763), .Q(I336215) );
not I_19618 (I336232,I336215);
nor I_19619 (I336249,I336232,I335913);
and I_19620 (I336266,I336139,I336249);
or I_19621 (I336283,I336060,I336266);
DFFARX1 I_19622  ( .D(I336283), .CLK(I2702), .RSTB(I335763), .Q(I335740) );
not I_19623 (I336314,I336232);
nor I_19624 (I336331,I336139,I336314);
nand I_19625 (I335743,I336232,I336331);
nand I_19626 (I335737,I335896,I336314);
not I_19627 (I336409,I2709);
not I_19628 (I336426,I1967);
nor I_19629 (I336443,I1431,I1655);
nand I_19630 (I336460,I336443,I1543);
nor I_19631 (I336477,I336426,I1431);
nand I_19632 (I336494,I336477,I2663);
DFFARX1 I_19633  ( .D(I336494), .CLK(I2702), .RSTB(I336409), .Q(I336511) );
not I_19634 (I336380,I336511);
not I_19635 (I336542,I1431);
not I_19636 (I336559,I336542);
not I_19637 (I336576,I1215);
nor I_19638 (I336593,I336576,I1719);
and I_19639 (I336610,I336593,I1623);
or I_19640 (I336627,I336610,I2575);
DFFARX1 I_19641  ( .D(I336627), .CLK(I2702), .RSTB(I336409), .Q(I336644) );
DFFARX1 I_19642  ( .D(I336644), .CLK(I2702), .RSTB(I336409), .Q(I336377) );
DFFARX1 I_19643  ( .D(I336644), .CLK(I2702), .RSTB(I336409), .Q(I336675) );
DFFARX1 I_19644  ( .D(I336644), .CLK(I2702), .RSTB(I336409), .Q(I336371) );
nand I_19645 (I336706,I336426,I1215);
nand I_19646 (I336723,I336706,I336460);
and I_19647 (I336740,I336542,I336723);
DFFARX1 I_19648  ( .D(I336740), .CLK(I2702), .RSTB(I336409), .Q(I336401) );
and I_19649 (I336374,I336706,I336675);
DFFARX1 I_19650  ( .D(I1927), .CLK(I2702), .RSTB(I336409), .Q(I336785) );
nor I_19651 (I336398,I336785,I336706);
nor I_19652 (I336816,I336785,I336460);
nand I_19653 (I336395,I336494,I336816);
not I_19654 (I336392,I336785);
DFFARX1 I_19655  ( .D(I1935), .CLK(I2702), .RSTB(I336409), .Q(I336861) );
not I_19656 (I336878,I336861);
nor I_19657 (I336895,I336878,I336559);
and I_19658 (I336912,I336785,I336895);
or I_19659 (I336929,I336706,I336912);
DFFARX1 I_19660  ( .D(I336929), .CLK(I2702), .RSTB(I336409), .Q(I336386) );
not I_19661 (I336960,I336878);
nor I_19662 (I336977,I336785,I336960);
nand I_19663 (I336389,I336878,I336977);
nand I_19664 (I336383,I336542,I336960);
not I_19665 (I337055,I2709);
not I_19666 (I337072,I87886);
nor I_19667 (I337089,I87877,I87868);
nand I_19668 (I337106,I337089,I87883);
nor I_19669 (I337123,I337072,I87877);
nand I_19670 (I337140,I337123,I87880);
DFFARX1 I_19671  ( .D(I337140), .CLK(I2702), .RSTB(I337055), .Q(I337157) );
not I_19672 (I337026,I337157);
not I_19673 (I337188,I87877);
not I_19674 (I337205,I337188);
not I_19675 (I337222,I87889);
nor I_19676 (I337239,I337222,I87874);
and I_19677 (I337256,I337239,I87892);
or I_19678 (I337273,I337256,I87865);
DFFARX1 I_19679  ( .D(I337273), .CLK(I2702), .RSTB(I337055), .Q(I337290) );
DFFARX1 I_19680  ( .D(I337290), .CLK(I2702), .RSTB(I337055), .Q(I337023) );
DFFARX1 I_19681  ( .D(I337290), .CLK(I2702), .RSTB(I337055), .Q(I337321) );
DFFARX1 I_19682  ( .D(I337290), .CLK(I2702), .RSTB(I337055), .Q(I337017) );
nand I_19683 (I337352,I337072,I87889);
nand I_19684 (I337369,I337352,I337106);
and I_19685 (I337386,I337188,I337369);
DFFARX1 I_19686  ( .D(I337386), .CLK(I2702), .RSTB(I337055), .Q(I337047) );
and I_19687 (I337020,I337352,I337321);
DFFARX1 I_19688  ( .D(I87895), .CLK(I2702), .RSTB(I337055), .Q(I337431) );
nor I_19689 (I337044,I337431,I337352);
nor I_19690 (I337462,I337431,I337106);
nand I_19691 (I337041,I337140,I337462);
not I_19692 (I337038,I337431);
DFFARX1 I_19693  ( .D(I87871), .CLK(I2702), .RSTB(I337055), .Q(I337507) );
not I_19694 (I337524,I337507);
nor I_19695 (I337541,I337524,I337205);
and I_19696 (I337558,I337431,I337541);
or I_19697 (I337575,I337352,I337558);
DFFARX1 I_19698  ( .D(I337575), .CLK(I2702), .RSTB(I337055), .Q(I337032) );
not I_19699 (I337606,I337524);
nor I_19700 (I337623,I337431,I337606);
nand I_19701 (I337035,I337524,I337623);
nand I_19702 (I337029,I337188,I337606);
not I_19703 (I337701,I2709);
not I_19704 (I337718,I17307);
nor I_19705 (I337735,I17322,I17316);
nand I_19706 (I337752,I337735,I17325);
nor I_19707 (I337769,I337718,I17322);
nand I_19708 (I337786,I337769,I17301);
DFFARX1 I_19709  ( .D(I337786), .CLK(I2702), .RSTB(I337701), .Q(I337803) );
not I_19710 (I337672,I337803);
not I_19711 (I337834,I17322);
not I_19712 (I337851,I337834);
not I_19713 (I337868,I17298);
nor I_19714 (I337885,I337868,I17313);
and I_19715 (I337902,I337885,I17319);
or I_19716 (I337919,I337902,I17328);
DFFARX1 I_19717  ( .D(I337919), .CLK(I2702), .RSTB(I337701), .Q(I337936) );
DFFARX1 I_19718  ( .D(I337936), .CLK(I2702), .RSTB(I337701), .Q(I337669) );
DFFARX1 I_19719  ( .D(I337936), .CLK(I2702), .RSTB(I337701), .Q(I337967) );
DFFARX1 I_19720  ( .D(I337936), .CLK(I2702), .RSTB(I337701), .Q(I337663) );
nand I_19721 (I337998,I337718,I17298);
nand I_19722 (I338015,I337998,I337752);
and I_19723 (I338032,I337834,I338015);
DFFARX1 I_19724  ( .D(I338032), .CLK(I2702), .RSTB(I337701), .Q(I337693) );
and I_19725 (I337666,I337998,I337967);
DFFARX1 I_19726  ( .D(I17310), .CLK(I2702), .RSTB(I337701), .Q(I338077) );
nor I_19727 (I337690,I338077,I337998);
nor I_19728 (I338108,I338077,I337752);
nand I_19729 (I337687,I337786,I338108);
not I_19730 (I337684,I338077);
DFFARX1 I_19731  ( .D(I17304), .CLK(I2702), .RSTB(I337701), .Q(I338153) );
not I_19732 (I338170,I338153);
nor I_19733 (I338187,I338170,I337851);
and I_19734 (I338204,I338077,I338187);
or I_19735 (I338221,I337998,I338204);
DFFARX1 I_19736  ( .D(I338221), .CLK(I2702), .RSTB(I337701), .Q(I337678) );
not I_19737 (I338252,I338170);
nor I_19738 (I338269,I338077,I338252);
nand I_19739 (I337681,I338170,I338269);
nand I_19740 (I337675,I337834,I338252);
not I_19741 (I338347,I2709);
not I_19742 (I338364,I561358);
nor I_19743 (I338381,I561370,I561364);
nand I_19744 (I338398,I338381,I561349);
nor I_19745 (I338415,I338364,I561370);
nand I_19746 (I338432,I338415,I561376);
DFFARX1 I_19747  ( .D(I338432), .CLK(I2702), .RSTB(I338347), .Q(I338449) );
not I_19748 (I338318,I338449);
not I_19749 (I338480,I561370);
not I_19750 (I338497,I338480);
not I_19751 (I338514,I561373);
nor I_19752 (I338531,I338514,I561355);
and I_19753 (I338548,I338531,I561352);
or I_19754 (I338565,I338548,I561379);
DFFARX1 I_19755  ( .D(I338565), .CLK(I2702), .RSTB(I338347), .Q(I338582) );
DFFARX1 I_19756  ( .D(I338582), .CLK(I2702), .RSTB(I338347), .Q(I338315) );
DFFARX1 I_19757  ( .D(I338582), .CLK(I2702), .RSTB(I338347), .Q(I338613) );
DFFARX1 I_19758  ( .D(I338582), .CLK(I2702), .RSTB(I338347), .Q(I338309) );
nand I_19759 (I338644,I338364,I561373);
nand I_19760 (I338661,I338644,I338398);
and I_19761 (I338678,I338480,I338661);
DFFARX1 I_19762  ( .D(I338678), .CLK(I2702), .RSTB(I338347), .Q(I338339) );
and I_19763 (I338312,I338644,I338613);
DFFARX1 I_19764  ( .D(I561367), .CLK(I2702), .RSTB(I338347), .Q(I338723) );
nor I_19765 (I338336,I338723,I338644);
nor I_19766 (I338754,I338723,I338398);
nand I_19767 (I338333,I338432,I338754);
not I_19768 (I338330,I338723);
DFFARX1 I_19769  ( .D(I561361), .CLK(I2702), .RSTB(I338347), .Q(I338799) );
not I_19770 (I338816,I338799);
nor I_19771 (I338833,I338816,I338497);
and I_19772 (I338850,I338723,I338833);
or I_19773 (I338867,I338644,I338850);
DFFARX1 I_19774  ( .D(I338867), .CLK(I2702), .RSTB(I338347), .Q(I338324) );
not I_19775 (I338898,I338816);
nor I_19776 (I338915,I338723,I338898);
nand I_19777 (I338327,I338816,I338915);
nand I_19778 (I338321,I338480,I338898);
not I_19779 (I338993,I2709);
not I_19780 (I339010,I13380);
nor I_19781 (I339027,I13395,I13389);
nand I_19782 (I339044,I339027,I13398);
nor I_19783 (I339061,I339010,I13395);
nand I_19784 (I339078,I339061,I13374);
DFFARX1 I_19785  ( .D(I339078), .CLK(I2702), .RSTB(I338993), .Q(I339095) );
not I_19786 (I338964,I339095);
not I_19787 (I339126,I13395);
not I_19788 (I339143,I339126);
not I_19789 (I339160,I13371);
nor I_19790 (I339177,I339160,I13386);
and I_19791 (I339194,I339177,I13392);
or I_19792 (I339211,I339194,I13401);
DFFARX1 I_19793  ( .D(I339211), .CLK(I2702), .RSTB(I338993), .Q(I339228) );
DFFARX1 I_19794  ( .D(I339228), .CLK(I2702), .RSTB(I338993), .Q(I338961) );
DFFARX1 I_19795  ( .D(I339228), .CLK(I2702), .RSTB(I338993), .Q(I339259) );
DFFARX1 I_19796  ( .D(I339228), .CLK(I2702), .RSTB(I338993), .Q(I338955) );
nand I_19797 (I339290,I339010,I13371);
nand I_19798 (I339307,I339290,I339044);
and I_19799 (I339324,I339126,I339307);
DFFARX1 I_19800  ( .D(I339324), .CLK(I2702), .RSTB(I338993), .Q(I338985) );
and I_19801 (I338958,I339290,I339259);
DFFARX1 I_19802  ( .D(I13383), .CLK(I2702), .RSTB(I338993), .Q(I339369) );
nor I_19803 (I338982,I339369,I339290);
nor I_19804 (I339400,I339369,I339044);
nand I_19805 (I338979,I339078,I339400);
not I_19806 (I338976,I339369);
DFFARX1 I_19807  ( .D(I13377), .CLK(I2702), .RSTB(I338993), .Q(I339445) );
not I_19808 (I339462,I339445);
nor I_19809 (I339479,I339462,I339143);
and I_19810 (I339496,I339369,I339479);
or I_19811 (I339513,I339290,I339496);
DFFARX1 I_19812  ( .D(I339513), .CLK(I2702), .RSTB(I338993), .Q(I338970) );
not I_19813 (I339544,I339462);
nor I_19814 (I339561,I339369,I339544);
nand I_19815 (I338973,I339462,I339561);
nand I_19816 (I338967,I339126,I339544);
not I_19817 (I339639,I2709);
not I_19818 (I339656,I558383);
nor I_19819 (I339673,I558395,I558389);
nand I_19820 (I339690,I339673,I558374);
nor I_19821 (I339707,I339656,I558395);
nand I_19822 (I339724,I339707,I558401);
DFFARX1 I_19823  ( .D(I339724), .CLK(I2702), .RSTB(I339639), .Q(I339741) );
not I_19824 (I339610,I339741);
not I_19825 (I339772,I558395);
not I_19826 (I339789,I339772);
not I_19827 (I339806,I558398);
nor I_19828 (I339823,I339806,I558380);
and I_19829 (I339840,I339823,I558377);
or I_19830 (I339857,I339840,I558404);
DFFARX1 I_19831  ( .D(I339857), .CLK(I2702), .RSTB(I339639), .Q(I339874) );
DFFARX1 I_19832  ( .D(I339874), .CLK(I2702), .RSTB(I339639), .Q(I339607) );
DFFARX1 I_19833  ( .D(I339874), .CLK(I2702), .RSTB(I339639), .Q(I339905) );
DFFARX1 I_19834  ( .D(I339874), .CLK(I2702), .RSTB(I339639), .Q(I339601) );
nand I_19835 (I339936,I339656,I558398);
nand I_19836 (I339953,I339936,I339690);
and I_19837 (I339970,I339772,I339953);
DFFARX1 I_19838  ( .D(I339970), .CLK(I2702), .RSTB(I339639), .Q(I339631) );
and I_19839 (I339604,I339936,I339905);
DFFARX1 I_19840  ( .D(I558392), .CLK(I2702), .RSTB(I339639), .Q(I340015) );
nor I_19841 (I339628,I340015,I339936);
nor I_19842 (I340046,I340015,I339690);
nand I_19843 (I339625,I339724,I340046);
not I_19844 (I339622,I340015);
DFFARX1 I_19845  ( .D(I558386), .CLK(I2702), .RSTB(I339639), .Q(I340091) );
not I_19846 (I340108,I340091);
nor I_19847 (I340125,I340108,I339789);
and I_19848 (I340142,I340015,I340125);
or I_19849 (I340159,I339936,I340142);
DFFARX1 I_19850  ( .D(I340159), .CLK(I2702), .RSTB(I339639), .Q(I339616) );
not I_19851 (I340190,I340108);
nor I_19852 (I340207,I340015,I340190);
nand I_19853 (I339619,I340108,I340207);
nand I_19854 (I339613,I339772,I340190);
not I_19855 (I340285,I2709);
not I_19856 (I340302,I123416);
nor I_19857 (I340319,I123407,I123398);
nand I_19858 (I340336,I340319,I123413);
nor I_19859 (I340353,I340302,I123407);
nand I_19860 (I340370,I340353,I123410);
DFFARX1 I_19861  ( .D(I340370), .CLK(I2702), .RSTB(I340285), .Q(I340387) );
not I_19862 (I340256,I340387);
not I_19863 (I340418,I123407);
not I_19864 (I340435,I340418);
not I_19865 (I340452,I123419);
nor I_19866 (I340469,I340452,I123404);
and I_19867 (I340486,I340469,I123422);
or I_19868 (I340503,I340486,I123395);
DFFARX1 I_19869  ( .D(I340503), .CLK(I2702), .RSTB(I340285), .Q(I340520) );
DFFARX1 I_19870  ( .D(I340520), .CLK(I2702), .RSTB(I340285), .Q(I340253) );
DFFARX1 I_19871  ( .D(I340520), .CLK(I2702), .RSTB(I340285), .Q(I340551) );
DFFARX1 I_19872  ( .D(I340520), .CLK(I2702), .RSTB(I340285), .Q(I340247) );
nand I_19873 (I340582,I340302,I123419);
nand I_19874 (I340599,I340582,I340336);
and I_19875 (I340616,I340418,I340599);
DFFARX1 I_19876  ( .D(I340616), .CLK(I2702), .RSTB(I340285), .Q(I340277) );
and I_19877 (I340250,I340582,I340551);
DFFARX1 I_19878  ( .D(I123425), .CLK(I2702), .RSTB(I340285), .Q(I340661) );
nor I_19879 (I340274,I340661,I340582);
nor I_19880 (I340692,I340661,I340336);
nand I_19881 (I340271,I340370,I340692);
not I_19882 (I340268,I340661);
DFFARX1 I_19883  ( .D(I123401), .CLK(I2702), .RSTB(I340285), .Q(I340737) );
not I_19884 (I340754,I340737);
nor I_19885 (I340771,I340754,I340435);
and I_19886 (I340788,I340661,I340771);
or I_19887 (I340805,I340582,I340788);
DFFARX1 I_19888  ( .D(I340805), .CLK(I2702), .RSTB(I340285), .Q(I340262) );
not I_19889 (I340836,I340754);
nor I_19890 (I340853,I340661,I340836);
nand I_19891 (I340265,I340754,I340853);
nand I_19892 (I340259,I340418,I340836);
not I_19893 (I340931,I2709);
not I_19894 (I340948,I116310);
nor I_19895 (I340965,I116301,I116292);
nand I_19896 (I340982,I340965,I116307);
nor I_19897 (I340999,I340948,I116301);
nand I_19898 (I341016,I340999,I116304);
DFFARX1 I_19899  ( .D(I341016), .CLK(I2702), .RSTB(I340931), .Q(I341033) );
not I_19900 (I340902,I341033);
not I_19901 (I341064,I116301);
not I_19902 (I341081,I341064);
not I_19903 (I341098,I116313);
nor I_19904 (I341115,I341098,I116298);
and I_19905 (I341132,I341115,I116316);
or I_19906 (I341149,I341132,I116289);
DFFARX1 I_19907  ( .D(I341149), .CLK(I2702), .RSTB(I340931), .Q(I341166) );
DFFARX1 I_19908  ( .D(I341166), .CLK(I2702), .RSTB(I340931), .Q(I340899) );
DFFARX1 I_19909  ( .D(I341166), .CLK(I2702), .RSTB(I340931), .Q(I341197) );
DFFARX1 I_19910  ( .D(I341166), .CLK(I2702), .RSTB(I340931), .Q(I340893) );
nand I_19911 (I341228,I340948,I116313);
nand I_19912 (I341245,I341228,I340982);
and I_19913 (I341262,I341064,I341245);
DFFARX1 I_19914  ( .D(I341262), .CLK(I2702), .RSTB(I340931), .Q(I340923) );
and I_19915 (I340896,I341228,I341197);
DFFARX1 I_19916  ( .D(I116319), .CLK(I2702), .RSTB(I340931), .Q(I341307) );
nor I_19917 (I340920,I341307,I341228);
nor I_19918 (I341338,I341307,I340982);
nand I_19919 (I340917,I341016,I341338);
not I_19920 (I340914,I341307);
DFFARX1 I_19921  ( .D(I116295), .CLK(I2702), .RSTB(I340931), .Q(I341383) );
not I_19922 (I341400,I341383);
nor I_19923 (I341417,I341400,I341081);
and I_19924 (I341434,I341307,I341417);
or I_19925 (I341451,I341228,I341434);
DFFARX1 I_19926  ( .D(I341451), .CLK(I2702), .RSTB(I340931), .Q(I340908) );
not I_19927 (I341482,I341400);
nor I_19928 (I341499,I341307,I341482);
nand I_19929 (I340911,I341400,I341499);
nand I_19930 (I340905,I341064,I341482);
not I_19931 (I341577,I2709);
not I_19932 (I341594,I52356);
nor I_19933 (I341611,I52347,I52338);
nand I_19934 (I341628,I341611,I52353);
nor I_19935 (I341645,I341594,I52347);
nand I_19936 (I341662,I341645,I52350);
DFFARX1 I_19937  ( .D(I341662), .CLK(I2702), .RSTB(I341577), .Q(I341679) );
not I_19938 (I341548,I341679);
not I_19939 (I341710,I52347);
not I_19940 (I341727,I341710);
not I_19941 (I341744,I52359);
nor I_19942 (I341761,I341744,I52344);
and I_19943 (I341778,I341761,I52362);
or I_19944 (I341795,I341778,I52335);
DFFARX1 I_19945  ( .D(I341795), .CLK(I2702), .RSTB(I341577), .Q(I341812) );
DFFARX1 I_19946  ( .D(I341812), .CLK(I2702), .RSTB(I341577), .Q(I341545) );
DFFARX1 I_19947  ( .D(I341812), .CLK(I2702), .RSTB(I341577), .Q(I341843) );
DFFARX1 I_19948  ( .D(I341812), .CLK(I2702), .RSTB(I341577), .Q(I341539) );
nand I_19949 (I341874,I341594,I52359);
nand I_19950 (I341891,I341874,I341628);
and I_19951 (I341908,I341710,I341891);
DFFARX1 I_19952  ( .D(I341908), .CLK(I2702), .RSTB(I341577), .Q(I341569) );
and I_19953 (I341542,I341874,I341843);
DFFARX1 I_19954  ( .D(I52365), .CLK(I2702), .RSTB(I341577), .Q(I341953) );
nor I_19955 (I341566,I341953,I341874);
nor I_19956 (I341984,I341953,I341628);
nand I_19957 (I341563,I341662,I341984);
not I_19958 (I341560,I341953);
DFFARX1 I_19959  ( .D(I52341), .CLK(I2702), .RSTB(I341577), .Q(I342029) );
not I_19960 (I342046,I342029);
nor I_19961 (I342063,I342046,I341727);
and I_19962 (I342080,I341953,I342063);
or I_19963 (I342097,I341874,I342080);
DFFARX1 I_19964  ( .D(I342097), .CLK(I2702), .RSTB(I341577), .Q(I341554) );
not I_19965 (I342128,I342046);
nor I_19966 (I342145,I341953,I342128);
nand I_19967 (I341557,I342046,I342145);
nand I_19968 (I341551,I341710,I342128);
not I_19969 (I342223,I2709);
not I_19970 (I342240,I620615);
nor I_19971 (I342257,I620612,I620597);
nand I_19972 (I342274,I342257,I620606);
nor I_19973 (I342291,I342240,I620612);
nand I_19974 (I342308,I342291,I620621);
DFFARX1 I_19975  ( .D(I342308), .CLK(I2702), .RSTB(I342223), .Q(I342325) );
not I_19976 (I342194,I342325);
not I_19977 (I342356,I620612);
not I_19978 (I342373,I342356);
not I_19979 (I342390,I620594);
nor I_19980 (I342407,I342390,I620600);
and I_19981 (I342424,I342407,I620624);
or I_19982 (I342441,I342424,I620618);
DFFARX1 I_19983  ( .D(I342441), .CLK(I2702), .RSTB(I342223), .Q(I342458) );
DFFARX1 I_19984  ( .D(I342458), .CLK(I2702), .RSTB(I342223), .Q(I342191) );
DFFARX1 I_19985  ( .D(I342458), .CLK(I2702), .RSTB(I342223), .Q(I342489) );
DFFARX1 I_19986  ( .D(I342458), .CLK(I2702), .RSTB(I342223), .Q(I342185) );
nand I_19987 (I342520,I342240,I620594);
nand I_19988 (I342537,I342520,I342274);
and I_19989 (I342554,I342356,I342537);
DFFARX1 I_19990  ( .D(I342554), .CLK(I2702), .RSTB(I342223), .Q(I342215) );
and I_19991 (I342188,I342520,I342489);
DFFARX1 I_19992  ( .D(I620603), .CLK(I2702), .RSTB(I342223), .Q(I342599) );
nor I_19993 (I342212,I342599,I342520);
nor I_19994 (I342630,I342599,I342274);
nand I_19995 (I342209,I342308,I342630);
not I_19996 (I342206,I342599);
DFFARX1 I_19997  ( .D(I620609), .CLK(I2702), .RSTB(I342223), .Q(I342675) );
not I_19998 (I342692,I342675);
nor I_19999 (I342709,I342692,I342373);
and I_20000 (I342726,I342599,I342709);
or I_20001 (I342743,I342520,I342726);
DFFARX1 I_20002  ( .D(I342743), .CLK(I2702), .RSTB(I342223), .Q(I342200) );
not I_20003 (I342774,I342692);
nor I_20004 (I342791,I342599,I342774);
nand I_20005 (I342203,I342692,I342791);
nand I_20006 (I342197,I342356,I342774);
not I_20007 (I342869,I2709);
not I_20008 (I342886,I41991);
nor I_20009 (I342903,I42006,I42000);
nand I_20010 (I342920,I342903,I42009);
nor I_20011 (I342937,I342886,I42006);
nand I_20012 (I342954,I342937,I41985);
DFFARX1 I_20013  ( .D(I342954), .CLK(I2702), .RSTB(I342869), .Q(I342971) );
not I_20014 (I342840,I342971);
not I_20015 (I343002,I42006);
not I_20016 (I343019,I343002);
not I_20017 (I343036,I41982);
nor I_20018 (I343053,I343036,I41997);
and I_20019 (I343070,I343053,I42003);
or I_20020 (I343087,I343070,I42012);
DFFARX1 I_20021  ( .D(I343087), .CLK(I2702), .RSTB(I342869), .Q(I343104) );
DFFARX1 I_20022  ( .D(I343104), .CLK(I2702), .RSTB(I342869), .Q(I342837) );
DFFARX1 I_20023  ( .D(I343104), .CLK(I2702), .RSTB(I342869), .Q(I343135) );
DFFARX1 I_20024  ( .D(I343104), .CLK(I2702), .RSTB(I342869), .Q(I342831) );
nand I_20025 (I343166,I342886,I41982);
nand I_20026 (I343183,I343166,I342920);
and I_20027 (I343200,I343002,I343183);
DFFARX1 I_20028  ( .D(I343200), .CLK(I2702), .RSTB(I342869), .Q(I342861) );
and I_20029 (I342834,I343166,I343135);
DFFARX1 I_20030  ( .D(I41994), .CLK(I2702), .RSTB(I342869), .Q(I343245) );
nor I_20031 (I342858,I343245,I343166);
nor I_20032 (I343276,I343245,I342920);
nand I_20033 (I342855,I342954,I343276);
not I_20034 (I342852,I343245);
DFFARX1 I_20035  ( .D(I41988), .CLK(I2702), .RSTB(I342869), .Q(I343321) );
not I_20036 (I343338,I343321);
nor I_20037 (I343355,I343338,I343019);
and I_20038 (I343372,I343245,I343355);
or I_20039 (I343389,I343166,I343372);
DFFARX1 I_20040  ( .D(I343389), .CLK(I2702), .RSTB(I342869), .Q(I342846) );
not I_20041 (I343420,I343338);
nor I_20042 (I343437,I343245,I343420);
nand I_20043 (I342849,I343338,I343437);
nand I_20044 (I342843,I343002,I343420);
not I_20045 (I343515,I2709);
not I_20046 (I343532,I582192);
nor I_20047 (I343549,I582180,I582189);
nand I_20048 (I343566,I343549,I582204);
nor I_20049 (I343583,I343532,I582180);
nand I_20050 (I343600,I343583,I582186);
DFFARX1 I_20051  ( .D(I343600), .CLK(I2702), .RSTB(I343515), .Q(I343617) );
not I_20052 (I343486,I343617);
not I_20053 (I343648,I582180);
not I_20054 (I343665,I343648);
not I_20055 (I343682,I582174);
nor I_20056 (I343699,I343682,I582195);
and I_20057 (I343716,I343699,I582177);
or I_20058 (I343733,I343716,I582183);
DFFARX1 I_20059  ( .D(I343733), .CLK(I2702), .RSTB(I343515), .Q(I343750) );
DFFARX1 I_20060  ( .D(I343750), .CLK(I2702), .RSTB(I343515), .Q(I343483) );
DFFARX1 I_20061  ( .D(I343750), .CLK(I2702), .RSTB(I343515), .Q(I343781) );
DFFARX1 I_20062  ( .D(I343750), .CLK(I2702), .RSTB(I343515), .Q(I343477) );
nand I_20063 (I343812,I343532,I582174);
nand I_20064 (I343829,I343812,I343566);
and I_20065 (I343846,I343648,I343829);
DFFARX1 I_20066  ( .D(I343846), .CLK(I2702), .RSTB(I343515), .Q(I343507) );
and I_20067 (I343480,I343812,I343781);
DFFARX1 I_20068  ( .D(I582201), .CLK(I2702), .RSTB(I343515), .Q(I343891) );
nor I_20069 (I343504,I343891,I343812);
nor I_20070 (I343922,I343891,I343566);
nand I_20071 (I343501,I343600,I343922);
not I_20072 (I343498,I343891);
DFFARX1 I_20073  ( .D(I582198), .CLK(I2702), .RSTB(I343515), .Q(I343967) );
not I_20074 (I343984,I343967);
nor I_20075 (I344001,I343984,I343665);
and I_20076 (I344018,I343891,I344001);
or I_20077 (I344035,I343812,I344018);
DFFARX1 I_20078  ( .D(I344035), .CLK(I2702), .RSTB(I343515), .Q(I343492) );
not I_20079 (I344066,I343984);
nor I_20080 (I344083,I343891,I344066);
nand I_20081 (I343495,I343984,I344083);
nand I_20082 (I343489,I343648,I344066);
not I_20083 (I344161,I2709);
not I_20084 (I344178,I328524);
nor I_20085 (I344195,I328503,I328515);
nand I_20086 (I344212,I344195,I328518);
nor I_20087 (I344229,I344178,I328503);
nand I_20088 (I344246,I344229,I328500);
DFFARX1 I_20089  ( .D(I344246), .CLK(I2702), .RSTB(I344161), .Q(I344263) );
not I_20090 (I344132,I344263);
not I_20091 (I344294,I328503);
not I_20092 (I344311,I344294);
not I_20093 (I344328,I328521);
nor I_20094 (I344345,I344328,I328512);
and I_20095 (I344362,I344345,I328506);
or I_20096 (I344379,I344362,I328530);
DFFARX1 I_20097  ( .D(I344379), .CLK(I2702), .RSTB(I344161), .Q(I344396) );
DFFARX1 I_20098  ( .D(I344396), .CLK(I2702), .RSTB(I344161), .Q(I344129) );
DFFARX1 I_20099  ( .D(I344396), .CLK(I2702), .RSTB(I344161), .Q(I344427) );
DFFARX1 I_20100  ( .D(I344396), .CLK(I2702), .RSTB(I344161), .Q(I344123) );
nand I_20101 (I344458,I344178,I328521);
nand I_20102 (I344475,I344458,I344212);
and I_20103 (I344492,I344294,I344475);
DFFARX1 I_20104  ( .D(I344492), .CLK(I2702), .RSTB(I344161), .Q(I344153) );
and I_20105 (I344126,I344458,I344427);
DFFARX1 I_20106  ( .D(I328527), .CLK(I2702), .RSTB(I344161), .Q(I344537) );
nor I_20107 (I344150,I344537,I344458);
nor I_20108 (I344568,I344537,I344212);
nand I_20109 (I344147,I344246,I344568);
not I_20110 (I344144,I344537);
DFFARX1 I_20111  ( .D(I328509), .CLK(I2702), .RSTB(I344161), .Q(I344613) );
not I_20112 (I344630,I344613);
nor I_20113 (I344647,I344630,I344311);
and I_20114 (I344664,I344537,I344647);
or I_20115 (I344681,I344458,I344664);
DFFARX1 I_20116  ( .D(I344681), .CLK(I2702), .RSTB(I344161), .Q(I344138) );
not I_20117 (I344712,I344630);
nor I_20118 (I344729,I344537,I344712);
nand I_20119 (I344141,I344630,I344729);
nand I_20120 (I344135,I344294,I344712);
not I_20121 (I344807,I2709);
not I_20122 (I344824,I531608);
nor I_20123 (I344841,I531620,I531614);
nand I_20124 (I344858,I344841,I531599);
nor I_20125 (I344875,I344824,I531620);
nand I_20126 (I344892,I344875,I531626);
DFFARX1 I_20127  ( .D(I344892), .CLK(I2702), .RSTB(I344807), .Q(I344909) );
not I_20128 (I344778,I344909);
not I_20129 (I344940,I531620);
not I_20130 (I344957,I344940);
not I_20131 (I344974,I531623);
nor I_20132 (I344991,I344974,I531605);
and I_20133 (I345008,I344991,I531602);
or I_20134 (I345025,I345008,I531629);
DFFARX1 I_20135  ( .D(I345025), .CLK(I2702), .RSTB(I344807), .Q(I345042) );
DFFARX1 I_20136  ( .D(I345042), .CLK(I2702), .RSTB(I344807), .Q(I344775) );
DFFARX1 I_20137  ( .D(I345042), .CLK(I2702), .RSTB(I344807), .Q(I345073) );
DFFARX1 I_20138  ( .D(I345042), .CLK(I2702), .RSTB(I344807), .Q(I344769) );
nand I_20139 (I345104,I344824,I531623);
nand I_20140 (I345121,I345104,I344858);
and I_20141 (I345138,I344940,I345121);
DFFARX1 I_20142  ( .D(I345138), .CLK(I2702), .RSTB(I344807), .Q(I344799) );
and I_20143 (I344772,I345104,I345073);
DFFARX1 I_20144  ( .D(I531617), .CLK(I2702), .RSTB(I344807), .Q(I345183) );
nor I_20145 (I344796,I345183,I345104);
nor I_20146 (I345214,I345183,I344858);
nand I_20147 (I344793,I344892,I345214);
not I_20148 (I344790,I345183);
DFFARX1 I_20149  ( .D(I531611), .CLK(I2702), .RSTB(I344807), .Q(I345259) );
not I_20150 (I345276,I345259);
nor I_20151 (I345293,I345276,I344957);
and I_20152 (I345310,I345183,I345293);
or I_20153 (I345327,I345104,I345310);
DFFARX1 I_20154  ( .D(I345327), .CLK(I2702), .RSTB(I344807), .Q(I344784) );
not I_20155 (I345358,I345276);
nor I_20156 (I345375,I345183,I345358);
nand I_20157 (I344787,I345276,I345375);
nand I_20158 (I344781,I344940,I345358);
not I_20159 (I345453,I2709);
not I_20160 (I345470,I295374);
nor I_20161 (I345487,I295353,I295365);
nand I_20162 (I345504,I345487,I295368);
nor I_20163 (I345521,I345470,I295353);
nand I_20164 (I345538,I345521,I295350);
DFFARX1 I_20165  ( .D(I345538), .CLK(I2702), .RSTB(I345453), .Q(I345555) );
not I_20166 (I345424,I345555);
not I_20167 (I345586,I295353);
not I_20168 (I345603,I345586);
not I_20169 (I345620,I295371);
nor I_20170 (I345637,I345620,I295362);
and I_20171 (I345654,I345637,I295356);
or I_20172 (I345671,I345654,I295380);
DFFARX1 I_20173  ( .D(I345671), .CLK(I2702), .RSTB(I345453), .Q(I345688) );
DFFARX1 I_20174  ( .D(I345688), .CLK(I2702), .RSTB(I345453), .Q(I345421) );
DFFARX1 I_20175  ( .D(I345688), .CLK(I2702), .RSTB(I345453), .Q(I345719) );
DFFARX1 I_20176  ( .D(I345688), .CLK(I2702), .RSTB(I345453), .Q(I345415) );
nand I_20177 (I345750,I345470,I295371);
nand I_20178 (I345767,I345750,I345504);
and I_20179 (I345784,I345586,I345767);
DFFARX1 I_20180  ( .D(I345784), .CLK(I2702), .RSTB(I345453), .Q(I345445) );
and I_20181 (I345418,I345750,I345719);
DFFARX1 I_20182  ( .D(I295377), .CLK(I2702), .RSTB(I345453), .Q(I345829) );
nor I_20183 (I345442,I345829,I345750);
nor I_20184 (I345860,I345829,I345504);
nand I_20185 (I345439,I345538,I345860);
not I_20186 (I345436,I345829);
DFFARX1 I_20187  ( .D(I295359), .CLK(I2702), .RSTB(I345453), .Q(I345905) );
not I_20188 (I345922,I345905);
nor I_20189 (I345939,I345922,I345603);
and I_20190 (I345956,I345829,I345939);
or I_20191 (I345973,I345750,I345956);
DFFARX1 I_20192  ( .D(I345973), .CLK(I2702), .RSTB(I345453), .Q(I345430) );
not I_20193 (I346004,I345922);
nor I_20194 (I346021,I345829,I346004);
nand I_20195 (I345433,I345922,I346021);
nand I_20196 (I345427,I345586,I346004);
not I_20197 (I346099,I2709);
not I_20198 (I346116,I307308);
nor I_20199 (I346133,I307287,I307299);
nand I_20200 (I346150,I346133,I307302);
nor I_20201 (I346167,I346116,I307287);
nand I_20202 (I346184,I346167,I307284);
DFFARX1 I_20203  ( .D(I346184), .CLK(I2702), .RSTB(I346099), .Q(I346201) );
not I_20204 (I346070,I346201);
not I_20205 (I346232,I307287);
not I_20206 (I346249,I346232);
not I_20207 (I346266,I307305);
nor I_20208 (I346283,I346266,I307296);
and I_20209 (I346300,I346283,I307290);
or I_20210 (I346317,I346300,I307314);
DFFARX1 I_20211  ( .D(I346317), .CLK(I2702), .RSTB(I346099), .Q(I346334) );
DFFARX1 I_20212  ( .D(I346334), .CLK(I2702), .RSTB(I346099), .Q(I346067) );
DFFARX1 I_20213  ( .D(I346334), .CLK(I2702), .RSTB(I346099), .Q(I346365) );
DFFARX1 I_20214  ( .D(I346334), .CLK(I2702), .RSTB(I346099), .Q(I346061) );
nand I_20215 (I346396,I346116,I307305);
nand I_20216 (I346413,I346396,I346150);
and I_20217 (I346430,I346232,I346413);
DFFARX1 I_20218  ( .D(I346430), .CLK(I2702), .RSTB(I346099), .Q(I346091) );
and I_20219 (I346064,I346396,I346365);
DFFARX1 I_20220  ( .D(I307311), .CLK(I2702), .RSTB(I346099), .Q(I346475) );
nor I_20221 (I346088,I346475,I346396);
nor I_20222 (I346506,I346475,I346150);
nand I_20223 (I346085,I346184,I346506);
not I_20224 (I346082,I346475);
DFFARX1 I_20225  ( .D(I307293), .CLK(I2702), .RSTB(I346099), .Q(I346551) );
not I_20226 (I346568,I346551);
nor I_20227 (I346585,I346568,I346249);
and I_20228 (I346602,I346475,I346585);
or I_20229 (I346619,I346396,I346602);
DFFARX1 I_20230  ( .D(I346619), .CLK(I2702), .RSTB(I346099), .Q(I346076) );
not I_20231 (I346650,I346568);
nor I_20232 (I346667,I346475,I346650);
nand I_20233 (I346079,I346568,I346667);
nand I_20234 (I346073,I346232,I346650);
not I_20235 (I346745,I2709);
not I_20236 (I346762,I556598);
nor I_20237 (I346779,I556610,I556604);
nand I_20238 (I346796,I346779,I556589);
nor I_20239 (I346813,I346762,I556610);
nand I_20240 (I346830,I346813,I556616);
DFFARX1 I_20241  ( .D(I346830), .CLK(I2702), .RSTB(I346745), .Q(I346847) );
not I_20242 (I346716,I346847);
not I_20243 (I346878,I556610);
not I_20244 (I346895,I346878);
not I_20245 (I346912,I556613);
nor I_20246 (I346929,I346912,I556595);
and I_20247 (I346946,I346929,I556592);
or I_20248 (I346963,I346946,I556619);
DFFARX1 I_20249  ( .D(I346963), .CLK(I2702), .RSTB(I346745), .Q(I346980) );
DFFARX1 I_20250  ( .D(I346980), .CLK(I2702), .RSTB(I346745), .Q(I346713) );
DFFARX1 I_20251  ( .D(I346980), .CLK(I2702), .RSTB(I346745), .Q(I347011) );
DFFARX1 I_20252  ( .D(I346980), .CLK(I2702), .RSTB(I346745), .Q(I346707) );
nand I_20253 (I347042,I346762,I556613);
nand I_20254 (I347059,I347042,I346796);
and I_20255 (I347076,I346878,I347059);
DFFARX1 I_20256  ( .D(I347076), .CLK(I2702), .RSTB(I346745), .Q(I346737) );
and I_20257 (I346710,I347042,I347011);
DFFARX1 I_20258  ( .D(I556607), .CLK(I2702), .RSTB(I346745), .Q(I347121) );
nor I_20259 (I346734,I347121,I347042);
nor I_20260 (I347152,I347121,I346796);
nand I_20261 (I346731,I346830,I347152);
not I_20262 (I346728,I347121);
DFFARX1 I_20263  ( .D(I556601), .CLK(I2702), .RSTB(I346745), .Q(I347197) );
not I_20264 (I347214,I347197);
nor I_20265 (I347231,I347214,I346895);
and I_20266 (I347248,I347121,I347231);
or I_20267 (I347265,I347042,I347248);
DFFARX1 I_20268  ( .D(I347265), .CLK(I2702), .RSTB(I346745), .Q(I346722) );
not I_20269 (I347296,I347214);
nor I_20270 (I347313,I347121,I347296);
nand I_20271 (I346725,I347214,I347313);
nand I_20272 (I346719,I346878,I347296);
not I_20273 (I347391,I2709);
not I_20274 (I347408,I27405);
nor I_20275 (I347425,I27420,I27414);
nand I_20276 (I347442,I347425,I27423);
nor I_20277 (I347459,I347408,I27420);
nand I_20278 (I347476,I347459,I27399);
DFFARX1 I_20279  ( .D(I347476), .CLK(I2702), .RSTB(I347391), .Q(I347493) );
not I_20280 (I347362,I347493);
not I_20281 (I347524,I27420);
not I_20282 (I347541,I347524);
not I_20283 (I347558,I27396);
nor I_20284 (I347575,I347558,I27411);
and I_20285 (I347592,I347575,I27417);
or I_20286 (I347609,I347592,I27426);
DFFARX1 I_20287  ( .D(I347609), .CLK(I2702), .RSTB(I347391), .Q(I347626) );
DFFARX1 I_20288  ( .D(I347626), .CLK(I2702), .RSTB(I347391), .Q(I347359) );
DFFARX1 I_20289  ( .D(I347626), .CLK(I2702), .RSTB(I347391), .Q(I347657) );
DFFARX1 I_20290  ( .D(I347626), .CLK(I2702), .RSTB(I347391), .Q(I347353) );
nand I_20291 (I347688,I347408,I27396);
nand I_20292 (I347705,I347688,I347442);
and I_20293 (I347722,I347524,I347705);
DFFARX1 I_20294  ( .D(I347722), .CLK(I2702), .RSTB(I347391), .Q(I347383) );
and I_20295 (I347356,I347688,I347657);
DFFARX1 I_20296  ( .D(I27408), .CLK(I2702), .RSTB(I347391), .Q(I347767) );
nor I_20297 (I347380,I347767,I347688);
nor I_20298 (I347798,I347767,I347442);
nand I_20299 (I347377,I347476,I347798);
not I_20300 (I347374,I347767);
DFFARX1 I_20301  ( .D(I27402), .CLK(I2702), .RSTB(I347391), .Q(I347843) );
not I_20302 (I347860,I347843);
nor I_20303 (I347877,I347860,I347541);
and I_20304 (I347894,I347767,I347877);
or I_20305 (I347911,I347688,I347894);
DFFARX1 I_20306  ( .D(I347911), .CLK(I2702), .RSTB(I347391), .Q(I347368) );
not I_20307 (I347942,I347860);
nor I_20308 (I347959,I347767,I347942);
nand I_20309 (I347371,I347860,I347959);
nand I_20310 (I347365,I347524,I347942);
not I_20311 (I348037,I2709);
not I_20312 (I348054,I133752);
nor I_20313 (I348071,I133743,I133734);
nand I_20314 (I348088,I348071,I133749);
nor I_20315 (I348105,I348054,I133743);
nand I_20316 (I348122,I348105,I133746);
DFFARX1 I_20317  ( .D(I348122), .CLK(I2702), .RSTB(I348037), .Q(I348139) );
not I_20318 (I348008,I348139);
not I_20319 (I348170,I133743);
not I_20320 (I348187,I348170);
not I_20321 (I348204,I133755);
nor I_20322 (I348221,I348204,I133740);
and I_20323 (I348238,I348221,I133758);
or I_20324 (I348255,I348238,I133731);
DFFARX1 I_20325  ( .D(I348255), .CLK(I2702), .RSTB(I348037), .Q(I348272) );
DFFARX1 I_20326  ( .D(I348272), .CLK(I2702), .RSTB(I348037), .Q(I348005) );
DFFARX1 I_20327  ( .D(I348272), .CLK(I2702), .RSTB(I348037), .Q(I348303) );
DFFARX1 I_20328  ( .D(I348272), .CLK(I2702), .RSTB(I348037), .Q(I347999) );
nand I_20329 (I348334,I348054,I133755);
nand I_20330 (I348351,I348334,I348088);
and I_20331 (I348368,I348170,I348351);
DFFARX1 I_20332  ( .D(I348368), .CLK(I2702), .RSTB(I348037), .Q(I348029) );
and I_20333 (I348002,I348334,I348303);
DFFARX1 I_20334  ( .D(I133761), .CLK(I2702), .RSTB(I348037), .Q(I348413) );
nor I_20335 (I348026,I348413,I348334);
nor I_20336 (I348444,I348413,I348088);
nand I_20337 (I348023,I348122,I348444);
not I_20338 (I348020,I348413);
DFFARX1 I_20339  ( .D(I133737), .CLK(I2702), .RSTB(I348037), .Q(I348489) );
not I_20340 (I348506,I348489);
nor I_20341 (I348523,I348506,I348187);
and I_20342 (I348540,I348413,I348523);
or I_20343 (I348557,I348334,I348540);
DFFARX1 I_20344  ( .D(I348557), .CLK(I2702), .RSTB(I348037), .Q(I348014) );
not I_20345 (I348588,I348506);
nor I_20346 (I348605,I348413,I348588);
nand I_20347 (I348017,I348506,I348605);
nand I_20348 (I348011,I348170,I348588);
not I_20349 (I348683,I2709);
not I_20350 (I348700,I64630);
nor I_20351 (I348717,I64621,I64612);
nand I_20352 (I348734,I348717,I64627);
nor I_20353 (I348751,I348700,I64621);
nand I_20354 (I348768,I348751,I64624);
DFFARX1 I_20355  ( .D(I348768), .CLK(I2702), .RSTB(I348683), .Q(I348785) );
not I_20356 (I348654,I348785);
not I_20357 (I348816,I64621);
not I_20358 (I348833,I348816);
not I_20359 (I348850,I64633);
nor I_20360 (I348867,I348850,I64618);
and I_20361 (I348884,I348867,I64636);
or I_20362 (I348901,I348884,I64609);
DFFARX1 I_20363  ( .D(I348901), .CLK(I2702), .RSTB(I348683), .Q(I348918) );
DFFARX1 I_20364  ( .D(I348918), .CLK(I2702), .RSTB(I348683), .Q(I348651) );
DFFARX1 I_20365  ( .D(I348918), .CLK(I2702), .RSTB(I348683), .Q(I348949) );
DFFARX1 I_20366  ( .D(I348918), .CLK(I2702), .RSTB(I348683), .Q(I348645) );
nand I_20367 (I348980,I348700,I64633);
nand I_20368 (I348997,I348980,I348734);
and I_20369 (I349014,I348816,I348997);
DFFARX1 I_20370  ( .D(I349014), .CLK(I2702), .RSTB(I348683), .Q(I348675) );
and I_20371 (I348648,I348980,I348949);
DFFARX1 I_20372  ( .D(I64639), .CLK(I2702), .RSTB(I348683), .Q(I349059) );
nor I_20373 (I348672,I349059,I348980);
nor I_20374 (I349090,I349059,I348734);
nand I_20375 (I348669,I348768,I349090);
not I_20376 (I348666,I349059);
DFFARX1 I_20377  ( .D(I64615), .CLK(I2702), .RSTB(I348683), .Q(I349135) );
not I_20378 (I349152,I349135);
nor I_20379 (I349169,I349152,I348833);
and I_20380 (I349186,I349059,I349169);
or I_20381 (I349203,I348980,I349186);
DFFARX1 I_20382  ( .D(I349203), .CLK(I2702), .RSTB(I348683), .Q(I348660) );
not I_20383 (I349234,I349152);
nor I_20384 (I349251,I349059,I349234);
nand I_20385 (I348663,I349152,I349251);
nand I_20386 (I348657,I348816,I349234);
not I_20387 (I349329,I2709);
not I_20388 (I349346,I24039);
nor I_20389 (I349363,I24054,I24048);
nand I_20390 (I349380,I349363,I24057);
nor I_20391 (I349397,I349346,I24054);
nand I_20392 (I349414,I349397,I24033);
DFFARX1 I_20393  ( .D(I349414), .CLK(I2702), .RSTB(I349329), .Q(I349431) );
not I_20394 (I349300,I349431);
not I_20395 (I349462,I24054);
not I_20396 (I349479,I349462);
not I_20397 (I349496,I24030);
nor I_20398 (I349513,I349496,I24045);
and I_20399 (I349530,I349513,I24051);
or I_20400 (I349547,I349530,I24060);
DFFARX1 I_20401  ( .D(I349547), .CLK(I2702), .RSTB(I349329), .Q(I349564) );
DFFARX1 I_20402  ( .D(I349564), .CLK(I2702), .RSTB(I349329), .Q(I349297) );
DFFARX1 I_20403  ( .D(I349564), .CLK(I2702), .RSTB(I349329), .Q(I349595) );
DFFARX1 I_20404  ( .D(I349564), .CLK(I2702), .RSTB(I349329), .Q(I349291) );
nand I_20405 (I349626,I349346,I24030);
nand I_20406 (I349643,I349626,I349380);
and I_20407 (I349660,I349462,I349643);
DFFARX1 I_20408  ( .D(I349660), .CLK(I2702), .RSTB(I349329), .Q(I349321) );
and I_20409 (I349294,I349626,I349595);
DFFARX1 I_20410  ( .D(I24042), .CLK(I2702), .RSTB(I349329), .Q(I349705) );
nor I_20411 (I349318,I349705,I349626);
nor I_20412 (I349736,I349705,I349380);
nand I_20413 (I349315,I349414,I349736);
not I_20414 (I349312,I349705);
DFFARX1 I_20415  ( .D(I24036), .CLK(I2702), .RSTB(I349329), .Q(I349781) );
not I_20416 (I349798,I349781);
nor I_20417 (I349815,I349798,I349479);
and I_20418 (I349832,I349705,I349815);
or I_20419 (I349849,I349626,I349832);
DFFARX1 I_20420  ( .D(I349849), .CLK(I2702), .RSTB(I349329), .Q(I349306) );
not I_20421 (I349880,I349798);
nor I_20422 (I349897,I349705,I349880);
nand I_20423 (I349309,I349798,I349897);
nand I_20424 (I349303,I349462,I349880);
not I_20425 (I349975,I2709);
not I_20426 (I349992,I423599);
nor I_20427 (I350009,I423608,I423593);
nand I_20428 (I350026,I350009,I423581);
nor I_20429 (I350043,I349992,I423608);
nand I_20430 (I350060,I350043,I423584);
DFFARX1 I_20431  ( .D(I350060), .CLK(I2702), .RSTB(I349975), .Q(I350077) );
not I_20432 (I349946,I350077);
not I_20433 (I350108,I423608);
not I_20434 (I350125,I350108);
not I_20435 (I350142,I423596);
nor I_20436 (I350159,I350142,I423590);
and I_20437 (I350176,I350159,I423587);
or I_20438 (I350193,I350176,I423602);
DFFARX1 I_20439  ( .D(I350193), .CLK(I2702), .RSTB(I349975), .Q(I350210) );
DFFARX1 I_20440  ( .D(I350210), .CLK(I2702), .RSTB(I349975), .Q(I349943) );
DFFARX1 I_20441  ( .D(I350210), .CLK(I2702), .RSTB(I349975), .Q(I350241) );
DFFARX1 I_20442  ( .D(I350210), .CLK(I2702), .RSTB(I349975), .Q(I349937) );
nand I_20443 (I350272,I349992,I423596);
nand I_20444 (I350289,I350272,I350026);
and I_20445 (I350306,I350108,I350289);
DFFARX1 I_20446  ( .D(I350306), .CLK(I2702), .RSTB(I349975), .Q(I349967) );
and I_20447 (I349940,I350272,I350241);
DFFARX1 I_20448  ( .D(I423611), .CLK(I2702), .RSTB(I349975), .Q(I350351) );
nor I_20449 (I349964,I350351,I350272);
nor I_20450 (I350382,I350351,I350026);
nand I_20451 (I349961,I350060,I350382);
not I_20452 (I349958,I350351);
DFFARX1 I_20453  ( .D(I423605), .CLK(I2702), .RSTB(I349975), .Q(I350427) );
not I_20454 (I350444,I350427);
nor I_20455 (I350461,I350444,I350125);
and I_20456 (I350478,I350351,I350461);
or I_20457 (I350495,I350272,I350478);
DFFARX1 I_20458  ( .D(I350495), .CLK(I2702), .RSTB(I349975), .Q(I349952) );
not I_20459 (I350526,I350444);
nor I_20460 (I350543,I350351,I350526);
nand I_20461 (I349955,I350444,I350543);
nand I_20462 (I349949,I350108,I350526);
not I_20463 (I350621,I2709);
not I_20464 (I350638,I719858);
nor I_20465 (I350655,I719843,I719849);
nand I_20466 (I350672,I350655,I719846);
nor I_20467 (I350689,I350638,I719843);
nand I_20468 (I350706,I350689,I719855);
DFFARX1 I_20469  ( .D(I350706), .CLK(I2702), .RSTB(I350621), .Q(I350723) );
not I_20470 (I350592,I350723);
not I_20471 (I350754,I719843);
not I_20472 (I350771,I350754);
not I_20473 (I350788,I719870);
nor I_20474 (I350805,I350788,I719864);
and I_20475 (I350822,I350805,I719861);
or I_20476 (I350839,I350822,I719840);
DFFARX1 I_20477  ( .D(I350839), .CLK(I2702), .RSTB(I350621), .Q(I350856) );
DFFARX1 I_20478  ( .D(I350856), .CLK(I2702), .RSTB(I350621), .Q(I350589) );
DFFARX1 I_20479  ( .D(I350856), .CLK(I2702), .RSTB(I350621), .Q(I350887) );
DFFARX1 I_20480  ( .D(I350856), .CLK(I2702), .RSTB(I350621), .Q(I350583) );
nand I_20481 (I350918,I350638,I719870);
nand I_20482 (I350935,I350918,I350672);
and I_20483 (I350952,I350754,I350935);
DFFARX1 I_20484  ( .D(I350952), .CLK(I2702), .RSTB(I350621), .Q(I350613) );
and I_20485 (I350586,I350918,I350887);
DFFARX1 I_20486  ( .D(I719867), .CLK(I2702), .RSTB(I350621), .Q(I350997) );
nor I_20487 (I350610,I350997,I350918);
nor I_20488 (I351028,I350997,I350672);
nand I_20489 (I350607,I350706,I351028);
not I_20490 (I350604,I350997);
DFFARX1 I_20491  ( .D(I719852), .CLK(I2702), .RSTB(I350621), .Q(I351073) );
not I_20492 (I351090,I351073);
nor I_20493 (I351107,I351090,I350771);
and I_20494 (I351124,I350997,I351107);
or I_20495 (I351141,I350918,I351124);
DFFARX1 I_20496  ( .D(I351141), .CLK(I2702), .RSTB(I350621), .Q(I350598) );
not I_20497 (I351172,I351090);
nor I_20498 (I351189,I350997,I351172);
nand I_20499 (I350601,I351090,I351189);
nand I_20500 (I350595,I350754,I351172);
not I_20501 (I351267,I2709);
not I_20502 (I351284,I18990);
nor I_20503 (I351301,I19005,I18999);
nand I_20504 (I351318,I351301,I19008);
nor I_20505 (I351335,I351284,I19005);
nand I_20506 (I351352,I351335,I18984);
DFFARX1 I_20507  ( .D(I351352), .CLK(I2702), .RSTB(I351267), .Q(I351369) );
not I_20508 (I351238,I351369);
not I_20509 (I351400,I19005);
not I_20510 (I351417,I351400);
not I_20511 (I351434,I18981);
nor I_20512 (I351451,I351434,I18996);
and I_20513 (I351468,I351451,I19002);
or I_20514 (I351485,I351468,I19011);
DFFARX1 I_20515  ( .D(I351485), .CLK(I2702), .RSTB(I351267), .Q(I351502) );
DFFARX1 I_20516  ( .D(I351502), .CLK(I2702), .RSTB(I351267), .Q(I351235) );
DFFARX1 I_20517  ( .D(I351502), .CLK(I2702), .RSTB(I351267), .Q(I351533) );
DFFARX1 I_20518  ( .D(I351502), .CLK(I2702), .RSTB(I351267), .Q(I351229) );
nand I_20519 (I351564,I351284,I18981);
nand I_20520 (I351581,I351564,I351318);
and I_20521 (I351598,I351400,I351581);
DFFARX1 I_20522  ( .D(I351598), .CLK(I2702), .RSTB(I351267), .Q(I351259) );
and I_20523 (I351232,I351564,I351533);
DFFARX1 I_20524  ( .D(I18993), .CLK(I2702), .RSTB(I351267), .Q(I351643) );
nor I_20525 (I351256,I351643,I351564);
nor I_20526 (I351674,I351643,I351318);
nand I_20527 (I351253,I351352,I351674);
not I_20528 (I351250,I351643);
DFFARX1 I_20529  ( .D(I18987), .CLK(I2702), .RSTB(I351267), .Q(I351719) );
not I_20530 (I351736,I351719);
nor I_20531 (I351753,I351736,I351417);
and I_20532 (I351770,I351643,I351753);
or I_20533 (I351787,I351564,I351770);
DFFARX1 I_20534  ( .D(I351787), .CLK(I2702), .RSTB(I351267), .Q(I351244) );
not I_20535 (I351818,I351736);
nor I_20536 (I351835,I351643,I351818);
nand I_20537 (I351247,I351736,I351835);
nand I_20538 (I351241,I351400,I351818);
not I_20539 (I351913,I2709);
not I_20540 (I351930,I704830);
nor I_20541 (I351947,I704815,I704821);
nand I_20542 (I351964,I351947,I704818);
nor I_20543 (I351981,I351930,I704815);
nand I_20544 (I351998,I351981,I704827);
DFFARX1 I_20545  ( .D(I351998), .CLK(I2702), .RSTB(I351913), .Q(I352015) );
not I_20546 (I351884,I352015);
not I_20547 (I352046,I704815);
not I_20548 (I352063,I352046);
not I_20549 (I352080,I704842);
nor I_20550 (I352097,I352080,I704836);
and I_20551 (I352114,I352097,I704833);
or I_20552 (I352131,I352114,I704812);
DFFARX1 I_20553  ( .D(I352131), .CLK(I2702), .RSTB(I351913), .Q(I352148) );
DFFARX1 I_20554  ( .D(I352148), .CLK(I2702), .RSTB(I351913), .Q(I351881) );
DFFARX1 I_20555  ( .D(I352148), .CLK(I2702), .RSTB(I351913), .Q(I352179) );
DFFARX1 I_20556  ( .D(I352148), .CLK(I2702), .RSTB(I351913), .Q(I351875) );
nand I_20557 (I352210,I351930,I704842);
nand I_20558 (I352227,I352210,I351964);
and I_20559 (I352244,I352046,I352227);
DFFARX1 I_20560  ( .D(I352244), .CLK(I2702), .RSTB(I351913), .Q(I351905) );
and I_20561 (I351878,I352210,I352179);
DFFARX1 I_20562  ( .D(I704839), .CLK(I2702), .RSTB(I351913), .Q(I352289) );
nor I_20563 (I351902,I352289,I352210);
nor I_20564 (I352320,I352289,I351964);
nand I_20565 (I351899,I351998,I352320);
not I_20566 (I351896,I352289);
DFFARX1 I_20567  ( .D(I704824), .CLK(I2702), .RSTB(I351913), .Q(I352365) );
not I_20568 (I352382,I352365);
nor I_20569 (I352399,I352382,I352063);
and I_20570 (I352416,I352289,I352399);
or I_20571 (I352433,I352210,I352416);
DFFARX1 I_20572  ( .D(I352433), .CLK(I2702), .RSTB(I351913), .Q(I351890) );
not I_20573 (I352464,I352382);
nor I_20574 (I352481,I352289,I352464);
nand I_20575 (I351893,I352382,I352481);
nand I_20576 (I351887,I352046,I352464);
not I_20577 (I352559,I2709);
not I_20578 (I352576,I471434);
nor I_20579 (I352593,I471437,I471419);
nand I_20580 (I352610,I352593,I471446);
nor I_20581 (I352627,I352576,I471437);
nand I_20582 (I352644,I352627,I471425);
DFFARX1 I_20583  ( .D(I352644), .CLK(I2702), .RSTB(I352559), .Q(I352661) );
not I_20584 (I352530,I352661);
not I_20585 (I352692,I471437);
not I_20586 (I352709,I352692);
not I_20587 (I352726,I471431);
nor I_20588 (I352743,I352726,I471443);
and I_20589 (I352760,I352743,I471449);
or I_20590 (I352777,I352760,I471428);
DFFARX1 I_20591  ( .D(I352777), .CLK(I2702), .RSTB(I352559), .Q(I352794) );
DFFARX1 I_20592  ( .D(I352794), .CLK(I2702), .RSTB(I352559), .Q(I352527) );
DFFARX1 I_20593  ( .D(I352794), .CLK(I2702), .RSTB(I352559), .Q(I352825) );
DFFARX1 I_20594  ( .D(I352794), .CLK(I2702), .RSTB(I352559), .Q(I352521) );
nand I_20595 (I352856,I352576,I471431);
nand I_20596 (I352873,I352856,I352610);
and I_20597 (I352890,I352692,I352873);
DFFARX1 I_20598  ( .D(I352890), .CLK(I2702), .RSTB(I352559), .Q(I352551) );
and I_20599 (I352524,I352856,I352825);
DFFARX1 I_20600  ( .D(I471440), .CLK(I2702), .RSTB(I352559), .Q(I352935) );
nor I_20601 (I352548,I352935,I352856);
nor I_20602 (I352966,I352935,I352610);
nand I_20603 (I352545,I352644,I352966);
not I_20604 (I352542,I352935);
DFFARX1 I_20605  ( .D(I471422), .CLK(I2702), .RSTB(I352559), .Q(I353011) );
not I_20606 (I353028,I353011);
nor I_20607 (I353045,I353028,I352709);
and I_20608 (I353062,I352935,I353045);
or I_20609 (I353079,I352856,I353062);
DFFARX1 I_20610  ( .D(I353079), .CLK(I2702), .RSTB(I352559), .Q(I352536) );
not I_20611 (I353110,I353028);
nor I_20612 (I353127,I352935,I353110);
nand I_20613 (I352539,I353028,I353127);
nand I_20614 (I352533,I352692,I353110);
not I_20615 (I353205,I2709);
not I_20616 (I353222,I120186);
nor I_20617 (I353239,I120177,I120168);
nand I_20618 (I353256,I353239,I120183);
nor I_20619 (I353273,I353222,I120177);
nand I_20620 (I353290,I353273,I120180);
DFFARX1 I_20621  ( .D(I353290), .CLK(I2702), .RSTB(I353205), .Q(I353307) );
not I_20622 (I353176,I353307);
not I_20623 (I353338,I120177);
not I_20624 (I353355,I353338);
not I_20625 (I353372,I120189);
nor I_20626 (I353389,I353372,I120174);
and I_20627 (I353406,I353389,I120192);
or I_20628 (I353423,I353406,I120165);
DFFARX1 I_20629  ( .D(I353423), .CLK(I2702), .RSTB(I353205), .Q(I353440) );
DFFARX1 I_20630  ( .D(I353440), .CLK(I2702), .RSTB(I353205), .Q(I353173) );
DFFARX1 I_20631  ( .D(I353440), .CLK(I2702), .RSTB(I353205), .Q(I353471) );
DFFARX1 I_20632  ( .D(I353440), .CLK(I2702), .RSTB(I353205), .Q(I353167) );
nand I_20633 (I353502,I353222,I120189);
nand I_20634 (I353519,I353502,I353256);
and I_20635 (I353536,I353338,I353519);
DFFARX1 I_20636  ( .D(I353536), .CLK(I2702), .RSTB(I353205), .Q(I353197) );
and I_20637 (I353170,I353502,I353471);
DFFARX1 I_20638  ( .D(I120195), .CLK(I2702), .RSTB(I353205), .Q(I353581) );
nor I_20639 (I353194,I353581,I353502);
nor I_20640 (I353612,I353581,I353256);
nand I_20641 (I353191,I353290,I353612);
not I_20642 (I353188,I353581);
DFFARX1 I_20643  ( .D(I120171), .CLK(I2702), .RSTB(I353205), .Q(I353657) );
not I_20644 (I353674,I353657);
nor I_20645 (I353691,I353674,I353355);
and I_20646 (I353708,I353581,I353691);
or I_20647 (I353725,I353502,I353708);
DFFARX1 I_20648  ( .D(I353725), .CLK(I2702), .RSTB(I353205), .Q(I353182) );
not I_20649 (I353756,I353674);
nor I_20650 (I353773,I353581,I353756);
nand I_20651 (I353185,I353674,I353773);
nand I_20652 (I353179,I353338,I353756);
not I_20653 (I353851,I2709);
not I_20654 (I353868,I215354);
nor I_20655 (I353885,I215360,I215357);
nand I_20656 (I353902,I353885,I215351);
nor I_20657 (I353919,I353868,I215360);
nand I_20658 (I353936,I353919,I215375);
DFFARX1 I_20659  ( .D(I353936), .CLK(I2702), .RSTB(I353851), .Q(I353953) );
not I_20660 (I353822,I353953);
not I_20661 (I353984,I215360);
not I_20662 (I354001,I353984);
not I_20663 (I354018,I215372);
nor I_20664 (I354035,I354018,I215363);
and I_20665 (I354052,I354035,I215348);
or I_20666 (I354069,I354052,I215369);
DFFARX1 I_20667  ( .D(I354069), .CLK(I2702), .RSTB(I353851), .Q(I354086) );
DFFARX1 I_20668  ( .D(I354086), .CLK(I2702), .RSTB(I353851), .Q(I353819) );
DFFARX1 I_20669  ( .D(I354086), .CLK(I2702), .RSTB(I353851), .Q(I354117) );
DFFARX1 I_20670  ( .D(I354086), .CLK(I2702), .RSTB(I353851), .Q(I353813) );
nand I_20671 (I354148,I353868,I215372);
nand I_20672 (I354165,I354148,I353902);
and I_20673 (I354182,I353984,I354165);
DFFARX1 I_20674  ( .D(I354182), .CLK(I2702), .RSTB(I353851), .Q(I353843) );
and I_20675 (I353816,I354148,I354117);
DFFARX1 I_20676  ( .D(I215366), .CLK(I2702), .RSTB(I353851), .Q(I354227) );
nor I_20677 (I353840,I354227,I354148);
nor I_20678 (I354258,I354227,I353902);
nand I_20679 (I353837,I353936,I354258);
not I_20680 (I353834,I354227);
DFFARX1 I_20681  ( .D(I215378), .CLK(I2702), .RSTB(I353851), .Q(I354303) );
not I_20682 (I354320,I354303);
nor I_20683 (I354337,I354320,I354001);
and I_20684 (I354354,I354227,I354337);
or I_20685 (I354371,I354148,I354354);
DFFARX1 I_20686  ( .D(I354371), .CLK(I2702), .RSTB(I353851), .Q(I353828) );
not I_20687 (I354402,I354320);
nor I_20688 (I354419,I354227,I354402);
nand I_20689 (I353831,I354320,I354419);
nand I_20690 (I353825,I353984,I354402);
not I_20691 (I354497,I2709);
not I_20692 (I354514,I308634);
nor I_20693 (I354531,I308613,I308625);
nand I_20694 (I354548,I354531,I308628);
nor I_20695 (I354565,I354514,I308613);
nand I_20696 (I354582,I354565,I308610);
DFFARX1 I_20697  ( .D(I354582), .CLK(I2702), .RSTB(I354497), .Q(I354599) );
not I_20698 (I354468,I354599);
not I_20699 (I354630,I308613);
not I_20700 (I354647,I354630);
not I_20701 (I354664,I308631);
nor I_20702 (I354681,I354664,I308622);
and I_20703 (I354698,I354681,I308616);
or I_20704 (I354715,I354698,I308640);
DFFARX1 I_20705  ( .D(I354715), .CLK(I2702), .RSTB(I354497), .Q(I354732) );
DFFARX1 I_20706  ( .D(I354732), .CLK(I2702), .RSTB(I354497), .Q(I354465) );
DFFARX1 I_20707  ( .D(I354732), .CLK(I2702), .RSTB(I354497), .Q(I354763) );
DFFARX1 I_20708  ( .D(I354732), .CLK(I2702), .RSTB(I354497), .Q(I354459) );
nand I_20709 (I354794,I354514,I308631);
nand I_20710 (I354811,I354794,I354548);
and I_20711 (I354828,I354630,I354811);
DFFARX1 I_20712  ( .D(I354828), .CLK(I2702), .RSTB(I354497), .Q(I354489) );
and I_20713 (I354462,I354794,I354763);
DFFARX1 I_20714  ( .D(I308637), .CLK(I2702), .RSTB(I354497), .Q(I354873) );
nor I_20715 (I354486,I354873,I354794);
nor I_20716 (I354904,I354873,I354548);
nand I_20717 (I354483,I354582,I354904);
not I_20718 (I354480,I354873);
DFFARX1 I_20719  ( .D(I308619), .CLK(I2702), .RSTB(I354497), .Q(I354949) );
not I_20720 (I354966,I354949);
nor I_20721 (I354983,I354966,I354647);
and I_20722 (I355000,I354873,I354983);
or I_20723 (I355017,I354794,I355000);
DFFARX1 I_20724  ( .D(I355017), .CLK(I2702), .RSTB(I354497), .Q(I354474) );
not I_20725 (I355048,I354966);
nor I_20726 (I355065,I354873,I355048);
nand I_20727 (I354477,I354966,I355065);
nand I_20728 (I354471,I354630,I355048);
not I_20729 (I355143,I2709);
not I_20730 (I355160,I206429);
nor I_20731 (I355177,I206435,I206432);
nand I_20732 (I355194,I355177,I206426);
nor I_20733 (I355211,I355160,I206435);
nand I_20734 (I355228,I355211,I206450);
DFFARX1 I_20735  ( .D(I355228), .CLK(I2702), .RSTB(I355143), .Q(I355245) );
not I_20736 (I355114,I355245);
not I_20737 (I355276,I206435);
not I_20738 (I355293,I355276);
not I_20739 (I355310,I206447);
nor I_20740 (I355327,I355310,I206438);
and I_20741 (I355344,I355327,I206423);
or I_20742 (I355361,I355344,I206444);
DFFARX1 I_20743  ( .D(I355361), .CLK(I2702), .RSTB(I355143), .Q(I355378) );
DFFARX1 I_20744  ( .D(I355378), .CLK(I2702), .RSTB(I355143), .Q(I355111) );
DFFARX1 I_20745  ( .D(I355378), .CLK(I2702), .RSTB(I355143), .Q(I355409) );
DFFARX1 I_20746  ( .D(I355378), .CLK(I2702), .RSTB(I355143), .Q(I355105) );
nand I_20747 (I355440,I355160,I206447);
nand I_20748 (I355457,I355440,I355194);
and I_20749 (I355474,I355276,I355457);
DFFARX1 I_20750  ( .D(I355474), .CLK(I2702), .RSTB(I355143), .Q(I355135) );
and I_20751 (I355108,I355440,I355409);
DFFARX1 I_20752  ( .D(I206441), .CLK(I2702), .RSTB(I355143), .Q(I355519) );
nor I_20753 (I355132,I355519,I355440);
nor I_20754 (I355550,I355519,I355194);
nand I_20755 (I355129,I355228,I355550);
not I_20756 (I355126,I355519);
DFFARX1 I_20757  ( .D(I206453), .CLK(I2702), .RSTB(I355143), .Q(I355595) );
not I_20758 (I355612,I355595);
nor I_20759 (I355629,I355612,I355293);
and I_20760 (I355646,I355519,I355629);
or I_20761 (I355663,I355440,I355646);
DFFARX1 I_20762  ( .D(I355663), .CLK(I2702), .RSTB(I355143), .Q(I355120) );
not I_20763 (I355694,I355612);
nor I_20764 (I355711,I355519,I355694);
nand I_20765 (I355123,I355612,I355711);
nand I_20766 (I355117,I355276,I355694);
not I_20767 (I355789,I2709);
not I_20768 (I355806,I67860);
nor I_20769 (I355823,I67851,I67842);
nand I_20770 (I355840,I355823,I67857);
nor I_20771 (I355857,I355806,I67851);
nand I_20772 (I355874,I355857,I67854);
DFFARX1 I_20773  ( .D(I355874), .CLK(I2702), .RSTB(I355789), .Q(I355891) );
not I_20774 (I355760,I355891);
not I_20775 (I355922,I67851);
not I_20776 (I355939,I355922);
not I_20777 (I355956,I67863);
nor I_20778 (I355973,I355956,I67848);
and I_20779 (I355990,I355973,I67866);
or I_20780 (I356007,I355990,I67839);
DFFARX1 I_20781  ( .D(I356007), .CLK(I2702), .RSTB(I355789), .Q(I356024) );
DFFARX1 I_20782  ( .D(I356024), .CLK(I2702), .RSTB(I355789), .Q(I355757) );
DFFARX1 I_20783  ( .D(I356024), .CLK(I2702), .RSTB(I355789), .Q(I356055) );
DFFARX1 I_20784  ( .D(I356024), .CLK(I2702), .RSTB(I355789), .Q(I355751) );
nand I_20785 (I356086,I355806,I67863);
nand I_20786 (I356103,I356086,I355840);
and I_20787 (I356120,I355922,I356103);
DFFARX1 I_20788  ( .D(I356120), .CLK(I2702), .RSTB(I355789), .Q(I355781) );
and I_20789 (I355754,I356086,I356055);
DFFARX1 I_20790  ( .D(I67869), .CLK(I2702), .RSTB(I355789), .Q(I356165) );
nor I_20791 (I355778,I356165,I356086);
nor I_20792 (I356196,I356165,I355840);
nand I_20793 (I355775,I355874,I356196);
not I_20794 (I355772,I356165);
DFFARX1 I_20795  ( .D(I67845), .CLK(I2702), .RSTB(I355789), .Q(I356241) );
not I_20796 (I356258,I356241);
nor I_20797 (I356275,I356258,I355939);
and I_20798 (I356292,I356165,I356275);
or I_20799 (I356309,I356086,I356292);
DFFARX1 I_20800  ( .D(I356309), .CLK(I2702), .RSTB(I355789), .Q(I355766) );
not I_20801 (I356340,I356258);
nor I_20802 (I356357,I356165,I356340);
nand I_20803 (I355769,I356258,I356357);
nand I_20804 (I355763,I355922,I356340);
not I_20805 (I356435,I2709);
not I_20806 (I356452,I309960);
nor I_20807 (I356469,I309939,I309951);
nand I_20808 (I356486,I356469,I309954);
nor I_20809 (I356503,I356452,I309939);
nand I_20810 (I356520,I356503,I309936);
DFFARX1 I_20811  ( .D(I356520), .CLK(I2702), .RSTB(I356435), .Q(I356537) );
not I_20812 (I356406,I356537);
not I_20813 (I356568,I309939);
not I_20814 (I356585,I356568);
not I_20815 (I356602,I309957);
nor I_20816 (I356619,I356602,I309948);
and I_20817 (I356636,I356619,I309942);
or I_20818 (I356653,I356636,I309966);
DFFARX1 I_20819  ( .D(I356653), .CLK(I2702), .RSTB(I356435), .Q(I356670) );
DFFARX1 I_20820  ( .D(I356670), .CLK(I2702), .RSTB(I356435), .Q(I356403) );
DFFARX1 I_20821  ( .D(I356670), .CLK(I2702), .RSTB(I356435), .Q(I356701) );
DFFARX1 I_20822  ( .D(I356670), .CLK(I2702), .RSTB(I356435), .Q(I356397) );
nand I_20823 (I356732,I356452,I309957);
nand I_20824 (I356749,I356732,I356486);
and I_20825 (I356766,I356568,I356749);
DFFARX1 I_20826  ( .D(I356766), .CLK(I2702), .RSTB(I356435), .Q(I356427) );
and I_20827 (I356400,I356732,I356701);
DFFARX1 I_20828  ( .D(I309963), .CLK(I2702), .RSTB(I356435), .Q(I356811) );
nor I_20829 (I356424,I356811,I356732);
nor I_20830 (I356842,I356811,I356486);
nand I_20831 (I356421,I356520,I356842);
not I_20832 (I356418,I356811);
DFFARX1 I_20833  ( .D(I309945), .CLK(I2702), .RSTB(I356435), .Q(I356887) );
not I_20834 (I356904,I356887);
nor I_20835 (I356921,I356904,I356585);
and I_20836 (I356938,I356811,I356921);
or I_20837 (I356955,I356732,I356938);
DFFARX1 I_20838  ( .D(I356955), .CLK(I2702), .RSTB(I356435), .Q(I356412) );
not I_20839 (I356986,I356904);
nor I_20840 (I357003,I356811,I356986);
nand I_20841 (I356415,I356904,I357003);
nand I_20842 (I356409,I356568,I356986);
not I_20843 (I357081,I2709);
not I_20844 (I357098,I557788);
nor I_20845 (I357115,I557800,I557794);
nand I_20846 (I357132,I357115,I557779);
nor I_20847 (I357149,I357098,I557800);
nand I_20848 (I357166,I357149,I557806);
DFFARX1 I_20849  ( .D(I357166), .CLK(I2702), .RSTB(I357081), .Q(I357183) );
not I_20850 (I357052,I357183);
not I_20851 (I357214,I557800);
not I_20852 (I357231,I357214);
not I_20853 (I357248,I557803);
nor I_20854 (I357265,I357248,I557785);
and I_20855 (I357282,I357265,I557782);
or I_20856 (I357299,I357282,I557809);
DFFARX1 I_20857  ( .D(I357299), .CLK(I2702), .RSTB(I357081), .Q(I357316) );
DFFARX1 I_20858  ( .D(I357316), .CLK(I2702), .RSTB(I357081), .Q(I357049) );
DFFARX1 I_20859  ( .D(I357316), .CLK(I2702), .RSTB(I357081), .Q(I357347) );
DFFARX1 I_20860  ( .D(I357316), .CLK(I2702), .RSTB(I357081), .Q(I357043) );
nand I_20861 (I357378,I357098,I557803);
nand I_20862 (I357395,I357378,I357132);
and I_20863 (I357412,I357214,I357395);
DFFARX1 I_20864  ( .D(I357412), .CLK(I2702), .RSTB(I357081), .Q(I357073) );
and I_20865 (I357046,I357378,I357347);
DFFARX1 I_20866  ( .D(I557797), .CLK(I2702), .RSTB(I357081), .Q(I357457) );
nor I_20867 (I357070,I357457,I357378);
nor I_20868 (I357488,I357457,I357132);
nand I_20869 (I357067,I357166,I357488);
not I_20870 (I357064,I357457);
DFFARX1 I_20871  ( .D(I557791), .CLK(I2702), .RSTB(I357081), .Q(I357533) );
not I_20872 (I357550,I357533);
nor I_20873 (I357567,I357550,I357231);
and I_20874 (I357584,I357457,I357567);
or I_20875 (I357601,I357378,I357584);
DFFARX1 I_20876  ( .D(I357601), .CLK(I2702), .RSTB(I357081), .Q(I357058) );
not I_20877 (I357632,I357550);
nor I_20878 (I357649,I357457,I357632);
nand I_20879 (I357061,I357550,I357649);
nand I_20880 (I357055,I357214,I357632);
not I_20881 (I357727,I2709);
not I_20882 (I357744,I175350);
nor I_20883 (I357761,I175371,I175353);
nand I_20884 (I357778,I357761,I175377);
nor I_20885 (I357795,I357744,I175371);
nand I_20886 (I357812,I357795,I175374);
DFFARX1 I_20887  ( .D(I357812), .CLK(I2702), .RSTB(I357727), .Q(I357829) );
not I_20888 (I357698,I357829);
not I_20889 (I357860,I175371);
not I_20890 (I357877,I357860);
not I_20891 (I357894,I175368);
nor I_20892 (I357911,I357894,I175347);
and I_20893 (I357928,I357911,I175359);
or I_20894 (I357945,I357928,I175356);
DFFARX1 I_20895  ( .D(I357945), .CLK(I2702), .RSTB(I357727), .Q(I357962) );
DFFARX1 I_20896  ( .D(I357962), .CLK(I2702), .RSTB(I357727), .Q(I357695) );
DFFARX1 I_20897  ( .D(I357962), .CLK(I2702), .RSTB(I357727), .Q(I357993) );
DFFARX1 I_20898  ( .D(I357962), .CLK(I2702), .RSTB(I357727), .Q(I357689) );
nand I_20899 (I358024,I357744,I175368);
nand I_20900 (I358041,I358024,I357778);
and I_20901 (I358058,I357860,I358041);
DFFARX1 I_20902  ( .D(I358058), .CLK(I2702), .RSTB(I357727), .Q(I357719) );
and I_20903 (I357692,I358024,I357993);
DFFARX1 I_20904  ( .D(I175362), .CLK(I2702), .RSTB(I357727), .Q(I358103) );
nor I_20905 (I357716,I358103,I358024);
nor I_20906 (I358134,I358103,I357778);
nand I_20907 (I357713,I357812,I358134);
not I_20908 (I357710,I358103);
DFFARX1 I_20909  ( .D(I175365), .CLK(I2702), .RSTB(I357727), .Q(I358179) );
not I_20910 (I358196,I358179);
nor I_20911 (I358213,I358196,I357877);
and I_20912 (I358230,I358103,I358213);
or I_20913 (I358247,I358024,I358230);
DFFARX1 I_20914  ( .D(I358247), .CLK(I2702), .RSTB(I357727), .Q(I357704) );
not I_20915 (I358278,I358196);
nor I_20916 (I358295,I358103,I358278);
nand I_20917 (I357707,I358196,I358295);
nand I_20918 (I357701,I357860,I358278);
not I_20919 (I358373,I2709);
not I_20920 (I358390,I74320);
nor I_20921 (I358407,I74311,I74302);
nand I_20922 (I358424,I358407,I74317);
nor I_20923 (I358441,I358390,I74311);
nand I_20924 (I358458,I358441,I74314);
DFFARX1 I_20925  ( .D(I358458), .CLK(I2702), .RSTB(I358373), .Q(I358475) );
not I_20926 (I358344,I358475);
not I_20927 (I358506,I74311);
not I_20928 (I358523,I358506);
not I_20929 (I358540,I74323);
nor I_20930 (I358557,I358540,I74308);
and I_20931 (I358574,I358557,I74326);
or I_20932 (I358591,I358574,I74299);
DFFARX1 I_20933  ( .D(I358591), .CLK(I2702), .RSTB(I358373), .Q(I358608) );
DFFARX1 I_20934  ( .D(I358608), .CLK(I2702), .RSTB(I358373), .Q(I358341) );
DFFARX1 I_20935  ( .D(I358608), .CLK(I2702), .RSTB(I358373), .Q(I358639) );
DFFARX1 I_20936  ( .D(I358608), .CLK(I2702), .RSTB(I358373), .Q(I358335) );
nand I_20937 (I358670,I358390,I74323);
nand I_20938 (I358687,I358670,I358424);
and I_20939 (I358704,I358506,I358687);
DFFARX1 I_20940  ( .D(I358704), .CLK(I2702), .RSTB(I358373), .Q(I358365) );
and I_20941 (I358338,I358670,I358639);
DFFARX1 I_20942  ( .D(I74329), .CLK(I2702), .RSTB(I358373), .Q(I358749) );
nor I_20943 (I358362,I358749,I358670);
nor I_20944 (I358780,I358749,I358424);
nand I_20945 (I358359,I358458,I358780);
not I_20946 (I358356,I358749);
DFFARX1 I_20947  ( .D(I74305), .CLK(I2702), .RSTB(I358373), .Q(I358825) );
not I_20948 (I358842,I358825);
nor I_20949 (I358859,I358842,I358523);
and I_20950 (I358876,I358749,I358859);
or I_20951 (I358893,I358670,I358876);
DFFARX1 I_20952  ( .D(I358893), .CLK(I2702), .RSTB(I358373), .Q(I358350) );
not I_20953 (I358924,I358842);
nor I_20954 (I358941,I358749,I358924);
nand I_20955 (I358353,I358842,I358941);
nand I_20956 (I358347,I358506,I358924);
not I_20957 (I359019,I2709);
not I_20958 (I359036,I674709);
nor I_20959 (I359053,I674706,I674691);
nand I_20960 (I359070,I359053,I674700);
nor I_20961 (I359087,I359036,I674706);
nand I_20962 (I359104,I359087,I674715);
DFFARX1 I_20963  ( .D(I359104), .CLK(I2702), .RSTB(I359019), .Q(I359121) );
not I_20964 (I358990,I359121);
not I_20965 (I359152,I674706);
not I_20966 (I359169,I359152);
not I_20967 (I359186,I674688);
nor I_20968 (I359203,I359186,I674694);
and I_20969 (I359220,I359203,I674718);
or I_20970 (I359237,I359220,I674712);
DFFARX1 I_20971  ( .D(I359237), .CLK(I2702), .RSTB(I359019), .Q(I359254) );
DFFARX1 I_20972  ( .D(I359254), .CLK(I2702), .RSTB(I359019), .Q(I358987) );
DFFARX1 I_20973  ( .D(I359254), .CLK(I2702), .RSTB(I359019), .Q(I359285) );
DFFARX1 I_20974  ( .D(I359254), .CLK(I2702), .RSTB(I359019), .Q(I358981) );
nand I_20975 (I359316,I359036,I674688);
nand I_20976 (I359333,I359316,I359070);
and I_20977 (I359350,I359152,I359333);
DFFARX1 I_20978  ( .D(I359350), .CLK(I2702), .RSTB(I359019), .Q(I359011) );
and I_20979 (I358984,I359316,I359285);
DFFARX1 I_20980  ( .D(I674697), .CLK(I2702), .RSTB(I359019), .Q(I359395) );
nor I_20981 (I359008,I359395,I359316);
nor I_20982 (I359426,I359395,I359070);
nand I_20983 (I359005,I359104,I359426);
not I_20984 (I359002,I359395);
DFFARX1 I_20985  ( .D(I674703), .CLK(I2702), .RSTB(I359019), .Q(I359471) );
not I_20986 (I359488,I359471);
nor I_20987 (I359505,I359488,I359169);
and I_20988 (I359522,I359395,I359505);
or I_20989 (I359539,I359316,I359522);
DFFARX1 I_20990  ( .D(I359539), .CLK(I2702), .RSTB(I359019), .Q(I358996) );
not I_20991 (I359570,I359488);
nor I_20992 (I359587,I359395,I359570);
nand I_20993 (I358999,I359488,I359587);
nand I_20994 (I358993,I359152,I359570);
not I_20995 (I359665,I2709);
not I_20996 (I359682,I502547);
nor I_20997 (I359699,I502553,I502538);
nand I_20998 (I359716,I359699,I502532);
nor I_20999 (I359733,I359682,I502553);
nand I_21000 (I359750,I359733,I502559);
DFFARX1 I_21001  ( .D(I359750), .CLK(I2702), .RSTB(I359665), .Q(I359767) );
not I_21002 (I359636,I359767);
not I_21003 (I359798,I502553);
not I_21004 (I359815,I359798);
not I_21005 (I359832,I502544);
nor I_21006 (I359849,I359832,I502550);
and I_21007 (I359866,I359849,I502556);
or I_21008 (I359883,I359866,I502529);
DFFARX1 I_21009  ( .D(I359883), .CLK(I2702), .RSTB(I359665), .Q(I359900) );
DFFARX1 I_21010  ( .D(I359900), .CLK(I2702), .RSTB(I359665), .Q(I359633) );
DFFARX1 I_21011  ( .D(I359900), .CLK(I2702), .RSTB(I359665), .Q(I359931) );
DFFARX1 I_21012  ( .D(I359900), .CLK(I2702), .RSTB(I359665), .Q(I359627) );
nand I_21013 (I359962,I359682,I502544);
nand I_21014 (I359979,I359962,I359716);
and I_21015 (I359996,I359798,I359979);
DFFARX1 I_21016  ( .D(I359996), .CLK(I2702), .RSTB(I359665), .Q(I359657) );
and I_21017 (I359630,I359962,I359931);
DFFARX1 I_21018  ( .D(I502535), .CLK(I2702), .RSTB(I359665), .Q(I360041) );
nor I_21019 (I359654,I360041,I359962);
nor I_21020 (I360072,I360041,I359716);
nand I_21021 (I359651,I359750,I360072);
not I_21022 (I359648,I360041);
DFFARX1 I_21023  ( .D(I502541), .CLK(I2702), .RSTB(I359665), .Q(I360117) );
not I_21024 (I360134,I360117);
nor I_21025 (I360151,I360134,I359815);
and I_21026 (I360168,I360041,I360151);
or I_21027 (I360185,I359962,I360168);
DFFARX1 I_21028  ( .D(I360185), .CLK(I2702), .RSTB(I359665), .Q(I359642) );
not I_21029 (I360216,I360134);
nor I_21030 (I360233,I360041,I360216);
nand I_21031 (I359645,I360134,I360233);
nand I_21032 (I359639,I359798,I360216);
not I_21033 (I360311,I2709);
not I_21034 (I360328,I35259);
nor I_21035 (I360345,I35274,I35268);
nand I_21036 (I360362,I360345,I35277);
nor I_21037 (I360379,I360328,I35274);
nand I_21038 (I360396,I360379,I35253);
DFFARX1 I_21039  ( .D(I360396), .CLK(I2702), .RSTB(I360311), .Q(I360413) );
not I_21040 (I360282,I360413);
not I_21041 (I360444,I35274);
not I_21042 (I360461,I360444);
not I_21043 (I360478,I35250);
nor I_21044 (I360495,I360478,I35265);
and I_21045 (I360512,I360495,I35271);
or I_21046 (I360529,I360512,I35280);
DFFARX1 I_21047  ( .D(I360529), .CLK(I2702), .RSTB(I360311), .Q(I360546) );
DFFARX1 I_21048  ( .D(I360546), .CLK(I2702), .RSTB(I360311), .Q(I360279) );
DFFARX1 I_21049  ( .D(I360546), .CLK(I2702), .RSTB(I360311), .Q(I360577) );
DFFARX1 I_21050  ( .D(I360546), .CLK(I2702), .RSTB(I360311), .Q(I360273) );
nand I_21051 (I360608,I360328,I35250);
nand I_21052 (I360625,I360608,I360362);
and I_21053 (I360642,I360444,I360625);
DFFARX1 I_21054  ( .D(I360642), .CLK(I2702), .RSTB(I360311), .Q(I360303) );
and I_21055 (I360276,I360608,I360577);
DFFARX1 I_21056  ( .D(I35262), .CLK(I2702), .RSTB(I360311), .Q(I360687) );
nor I_21057 (I360300,I360687,I360608);
nor I_21058 (I360718,I360687,I360362);
nand I_21059 (I360297,I360396,I360718);
not I_21060 (I360294,I360687);
DFFARX1 I_21061  ( .D(I35256), .CLK(I2702), .RSTB(I360311), .Q(I360763) );
not I_21062 (I360780,I360763);
nor I_21063 (I360797,I360780,I360461);
and I_21064 (I360814,I360687,I360797);
or I_21065 (I360831,I360608,I360814);
DFFARX1 I_21066  ( .D(I360831), .CLK(I2702), .RSTB(I360311), .Q(I360288) );
not I_21067 (I360862,I360780);
nor I_21068 (I360879,I360687,I360862);
nand I_21069 (I360291,I360780,I360879);
nand I_21070 (I360285,I360444,I360862);
not I_21071 (I360957,I2709);
not I_21072 (I360974,I456406);
nor I_21073 (I360991,I456409,I456391);
nand I_21074 (I361008,I360991,I456418);
nor I_21075 (I361025,I360974,I456409);
nand I_21076 (I361042,I361025,I456397);
DFFARX1 I_21077  ( .D(I361042), .CLK(I2702), .RSTB(I360957), .Q(I361059) );
not I_21078 (I360928,I361059);
not I_21079 (I361090,I456409);
not I_21080 (I361107,I361090);
not I_21081 (I361124,I456403);
nor I_21082 (I361141,I361124,I456415);
and I_21083 (I361158,I361141,I456421);
or I_21084 (I361175,I361158,I456400);
DFFARX1 I_21085  ( .D(I361175), .CLK(I2702), .RSTB(I360957), .Q(I361192) );
DFFARX1 I_21086  ( .D(I361192), .CLK(I2702), .RSTB(I360957), .Q(I360925) );
DFFARX1 I_21087  ( .D(I361192), .CLK(I2702), .RSTB(I360957), .Q(I361223) );
DFFARX1 I_21088  ( .D(I361192), .CLK(I2702), .RSTB(I360957), .Q(I360919) );
nand I_21089 (I361254,I360974,I456403);
nand I_21090 (I361271,I361254,I361008);
and I_21091 (I361288,I361090,I361271);
DFFARX1 I_21092  ( .D(I361288), .CLK(I2702), .RSTB(I360957), .Q(I360949) );
and I_21093 (I360922,I361254,I361223);
DFFARX1 I_21094  ( .D(I456412), .CLK(I2702), .RSTB(I360957), .Q(I361333) );
nor I_21095 (I360946,I361333,I361254);
nor I_21096 (I361364,I361333,I361008);
nand I_21097 (I360943,I361042,I361364);
not I_21098 (I360940,I361333);
DFFARX1 I_21099  ( .D(I456394), .CLK(I2702), .RSTB(I360957), .Q(I361409) );
not I_21100 (I361426,I361409);
nor I_21101 (I361443,I361426,I361107);
and I_21102 (I361460,I361333,I361443);
or I_21103 (I361477,I361254,I361460);
DFFARX1 I_21104  ( .D(I361477), .CLK(I2702), .RSTB(I360957), .Q(I360934) );
not I_21105 (I361508,I361426);
nor I_21106 (I361525,I361333,I361508);
nand I_21107 (I360937,I361426,I361525);
nand I_21108 (I360931,I361090,I361508);
not I_21109 (I361603,I2709);
not I_21110 (I361620,I508998);
nor I_21111 (I361637,I509010,I509004);
nand I_21112 (I361654,I361637,I508989);
nor I_21113 (I361671,I361620,I509010);
nand I_21114 (I361688,I361671,I509016);
DFFARX1 I_21115  ( .D(I361688), .CLK(I2702), .RSTB(I361603), .Q(I361705) );
not I_21116 (I361574,I361705);
not I_21117 (I361736,I509010);
not I_21118 (I361753,I361736);
not I_21119 (I361770,I509013);
nor I_21120 (I361787,I361770,I508995);
and I_21121 (I361804,I361787,I508992);
or I_21122 (I361821,I361804,I509019);
DFFARX1 I_21123  ( .D(I361821), .CLK(I2702), .RSTB(I361603), .Q(I361838) );
DFFARX1 I_21124  ( .D(I361838), .CLK(I2702), .RSTB(I361603), .Q(I361571) );
DFFARX1 I_21125  ( .D(I361838), .CLK(I2702), .RSTB(I361603), .Q(I361869) );
DFFARX1 I_21126  ( .D(I361838), .CLK(I2702), .RSTB(I361603), .Q(I361565) );
nand I_21127 (I361900,I361620,I509013);
nand I_21128 (I361917,I361900,I361654);
and I_21129 (I361934,I361736,I361917);
DFFARX1 I_21130  ( .D(I361934), .CLK(I2702), .RSTB(I361603), .Q(I361595) );
and I_21131 (I361568,I361900,I361869);
DFFARX1 I_21132  ( .D(I509007), .CLK(I2702), .RSTB(I361603), .Q(I361979) );
nor I_21133 (I361592,I361979,I361900);
nor I_21134 (I362010,I361979,I361654);
nand I_21135 (I361589,I361688,I362010);
not I_21136 (I361586,I361979);
DFFARX1 I_21137  ( .D(I509001), .CLK(I2702), .RSTB(I361603), .Q(I362055) );
not I_21138 (I362072,I362055);
nor I_21139 (I362089,I362072,I361753);
and I_21140 (I362106,I361979,I362089);
or I_21141 (I362123,I361900,I362106);
DFFARX1 I_21142  ( .D(I362123), .CLK(I2702), .RSTB(I361603), .Q(I361580) );
not I_21143 (I362154,I362072);
nor I_21144 (I362171,I361979,I362154);
nand I_21145 (I361583,I362072,I362171);
nand I_21146 (I361577,I361736,I362154);
not I_21147 (I362249,I2709);
not I_21148 (I362266,I168720);
nor I_21149 (I362283,I168741,I168723);
nand I_21150 (I362300,I362283,I168747);
nor I_21151 (I362317,I362266,I168741);
nand I_21152 (I362334,I362317,I168744);
DFFARX1 I_21153  ( .D(I362334), .CLK(I2702), .RSTB(I362249), .Q(I362351) );
not I_21154 (I362220,I362351);
not I_21155 (I362382,I168741);
not I_21156 (I362399,I362382);
not I_21157 (I362416,I168738);
nor I_21158 (I362433,I362416,I168717);
and I_21159 (I362450,I362433,I168729);
or I_21160 (I362467,I362450,I168726);
DFFARX1 I_21161  ( .D(I362467), .CLK(I2702), .RSTB(I362249), .Q(I362484) );
DFFARX1 I_21162  ( .D(I362484), .CLK(I2702), .RSTB(I362249), .Q(I362217) );
DFFARX1 I_21163  ( .D(I362484), .CLK(I2702), .RSTB(I362249), .Q(I362515) );
DFFARX1 I_21164  ( .D(I362484), .CLK(I2702), .RSTB(I362249), .Q(I362211) );
nand I_21165 (I362546,I362266,I168738);
nand I_21166 (I362563,I362546,I362300);
and I_21167 (I362580,I362382,I362563);
DFFARX1 I_21168  ( .D(I362580), .CLK(I2702), .RSTB(I362249), .Q(I362241) );
and I_21169 (I362214,I362546,I362515);
DFFARX1 I_21170  ( .D(I168732), .CLK(I2702), .RSTB(I362249), .Q(I362625) );
nor I_21171 (I362238,I362625,I362546);
nor I_21172 (I362656,I362625,I362300);
nand I_21173 (I362235,I362334,I362656);
not I_21174 (I362232,I362625);
DFFARX1 I_21175  ( .D(I168735), .CLK(I2702), .RSTB(I362249), .Q(I362701) );
not I_21176 (I362718,I362701);
nor I_21177 (I362735,I362718,I362399);
and I_21178 (I362752,I362625,I362735);
or I_21179 (I362769,I362546,I362752);
DFFARX1 I_21180  ( .D(I362769), .CLK(I2702), .RSTB(I362249), .Q(I362226) );
not I_21181 (I362800,I362718);
nor I_21182 (I362817,I362625,I362800);
nand I_21183 (I362229,I362718,I362817);
nand I_21184 (I362223,I362382,I362800);
not I_21185 (I362895,I2709);
not I_21186 (I362912,I292722);
nor I_21187 (I362929,I292701,I292713);
nand I_21188 (I362946,I362929,I292716);
nor I_21189 (I362963,I362912,I292701);
nand I_21190 (I362980,I362963,I292698);
DFFARX1 I_21191  ( .D(I362980), .CLK(I2702), .RSTB(I362895), .Q(I362997) );
not I_21192 (I362866,I362997);
not I_21193 (I363028,I292701);
not I_21194 (I363045,I363028);
not I_21195 (I363062,I292719);
nor I_21196 (I363079,I363062,I292710);
and I_21197 (I363096,I363079,I292704);
or I_21198 (I363113,I363096,I292728);
DFFARX1 I_21199  ( .D(I363113), .CLK(I2702), .RSTB(I362895), .Q(I363130) );
DFFARX1 I_21200  ( .D(I363130), .CLK(I2702), .RSTB(I362895), .Q(I362863) );
DFFARX1 I_21201  ( .D(I363130), .CLK(I2702), .RSTB(I362895), .Q(I363161) );
DFFARX1 I_21202  ( .D(I363130), .CLK(I2702), .RSTB(I362895), .Q(I362857) );
nand I_21203 (I363192,I362912,I292719);
nand I_21204 (I363209,I363192,I362946);
and I_21205 (I363226,I363028,I363209);
DFFARX1 I_21206  ( .D(I363226), .CLK(I2702), .RSTB(I362895), .Q(I362887) );
and I_21207 (I362860,I363192,I363161);
DFFARX1 I_21208  ( .D(I292725), .CLK(I2702), .RSTB(I362895), .Q(I363271) );
nor I_21209 (I362884,I363271,I363192);
nor I_21210 (I363302,I363271,I362946);
nand I_21211 (I362881,I362980,I363302);
not I_21212 (I362878,I363271);
DFFARX1 I_21213  ( .D(I292707), .CLK(I2702), .RSTB(I362895), .Q(I363347) );
not I_21214 (I363364,I363347);
nor I_21215 (I363381,I363364,I363045);
and I_21216 (I363398,I363271,I363381);
or I_21217 (I363415,I363192,I363398);
DFFARX1 I_21218  ( .D(I363415), .CLK(I2702), .RSTB(I362895), .Q(I362872) );
not I_21219 (I363446,I363364);
nor I_21220 (I363463,I363271,I363446);
nand I_21221 (I362875,I363364,I363463);
nand I_21222 (I362869,I363028,I363446);
not I_21223 (I363541,I2709);
not I_21224 (I363558,I298689);
nor I_21225 (I363575,I298668,I298680);
nand I_21226 (I363592,I363575,I298683);
nor I_21227 (I363609,I363558,I298668);
nand I_21228 (I363626,I363609,I298665);
DFFARX1 I_21229  ( .D(I363626), .CLK(I2702), .RSTB(I363541), .Q(I363643) );
not I_21230 (I363512,I363643);
not I_21231 (I363674,I298668);
not I_21232 (I363691,I363674);
not I_21233 (I363708,I298686);
nor I_21234 (I363725,I363708,I298677);
and I_21235 (I363742,I363725,I298671);
or I_21236 (I363759,I363742,I298695);
DFFARX1 I_21237  ( .D(I363759), .CLK(I2702), .RSTB(I363541), .Q(I363776) );
DFFARX1 I_21238  ( .D(I363776), .CLK(I2702), .RSTB(I363541), .Q(I363509) );
DFFARX1 I_21239  ( .D(I363776), .CLK(I2702), .RSTB(I363541), .Q(I363807) );
DFFARX1 I_21240  ( .D(I363776), .CLK(I2702), .RSTB(I363541), .Q(I363503) );
nand I_21241 (I363838,I363558,I298686);
nand I_21242 (I363855,I363838,I363592);
and I_21243 (I363872,I363674,I363855);
DFFARX1 I_21244  ( .D(I363872), .CLK(I2702), .RSTB(I363541), .Q(I363533) );
and I_21245 (I363506,I363838,I363807);
DFFARX1 I_21246  ( .D(I298692), .CLK(I2702), .RSTB(I363541), .Q(I363917) );
nor I_21247 (I363530,I363917,I363838);
nor I_21248 (I363948,I363917,I363592);
nand I_21249 (I363527,I363626,I363948);
not I_21250 (I363524,I363917);
DFFARX1 I_21251  ( .D(I298674), .CLK(I2702), .RSTB(I363541), .Q(I363993) );
not I_21252 (I364010,I363993);
nor I_21253 (I364027,I364010,I363691);
and I_21254 (I364044,I363917,I364027);
or I_21255 (I364061,I363838,I364044);
DFFARX1 I_21256  ( .D(I364061), .CLK(I2702), .RSTB(I363541), .Q(I363518) );
not I_21257 (I364092,I364010);
nor I_21258 (I364109,I363917,I364092);
nand I_21259 (I363521,I364010,I364109);
nand I_21260 (I363515,I363674,I364092);
not I_21261 (I364187,I2709);
not I_21262 (I364204,I174024);
nor I_21263 (I364221,I174045,I174027);
nand I_21264 (I364238,I364221,I174051);
nor I_21265 (I364255,I364204,I174045);
nand I_21266 (I364272,I364255,I174048);
DFFARX1 I_21267  ( .D(I364272), .CLK(I2702), .RSTB(I364187), .Q(I364289) );
not I_21268 (I364158,I364289);
not I_21269 (I364320,I174045);
not I_21270 (I364337,I364320);
not I_21271 (I364354,I174042);
nor I_21272 (I364371,I364354,I174021);
and I_21273 (I364388,I364371,I174033);
or I_21274 (I364405,I364388,I174030);
DFFARX1 I_21275  ( .D(I364405), .CLK(I2702), .RSTB(I364187), .Q(I364422) );
DFFARX1 I_21276  ( .D(I364422), .CLK(I2702), .RSTB(I364187), .Q(I364155) );
DFFARX1 I_21277  ( .D(I364422), .CLK(I2702), .RSTB(I364187), .Q(I364453) );
DFFARX1 I_21278  ( .D(I364422), .CLK(I2702), .RSTB(I364187), .Q(I364149) );
nand I_21279 (I364484,I364204,I174042);
nand I_21280 (I364501,I364484,I364238);
and I_21281 (I364518,I364320,I364501);
DFFARX1 I_21282  ( .D(I364518), .CLK(I2702), .RSTB(I364187), .Q(I364179) );
and I_21283 (I364152,I364484,I364453);
DFFARX1 I_21284  ( .D(I174036), .CLK(I2702), .RSTB(I364187), .Q(I364563) );
nor I_21285 (I364176,I364563,I364484);
nor I_21286 (I364594,I364563,I364238);
nand I_21287 (I364173,I364272,I364594);
not I_21288 (I364170,I364563);
DFFARX1 I_21289  ( .D(I174039), .CLK(I2702), .RSTB(I364187), .Q(I364639) );
not I_21290 (I364656,I364639);
nor I_21291 (I364673,I364656,I364337);
and I_21292 (I364690,I364563,I364673);
or I_21293 (I364707,I364484,I364690);
DFFARX1 I_21294  ( .D(I364707), .CLK(I2702), .RSTB(I364187), .Q(I364164) );
not I_21295 (I364738,I364656);
nor I_21296 (I364755,I364563,I364738);
nand I_21297 (I364167,I364656,I364755);
nand I_21298 (I364161,I364320,I364738);
not I_21299 (I364833,I2709);
not I_21300 (I364850,I599447);
nor I_21301 (I364867,I599435,I599444);
nand I_21302 (I364884,I364867,I599459);
nor I_21303 (I364901,I364850,I599435);
nand I_21304 (I364918,I364901,I599441);
DFFARX1 I_21305  ( .D(I364918), .CLK(I2702), .RSTB(I364833), .Q(I364935) );
not I_21306 (I364804,I364935);
not I_21307 (I364966,I599435);
not I_21308 (I364983,I364966);
not I_21309 (I365000,I599429);
nor I_21310 (I365017,I365000,I599450);
and I_21311 (I365034,I365017,I599432);
or I_21312 (I365051,I365034,I599438);
DFFARX1 I_21313  ( .D(I365051), .CLK(I2702), .RSTB(I364833), .Q(I365068) );
DFFARX1 I_21314  ( .D(I365068), .CLK(I2702), .RSTB(I364833), .Q(I364801) );
DFFARX1 I_21315  ( .D(I365068), .CLK(I2702), .RSTB(I364833), .Q(I365099) );
DFFARX1 I_21316  ( .D(I365068), .CLK(I2702), .RSTB(I364833), .Q(I364795) );
nand I_21317 (I365130,I364850,I599429);
nand I_21318 (I365147,I365130,I364884);
and I_21319 (I365164,I364966,I365147);
DFFARX1 I_21320  ( .D(I365164), .CLK(I2702), .RSTB(I364833), .Q(I364825) );
and I_21321 (I364798,I365130,I365099);
DFFARX1 I_21322  ( .D(I599456), .CLK(I2702), .RSTB(I364833), .Q(I365209) );
nor I_21323 (I364822,I365209,I365130);
nor I_21324 (I365240,I365209,I364884);
nand I_21325 (I364819,I364918,I365240);
not I_21326 (I364816,I365209);
DFFARX1 I_21327  ( .D(I599453), .CLK(I2702), .RSTB(I364833), .Q(I365285) );
not I_21328 (I365302,I365285);
nor I_21329 (I365319,I365302,I364983);
and I_21330 (I365336,I365209,I365319);
or I_21331 (I365353,I365130,I365336);
DFFARX1 I_21332  ( .D(I365353), .CLK(I2702), .RSTB(I364833), .Q(I364810) );
not I_21333 (I365384,I365302);
nor I_21334 (I365401,I365209,I365384);
nand I_21335 (I364813,I365302,I365401);
nand I_21336 (I364807,I364966,I365384);
not I_21337 (I365479,I2709);
not I_21338 (I365496,I174687);
nor I_21339 (I365513,I174708,I174690);
nand I_21340 (I365530,I365513,I174714);
nor I_21341 (I365547,I365496,I174708);
nand I_21342 (I365564,I365547,I174711);
DFFARX1 I_21343  ( .D(I365564), .CLK(I2702), .RSTB(I365479), .Q(I365581) );
not I_21344 (I365450,I365581);
not I_21345 (I365612,I174708);
not I_21346 (I365629,I365612);
not I_21347 (I365646,I174705);
nor I_21348 (I365663,I365646,I174684);
and I_21349 (I365680,I365663,I174696);
or I_21350 (I365697,I365680,I174693);
DFFARX1 I_21351  ( .D(I365697), .CLK(I2702), .RSTB(I365479), .Q(I365714) );
DFFARX1 I_21352  ( .D(I365714), .CLK(I2702), .RSTB(I365479), .Q(I365447) );
DFFARX1 I_21353  ( .D(I365714), .CLK(I2702), .RSTB(I365479), .Q(I365745) );
DFFARX1 I_21354  ( .D(I365714), .CLK(I2702), .RSTB(I365479), .Q(I365441) );
nand I_21355 (I365776,I365496,I174705);
nand I_21356 (I365793,I365776,I365530);
and I_21357 (I365810,I365612,I365793);
DFFARX1 I_21358  ( .D(I365810), .CLK(I2702), .RSTB(I365479), .Q(I365471) );
and I_21359 (I365444,I365776,I365745);
DFFARX1 I_21360  ( .D(I174699), .CLK(I2702), .RSTB(I365479), .Q(I365855) );
nor I_21361 (I365468,I365855,I365776);
nor I_21362 (I365886,I365855,I365530);
nand I_21363 (I365465,I365564,I365886);
not I_21364 (I365462,I365855);
DFFARX1 I_21365  ( .D(I174702), .CLK(I2702), .RSTB(I365479), .Q(I365931) );
not I_21366 (I365948,I365931);
nor I_21367 (I365965,I365948,I365629);
and I_21368 (I365982,I365855,I365965);
or I_21369 (I365999,I365776,I365982);
DFFARX1 I_21370  ( .D(I365999), .CLK(I2702), .RSTB(I365479), .Q(I365456) );
not I_21371 (I366030,I365948);
nor I_21372 (I366047,I365855,I366030);
nand I_21373 (I365459,I365948,I366047);
nand I_21374 (I365453,I365612,I366030);
not I_21375 (I366125,I2709);
not I_21376 (I366142,I416867);
nor I_21377 (I366159,I416876,I416861);
nand I_21378 (I366176,I366159,I416849);
nor I_21379 (I366193,I366142,I416876);
nand I_21380 (I366210,I366193,I416852);
DFFARX1 I_21381  ( .D(I366210), .CLK(I2702), .RSTB(I366125), .Q(I366227) );
not I_21382 (I366096,I366227);
not I_21383 (I366258,I416876);
not I_21384 (I366275,I366258);
not I_21385 (I366292,I416864);
nor I_21386 (I366309,I366292,I416858);
and I_21387 (I366326,I366309,I416855);
or I_21388 (I366343,I366326,I416870);
DFFARX1 I_21389  ( .D(I366343), .CLK(I2702), .RSTB(I366125), .Q(I366360) );
DFFARX1 I_21390  ( .D(I366360), .CLK(I2702), .RSTB(I366125), .Q(I366093) );
DFFARX1 I_21391  ( .D(I366360), .CLK(I2702), .RSTB(I366125), .Q(I366391) );
DFFARX1 I_21392  ( .D(I366360), .CLK(I2702), .RSTB(I366125), .Q(I366087) );
nand I_21393 (I366422,I366142,I416864);
nand I_21394 (I366439,I366422,I366176);
and I_21395 (I366456,I366258,I366439);
DFFARX1 I_21396  ( .D(I366456), .CLK(I2702), .RSTB(I366125), .Q(I366117) );
and I_21397 (I366090,I366422,I366391);
DFFARX1 I_21398  ( .D(I416879), .CLK(I2702), .RSTB(I366125), .Q(I366501) );
nor I_21399 (I366114,I366501,I366422);
nor I_21400 (I366532,I366501,I366176);
nand I_21401 (I366111,I366210,I366532);
not I_21402 (I366108,I366501);
DFFARX1 I_21403  ( .D(I416873), .CLK(I2702), .RSTB(I366125), .Q(I366577) );
not I_21404 (I366594,I366577);
nor I_21405 (I366611,I366594,I366275);
and I_21406 (I366628,I366501,I366611);
or I_21407 (I366645,I366422,I366628);
DFFARX1 I_21408  ( .D(I366645), .CLK(I2702), .RSTB(I366125), .Q(I366102) );
not I_21409 (I366676,I366594);
nor I_21410 (I366693,I366501,I366676);
nand I_21411 (I366105,I366594,I366693);
nand I_21412 (I366099,I366258,I366676);
not I_21413 (I366771,I2709);
not I_21414 (I366788,I725638);
nor I_21415 (I366805,I725623,I725629);
nand I_21416 (I366822,I366805,I725626);
nor I_21417 (I366839,I366788,I725623);
nand I_21418 (I366856,I366839,I725635);
DFFARX1 I_21419  ( .D(I366856), .CLK(I2702), .RSTB(I366771), .Q(I366873) );
not I_21420 (I366742,I366873);
not I_21421 (I366904,I725623);
not I_21422 (I366921,I366904);
not I_21423 (I366938,I725650);
nor I_21424 (I366955,I366938,I725644);
and I_21425 (I366972,I366955,I725641);
or I_21426 (I366989,I366972,I725620);
DFFARX1 I_21427  ( .D(I366989), .CLK(I2702), .RSTB(I366771), .Q(I367006) );
DFFARX1 I_21428  ( .D(I367006), .CLK(I2702), .RSTB(I366771), .Q(I366739) );
DFFARX1 I_21429  ( .D(I367006), .CLK(I2702), .RSTB(I366771), .Q(I367037) );
DFFARX1 I_21430  ( .D(I367006), .CLK(I2702), .RSTB(I366771), .Q(I366733) );
nand I_21431 (I367068,I366788,I725650);
nand I_21432 (I367085,I367068,I366822);
and I_21433 (I367102,I366904,I367085);
DFFARX1 I_21434  ( .D(I367102), .CLK(I2702), .RSTB(I366771), .Q(I366763) );
and I_21435 (I366736,I367068,I367037);
DFFARX1 I_21436  ( .D(I725647), .CLK(I2702), .RSTB(I366771), .Q(I367147) );
nor I_21437 (I366760,I367147,I367068);
nor I_21438 (I367178,I367147,I366822);
nand I_21439 (I366757,I366856,I367178);
not I_21440 (I366754,I367147);
DFFARX1 I_21441  ( .D(I725632), .CLK(I2702), .RSTB(I366771), .Q(I367223) );
not I_21442 (I367240,I367223);
nor I_21443 (I367257,I367240,I366921);
and I_21444 (I367274,I367147,I367257);
or I_21445 (I367291,I367068,I367274);
DFFARX1 I_21446  ( .D(I367291), .CLK(I2702), .RSTB(I366771), .Q(I366748) );
not I_21447 (I367322,I367240);
nor I_21448 (I367339,I367147,I367322);
nand I_21449 (I366751,I367240,I367339);
nand I_21450 (I366745,I366904,I367322);
not I_21451 (I367417,I2709);
not I_21452 (I367434,I526253);
nor I_21453 (I367451,I526265,I526259);
nand I_21454 (I367468,I367451,I526244);
nor I_21455 (I367485,I367434,I526265);
nand I_21456 (I367502,I367485,I526271);
DFFARX1 I_21457  ( .D(I367502), .CLK(I2702), .RSTB(I367417), .Q(I367519) );
not I_21458 (I367388,I367519);
not I_21459 (I367550,I526265);
not I_21460 (I367567,I367550);
not I_21461 (I367584,I526268);
nor I_21462 (I367601,I367584,I526250);
and I_21463 (I367618,I367601,I526247);
or I_21464 (I367635,I367618,I526274);
DFFARX1 I_21465  ( .D(I367635), .CLK(I2702), .RSTB(I367417), .Q(I367652) );
DFFARX1 I_21466  ( .D(I367652), .CLK(I2702), .RSTB(I367417), .Q(I367385) );
DFFARX1 I_21467  ( .D(I367652), .CLK(I2702), .RSTB(I367417), .Q(I367683) );
DFFARX1 I_21468  ( .D(I367652), .CLK(I2702), .RSTB(I367417), .Q(I367379) );
nand I_21469 (I367714,I367434,I526268);
nand I_21470 (I367731,I367714,I367468);
and I_21471 (I367748,I367550,I367731);
DFFARX1 I_21472  ( .D(I367748), .CLK(I2702), .RSTB(I367417), .Q(I367409) );
and I_21473 (I367382,I367714,I367683);
DFFARX1 I_21474  ( .D(I526262), .CLK(I2702), .RSTB(I367417), .Q(I367793) );
nor I_21475 (I367406,I367793,I367714);
nor I_21476 (I367824,I367793,I367468);
nand I_21477 (I367403,I367502,I367824);
not I_21478 (I367400,I367793);
DFFARX1 I_21479  ( .D(I526256), .CLK(I2702), .RSTB(I367417), .Q(I367869) );
not I_21480 (I367886,I367869);
nor I_21481 (I367903,I367886,I367567);
and I_21482 (I367920,I367793,I367903);
or I_21483 (I367937,I367714,I367920);
DFFARX1 I_21484  ( .D(I367937), .CLK(I2702), .RSTB(I367417), .Q(I367394) );
not I_21485 (I367968,I367886);
nor I_21486 (I367985,I367793,I367968);
nand I_21487 (I367397,I367886,I367985);
nand I_21488 (I367391,I367550,I367968);
not I_21489 (I368063,I2709);
not I_21490 (I368080,I452360);
nor I_21491 (I368097,I452363,I452345);
nand I_21492 (I368114,I368097,I452372);
nor I_21493 (I368131,I368080,I452363);
nand I_21494 (I368148,I368131,I452351);
DFFARX1 I_21495  ( .D(I368148), .CLK(I2702), .RSTB(I368063), .Q(I368165) );
not I_21496 (I368034,I368165);
not I_21497 (I368196,I452363);
not I_21498 (I368213,I368196);
not I_21499 (I368230,I452357);
nor I_21500 (I368247,I368230,I452369);
and I_21501 (I368264,I368247,I452375);
or I_21502 (I368281,I368264,I452354);
DFFARX1 I_21503  ( .D(I368281), .CLK(I2702), .RSTB(I368063), .Q(I368298) );
DFFARX1 I_21504  ( .D(I368298), .CLK(I2702), .RSTB(I368063), .Q(I368031) );
DFFARX1 I_21505  ( .D(I368298), .CLK(I2702), .RSTB(I368063), .Q(I368329) );
DFFARX1 I_21506  ( .D(I368298), .CLK(I2702), .RSTB(I368063), .Q(I368025) );
nand I_21507 (I368360,I368080,I452357);
nand I_21508 (I368377,I368360,I368114);
and I_21509 (I368394,I368196,I368377);
DFFARX1 I_21510  ( .D(I368394), .CLK(I2702), .RSTB(I368063), .Q(I368055) );
and I_21511 (I368028,I368360,I368329);
DFFARX1 I_21512  ( .D(I452366), .CLK(I2702), .RSTB(I368063), .Q(I368439) );
nor I_21513 (I368052,I368439,I368360);
nor I_21514 (I368470,I368439,I368114);
nand I_21515 (I368049,I368148,I368470);
not I_21516 (I368046,I368439);
DFFARX1 I_21517  ( .D(I452348), .CLK(I2702), .RSTB(I368063), .Q(I368515) );
not I_21518 (I368532,I368515);
nor I_21519 (I368549,I368532,I368213);
and I_21520 (I368566,I368439,I368549);
or I_21521 (I368583,I368360,I368566);
DFFARX1 I_21522  ( .D(I368583), .CLK(I2702), .RSTB(I368063), .Q(I368040) );
not I_21523 (I368614,I368532);
nor I_21524 (I368631,I368439,I368614);
nand I_21525 (I368043,I368532,I368631);
nand I_21526 (I368037,I368196,I368614);
not I_21527 (I368709,I2709);
not I_21528 (I368726,I676596);
nor I_21529 (I368743,I676593,I676578);
nand I_21530 (I368760,I368743,I676587);
nor I_21531 (I368777,I368726,I676593);
nand I_21532 (I368794,I368777,I676602);
DFFARX1 I_21533  ( .D(I368794), .CLK(I2702), .RSTB(I368709), .Q(I368811) );
not I_21534 (I368680,I368811);
not I_21535 (I368842,I676593);
not I_21536 (I368859,I368842);
not I_21537 (I368876,I676575);
nor I_21538 (I368893,I368876,I676581);
and I_21539 (I368910,I368893,I676605);
or I_21540 (I368927,I368910,I676599);
DFFARX1 I_21541  ( .D(I368927), .CLK(I2702), .RSTB(I368709), .Q(I368944) );
DFFARX1 I_21542  ( .D(I368944), .CLK(I2702), .RSTB(I368709), .Q(I368677) );
DFFARX1 I_21543  ( .D(I368944), .CLK(I2702), .RSTB(I368709), .Q(I368975) );
DFFARX1 I_21544  ( .D(I368944), .CLK(I2702), .RSTB(I368709), .Q(I368671) );
nand I_21545 (I369006,I368726,I676575);
nand I_21546 (I369023,I369006,I368760);
and I_21547 (I369040,I368842,I369023);
DFFARX1 I_21548  ( .D(I369040), .CLK(I2702), .RSTB(I368709), .Q(I368701) );
and I_21549 (I368674,I369006,I368975);
DFFARX1 I_21550  ( .D(I676584), .CLK(I2702), .RSTB(I368709), .Q(I369085) );
nor I_21551 (I368698,I369085,I369006);
nor I_21552 (I369116,I369085,I368760);
nand I_21553 (I368695,I368794,I369116);
not I_21554 (I368692,I369085);
DFFARX1 I_21555  ( .D(I676590), .CLK(I2702), .RSTB(I368709), .Q(I369161) );
not I_21556 (I369178,I369161);
nor I_21557 (I369195,I369178,I368859);
and I_21558 (I369212,I369085,I369195);
or I_21559 (I369229,I369006,I369212);
DFFARX1 I_21560  ( .D(I369229), .CLK(I2702), .RSTB(I368709), .Q(I368686) );
not I_21561 (I369260,I369178);
nor I_21562 (I369277,I369085,I369260);
nand I_21563 (I368689,I369178,I369277);
nand I_21564 (I368683,I368842,I369260);
not I_21565 (I369355,I2709);
not I_21566 (I369372,I551838);
nor I_21567 (I369389,I551850,I551844);
nand I_21568 (I369406,I369389,I551829);
nor I_21569 (I369423,I369372,I551850);
nand I_21570 (I369440,I369423,I551856);
DFFARX1 I_21571  ( .D(I369440), .CLK(I2702), .RSTB(I369355), .Q(I369457) );
not I_21572 (I369326,I369457);
not I_21573 (I369488,I551850);
not I_21574 (I369505,I369488);
not I_21575 (I369522,I551853);
nor I_21576 (I369539,I369522,I551835);
and I_21577 (I369556,I369539,I551832);
or I_21578 (I369573,I369556,I551859);
DFFARX1 I_21579  ( .D(I369573), .CLK(I2702), .RSTB(I369355), .Q(I369590) );
DFFARX1 I_21580  ( .D(I369590), .CLK(I2702), .RSTB(I369355), .Q(I369323) );
DFFARX1 I_21581  ( .D(I369590), .CLK(I2702), .RSTB(I369355), .Q(I369621) );
DFFARX1 I_21582  ( .D(I369590), .CLK(I2702), .RSTB(I369355), .Q(I369317) );
nand I_21583 (I369652,I369372,I551853);
nand I_21584 (I369669,I369652,I369406);
and I_21585 (I369686,I369488,I369669);
DFFARX1 I_21586  ( .D(I369686), .CLK(I2702), .RSTB(I369355), .Q(I369347) );
and I_21587 (I369320,I369652,I369621);
DFFARX1 I_21588  ( .D(I551847), .CLK(I2702), .RSTB(I369355), .Q(I369731) );
nor I_21589 (I369344,I369731,I369652);
nor I_21590 (I369762,I369731,I369406);
nand I_21591 (I369341,I369440,I369762);
not I_21592 (I369338,I369731);
DFFARX1 I_21593  ( .D(I551841), .CLK(I2702), .RSTB(I369355), .Q(I369807) );
not I_21594 (I369824,I369807);
nor I_21595 (I369841,I369824,I369505);
and I_21596 (I369858,I369731,I369841);
or I_21597 (I369875,I369652,I369858);
DFFARX1 I_21598  ( .D(I369875), .CLK(I2702), .RSTB(I369355), .Q(I369332) );
not I_21599 (I369906,I369824);
nor I_21600 (I369923,I369731,I369906);
nand I_21601 (I369335,I369824,I369923);
nand I_21602 (I369329,I369488,I369906);
not I_21603 (I370001,I2709);
not I_21604 (I370018,I233213);
nor I_21605 (I370035,I233201,I233204);
nand I_21606 (I370052,I370035,I233228);
nor I_21607 (I370069,I370018,I233201);
nand I_21608 (I370086,I370069,I233210);
DFFARX1 I_21609  ( .D(I370086), .CLK(I2702), .RSTB(I370001), .Q(I370103) );
not I_21610 (I369972,I370103);
not I_21611 (I370134,I233201);
not I_21612 (I370151,I370134);
not I_21613 (I370168,I233207);
nor I_21614 (I370185,I370168,I233222);
and I_21615 (I370202,I370185,I233198);
or I_21616 (I370219,I370202,I233225);
DFFARX1 I_21617  ( .D(I370219), .CLK(I2702), .RSTB(I370001), .Q(I370236) );
DFFARX1 I_21618  ( .D(I370236), .CLK(I2702), .RSTB(I370001), .Q(I369969) );
DFFARX1 I_21619  ( .D(I370236), .CLK(I2702), .RSTB(I370001), .Q(I370267) );
DFFARX1 I_21620  ( .D(I370236), .CLK(I2702), .RSTB(I370001), .Q(I369963) );
nand I_21621 (I370298,I370018,I233207);
nand I_21622 (I370315,I370298,I370052);
and I_21623 (I370332,I370134,I370315);
DFFARX1 I_21624  ( .D(I370332), .CLK(I2702), .RSTB(I370001), .Q(I369993) );
and I_21625 (I369966,I370298,I370267);
DFFARX1 I_21626  ( .D(I233216), .CLK(I2702), .RSTB(I370001), .Q(I370377) );
nor I_21627 (I369990,I370377,I370298);
nor I_21628 (I370408,I370377,I370052);
nand I_21629 (I369987,I370086,I370408);
not I_21630 (I369984,I370377);
DFFARX1 I_21631  ( .D(I233219), .CLK(I2702), .RSTB(I370001), .Q(I370453) );
not I_21632 (I370470,I370453);
nor I_21633 (I370487,I370470,I370151);
and I_21634 (I370504,I370377,I370487);
or I_21635 (I370521,I370298,I370504);
DFFARX1 I_21636  ( .D(I370521), .CLK(I2702), .RSTB(I370001), .Q(I369978) );
not I_21637 (I370552,I370470);
nor I_21638 (I370569,I370377,I370552);
nand I_21639 (I369981,I370470,I370569);
nand I_21640 (I369975,I370134,I370552);
not I_21641 (I370647,I2709);
not I_21642 (I370664,I183306);
nor I_21643 (I370681,I183327,I183309);
nand I_21644 (I370698,I370681,I183333);
nor I_21645 (I370715,I370664,I183327);
nand I_21646 (I370732,I370715,I183330);
DFFARX1 I_21647  ( .D(I370732), .CLK(I2702), .RSTB(I370647), .Q(I370749) );
not I_21648 (I370618,I370749);
not I_21649 (I370780,I183327);
not I_21650 (I370797,I370780);
not I_21651 (I370814,I183324);
nor I_21652 (I370831,I370814,I183303);
and I_21653 (I370848,I370831,I183315);
or I_21654 (I370865,I370848,I183312);
DFFARX1 I_21655  ( .D(I370865), .CLK(I2702), .RSTB(I370647), .Q(I370882) );
DFFARX1 I_21656  ( .D(I370882), .CLK(I2702), .RSTB(I370647), .Q(I370615) );
DFFARX1 I_21657  ( .D(I370882), .CLK(I2702), .RSTB(I370647), .Q(I370913) );
DFFARX1 I_21658  ( .D(I370882), .CLK(I2702), .RSTB(I370647), .Q(I370609) );
nand I_21659 (I370944,I370664,I183324);
nand I_21660 (I370961,I370944,I370698);
and I_21661 (I370978,I370780,I370961);
DFFARX1 I_21662  ( .D(I370978), .CLK(I2702), .RSTB(I370647), .Q(I370639) );
and I_21663 (I370612,I370944,I370913);
DFFARX1 I_21664  ( .D(I183318), .CLK(I2702), .RSTB(I370647), .Q(I371023) );
nor I_21665 (I370636,I371023,I370944);
nor I_21666 (I371054,I371023,I370698);
nand I_21667 (I370633,I370732,I371054);
not I_21668 (I370630,I371023);
DFFARX1 I_21669  ( .D(I183321), .CLK(I2702), .RSTB(I370647), .Q(I371099) );
not I_21670 (I371116,I371099);
nor I_21671 (I371133,I371116,I370797);
and I_21672 (I371150,I371023,I371133);
or I_21673 (I371167,I370944,I371150);
DFFARX1 I_21674  ( .D(I371167), .CLK(I2702), .RSTB(I370647), .Q(I370624) );
not I_21675 (I371198,I371116);
nor I_21676 (I371215,I371023,I371198);
nand I_21677 (I370627,I371116,I371215);
nand I_21678 (I370621,I370780,I371198);
not I_21679 (I371293,I2709);
not I_21680 (I371310,I669048);
nor I_21681 (I371327,I669045,I669030);
nand I_21682 (I371344,I371327,I669039);
nor I_21683 (I371361,I371310,I669045);
nand I_21684 (I371378,I371361,I669054);
DFFARX1 I_21685  ( .D(I371378), .CLK(I2702), .RSTB(I371293), .Q(I371395) );
not I_21686 (I371264,I371395);
not I_21687 (I371426,I669045);
not I_21688 (I371443,I371426);
not I_21689 (I371460,I669027);
nor I_21690 (I371477,I371460,I669033);
and I_21691 (I371494,I371477,I669057);
or I_21692 (I371511,I371494,I669051);
DFFARX1 I_21693  ( .D(I371511), .CLK(I2702), .RSTB(I371293), .Q(I371528) );
DFFARX1 I_21694  ( .D(I371528), .CLK(I2702), .RSTB(I371293), .Q(I371261) );
DFFARX1 I_21695  ( .D(I371528), .CLK(I2702), .RSTB(I371293), .Q(I371559) );
DFFARX1 I_21696  ( .D(I371528), .CLK(I2702), .RSTB(I371293), .Q(I371255) );
nand I_21697 (I371590,I371310,I669027);
nand I_21698 (I371607,I371590,I371344);
and I_21699 (I371624,I371426,I371607);
DFFARX1 I_21700  ( .D(I371624), .CLK(I2702), .RSTB(I371293), .Q(I371285) );
and I_21701 (I371258,I371590,I371559);
DFFARX1 I_21702  ( .D(I669036), .CLK(I2702), .RSTB(I371293), .Q(I371669) );
nor I_21703 (I371282,I371669,I371590);
nor I_21704 (I371700,I371669,I371344);
nand I_21705 (I371279,I371378,I371700);
not I_21706 (I371276,I371669);
DFFARX1 I_21707  ( .D(I669042), .CLK(I2702), .RSTB(I371293), .Q(I371745) );
not I_21708 (I371762,I371745);
nor I_21709 (I371779,I371762,I371443);
and I_21710 (I371796,I371669,I371779);
or I_21711 (I371813,I371590,I371796);
DFFARX1 I_21712  ( .D(I371813), .CLK(I2702), .RSTB(I371293), .Q(I371270) );
not I_21713 (I371844,I371762);
nor I_21714 (I371861,I371669,I371844);
nand I_21715 (I371273,I371762,I371861);
nand I_21716 (I371267,I371426,I371844);
not I_21717 (I371939,I2709);
not I_21718 (I371956,I619357);
nor I_21719 (I371973,I619354,I619339);
nand I_21720 (I371990,I371973,I619348);
nor I_21721 (I372007,I371956,I619354);
nand I_21722 (I372024,I372007,I619363);
DFFARX1 I_21723  ( .D(I372024), .CLK(I2702), .RSTB(I371939), .Q(I372041) );
not I_21724 (I371910,I372041);
not I_21725 (I372072,I619354);
not I_21726 (I372089,I372072);
not I_21727 (I372106,I619336);
nor I_21728 (I372123,I372106,I619342);
and I_21729 (I372140,I372123,I619366);
or I_21730 (I372157,I372140,I619360);
DFFARX1 I_21731  ( .D(I372157), .CLK(I2702), .RSTB(I371939), .Q(I372174) );
DFFARX1 I_21732  ( .D(I372174), .CLK(I2702), .RSTB(I371939), .Q(I371907) );
DFFARX1 I_21733  ( .D(I372174), .CLK(I2702), .RSTB(I371939), .Q(I372205) );
DFFARX1 I_21734  ( .D(I372174), .CLK(I2702), .RSTB(I371939), .Q(I371901) );
nand I_21735 (I372236,I371956,I619336);
nand I_21736 (I372253,I372236,I371990);
and I_21737 (I372270,I372072,I372253);
DFFARX1 I_21738  ( .D(I372270), .CLK(I2702), .RSTB(I371939), .Q(I371931) );
and I_21739 (I371904,I372236,I372205);
DFFARX1 I_21740  ( .D(I619345), .CLK(I2702), .RSTB(I371939), .Q(I372315) );
nor I_21741 (I371928,I372315,I372236);
nor I_21742 (I372346,I372315,I371990);
nand I_21743 (I371925,I372024,I372346);
not I_21744 (I371922,I372315);
DFFARX1 I_21745  ( .D(I619351), .CLK(I2702), .RSTB(I371939), .Q(I372391) );
not I_21746 (I372408,I372391);
nor I_21747 (I372425,I372408,I372089);
and I_21748 (I372442,I372315,I372425);
or I_21749 (I372459,I372236,I372442);
DFFARX1 I_21750  ( .D(I372459), .CLK(I2702), .RSTB(I371939), .Q(I371916) );
not I_21751 (I372490,I372408);
nor I_21752 (I372507,I372315,I372490);
nand I_21753 (I371919,I372408,I372507);
nand I_21754 (I371913,I372072,I372490);
not I_21755 (I372585,I2709);
not I_21756 (I372602,I16185);
nor I_21757 (I372619,I16200,I16194);
nand I_21758 (I372636,I372619,I16203);
nor I_21759 (I372653,I372602,I16200);
nand I_21760 (I372670,I372653,I16179);
DFFARX1 I_21761  ( .D(I372670), .CLK(I2702), .RSTB(I372585), .Q(I372687) );
not I_21762 (I372556,I372687);
not I_21763 (I372718,I16200);
not I_21764 (I372735,I372718);
not I_21765 (I372752,I16176);
nor I_21766 (I372769,I372752,I16191);
and I_21767 (I372786,I372769,I16197);
or I_21768 (I372803,I372786,I16206);
DFFARX1 I_21769  ( .D(I372803), .CLK(I2702), .RSTB(I372585), .Q(I372820) );
DFFARX1 I_21770  ( .D(I372820), .CLK(I2702), .RSTB(I372585), .Q(I372553) );
DFFARX1 I_21771  ( .D(I372820), .CLK(I2702), .RSTB(I372585), .Q(I372851) );
DFFARX1 I_21772  ( .D(I372820), .CLK(I2702), .RSTB(I372585), .Q(I372547) );
nand I_21773 (I372882,I372602,I16176);
nand I_21774 (I372899,I372882,I372636);
and I_21775 (I372916,I372718,I372899);
DFFARX1 I_21776  ( .D(I372916), .CLK(I2702), .RSTB(I372585), .Q(I372577) );
and I_21777 (I372550,I372882,I372851);
DFFARX1 I_21778  ( .D(I16188), .CLK(I2702), .RSTB(I372585), .Q(I372961) );
nor I_21779 (I372574,I372961,I372882);
nor I_21780 (I372992,I372961,I372636);
nand I_21781 (I372571,I372670,I372992);
not I_21782 (I372568,I372961);
DFFARX1 I_21783  ( .D(I16182), .CLK(I2702), .RSTB(I372585), .Q(I373037) );
not I_21784 (I373054,I373037);
nor I_21785 (I373071,I373054,I372735);
and I_21786 (I373088,I372961,I373071);
or I_21787 (I373105,I372882,I373088);
DFFARX1 I_21788  ( .D(I373105), .CLK(I2702), .RSTB(I372585), .Q(I372562) );
not I_21789 (I373136,I373054);
nor I_21790 (I373153,I372961,I373136);
nand I_21791 (I372565,I373054,I373153);
nand I_21792 (I372559,I372718,I373136);
not I_21793 (I373231,I2709);
not I_21794 (I373248,I588142);
nor I_21795 (I373265,I588130,I588139);
nand I_21796 (I373282,I373265,I588154);
nor I_21797 (I373299,I373248,I588130);
nand I_21798 (I373316,I373299,I588136);
DFFARX1 I_21799  ( .D(I373316), .CLK(I2702), .RSTB(I373231), .Q(I373333) );
not I_21800 (I373202,I373333);
not I_21801 (I373364,I588130);
not I_21802 (I373381,I373364);
not I_21803 (I373398,I588124);
nor I_21804 (I373415,I373398,I588145);
and I_21805 (I373432,I373415,I588127);
or I_21806 (I373449,I373432,I588133);
DFFARX1 I_21807  ( .D(I373449), .CLK(I2702), .RSTB(I373231), .Q(I373466) );
DFFARX1 I_21808  ( .D(I373466), .CLK(I2702), .RSTB(I373231), .Q(I373199) );
DFFARX1 I_21809  ( .D(I373466), .CLK(I2702), .RSTB(I373231), .Q(I373497) );
DFFARX1 I_21810  ( .D(I373466), .CLK(I2702), .RSTB(I373231), .Q(I373193) );
nand I_21811 (I373528,I373248,I588124);
nand I_21812 (I373545,I373528,I373282);
and I_21813 (I373562,I373364,I373545);
DFFARX1 I_21814  ( .D(I373562), .CLK(I2702), .RSTB(I373231), .Q(I373223) );
and I_21815 (I373196,I373528,I373497);
DFFARX1 I_21816  ( .D(I588151), .CLK(I2702), .RSTB(I373231), .Q(I373607) );
nor I_21817 (I373220,I373607,I373528);
nor I_21818 (I373638,I373607,I373282);
nand I_21819 (I373217,I373316,I373638);
not I_21820 (I373214,I373607);
DFFARX1 I_21821  ( .D(I588148), .CLK(I2702), .RSTB(I373231), .Q(I373683) );
not I_21822 (I373700,I373683);
nor I_21823 (I373717,I373700,I373381);
and I_21824 (I373734,I373607,I373717);
or I_21825 (I373751,I373528,I373734);
DFFARX1 I_21826  ( .D(I373751), .CLK(I2702), .RSTB(I373231), .Q(I373208) );
not I_21827 (I373782,I373700);
nor I_21828 (I373799,I373607,I373782);
nand I_21829 (I373211,I373700,I373799);
nand I_21830 (I373205,I373364,I373782);
not I_21831 (I373877,I2709);
not I_21832 (I373894,I578027);
nor I_21833 (I373911,I578015,I578024);
nand I_21834 (I373928,I373911,I578039);
nor I_21835 (I373945,I373894,I578015);
nand I_21836 (I373962,I373945,I578021);
DFFARX1 I_21837  ( .D(I373962), .CLK(I2702), .RSTB(I373877), .Q(I373979) );
not I_21838 (I373848,I373979);
not I_21839 (I374010,I578015);
not I_21840 (I374027,I374010);
not I_21841 (I374044,I578009);
nor I_21842 (I374061,I374044,I578030);
and I_21843 (I374078,I374061,I578012);
or I_21844 (I374095,I374078,I578018);
DFFARX1 I_21845  ( .D(I374095), .CLK(I2702), .RSTB(I373877), .Q(I374112) );
DFFARX1 I_21846  ( .D(I374112), .CLK(I2702), .RSTB(I373877), .Q(I373845) );
DFFARX1 I_21847  ( .D(I374112), .CLK(I2702), .RSTB(I373877), .Q(I374143) );
DFFARX1 I_21848  ( .D(I374112), .CLK(I2702), .RSTB(I373877), .Q(I373839) );
nand I_21849 (I374174,I373894,I578009);
nand I_21850 (I374191,I374174,I373928);
and I_21851 (I374208,I374010,I374191);
DFFARX1 I_21852  ( .D(I374208), .CLK(I2702), .RSTB(I373877), .Q(I373869) );
and I_21853 (I373842,I374174,I374143);
DFFARX1 I_21854  ( .D(I578036), .CLK(I2702), .RSTB(I373877), .Q(I374253) );
nor I_21855 (I373866,I374253,I374174);
nor I_21856 (I374284,I374253,I373928);
nand I_21857 (I373863,I373962,I374284);
not I_21858 (I373860,I374253);
DFFARX1 I_21859  ( .D(I578033), .CLK(I2702), .RSTB(I373877), .Q(I374329) );
not I_21860 (I374346,I374329);
nor I_21861 (I374363,I374346,I374027);
and I_21862 (I374380,I374253,I374363);
or I_21863 (I374397,I374174,I374380);
DFFARX1 I_21864  ( .D(I374397), .CLK(I2702), .RSTB(I373877), .Q(I373854) );
not I_21865 (I374428,I374346);
nor I_21866 (I374445,I374253,I374428);
nand I_21867 (I373857,I374346,I374445);
nand I_21868 (I373851,I374010,I374428);
not I_21869 (I374523,I2709);
not I_21870 (I374540,I176013);
nor I_21871 (I374557,I176034,I176016);
nand I_21872 (I374574,I374557,I176040);
nor I_21873 (I374591,I374540,I176034);
nand I_21874 (I374608,I374591,I176037);
DFFARX1 I_21875  ( .D(I374608), .CLK(I2702), .RSTB(I374523), .Q(I374625) );
not I_21876 (I374494,I374625);
not I_21877 (I374656,I176034);
not I_21878 (I374673,I374656);
not I_21879 (I374690,I176031);
nor I_21880 (I374707,I374690,I176010);
and I_21881 (I374724,I374707,I176022);
or I_21882 (I374741,I374724,I176019);
DFFARX1 I_21883  ( .D(I374741), .CLK(I2702), .RSTB(I374523), .Q(I374758) );
DFFARX1 I_21884  ( .D(I374758), .CLK(I2702), .RSTB(I374523), .Q(I374491) );
DFFARX1 I_21885  ( .D(I374758), .CLK(I2702), .RSTB(I374523), .Q(I374789) );
DFFARX1 I_21886  ( .D(I374758), .CLK(I2702), .RSTB(I374523), .Q(I374485) );
nand I_21887 (I374820,I374540,I176031);
nand I_21888 (I374837,I374820,I374574);
and I_21889 (I374854,I374656,I374837);
DFFARX1 I_21890  ( .D(I374854), .CLK(I2702), .RSTB(I374523), .Q(I374515) );
and I_21891 (I374488,I374820,I374789);
DFFARX1 I_21892  ( .D(I176025), .CLK(I2702), .RSTB(I374523), .Q(I374899) );
nor I_21893 (I374512,I374899,I374820);
nor I_21894 (I374930,I374899,I374574);
nand I_21895 (I374509,I374608,I374930);
not I_21896 (I374506,I374899);
DFFARX1 I_21897  ( .D(I176028), .CLK(I2702), .RSTB(I374523), .Q(I374975) );
not I_21898 (I374992,I374975);
nor I_21899 (I375009,I374992,I374673);
and I_21900 (I375026,I374899,I375009);
or I_21901 (I375043,I374820,I375026);
DFFARX1 I_21902  ( .D(I375043), .CLK(I2702), .RSTB(I374523), .Q(I374500) );
not I_21903 (I375074,I374992);
nor I_21904 (I375091,I374899,I375074);
nand I_21905 (I374503,I374992,I375091);
nand I_21906 (I374497,I374656,I375074);
not I_21907 (I375169,I2709);
not I_21908 (I375186,I124708);
nor I_21909 (I375203,I124699,I124690);
nand I_21910 (I375220,I375203,I124705);
nor I_21911 (I375237,I375186,I124699);
nand I_21912 (I375254,I375237,I124702);
DFFARX1 I_21913  ( .D(I375254), .CLK(I2702), .RSTB(I375169), .Q(I375271) );
not I_21914 (I375140,I375271);
not I_21915 (I375302,I124699);
not I_21916 (I375319,I375302);
not I_21917 (I375336,I124711);
nor I_21918 (I375353,I375336,I124696);
and I_21919 (I375370,I375353,I124714);
or I_21920 (I375387,I375370,I124687);
DFFARX1 I_21921  ( .D(I375387), .CLK(I2702), .RSTB(I375169), .Q(I375404) );
DFFARX1 I_21922  ( .D(I375404), .CLK(I2702), .RSTB(I375169), .Q(I375137) );
DFFARX1 I_21923  ( .D(I375404), .CLK(I2702), .RSTB(I375169), .Q(I375435) );
DFFARX1 I_21924  ( .D(I375404), .CLK(I2702), .RSTB(I375169), .Q(I375131) );
nand I_21925 (I375466,I375186,I124711);
nand I_21926 (I375483,I375466,I375220);
and I_21927 (I375500,I375302,I375483);
DFFARX1 I_21928  ( .D(I375500), .CLK(I2702), .RSTB(I375169), .Q(I375161) );
and I_21929 (I375134,I375466,I375435);
DFFARX1 I_21930  ( .D(I124717), .CLK(I2702), .RSTB(I375169), .Q(I375545) );
nor I_21931 (I375158,I375545,I375466);
nor I_21932 (I375576,I375545,I375220);
nand I_21933 (I375155,I375254,I375576);
not I_21934 (I375152,I375545);
DFFARX1 I_21935  ( .D(I124693), .CLK(I2702), .RSTB(I375169), .Q(I375621) );
not I_21936 (I375638,I375621);
nor I_21937 (I375655,I375638,I375319);
and I_21938 (I375672,I375545,I375655);
or I_21939 (I375689,I375466,I375672);
DFFARX1 I_21940  ( .D(I375689), .CLK(I2702), .RSTB(I375169), .Q(I375146) );
not I_21941 (I375720,I375638);
nor I_21942 (I375737,I375545,I375720);
nand I_21943 (I375149,I375638,I375737);
nand I_21944 (I375143,I375302,I375720);
not I_21945 (I375815,I2709);
not I_21946 (I375832,I185958);
nor I_21947 (I375849,I185979,I185961);
nand I_21948 (I375866,I375849,I185985);
nor I_21949 (I375883,I375832,I185979);
nand I_21950 (I375900,I375883,I185982);
DFFARX1 I_21951  ( .D(I375900), .CLK(I2702), .RSTB(I375815), .Q(I375917) );
not I_21952 (I375786,I375917);
not I_21953 (I375948,I185979);
not I_21954 (I375965,I375948);
not I_21955 (I375982,I185976);
nor I_21956 (I375999,I375982,I185955);
and I_21957 (I376016,I375999,I185967);
or I_21958 (I376033,I376016,I185964);
DFFARX1 I_21959  ( .D(I376033), .CLK(I2702), .RSTB(I375815), .Q(I376050) );
DFFARX1 I_21960  ( .D(I376050), .CLK(I2702), .RSTB(I375815), .Q(I375783) );
DFFARX1 I_21961  ( .D(I376050), .CLK(I2702), .RSTB(I375815), .Q(I376081) );
DFFARX1 I_21962  ( .D(I376050), .CLK(I2702), .RSTB(I375815), .Q(I375777) );
nand I_21963 (I376112,I375832,I185976);
nand I_21964 (I376129,I376112,I375866);
and I_21965 (I376146,I375948,I376129);
DFFARX1 I_21966  ( .D(I376146), .CLK(I2702), .RSTB(I375815), .Q(I375807) );
and I_21967 (I375780,I376112,I376081);
DFFARX1 I_21968  ( .D(I185970), .CLK(I2702), .RSTB(I375815), .Q(I376191) );
nor I_21969 (I375804,I376191,I376112);
nor I_21970 (I376222,I376191,I375866);
nand I_21971 (I375801,I375900,I376222);
not I_21972 (I375798,I376191);
DFFARX1 I_21973  ( .D(I185973), .CLK(I2702), .RSTB(I375815), .Q(I376267) );
not I_21974 (I376284,I376267);
nor I_21975 (I376301,I376284,I375965);
and I_21976 (I376318,I376191,I376301);
or I_21977 (I376335,I376112,I376318);
DFFARX1 I_21978  ( .D(I376335), .CLK(I2702), .RSTB(I375815), .Q(I375792) );
not I_21979 (I376366,I376284);
nor I_21980 (I376383,I376191,I376366);
nand I_21981 (I375795,I376284,I376383);
nand I_21982 (I375789,I375948,I376366);
not I_21983 (I376461,I2709);
not I_21984 (I376478,I95638);
nor I_21985 (I376495,I95629,I95620);
nand I_21986 (I376512,I376495,I95635);
nor I_21987 (I376529,I376478,I95629);
nand I_21988 (I376546,I376529,I95632);
DFFARX1 I_21989  ( .D(I376546), .CLK(I2702), .RSTB(I376461), .Q(I376563) );
not I_21990 (I376432,I376563);
not I_21991 (I376594,I95629);
not I_21992 (I376611,I376594);
not I_21993 (I376628,I95641);
nor I_21994 (I376645,I376628,I95626);
and I_21995 (I376662,I376645,I95644);
or I_21996 (I376679,I376662,I95617);
DFFARX1 I_21997  ( .D(I376679), .CLK(I2702), .RSTB(I376461), .Q(I376696) );
DFFARX1 I_21998  ( .D(I376696), .CLK(I2702), .RSTB(I376461), .Q(I376429) );
DFFARX1 I_21999  ( .D(I376696), .CLK(I2702), .RSTB(I376461), .Q(I376727) );
DFFARX1 I_22000  ( .D(I376696), .CLK(I2702), .RSTB(I376461), .Q(I376423) );
nand I_22001 (I376758,I376478,I95641);
nand I_22002 (I376775,I376758,I376512);
and I_22003 (I376792,I376594,I376775);
DFFARX1 I_22004  ( .D(I376792), .CLK(I2702), .RSTB(I376461), .Q(I376453) );
and I_22005 (I376426,I376758,I376727);
DFFARX1 I_22006  ( .D(I95647), .CLK(I2702), .RSTB(I376461), .Q(I376837) );
nor I_22007 (I376450,I376837,I376758);
nor I_22008 (I376868,I376837,I376512);
nand I_22009 (I376447,I376546,I376868);
not I_22010 (I376444,I376837);
DFFARX1 I_22011  ( .D(I95623), .CLK(I2702), .RSTB(I376461), .Q(I376913) );
not I_22012 (I376930,I376913);
nor I_22013 (I376947,I376930,I376611);
and I_22014 (I376964,I376837,I376947);
or I_22015 (I376981,I376758,I376964);
DFFARX1 I_22016  ( .D(I376981), .CLK(I2702), .RSTB(I376461), .Q(I376438) );
not I_22017 (I377012,I376930);
nor I_22018 (I377029,I376837,I377012);
nand I_22019 (I376441,I376930,I377029);
nand I_22020 (I376435,I376594,I377012);
not I_22021 (I377107,I2709);
not I_22022 (I377124,I697894);
nor I_22023 (I377141,I697879,I697885);
nand I_22024 (I377158,I377141,I697882);
nor I_22025 (I377175,I377124,I697879);
nand I_22026 (I377192,I377175,I697891);
DFFARX1 I_22027  ( .D(I377192), .CLK(I2702), .RSTB(I377107), .Q(I377209) );
not I_22028 (I377078,I377209);
not I_22029 (I377240,I697879);
not I_22030 (I377257,I377240);
not I_22031 (I377274,I697906);
nor I_22032 (I377291,I377274,I697900);
and I_22033 (I377308,I377291,I697897);
or I_22034 (I377325,I377308,I697876);
DFFARX1 I_22035  ( .D(I377325), .CLK(I2702), .RSTB(I377107), .Q(I377342) );
DFFARX1 I_22036  ( .D(I377342), .CLK(I2702), .RSTB(I377107), .Q(I377075) );
DFFARX1 I_22037  ( .D(I377342), .CLK(I2702), .RSTB(I377107), .Q(I377373) );
DFFARX1 I_22038  ( .D(I377342), .CLK(I2702), .RSTB(I377107), .Q(I377069) );
nand I_22039 (I377404,I377124,I697906);
nand I_22040 (I377421,I377404,I377158);
and I_22041 (I377438,I377240,I377421);
DFFARX1 I_22042  ( .D(I377438), .CLK(I2702), .RSTB(I377107), .Q(I377099) );
and I_22043 (I377072,I377404,I377373);
DFFARX1 I_22044  ( .D(I697903), .CLK(I2702), .RSTB(I377107), .Q(I377483) );
nor I_22045 (I377096,I377483,I377404);
nor I_22046 (I377514,I377483,I377158);
nand I_22047 (I377093,I377192,I377514);
not I_22048 (I377090,I377483);
DFFARX1 I_22049  ( .D(I697888), .CLK(I2702), .RSTB(I377107), .Q(I377559) );
not I_22050 (I377576,I377559);
nor I_22051 (I377593,I377576,I377257);
and I_22052 (I377610,I377483,I377593);
or I_22053 (I377627,I377404,I377610);
DFFARX1 I_22054  ( .D(I377627), .CLK(I2702), .RSTB(I377107), .Q(I377084) );
not I_22055 (I377658,I377576);
nor I_22056 (I377675,I377483,I377658);
nand I_22057 (I377087,I377576,I377675);
nand I_22058 (I377081,I377240,I377658);
not I_22059 (I377753,I2709);
not I_22060 (I377770,I269517);
nor I_22061 (I377787,I269496,I269508);
nand I_22062 (I377804,I377787,I269511);
nor I_22063 (I377821,I377770,I269496);
nand I_22064 (I377838,I377821,I269493);
DFFARX1 I_22065  ( .D(I377838), .CLK(I2702), .RSTB(I377753), .Q(I377855) );
not I_22066 (I377724,I377855);
not I_22067 (I377886,I269496);
not I_22068 (I377903,I377886);
not I_22069 (I377920,I269514);
nor I_22070 (I377937,I377920,I269505);
and I_22071 (I377954,I377937,I269499);
or I_22072 (I377971,I377954,I269523);
DFFARX1 I_22073  ( .D(I377971), .CLK(I2702), .RSTB(I377753), .Q(I377988) );
DFFARX1 I_22074  ( .D(I377988), .CLK(I2702), .RSTB(I377753), .Q(I377721) );
DFFARX1 I_22075  ( .D(I377988), .CLK(I2702), .RSTB(I377753), .Q(I378019) );
DFFARX1 I_22076  ( .D(I377988), .CLK(I2702), .RSTB(I377753), .Q(I377715) );
nand I_22077 (I378050,I377770,I269514);
nand I_22078 (I378067,I378050,I377804);
and I_22079 (I378084,I377886,I378067);
DFFARX1 I_22080  ( .D(I378084), .CLK(I2702), .RSTB(I377753), .Q(I377745) );
and I_22081 (I377718,I378050,I378019);
DFFARX1 I_22082  ( .D(I269520), .CLK(I2702), .RSTB(I377753), .Q(I378129) );
nor I_22083 (I377742,I378129,I378050);
nor I_22084 (I378160,I378129,I377804);
nand I_22085 (I377739,I377838,I378160);
not I_22086 (I377736,I378129);
DFFARX1 I_22087  ( .D(I269502), .CLK(I2702), .RSTB(I377753), .Q(I378205) );
not I_22088 (I378222,I378205);
nor I_22089 (I378239,I378222,I377903);
and I_22090 (I378256,I378129,I378239);
or I_22091 (I378273,I378050,I378256);
DFFARX1 I_22092  ( .D(I378273), .CLK(I2702), .RSTB(I377753), .Q(I377730) );
not I_22093 (I378304,I378222);
nor I_22094 (I378321,I378129,I378304);
nand I_22095 (I377733,I378222,I378321);
nand I_22096 (I377727,I377886,I378304);
not I_22097 (I378399,I2709);
not I_22098 (I378416,I441378);
nor I_22099 (I378433,I441381,I441363);
nand I_22100 (I378450,I378433,I441390);
nor I_22101 (I378467,I378416,I441381);
nand I_22102 (I378484,I378467,I441369);
DFFARX1 I_22103  ( .D(I378484), .CLK(I2702), .RSTB(I378399), .Q(I378501) );
not I_22104 (I378370,I378501);
not I_22105 (I378532,I441381);
not I_22106 (I378549,I378532);
not I_22107 (I378566,I441375);
nor I_22108 (I378583,I378566,I441387);
and I_22109 (I378600,I378583,I441393);
or I_22110 (I378617,I378600,I441372);
DFFARX1 I_22111  ( .D(I378617), .CLK(I2702), .RSTB(I378399), .Q(I378634) );
DFFARX1 I_22112  ( .D(I378634), .CLK(I2702), .RSTB(I378399), .Q(I378367) );
DFFARX1 I_22113  ( .D(I378634), .CLK(I2702), .RSTB(I378399), .Q(I378665) );
DFFARX1 I_22114  ( .D(I378634), .CLK(I2702), .RSTB(I378399), .Q(I378361) );
nand I_22115 (I378696,I378416,I441375);
nand I_22116 (I378713,I378696,I378450);
and I_22117 (I378730,I378532,I378713);
DFFARX1 I_22118  ( .D(I378730), .CLK(I2702), .RSTB(I378399), .Q(I378391) );
and I_22119 (I378364,I378696,I378665);
DFFARX1 I_22120  ( .D(I441384), .CLK(I2702), .RSTB(I378399), .Q(I378775) );
nor I_22121 (I378388,I378775,I378696);
nor I_22122 (I378806,I378775,I378450);
nand I_22123 (I378385,I378484,I378806);
not I_22124 (I378382,I378775);
DFFARX1 I_22125  ( .D(I441366), .CLK(I2702), .RSTB(I378399), .Q(I378851) );
not I_22126 (I378868,I378851);
nor I_22127 (I378885,I378868,I378549);
and I_22128 (I378902,I378775,I378885);
or I_22129 (I378919,I378696,I378902);
DFFARX1 I_22130  ( .D(I378919), .CLK(I2702), .RSTB(I378399), .Q(I378376) );
not I_22131 (I378950,I378868);
nor I_22132 (I378967,I378775,I378950);
nand I_22133 (I378379,I378868,I378967);
nand I_22134 (I378373,I378532,I378950);
not I_22135 (I379045,I2709);
not I_22136 (I379062,I9453);
nor I_22137 (I379079,I9468,I9462);
nand I_22138 (I379096,I379079,I9471);
nor I_22139 (I379113,I379062,I9468);
nand I_22140 (I379130,I379113,I9447);
DFFARX1 I_22141  ( .D(I379130), .CLK(I2702), .RSTB(I379045), .Q(I379147) );
not I_22142 (I379016,I379147);
not I_22143 (I379178,I9468);
not I_22144 (I379195,I379178);
not I_22145 (I379212,I9444);
nor I_22146 (I379229,I379212,I9459);
and I_22147 (I379246,I379229,I9465);
or I_22148 (I379263,I379246,I9474);
DFFARX1 I_22149  ( .D(I379263), .CLK(I2702), .RSTB(I379045), .Q(I379280) );
DFFARX1 I_22150  ( .D(I379280), .CLK(I2702), .RSTB(I379045), .Q(I379013) );
DFFARX1 I_22151  ( .D(I379280), .CLK(I2702), .RSTB(I379045), .Q(I379311) );
DFFARX1 I_22152  ( .D(I379280), .CLK(I2702), .RSTB(I379045), .Q(I379007) );
nand I_22153 (I379342,I379062,I9444);
nand I_22154 (I379359,I379342,I379096);
and I_22155 (I379376,I379178,I379359);
DFFARX1 I_22156  ( .D(I379376), .CLK(I2702), .RSTB(I379045), .Q(I379037) );
and I_22157 (I379010,I379342,I379311);
DFFARX1 I_22158  ( .D(I9456), .CLK(I2702), .RSTB(I379045), .Q(I379421) );
nor I_22159 (I379034,I379421,I379342);
nor I_22160 (I379452,I379421,I379096);
nand I_22161 (I379031,I379130,I379452);
not I_22162 (I379028,I379421);
DFFARX1 I_22163  ( .D(I9450), .CLK(I2702), .RSTB(I379045), .Q(I379497) );
not I_22164 (I379514,I379497);
nor I_22165 (I379531,I379514,I379195);
and I_22166 (I379548,I379421,I379531);
or I_22167 (I379565,I379342,I379548);
DFFARX1 I_22168  ( .D(I379565), .CLK(I2702), .RSTB(I379045), .Q(I379022) );
not I_22169 (I379596,I379514);
nor I_22170 (I379613,I379421,I379596);
nand I_22171 (I379025,I379514,I379613);
nand I_22172 (I379019,I379178,I379596);
not I_22173 (I379691,I2709);
not I_22174 (I379708,I653952);
nor I_22175 (I379725,I653949,I653934);
nand I_22176 (I379742,I379725,I653943);
nor I_22177 (I379759,I379708,I653949);
nand I_22178 (I379776,I379759,I653958);
DFFARX1 I_22179  ( .D(I379776), .CLK(I2702), .RSTB(I379691), .Q(I379793) );
not I_22180 (I379662,I379793);
not I_22181 (I379824,I653949);
not I_22182 (I379841,I379824);
not I_22183 (I379858,I653931);
nor I_22184 (I379875,I379858,I653937);
and I_22185 (I379892,I379875,I653961);
or I_22186 (I379909,I379892,I653955);
DFFARX1 I_22187  ( .D(I379909), .CLK(I2702), .RSTB(I379691), .Q(I379926) );
DFFARX1 I_22188  ( .D(I379926), .CLK(I2702), .RSTB(I379691), .Q(I379659) );
DFFARX1 I_22189  ( .D(I379926), .CLK(I2702), .RSTB(I379691), .Q(I379957) );
DFFARX1 I_22190  ( .D(I379926), .CLK(I2702), .RSTB(I379691), .Q(I379653) );
nand I_22191 (I379988,I379708,I653931);
nand I_22192 (I380005,I379988,I379742);
and I_22193 (I380022,I379824,I380005);
DFFARX1 I_22194  ( .D(I380022), .CLK(I2702), .RSTB(I379691), .Q(I379683) );
and I_22195 (I379656,I379988,I379957);
DFFARX1 I_22196  ( .D(I653940), .CLK(I2702), .RSTB(I379691), .Q(I380067) );
nor I_22197 (I379680,I380067,I379988);
nor I_22198 (I380098,I380067,I379742);
nand I_22199 (I379677,I379776,I380098);
not I_22200 (I379674,I380067);
DFFARX1 I_22201  ( .D(I653946), .CLK(I2702), .RSTB(I379691), .Q(I380143) );
not I_22202 (I380160,I380143);
nor I_22203 (I380177,I380160,I379841);
and I_22204 (I380194,I380067,I380177);
or I_22205 (I380211,I379988,I380194);
DFFARX1 I_22206  ( .D(I380211), .CLK(I2702), .RSTB(I379691), .Q(I379668) );
not I_22207 (I380242,I380160);
nor I_22208 (I380259,I380067,I380242);
nand I_22209 (I379671,I380160,I380259);
nand I_22210 (I379665,I379824,I380242);
not I_22211 (I380337,I2709);
not I_22212 (I380354,I50418);
nor I_22213 (I380371,I50409,I50400);
nand I_22214 (I380388,I380371,I50415);
nor I_22215 (I380405,I380354,I50409);
nand I_22216 (I380422,I380405,I50412);
DFFARX1 I_22217  ( .D(I380422), .CLK(I2702), .RSTB(I380337), .Q(I380439) );
not I_22218 (I380308,I380439);
not I_22219 (I380470,I50409);
not I_22220 (I380487,I380470);
not I_22221 (I380504,I50421);
nor I_22222 (I380521,I380504,I50406);
and I_22223 (I380538,I380521,I50424);
or I_22224 (I380555,I380538,I50397);
DFFARX1 I_22225  ( .D(I380555), .CLK(I2702), .RSTB(I380337), .Q(I380572) );
DFFARX1 I_22226  ( .D(I380572), .CLK(I2702), .RSTB(I380337), .Q(I380305) );
DFFARX1 I_22227  ( .D(I380572), .CLK(I2702), .RSTB(I380337), .Q(I380603) );
DFFARX1 I_22228  ( .D(I380572), .CLK(I2702), .RSTB(I380337), .Q(I380299) );
nand I_22229 (I380634,I380354,I50421);
nand I_22230 (I380651,I380634,I380388);
and I_22231 (I380668,I380470,I380651);
DFFARX1 I_22232  ( .D(I380668), .CLK(I2702), .RSTB(I380337), .Q(I380329) );
and I_22233 (I380302,I380634,I380603);
DFFARX1 I_22234  ( .D(I50427), .CLK(I2702), .RSTB(I380337), .Q(I380713) );
nor I_22235 (I380326,I380713,I380634);
nor I_22236 (I380744,I380713,I380388);
nand I_22237 (I380323,I380422,I380744);
not I_22238 (I380320,I380713);
DFFARX1 I_22239  ( .D(I50403), .CLK(I2702), .RSTB(I380337), .Q(I380789) );
not I_22240 (I380806,I380789);
nor I_22241 (I380823,I380806,I380487);
and I_22242 (I380840,I380713,I380823);
or I_22243 (I380857,I380634,I380840);
DFFARX1 I_22244  ( .D(I380857), .CLK(I2702), .RSTB(I380337), .Q(I380314) );
not I_22245 (I380888,I380806);
nor I_22246 (I380905,I380713,I380888);
nand I_22247 (I380317,I380806,I380905);
nand I_22248 (I380311,I380470,I380888);
not I_22249 (I380983,I2709);
not I_22250 (I381000,I33576);
nor I_22251 (I381017,I33591,I33585);
nand I_22252 (I381034,I381017,I33594);
nor I_22253 (I381051,I381000,I33591);
nand I_22254 (I381068,I381051,I33570);
DFFARX1 I_22255  ( .D(I381068), .CLK(I2702), .RSTB(I380983), .Q(I381085) );
not I_22256 (I380954,I381085);
not I_22257 (I381116,I33591);
not I_22258 (I381133,I381116);
not I_22259 (I381150,I33567);
nor I_22260 (I381167,I381150,I33582);
and I_22261 (I381184,I381167,I33588);
or I_22262 (I381201,I381184,I33597);
DFFARX1 I_22263  ( .D(I381201), .CLK(I2702), .RSTB(I380983), .Q(I381218) );
DFFARX1 I_22264  ( .D(I381218), .CLK(I2702), .RSTB(I380983), .Q(I380951) );
DFFARX1 I_22265  ( .D(I381218), .CLK(I2702), .RSTB(I380983), .Q(I381249) );
DFFARX1 I_22266  ( .D(I381218), .CLK(I2702), .RSTB(I380983), .Q(I380945) );
nand I_22267 (I381280,I381000,I33567);
nand I_22268 (I381297,I381280,I381034);
and I_22269 (I381314,I381116,I381297);
DFFARX1 I_22270  ( .D(I381314), .CLK(I2702), .RSTB(I380983), .Q(I380975) );
and I_22271 (I380948,I381280,I381249);
DFFARX1 I_22272  ( .D(I33579), .CLK(I2702), .RSTB(I380983), .Q(I381359) );
nor I_22273 (I380972,I381359,I381280);
nor I_22274 (I381390,I381359,I381034);
nand I_22275 (I380969,I381068,I381390);
not I_22276 (I380966,I381359);
DFFARX1 I_22277  ( .D(I33573), .CLK(I2702), .RSTB(I380983), .Q(I381435) );
not I_22278 (I381452,I381435);
nor I_22279 (I381469,I381452,I381133);
and I_22280 (I381486,I381359,I381469);
or I_22281 (I381503,I381280,I381486);
DFFARX1 I_22282  ( .D(I381503), .CLK(I2702), .RSTB(I380983), .Q(I380960) );
not I_22283 (I381534,I381452);
nor I_22284 (I381551,I381359,I381534);
nand I_22285 (I380963,I381452,I381551);
nand I_22286 (I380957,I381116,I381534);
not I_22287 (I381629,I2709);
not I_22288 (I381646,I414419);
nor I_22289 (I381663,I414428,I414413);
nand I_22290 (I381680,I381663,I414401);
nor I_22291 (I381697,I381646,I414428);
nand I_22292 (I381714,I381697,I414404);
DFFARX1 I_22293  ( .D(I381714), .CLK(I2702), .RSTB(I381629), .Q(I381731) );
not I_22294 (I381600,I381731);
not I_22295 (I381762,I414428);
not I_22296 (I381779,I381762);
not I_22297 (I381796,I414416);
nor I_22298 (I381813,I381796,I414410);
and I_22299 (I381830,I381813,I414407);
or I_22300 (I381847,I381830,I414422);
DFFARX1 I_22301  ( .D(I381847), .CLK(I2702), .RSTB(I381629), .Q(I381864) );
DFFARX1 I_22302  ( .D(I381864), .CLK(I2702), .RSTB(I381629), .Q(I381597) );
DFFARX1 I_22303  ( .D(I381864), .CLK(I2702), .RSTB(I381629), .Q(I381895) );
DFFARX1 I_22304  ( .D(I381864), .CLK(I2702), .RSTB(I381629), .Q(I381591) );
nand I_22305 (I381926,I381646,I414416);
nand I_22306 (I381943,I381926,I381680);
and I_22307 (I381960,I381762,I381943);
DFFARX1 I_22308  ( .D(I381960), .CLK(I2702), .RSTB(I381629), .Q(I381621) );
and I_22309 (I381594,I381926,I381895);
DFFARX1 I_22310  ( .D(I414431), .CLK(I2702), .RSTB(I381629), .Q(I382005) );
nor I_22311 (I381618,I382005,I381926);
nor I_22312 (I382036,I382005,I381680);
nand I_22313 (I381615,I381714,I382036);
not I_22314 (I381612,I382005);
DFFARX1 I_22315  ( .D(I414425), .CLK(I2702), .RSTB(I381629), .Q(I382081) );
not I_22316 (I382098,I382081);
nor I_22317 (I382115,I382098,I381779);
and I_22318 (I382132,I382005,I382115);
or I_22319 (I382149,I381926,I382132);
DFFARX1 I_22320  ( .D(I382149), .CLK(I2702), .RSTB(I381629), .Q(I381606) );
not I_22321 (I382180,I382098);
nor I_22322 (I382197,I382005,I382180);
nand I_22323 (I381609,I382098,I382197);
nand I_22324 (I381603,I381762,I382180);
not I_22325 (I382275,I2709);
not I_22326 (I382292,I11697);
nor I_22327 (I382309,I11712,I11706);
nand I_22328 (I382326,I382309,I11715);
nor I_22329 (I382343,I382292,I11712);
nand I_22330 (I382360,I382343,I11691);
DFFARX1 I_22331  ( .D(I382360), .CLK(I2702), .RSTB(I382275), .Q(I382377) );
not I_22332 (I382246,I382377);
not I_22333 (I382408,I11712);
not I_22334 (I382425,I382408);
not I_22335 (I382442,I11688);
nor I_22336 (I382459,I382442,I11703);
and I_22337 (I382476,I382459,I11709);
or I_22338 (I382493,I382476,I11718);
DFFARX1 I_22339  ( .D(I382493), .CLK(I2702), .RSTB(I382275), .Q(I382510) );
DFFARX1 I_22340  ( .D(I382510), .CLK(I2702), .RSTB(I382275), .Q(I382243) );
DFFARX1 I_22341  ( .D(I382510), .CLK(I2702), .RSTB(I382275), .Q(I382541) );
DFFARX1 I_22342  ( .D(I382510), .CLK(I2702), .RSTB(I382275), .Q(I382237) );
nand I_22343 (I382572,I382292,I11688);
nand I_22344 (I382589,I382572,I382326);
and I_22345 (I382606,I382408,I382589);
DFFARX1 I_22346  ( .D(I382606), .CLK(I2702), .RSTB(I382275), .Q(I382267) );
and I_22347 (I382240,I382572,I382541);
DFFARX1 I_22348  ( .D(I11700), .CLK(I2702), .RSTB(I382275), .Q(I382651) );
nor I_22349 (I382264,I382651,I382572);
nor I_22350 (I382682,I382651,I382326);
nand I_22351 (I382261,I382360,I382682);
not I_22352 (I382258,I382651);
DFFARX1 I_22353  ( .D(I11694), .CLK(I2702), .RSTB(I382275), .Q(I382727) );
not I_22354 (I382744,I382727);
nor I_22355 (I382761,I382744,I382425);
and I_22356 (I382778,I382651,I382761);
or I_22357 (I382795,I382572,I382778);
DFFARX1 I_22358  ( .D(I382795), .CLK(I2702), .RSTB(I382275), .Q(I382252) );
not I_22359 (I382826,I382744);
nor I_22360 (I382843,I382651,I382826);
nand I_22361 (I382255,I382744,I382843);
nand I_22362 (I382249,I382408,I382826);
not I_22363 (I382921,I2709);
not I_22364 (I382938,I19551);
nor I_22365 (I382955,I19566,I19560);
nand I_22366 (I382972,I382955,I19569);
nor I_22367 (I382989,I382938,I19566);
nand I_22368 (I383006,I382989,I19545);
DFFARX1 I_22369  ( .D(I383006), .CLK(I2702), .RSTB(I382921), .Q(I383023) );
not I_22370 (I382892,I383023);
not I_22371 (I383054,I19566);
not I_22372 (I383071,I383054);
not I_22373 (I383088,I19542);
nor I_22374 (I383105,I383088,I19557);
and I_22375 (I383122,I383105,I19563);
or I_22376 (I383139,I383122,I19572);
DFFARX1 I_22377  ( .D(I383139), .CLK(I2702), .RSTB(I382921), .Q(I383156) );
DFFARX1 I_22378  ( .D(I383156), .CLK(I2702), .RSTB(I382921), .Q(I382889) );
DFFARX1 I_22379  ( .D(I383156), .CLK(I2702), .RSTB(I382921), .Q(I383187) );
DFFARX1 I_22380  ( .D(I383156), .CLK(I2702), .RSTB(I382921), .Q(I382883) );
nand I_22381 (I383218,I382938,I19542);
nand I_22382 (I383235,I383218,I382972);
and I_22383 (I383252,I383054,I383235);
DFFARX1 I_22384  ( .D(I383252), .CLK(I2702), .RSTB(I382921), .Q(I382913) );
and I_22385 (I382886,I383218,I383187);
DFFARX1 I_22386  ( .D(I19554), .CLK(I2702), .RSTB(I382921), .Q(I383297) );
nor I_22387 (I382910,I383297,I383218);
nor I_22388 (I383328,I383297,I382972);
nand I_22389 (I382907,I383006,I383328);
not I_22390 (I382904,I383297);
DFFARX1 I_22391  ( .D(I19548), .CLK(I2702), .RSTB(I382921), .Q(I383373) );
not I_22392 (I383390,I383373);
nor I_22393 (I383407,I383390,I383071);
and I_22394 (I383424,I383297,I383407);
or I_22395 (I383441,I383218,I383424);
DFFARX1 I_22396  ( .D(I383441), .CLK(I2702), .RSTB(I382921), .Q(I382898) );
not I_22397 (I383472,I383390);
nor I_22398 (I383489,I383297,I383472);
nand I_22399 (I382901,I383390,I383489);
nand I_22400 (I382895,I383054,I383472);
not I_22401 (I383567,I2709);
not I_22402 (I383584,I623131);
nor I_22403 (I383601,I623128,I623113);
nand I_22404 (I383618,I383601,I623122);
nor I_22405 (I383635,I383584,I623128);
nand I_22406 (I383652,I383635,I623137);
DFFARX1 I_22407  ( .D(I383652), .CLK(I2702), .RSTB(I383567), .Q(I383669) );
not I_22408 (I383538,I383669);
not I_22409 (I383700,I623128);
not I_22410 (I383717,I383700);
not I_22411 (I383734,I623110);
nor I_22412 (I383751,I383734,I623116);
and I_22413 (I383768,I383751,I623140);
or I_22414 (I383785,I383768,I623134);
DFFARX1 I_22415  ( .D(I383785), .CLK(I2702), .RSTB(I383567), .Q(I383802) );
DFFARX1 I_22416  ( .D(I383802), .CLK(I2702), .RSTB(I383567), .Q(I383535) );
DFFARX1 I_22417  ( .D(I383802), .CLK(I2702), .RSTB(I383567), .Q(I383833) );
DFFARX1 I_22418  ( .D(I383802), .CLK(I2702), .RSTB(I383567), .Q(I383529) );
nand I_22419 (I383864,I383584,I623110);
nand I_22420 (I383881,I383864,I383618);
and I_22421 (I383898,I383700,I383881);
DFFARX1 I_22422  ( .D(I383898), .CLK(I2702), .RSTB(I383567), .Q(I383559) );
and I_22423 (I383532,I383864,I383833);
DFFARX1 I_22424  ( .D(I623119), .CLK(I2702), .RSTB(I383567), .Q(I383943) );
nor I_22425 (I383556,I383943,I383864);
nor I_22426 (I383974,I383943,I383618);
nand I_22427 (I383553,I383652,I383974);
not I_22428 (I383550,I383943);
DFFARX1 I_22429  ( .D(I623125), .CLK(I2702), .RSTB(I383567), .Q(I384019) );
not I_22430 (I384036,I384019);
nor I_22431 (I384053,I384036,I383717);
and I_22432 (I384070,I383943,I384053);
or I_22433 (I384087,I383864,I384070);
DFFARX1 I_22434  ( .D(I384087), .CLK(I2702), .RSTB(I383567), .Q(I383544) );
not I_22435 (I384118,I384036);
nor I_22436 (I384135,I383943,I384118);
nand I_22437 (I383547,I384036,I384135);
nand I_22438 (I383541,I383700,I384118);
not I_22439 (I384213,I2709);
not I_22440 (I384230,I301341);
nor I_22441 (I384247,I301320,I301332);
nand I_22442 (I384264,I384247,I301335);
nor I_22443 (I384281,I384230,I301320);
nand I_22444 (I384298,I384281,I301317);
DFFARX1 I_22445  ( .D(I384298), .CLK(I2702), .RSTB(I384213), .Q(I384315) );
not I_22446 (I384184,I384315);
not I_22447 (I384346,I301320);
not I_22448 (I384363,I384346);
not I_22449 (I384380,I301338);
nor I_22450 (I384397,I384380,I301329);
and I_22451 (I384414,I384397,I301323);
or I_22452 (I384431,I384414,I301347);
DFFARX1 I_22453  ( .D(I384431), .CLK(I2702), .RSTB(I384213), .Q(I384448) );
DFFARX1 I_22454  ( .D(I384448), .CLK(I2702), .RSTB(I384213), .Q(I384181) );
DFFARX1 I_22455  ( .D(I384448), .CLK(I2702), .RSTB(I384213), .Q(I384479) );
DFFARX1 I_22456  ( .D(I384448), .CLK(I2702), .RSTB(I384213), .Q(I384175) );
nand I_22457 (I384510,I384230,I301338);
nand I_22458 (I384527,I384510,I384264);
and I_22459 (I384544,I384346,I384527);
DFFARX1 I_22460  ( .D(I384544), .CLK(I2702), .RSTB(I384213), .Q(I384205) );
and I_22461 (I384178,I384510,I384479);
DFFARX1 I_22462  ( .D(I301344), .CLK(I2702), .RSTB(I384213), .Q(I384589) );
nor I_22463 (I384202,I384589,I384510);
nor I_22464 (I384620,I384589,I384264);
nand I_22465 (I384199,I384298,I384620);
not I_22466 (I384196,I384589);
DFFARX1 I_22467  ( .D(I301326), .CLK(I2702), .RSTB(I384213), .Q(I384665) );
not I_22468 (I384682,I384665);
nor I_22469 (I384699,I384682,I384363);
and I_22470 (I384716,I384589,I384699);
or I_22471 (I384733,I384510,I384716);
DFFARX1 I_22472  ( .D(I384733), .CLK(I2702), .RSTB(I384213), .Q(I384190) );
not I_22473 (I384764,I384682);
nor I_22474 (I384781,I384589,I384764);
nand I_22475 (I384193,I384682,I384781);
nand I_22476 (I384187,I384346,I384764);
not I_22477 (I384859,I2709);
not I_22478 (I384876,I597662);
nor I_22479 (I384893,I597650,I597659);
nand I_22480 (I384910,I384893,I597674);
nor I_22481 (I384927,I384876,I597650);
nand I_22482 (I384944,I384927,I597656);
DFFARX1 I_22483  ( .D(I384944), .CLK(I2702), .RSTB(I384859), .Q(I384961) );
not I_22484 (I384830,I384961);
not I_22485 (I384992,I597650);
not I_22486 (I385009,I384992);
not I_22487 (I385026,I597644);
nor I_22488 (I385043,I385026,I597665);
and I_22489 (I385060,I385043,I597647);
or I_22490 (I385077,I385060,I597653);
DFFARX1 I_22491  ( .D(I385077), .CLK(I2702), .RSTB(I384859), .Q(I385094) );
DFFARX1 I_22492  ( .D(I385094), .CLK(I2702), .RSTB(I384859), .Q(I384827) );
DFFARX1 I_22493  ( .D(I385094), .CLK(I2702), .RSTB(I384859), .Q(I385125) );
DFFARX1 I_22494  ( .D(I385094), .CLK(I2702), .RSTB(I384859), .Q(I384821) );
nand I_22495 (I385156,I384876,I597644);
nand I_22496 (I385173,I385156,I384910);
and I_22497 (I385190,I384992,I385173);
DFFARX1 I_22498  ( .D(I385190), .CLK(I2702), .RSTB(I384859), .Q(I384851) );
and I_22499 (I384824,I385156,I385125);
DFFARX1 I_22500  ( .D(I597671), .CLK(I2702), .RSTB(I384859), .Q(I385235) );
nor I_22501 (I384848,I385235,I385156);
nor I_22502 (I385266,I385235,I384910);
nand I_22503 (I384845,I384944,I385266);
not I_22504 (I384842,I385235);
DFFARX1 I_22505  ( .D(I597668), .CLK(I2702), .RSTB(I384859), .Q(I385311) );
not I_22506 (I385328,I385311);
nor I_22507 (I385345,I385328,I385009);
and I_22508 (I385362,I385235,I385345);
or I_22509 (I385379,I385156,I385362);
DFFARX1 I_22510  ( .D(I385379), .CLK(I2702), .RSTB(I384859), .Q(I384836) );
not I_22511 (I385410,I385328);
nor I_22512 (I385427,I385235,I385410);
nand I_22513 (I384839,I385328,I385427);
nand I_22514 (I384833,I384992,I385410);
not I_22515 (I385505,I2709);
not I_22516 (I385522,I315264);
nor I_22517 (I385539,I315243,I315255);
nand I_22518 (I385556,I385539,I315258);
nor I_22519 (I385573,I385522,I315243);
nand I_22520 (I385590,I385573,I315240);
DFFARX1 I_22521  ( .D(I385590), .CLK(I2702), .RSTB(I385505), .Q(I385607) );
not I_22522 (I385476,I385607);
not I_22523 (I385638,I315243);
not I_22524 (I385655,I385638);
not I_22525 (I385672,I315261);
nor I_22526 (I385689,I385672,I315252);
and I_22527 (I385706,I385689,I315246);
or I_22528 (I385723,I385706,I315270);
DFFARX1 I_22529  ( .D(I385723), .CLK(I2702), .RSTB(I385505), .Q(I385740) );
DFFARX1 I_22530  ( .D(I385740), .CLK(I2702), .RSTB(I385505), .Q(I385473) );
DFFARX1 I_22531  ( .D(I385740), .CLK(I2702), .RSTB(I385505), .Q(I385771) );
DFFARX1 I_22532  ( .D(I385740), .CLK(I2702), .RSTB(I385505), .Q(I385467) );
nand I_22533 (I385802,I385522,I315261);
nand I_22534 (I385819,I385802,I385556);
and I_22535 (I385836,I385638,I385819);
DFFARX1 I_22536  ( .D(I385836), .CLK(I2702), .RSTB(I385505), .Q(I385497) );
and I_22537 (I385470,I385802,I385771);
DFFARX1 I_22538  ( .D(I315267), .CLK(I2702), .RSTB(I385505), .Q(I385881) );
nor I_22539 (I385494,I385881,I385802);
nor I_22540 (I385912,I385881,I385556);
nand I_22541 (I385491,I385590,I385912);
not I_22542 (I385488,I385881);
DFFARX1 I_22543  ( .D(I315249), .CLK(I2702), .RSTB(I385505), .Q(I385957) );
not I_22544 (I385974,I385957);
nor I_22545 (I385991,I385974,I385655);
and I_22546 (I386008,I385881,I385991);
or I_22547 (I386025,I385802,I386008);
DFFARX1 I_22548  ( .D(I386025), .CLK(I2702), .RSTB(I385505), .Q(I385482) );
not I_22549 (I386056,I385974);
nor I_22550 (I386073,I385881,I386056);
nand I_22551 (I385485,I385974,I386073);
nand I_22552 (I385479,I385638,I386056);
not I_22553 (I386151,I2709);
not I_22554 (I386168,I690958);
nor I_22555 (I386185,I690943,I690949);
nand I_22556 (I386202,I386185,I690946);
nor I_22557 (I386219,I386168,I690943);
nand I_22558 (I386236,I386219,I690955);
DFFARX1 I_22559  ( .D(I386236), .CLK(I2702), .RSTB(I386151), .Q(I386253) );
not I_22560 (I386122,I386253);
not I_22561 (I386284,I690943);
not I_22562 (I386301,I386284);
not I_22563 (I386318,I690970);
nor I_22564 (I386335,I386318,I690964);
and I_22565 (I386352,I386335,I690961);
or I_22566 (I386369,I386352,I690940);
DFFARX1 I_22567  ( .D(I386369), .CLK(I2702), .RSTB(I386151), .Q(I386386) );
DFFARX1 I_22568  ( .D(I386386), .CLK(I2702), .RSTB(I386151), .Q(I386119) );
DFFARX1 I_22569  ( .D(I386386), .CLK(I2702), .RSTB(I386151), .Q(I386417) );
DFFARX1 I_22570  ( .D(I386386), .CLK(I2702), .RSTB(I386151), .Q(I386113) );
nand I_22571 (I386448,I386168,I690970);
nand I_22572 (I386465,I386448,I386202);
and I_22573 (I386482,I386284,I386465);
DFFARX1 I_22574  ( .D(I386482), .CLK(I2702), .RSTB(I386151), .Q(I386143) );
and I_22575 (I386116,I386448,I386417);
DFFARX1 I_22576  ( .D(I690967), .CLK(I2702), .RSTB(I386151), .Q(I386527) );
nor I_22577 (I386140,I386527,I386448);
nor I_22578 (I386558,I386527,I386202);
nand I_22579 (I386137,I386236,I386558);
not I_22580 (I386134,I386527);
DFFARX1 I_22581  ( .D(I690952), .CLK(I2702), .RSTB(I386151), .Q(I386603) );
not I_22582 (I386620,I386603);
nor I_22583 (I386637,I386620,I386301);
and I_22584 (I386654,I386527,I386637);
or I_22585 (I386671,I386448,I386654);
DFFARX1 I_22586  ( .D(I386671), .CLK(I2702), .RSTB(I386151), .Q(I386128) );
not I_22587 (I386702,I386620);
nor I_22588 (I386719,I386527,I386702);
nand I_22589 (I386131,I386620,I386719);
nand I_22590 (I386125,I386284,I386702);
not I_22591 (I386797,I2709);
not I_22592 (I386814,I253605);
nor I_22593 (I386831,I253584,I253596);
nand I_22594 (I386848,I386831,I253599);
nor I_22595 (I386865,I386814,I253584);
nand I_22596 (I386882,I386865,I253581);
DFFARX1 I_22597  ( .D(I386882), .CLK(I2702), .RSTB(I386797), .Q(I386899) );
not I_22598 (I386768,I386899);
not I_22599 (I386930,I253584);
not I_22600 (I386947,I386930);
not I_22601 (I386964,I253602);
nor I_22602 (I386981,I386964,I253593);
and I_22603 (I386998,I386981,I253587);
or I_22604 (I387015,I386998,I253611);
DFFARX1 I_22605  ( .D(I387015), .CLK(I2702), .RSTB(I386797), .Q(I387032) );
DFFARX1 I_22606  ( .D(I387032), .CLK(I2702), .RSTB(I386797), .Q(I386765) );
DFFARX1 I_22607  ( .D(I387032), .CLK(I2702), .RSTB(I386797), .Q(I387063) );
DFFARX1 I_22608  ( .D(I387032), .CLK(I2702), .RSTB(I386797), .Q(I386759) );
nand I_22609 (I387094,I386814,I253602);
nand I_22610 (I387111,I387094,I386848);
and I_22611 (I387128,I386930,I387111);
DFFARX1 I_22612  ( .D(I387128), .CLK(I2702), .RSTB(I386797), .Q(I386789) );
and I_22613 (I386762,I387094,I387063);
DFFARX1 I_22614  ( .D(I253608), .CLK(I2702), .RSTB(I386797), .Q(I387173) );
nor I_22615 (I386786,I387173,I387094);
nor I_22616 (I387204,I387173,I386848);
nand I_22617 (I386783,I386882,I387204);
not I_22618 (I386780,I387173);
DFFARX1 I_22619  ( .D(I253590), .CLK(I2702), .RSTB(I386797), .Q(I387249) );
not I_22620 (I387266,I387249);
nor I_22621 (I387283,I387266,I386947);
and I_22622 (I387300,I387173,I387283);
or I_22623 (I387317,I387094,I387300);
DFFARX1 I_22624  ( .D(I387317), .CLK(I2702), .RSTB(I386797), .Q(I386774) );
not I_22625 (I387348,I387266);
nor I_22626 (I387365,I387173,I387348);
nand I_22627 (I386777,I387266,I387365);
nand I_22628 (I386771,I386930,I387348);
not I_22629 (I387443,I2709);
not I_22630 (I387460,I547673);
nor I_22631 (I387477,I547685,I547679);
nand I_22632 (I387494,I387477,I547664);
nor I_22633 (I387511,I387460,I547685);
nand I_22634 (I387528,I387511,I547691);
DFFARX1 I_22635  ( .D(I387528), .CLK(I2702), .RSTB(I387443), .Q(I387545) );
not I_22636 (I387414,I387545);
not I_22637 (I387576,I547685);
not I_22638 (I387593,I387576);
not I_22639 (I387610,I547688);
nor I_22640 (I387627,I387610,I547670);
and I_22641 (I387644,I387627,I547667);
or I_22642 (I387661,I387644,I547694);
DFFARX1 I_22643  ( .D(I387661), .CLK(I2702), .RSTB(I387443), .Q(I387678) );
DFFARX1 I_22644  ( .D(I387678), .CLK(I2702), .RSTB(I387443), .Q(I387411) );
DFFARX1 I_22645  ( .D(I387678), .CLK(I2702), .RSTB(I387443), .Q(I387709) );
DFFARX1 I_22646  ( .D(I387678), .CLK(I2702), .RSTB(I387443), .Q(I387405) );
nand I_22647 (I387740,I387460,I547688);
nand I_22648 (I387757,I387740,I387494);
and I_22649 (I387774,I387576,I387757);
DFFARX1 I_22650  ( .D(I387774), .CLK(I2702), .RSTB(I387443), .Q(I387435) );
and I_22651 (I387408,I387740,I387709);
DFFARX1 I_22652  ( .D(I547682), .CLK(I2702), .RSTB(I387443), .Q(I387819) );
nor I_22653 (I387432,I387819,I387740);
nor I_22654 (I387850,I387819,I387494);
nand I_22655 (I387429,I387528,I387850);
not I_22656 (I387426,I387819);
DFFARX1 I_22657  ( .D(I547676), .CLK(I2702), .RSTB(I387443), .Q(I387895) );
not I_22658 (I387912,I387895);
nor I_22659 (I387929,I387912,I387593);
and I_22660 (I387946,I387819,I387929);
or I_22661 (I387963,I387740,I387946);
DFFARX1 I_22662  ( .D(I387963), .CLK(I2702), .RSTB(I387443), .Q(I387420) );
not I_22663 (I387994,I387912);
nor I_22664 (I388011,I387819,I387994);
nand I_22665 (I387423,I387912,I388011);
nand I_22666 (I387417,I387576,I387994);
not I_22667 (I388089,I2709);
not I_22668 (I388106,I701940);
nor I_22669 (I388123,I701925,I701931);
nand I_22670 (I388140,I388123,I701928);
nor I_22671 (I388157,I388106,I701925);
nand I_22672 (I388174,I388157,I701937);
DFFARX1 I_22673  ( .D(I388174), .CLK(I2702), .RSTB(I388089), .Q(I388191) );
not I_22674 (I388060,I388191);
not I_22675 (I388222,I701925);
not I_22676 (I388239,I388222);
not I_22677 (I388256,I701952);
nor I_22678 (I388273,I388256,I701946);
and I_22679 (I388290,I388273,I701943);
or I_22680 (I388307,I388290,I701922);
DFFARX1 I_22681  ( .D(I388307), .CLK(I2702), .RSTB(I388089), .Q(I388324) );
DFFARX1 I_22682  ( .D(I388324), .CLK(I2702), .RSTB(I388089), .Q(I388057) );
DFFARX1 I_22683  ( .D(I388324), .CLK(I2702), .RSTB(I388089), .Q(I388355) );
DFFARX1 I_22684  ( .D(I388324), .CLK(I2702), .RSTB(I388089), .Q(I388051) );
nand I_22685 (I388386,I388106,I701952);
nand I_22686 (I388403,I388386,I388140);
and I_22687 (I388420,I388222,I388403);
DFFARX1 I_22688  ( .D(I388420), .CLK(I2702), .RSTB(I388089), .Q(I388081) );
and I_22689 (I388054,I388386,I388355);
DFFARX1 I_22690  ( .D(I701949), .CLK(I2702), .RSTB(I388089), .Q(I388465) );
nor I_22691 (I388078,I388465,I388386);
nor I_22692 (I388496,I388465,I388140);
nand I_22693 (I388075,I388174,I388496);
not I_22694 (I388072,I388465);
DFFARX1 I_22695  ( .D(I701934), .CLK(I2702), .RSTB(I388089), .Q(I388541) );
not I_22696 (I388558,I388541);
nor I_22697 (I388575,I388558,I388239);
and I_22698 (I388592,I388465,I388575);
or I_22699 (I388609,I388386,I388592);
DFFARX1 I_22700  ( .D(I388609), .CLK(I2702), .RSTB(I388089), .Q(I388066) );
not I_22701 (I388640,I388558);
nor I_22702 (I388657,I388465,I388640);
nand I_22703 (I388069,I388558,I388657);
nand I_22704 (I388063,I388222,I388640);
not I_22705 (I388735,I2709);
not I_22706 (I388752,I523278);
nor I_22707 (I388769,I523290,I523284);
nand I_22708 (I388786,I388769,I523269);
nor I_22709 (I388803,I388752,I523290);
nand I_22710 (I388820,I388803,I523296);
DFFARX1 I_22711  ( .D(I388820), .CLK(I2702), .RSTB(I388735), .Q(I388837) );
not I_22712 (I388706,I388837);
not I_22713 (I388868,I523290);
not I_22714 (I388885,I388868);
not I_22715 (I388902,I523293);
nor I_22716 (I388919,I388902,I523275);
and I_22717 (I388936,I388919,I523272);
or I_22718 (I388953,I388936,I523299);
DFFARX1 I_22719  ( .D(I388953), .CLK(I2702), .RSTB(I388735), .Q(I388970) );
DFFARX1 I_22720  ( .D(I388970), .CLK(I2702), .RSTB(I388735), .Q(I388703) );
DFFARX1 I_22721  ( .D(I388970), .CLK(I2702), .RSTB(I388735), .Q(I389001) );
DFFARX1 I_22722  ( .D(I388970), .CLK(I2702), .RSTB(I388735), .Q(I388697) );
nand I_22723 (I389032,I388752,I523293);
nand I_22724 (I389049,I389032,I388786);
and I_22725 (I389066,I388868,I389049);
DFFARX1 I_22726  ( .D(I389066), .CLK(I2702), .RSTB(I388735), .Q(I388727) );
and I_22727 (I388700,I389032,I389001);
DFFARX1 I_22728  ( .D(I523287), .CLK(I2702), .RSTB(I388735), .Q(I389111) );
nor I_22729 (I388724,I389111,I389032);
nor I_22730 (I389142,I389111,I388786);
nand I_22731 (I388721,I388820,I389142);
not I_22732 (I388718,I389111);
DFFARX1 I_22733  ( .D(I523281), .CLK(I2702), .RSTB(I388735), .Q(I389187) );
not I_22734 (I389204,I389187);
nor I_22735 (I389221,I389204,I388885);
and I_22736 (I389238,I389111,I389221);
or I_22737 (I389255,I389032,I389238);
DFFARX1 I_22738  ( .D(I389255), .CLK(I2702), .RSTB(I388735), .Q(I388712) );
not I_22739 (I389286,I389204);
nor I_22740 (I389303,I389111,I389286);
nand I_22741 (I388715,I389204,I389303);
nand I_22742 (I388709,I388868,I389286);
not I_22743 (I389381,I2709);
not I_22744 (I389398,I92408);
nor I_22745 (I389415,I92399,I92390);
nand I_22746 (I389432,I389415,I92405);
nor I_22747 (I389449,I389398,I92399);
nand I_22748 (I389466,I389449,I92402);
DFFARX1 I_22749  ( .D(I389466), .CLK(I2702), .RSTB(I389381), .Q(I389483) );
not I_22750 (I389352,I389483);
not I_22751 (I389514,I92399);
not I_22752 (I389531,I389514);
not I_22753 (I389548,I92411);
nor I_22754 (I389565,I389548,I92396);
and I_22755 (I389582,I389565,I92414);
or I_22756 (I389599,I389582,I92387);
DFFARX1 I_22757  ( .D(I389599), .CLK(I2702), .RSTB(I389381), .Q(I389616) );
DFFARX1 I_22758  ( .D(I389616), .CLK(I2702), .RSTB(I389381), .Q(I389349) );
DFFARX1 I_22759  ( .D(I389616), .CLK(I2702), .RSTB(I389381), .Q(I389647) );
DFFARX1 I_22760  ( .D(I389616), .CLK(I2702), .RSTB(I389381), .Q(I389343) );
nand I_22761 (I389678,I389398,I92411);
nand I_22762 (I389695,I389678,I389432);
and I_22763 (I389712,I389514,I389695);
DFFARX1 I_22764  ( .D(I389712), .CLK(I2702), .RSTB(I389381), .Q(I389373) );
and I_22765 (I389346,I389678,I389647);
DFFARX1 I_22766  ( .D(I92417), .CLK(I2702), .RSTB(I389381), .Q(I389757) );
nor I_22767 (I389370,I389757,I389678);
nor I_22768 (I389788,I389757,I389432);
nand I_22769 (I389367,I389466,I389788);
not I_22770 (I389364,I389757);
DFFARX1 I_22771  ( .D(I92393), .CLK(I2702), .RSTB(I389381), .Q(I389833) );
not I_22772 (I389850,I389833);
nor I_22773 (I389867,I389850,I389531);
and I_22774 (I389884,I389757,I389867);
or I_22775 (I389901,I389678,I389884);
DFFARX1 I_22776  ( .D(I389901), .CLK(I2702), .RSTB(I389381), .Q(I389358) );
not I_22777 (I389932,I389850);
nor I_22778 (I389949,I389757,I389932);
nand I_22779 (I389361,I389850,I389949);
nand I_22780 (I389355,I389514,I389932);
not I_22781 (I390027,I2709);
not I_22782 (I390044,I225469);
nor I_22783 (I390061,I225475,I225472);
nand I_22784 (I390078,I390061,I225466);
nor I_22785 (I390095,I390044,I225475);
nand I_22786 (I390112,I390095,I225490);
DFFARX1 I_22787  ( .D(I390112), .CLK(I2702), .RSTB(I390027), .Q(I390129) );
not I_22788 (I389998,I390129);
not I_22789 (I390160,I225475);
not I_22790 (I390177,I390160);
not I_22791 (I390194,I225487);
nor I_22792 (I390211,I390194,I225478);
and I_22793 (I390228,I390211,I225463);
or I_22794 (I390245,I390228,I225484);
DFFARX1 I_22795  ( .D(I390245), .CLK(I2702), .RSTB(I390027), .Q(I390262) );
DFFARX1 I_22796  ( .D(I390262), .CLK(I2702), .RSTB(I390027), .Q(I389995) );
DFFARX1 I_22797  ( .D(I390262), .CLK(I2702), .RSTB(I390027), .Q(I390293) );
DFFARX1 I_22798  ( .D(I390262), .CLK(I2702), .RSTB(I390027), .Q(I389989) );
nand I_22799 (I390324,I390044,I225487);
nand I_22800 (I390341,I390324,I390078);
and I_22801 (I390358,I390160,I390341);
DFFARX1 I_22802  ( .D(I390358), .CLK(I2702), .RSTB(I390027), .Q(I390019) );
and I_22803 (I389992,I390324,I390293);
DFFARX1 I_22804  ( .D(I225481), .CLK(I2702), .RSTB(I390027), .Q(I390403) );
nor I_22805 (I390016,I390403,I390324);
nor I_22806 (I390434,I390403,I390078);
nand I_22807 (I390013,I390112,I390434);
not I_22808 (I390010,I390403);
DFFARX1 I_22809  ( .D(I225493), .CLK(I2702), .RSTB(I390027), .Q(I390479) );
not I_22810 (I390496,I390479);
nor I_22811 (I390513,I390496,I390177);
and I_22812 (I390530,I390403,I390513);
or I_22813 (I390547,I390324,I390530);
DFFARX1 I_22814  ( .D(I390547), .CLK(I2702), .RSTB(I390027), .Q(I390004) );
not I_22815 (I390578,I390496);
nor I_22816 (I390595,I390403,I390578);
nand I_22817 (I390007,I390496,I390595);
nand I_22818 (I390001,I390160,I390578);
not I_22819 (I390673,I2709);
not I_22820 (I390690,I472590);
nor I_22821 (I390707,I472593,I472575);
nand I_22822 (I390724,I390707,I472602);
nor I_22823 (I390741,I390690,I472593);
nand I_22824 (I390758,I390741,I472581);
DFFARX1 I_22825  ( .D(I390758), .CLK(I2702), .RSTB(I390673), .Q(I390775) );
not I_22826 (I390644,I390775);
not I_22827 (I390806,I472593);
not I_22828 (I390823,I390806);
not I_22829 (I390840,I472587);
nor I_22830 (I390857,I390840,I472599);
and I_22831 (I390874,I390857,I472605);
or I_22832 (I390891,I390874,I472584);
DFFARX1 I_22833  ( .D(I390891), .CLK(I2702), .RSTB(I390673), .Q(I390908) );
DFFARX1 I_22834  ( .D(I390908), .CLK(I2702), .RSTB(I390673), .Q(I390641) );
DFFARX1 I_22835  ( .D(I390908), .CLK(I2702), .RSTB(I390673), .Q(I390939) );
DFFARX1 I_22836  ( .D(I390908), .CLK(I2702), .RSTB(I390673), .Q(I390635) );
nand I_22837 (I390970,I390690,I472587);
nand I_22838 (I390987,I390970,I390724);
and I_22839 (I391004,I390806,I390987);
DFFARX1 I_22840  ( .D(I391004), .CLK(I2702), .RSTB(I390673), .Q(I390665) );
and I_22841 (I390638,I390970,I390939);
DFFARX1 I_22842  ( .D(I472596), .CLK(I2702), .RSTB(I390673), .Q(I391049) );
nor I_22843 (I390662,I391049,I390970);
nor I_22844 (I391080,I391049,I390724);
nand I_22845 (I390659,I390758,I391080);
not I_22846 (I390656,I391049);
DFFARX1 I_22847  ( .D(I472578), .CLK(I2702), .RSTB(I390673), .Q(I391125) );
not I_22848 (I391142,I391125);
nor I_22849 (I391159,I391142,I390823);
and I_22850 (I391176,I391049,I391159);
or I_22851 (I391193,I390970,I391176);
DFFARX1 I_22852  ( .D(I391193), .CLK(I2702), .RSTB(I390673), .Q(I390650) );
not I_22853 (I391224,I391142);
nor I_22854 (I391241,I391049,I391224);
nand I_22855 (I390653,I391142,I391241);
nand I_22856 (I390647,I390806,I391224);
not I_22857 (I391319,I2709);
not I_22858 (I391336,I144189);
nor I_22859 (I391353,I144210,I144192);
nand I_22860 (I391370,I391353,I144216);
nor I_22861 (I391387,I391336,I144210);
nand I_22862 (I391404,I391387,I144213);
DFFARX1 I_22863  ( .D(I391404), .CLK(I2702), .RSTB(I391319), .Q(I391421) );
not I_22864 (I391290,I391421);
not I_22865 (I391452,I144210);
not I_22866 (I391469,I391452);
not I_22867 (I391486,I144207);
nor I_22868 (I391503,I391486,I144186);
and I_22869 (I391520,I391503,I144198);
or I_22870 (I391537,I391520,I144195);
DFFARX1 I_22871  ( .D(I391537), .CLK(I2702), .RSTB(I391319), .Q(I391554) );
DFFARX1 I_22872  ( .D(I391554), .CLK(I2702), .RSTB(I391319), .Q(I391287) );
DFFARX1 I_22873  ( .D(I391554), .CLK(I2702), .RSTB(I391319), .Q(I391585) );
DFFARX1 I_22874  ( .D(I391554), .CLK(I2702), .RSTB(I391319), .Q(I391281) );
nand I_22875 (I391616,I391336,I144207);
nand I_22876 (I391633,I391616,I391370);
and I_22877 (I391650,I391452,I391633);
DFFARX1 I_22878  ( .D(I391650), .CLK(I2702), .RSTB(I391319), .Q(I391311) );
and I_22879 (I391284,I391616,I391585);
DFFARX1 I_22880  ( .D(I144201), .CLK(I2702), .RSTB(I391319), .Q(I391695) );
nor I_22881 (I391308,I391695,I391616);
nor I_22882 (I391726,I391695,I391370);
nand I_22883 (I391305,I391404,I391726);
not I_22884 (I391302,I391695);
DFFARX1 I_22885  ( .D(I144204), .CLK(I2702), .RSTB(I391319), .Q(I391771) );
not I_22886 (I391788,I391771);
nor I_22887 (I391805,I391788,I391469);
and I_22888 (I391822,I391695,I391805);
or I_22889 (I391839,I391616,I391822);
DFFARX1 I_22890  ( .D(I391839), .CLK(I2702), .RSTB(I391319), .Q(I391296) );
not I_22891 (I391870,I391788);
nor I_22892 (I391887,I391695,I391870);
nand I_22893 (I391299,I391788,I391887);
nand I_22894 (I391293,I391452,I391870);
not I_22895 (I391965,I2709);
not I_22896 (I391982,I298026);
nor I_22897 (I391999,I298005,I298017);
nand I_22898 (I392016,I391999,I298020);
nor I_22899 (I392033,I391982,I298005);
nand I_22900 (I392050,I392033,I298002);
DFFARX1 I_22901  ( .D(I392050), .CLK(I2702), .RSTB(I391965), .Q(I392067) );
not I_22902 (I391936,I392067);
not I_22903 (I392098,I298005);
not I_22904 (I392115,I392098);
not I_22905 (I392132,I298023);
nor I_22906 (I392149,I392132,I298014);
and I_22907 (I392166,I392149,I298008);
or I_22908 (I392183,I392166,I298032);
DFFARX1 I_22909  ( .D(I392183), .CLK(I2702), .RSTB(I391965), .Q(I392200) );
DFFARX1 I_22910  ( .D(I392200), .CLK(I2702), .RSTB(I391965), .Q(I391933) );
DFFARX1 I_22911  ( .D(I392200), .CLK(I2702), .RSTB(I391965), .Q(I392231) );
DFFARX1 I_22912  ( .D(I392200), .CLK(I2702), .RSTB(I391965), .Q(I391927) );
nand I_22913 (I392262,I391982,I298023);
nand I_22914 (I392279,I392262,I392016);
and I_22915 (I392296,I392098,I392279);
DFFARX1 I_22916  ( .D(I392296), .CLK(I2702), .RSTB(I391965), .Q(I391957) );
and I_22917 (I391930,I392262,I392231);
DFFARX1 I_22918  ( .D(I298029), .CLK(I2702), .RSTB(I391965), .Q(I392341) );
nor I_22919 (I391954,I392341,I392262);
nor I_22920 (I392372,I392341,I392016);
nand I_22921 (I391951,I392050,I392372);
not I_22922 (I391948,I392341);
DFFARX1 I_22923  ( .D(I298011), .CLK(I2702), .RSTB(I391965), .Q(I392417) );
not I_22924 (I392434,I392417);
nor I_22925 (I392451,I392434,I392115);
and I_22926 (I392468,I392341,I392451);
or I_22927 (I392485,I392262,I392468);
DFFARX1 I_22928  ( .D(I392485), .CLK(I2702), .RSTB(I391965), .Q(I391942) );
not I_22929 (I392516,I392434);
nor I_22930 (I392533,I392341,I392516);
nand I_22931 (I391945,I392434,I392533);
nand I_22932 (I391939,I392098,I392516);
not I_22933 (I392611,I2709);
not I_22934 (I392628,I463920);
nor I_22935 (I392645,I463923,I463905);
nand I_22936 (I392662,I392645,I463932);
nor I_22937 (I392679,I392628,I463923);
nand I_22938 (I392696,I392679,I463911);
DFFARX1 I_22939  ( .D(I392696), .CLK(I2702), .RSTB(I392611), .Q(I392713) );
not I_22940 (I392582,I392713);
not I_22941 (I392744,I463923);
not I_22942 (I392761,I392744);
not I_22943 (I392778,I463917);
nor I_22944 (I392795,I392778,I463929);
and I_22945 (I392812,I392795,I463935);
or I_22946 (I392829,I392812,I463914);
DFFARX1 I_22947  ( .D(I392829), .CLK(I2702), .RSTB(I392611), .Q(I392846) );
DFFARX1 I_22948  ( .D(I392846), .CLK(I2702), .RSTB(I392611), .Q(I392579) );
DFFARX1 I_22949  ( .D(I392846), .CLK(I2702), .RSTB(I392611), .Q(I392877) );
DFFARX1 I_22950  ( .D(I392846), .CLK(I2702), .RSTB(I392611), .Q(I392573) );
nand I_22951 (I392908,I392628,I463917);
nand I_22952 (I392925,I392908,I392662);
and I_22953 (I392942,I392744,I392925);
DFFARX1 I_22954  ( .D(I392942), .CLK(I2702), .RSTB(I392611), .Q(I392603) );
and I_22955 (I392576,I392908,I392877);
DFFARX1 I_22956  ( .D(I463926), .CLK(I2702), .RSTB(I392611), .Q(I392987) );
nor I_22957 (I392600,I392987,I392908);
nor I_22958 (I393018,I392987,I392662);
nand I_22959 (I392597,I392696,I393018);
not I_22960 (I392594,I392987);
DFFARX1 I_22961  ( .D(I463908), .CLK(I2702), .RSTB(I392611), .Q(I393063) );
not I_22962 (I393080,I393063);
nor I_22963 (I393097,I393080,I392761);
and I_22964 (I393114,I392987,I393097);
or I_22965 (I393131,I392908,I393114);
DFFARX1 I_22966  ( .D(I393131), .CLK(I2702), .RSTB(I392611), .Q(I392588) );
not I_22967 (I393162,I393080);
nor I_22968 (I393179,I392987,I393162);
nand I_22969 (I392591,I393080,I393179);
nand I_22970 (I392585,I392744,I393162);
not I_22971 (I393257,I2709);
not I_22972 (I393274,I125354);
nor I_22973 (I393291,I125345,I125336);
nand I_22974 (I393308,I393291,I125351);
nor I_22975 (I393325,I393274,I125345);
nand I_22976 (I393342,I393325,I125348);
DFFARX1 I_22977  ( .D(I393342), .CLK(I2702), .RSTB(I393257), .Q(I393359) );
not I_22978 (I393228,I393359);
not I_22979 (I393390,I125345);
not I_22980 (I393407,I393390);
not I_22981 (I393424,I125357);
nor I_22982 (I393441,I393424,I125342);
and I_22983 (I393458,I393441,I125360);
or I_22984 (I393475,I393458,I125333);
DFFARX1 I_22985  ( .D(I393475), .CLK(I2702), .RSTB(I393257), .Q(I393492) );
DFFARX1 I_22986  ( .D(I393492), .CLK(I2702), .RSTB(I393257), .Q(I393225) );
DFFARX1 I_22987  ( .D(I393492), .CLK(I2702), .RSTB(I393257), .Q(I393523) );
DFFARX1 I_22988  ( .D(I393492), .CLK(I2702), .RSTB(I393257), .Q(I393219) );
nand I_22989 (I393554,I393274,I125357);
nand I_22990 (I393571,I393554,I393308);
and I_22991 (I393588,I393390,I393571);
DFFARX1 I_22992  ( .D(I393588), .CLK(I2702), .RSTB(I393257), .Q(I393249) );
and I_22993 (I393222,I393554,I393523);
DFFARX1 I_22994  ( .D(I125363), .CLK(I2702), .RSTB(I393257), .Q(I393633) );
nor I_22995 (I393246,I393633,I393554);
nor I_22996 (I393664,I393633,I393308);
nand I_22997 (I393243,I393342,I393664);
not I_22998 (I393240,I393633);
DFFARX1 I_22999  ( .D(I125339), .CLK(I2702), .RSTB(I393257), .Q(I393709) );
not I_23000 (I393726,I393709);
nor I_23001 (I393743,I393726,I393407);
and I_23002 (I393760,I393633,I393743);
or I_23003 (I393777,I393554,I393760);
DFFARX1 I_23004  ( .D(I393777), .CLK(I2702), .RSTB(I393257), .Q(I393234) );
not I_23005 (I393808,I393726);
nor I_23006 (I393825,I393633,I393808);
nand I_23007 (I393237,I393726,I393825);
nand I_23008 (I393231,I393390,I393808);
not I_23009 (I393903,I2709);
not I_23010 (I393920,I258909);
nor I_23011 (I393937,I258888,I258900);
nand I_23012 (I393954,I393937,I258903);
nor I_23013 (I393971,I393920,I258888);
nand I_23014 (I393988,I393971,I258885);
DFFARX1 I_23015  ( .D(I393988), .CLK(I2702), .RSTB(I393903), .Q(I394005) );
not I_23016 (I393874,I394005);
not I_23017 (I394036,I258888);
not I_23018 (I394053,I394036);
not I_23019 (I394070,I258906);
nor I_23020 (I394087,I394070,I258897);
and I_23021 (I394104,I394087,I258891);
or I_23022 (I394121,I394104,I258915);
DFFARX1 I_23023  ( .D(I394121), .CLK(I2702), .RSTB(I393903), .Q(I394138) );
DFFARX1 I_23024  ( .D(I394138), .CLK(I2702), .RSTB(I393903), .Q(I393871) );
DFFARX1 I_23025  ( .D(I394138), .CLK(I2702), .RSTB(I393903), .Q(I394169) );
DFFARX1 I_23026  ( .D(I394138), .CLK(I2702), .RSTB(I393903), .Q(I393865) );
nand I_23027 (I394200,I393920,I258906);
nand I_23028 (I394217,I394200,I393954);
and I_23029 (I394234,I394036,I394217);
DFFARX1 I_23030  ( .D(I394234), .CLK(I2702), .RSTB(I393903), .Q(I393895) );
and I_23031 (I393868,I394200,I394169);
DFFARX1 I_23032  ( .D(I258912), .CLK(I2702), .RSTB(I393903), .Q(I394279) );
nor I_23033 (I393892,I394279,I394200);
nor I_23034 (I394310,I394279,I393954);
nand I_23035 (I393889,I393988,I394310);
not I_23036 (I393886,I394279);
DFFARX1 I_23037  ( .D(I258894), .CLK(I2702), .RSTB(I393903), .Q(I394355) );
not I_23038 (I394372,I394355);
nor I_23039 (I394389,I394372,I394053);
and I_23040 (I394406,I394279,I394389);
or I_23041 (I394423,I394200,I394406);
DFFARX1 I_23042  ( .D(I394423), .CLK(I2702), .RSTB(I393903), .Q(I393880) );
not I_23043 (I394454,I394372);
nor I_23044 (I394471,I394279,I394454);
nand I_23045 (I393883,I394372,I394471);
nand I_23046 (I393877,I394036,I394454);
not I_23047 (I394549,I2709);
not I_23048 (I394566,I317253);
nor I_23049 (I394583,I317232,I317244);
nand I_23050 (I394600,I394583,I317247);
nor I_23051 (I394617,I394566,I317232);
nand I_23052 (I394634,I394617,I317229);
DFFARX1 I_23053  ( .D(I394634), .CLK(I2702), .RSTB(I394549), .Q(I394651) );
not I_23054 (I394520,I394651);
not I_23055 (I394682,I317232);
not I_23056 (I394699,I394682);
not I_23057 (I394716,I317250);
nor I_23058 (I394733,I394716,I317241);
and I_23059 (I394750,I394733,I317235);
or I_23060 (I394767,I394750,I317259);
DFFARX1 I_23061  ( .D(I394767), .CLK(I2702), .RSTB(I394549), .Q(I394784) );
DFFARX1 I_23062  ( .D(I394784), .CLK(I2702), .RSTB(I394549), .Q(I394517) );
DFFARX1 I_23063  ( .D(I394784), .CLK(I2702), .RSTB(I394549), .Q(I394815) );
DFFARX1 I_23064  ( .D(I394784), .CLK(I2702), .RSTB(I394549), .Q(I394511) );
nand I_23065 (I394846,I394566,I317250);
nand I_23066 (I394863,I394846,I394600);
and I_23067 (I394880,I394682,I394863);
DFFARX1 I_23068  ( .D(I394880), .CLK(I2702), .RSTB(I394549), .Q(I394541) );
and I_23069 (I394514,I394846,I394815);
DFFARX1 I_23070  ( .D(I317256), .CLK(I2702), .RSTB(I394549), .Q(I394925) );
nor I_23071 (I394538,I394925,I394846);
nor I_23072 (I394956,I394925,I394600);
nand I_23073 (I394535,I394634,I394956);
not I_23074 (I394532,I394925);
DFFARX1 I_23075  ( .D(I317238), .CLK(I2702), .RSTB(I394549), .Q(I395001) );
not I_23076 (I395018,I395001);
nor I_23077 (I395035,I395018,I394699);
and I_23078 (I395052,I394925,I395035);
or I_23079 (I395069,I394846,I395052);
DFFARX1 I_23080  ( .D(I395069), .CLK(I2702), .RSTB(I394549), .Q(I394526) );
not I_23081 (I395100,I395018);
nor I_23082 (I395117,I394925,I395100);
nand I_23083 (I394529,I395018,I395117);
nand I_23084 (I394523,I394682,I395100);
not I_23085 (I395195,I2709);
not I_23086 (I395212,I329850);
nor I_23087 (I395229,I329829,I329841);
nand I_23088 (I395246,I395229,I329844);
nor I_23089 (I395263,I395212,I329829);
nand I_23090 (I395280,I395263,I329826);
DFFARX1 I_23091  ( .D(I395280), .CLK(I2702), .RSTB(I395195), .Q(I395297) );
not I_23092 (I395166,I395297);
not I_23093 (I395328,I329829);
not I_23094 (I395345,I395328);
not I_23095 (I395362,I329847);
nor I_23096 (I395379,I395362,I329838);
and I_23097 (I395396,I395379,I329832);
or I_23098 (I395413,I395396,I329856);
DFFARX1 I_23099  ( .D(I395413), .CLK(I2702), .RSTB(I395195), .Q(I395430) );
DFFARX1 I_23100  ( .D(I395430), .CLK(I2702), .RSTB(I395195), .Q(I395163) );
DFFARX1 I_23101  ( .D(I395430), .CLK(I2702), .RSTB(I395195), .Q(I395461) );
DFFARX1 I_23102  ( .D(I395430), .CLK(I2702), .RSTB(I395195), .Q(I395157) );
nand I_23103 (I395492,I395212,I329847);
nand I_23104 (I395509,I395492,I395246);
and I_23105 (I395526,I395328,I395509);
DFFARX1 I_23106  ( .D(I395526), .CLK(I2702), .RSTB(I395195), .Q(I395187) );
and I_23107 (I395160,I395492,I395461);
DFFARX1 I_23108  ( .D(I329853), .CLK(I2702), .RSTB(I395195), .Q(I395571) );
nor I_23109 (I395184,I395571,I395492);
nor I_23110 (I395602,I395571,I395246);
nand I_23111 (I395181,I395280,I395602);
not I_23112 (I395178,I395571);
DFFARX1 I_23113  ( .D(I329835), .CLK(I2702), .RSTB(I395195), .Q(I395647) );
not I_23114 (I395664,I395647);
nor I_23115 (I395681,I395664,I395345);
and I_23116 (I395698,I395571,I395681);
or I_23117 (I395715,I395492,I395698);
DFFARX1 I_23118  ( .D(I395715), .CLK(I2702), .RSTB(I395195), .Q(I395172) );
not I_23119 (I395746,I395664);
nor I_23120 (I395763,I395571,I395746);
nand I_23121 (I395175,I395664,I395763);
nand I_23122 (I395169,I395328,I395746);
not I_23123 (I395841,I2709);
not I_23124 (I395858,I548863);
nor I_23125 (I395875,I548875,I548869);
nand I_23126 (I395892,I395875,I548854);
nor I_23127 (I395909,I395858,I548875);
nand I_23128 (I395926,I395909,I548881);
DFFARX1 I_23129  ( .D(I395926), .CLK(I2702), .RSTB(I395841), .Q(I395943) );
not I_23130 (I395812,I395943);
not I_23131 (I395974,I548875);
not I_23132 (I395991,I395974);
not I_23133 (I396008,I548878);
nor I_23134 (I396025,I396008,I548860);
and I_23135 (I396042,I396025,I548857);
or I_23136 (I396059,I396042,I548884);
DFFARX1 I_23137  ( .D(I396059), .CLK(I2702), .RSTB(I395841), .Q(I396076) );
DFFARX1 I_23138  ( .D(I396076), .CLK(I2702), .RSTB(I395841), .Q(I395809) );
DFFARX1 I_23139  ( .D(I396076), .CLK(I2702), .RSTB(I395841), .Q(I396107) );
DFFARX1 I_23140  ( .D(I396076), .CLK(I2702), .RSTB(I395841), .Q(I395803) );
nand I_23141 (I396138,I395858,I548878);
nand I_23142 (I396155,I396138,I395892);
and I_23143 (I396172,I395974,I396155);
DFFARX1 I_23144  ( .D(I396172), .CLK(I2702), .RSTB(I395841), .Q(I395833) );
and I_23145 (I395806,I396138,I396107);
DFFARX1 I_23146  ( .D(I548872), .CLK(I2702), .RSTB(I395841), .Q(I396217) );
nor I_23147 (I395830,I396217,I396138);
nor I_23148 (I396248,I396217,I395892);
nand I_23149 (I395827,I395926,I396248);
not I_23150 (I395824,I396217);
DFFARX1 I_23151  ( .D(I548866), .CLK(I2702), .RSTB(I395841), .Q(I396293) );
not I_23152 (I396310,I396293);
nor I_23153 (I396327,I396310,I395991);
and I_23154 (I396344,I396217,I396327);
or I_23155 (I396361,I396138,I396344);
DFFARX1 I_23156  ( .D(I396361), .CLK(I2702), .RSTB(I395841), .Q(I395818) );
not I_23157 (I396392,I396310);
nor I_23158 (I396409,I396217,I396392);
nand I_23159 (I395821,I396310,I396409);
nand I_23160 (I395815,I395974,I396392);
not I_23161 (I396487,I2709);
not I_23162 (I396504,I321231);
nor I_23163 (I396521,I321210,I321222);
nand I_23164 (I396538,I396521,I321225);
nor I_23165 (I396555,I396504,I321210);
nand I_23166 (I396572,I396555,I321207);
DFFARX1 I_23167  ( .D(I396572), .CLK(I2702), .RSTB(I396487), .Q(I396589) );
not I_23168 (I396458,I396589);
not I_23169 (I396620,I321210);
not I_23170 (I396637,I396620);
not I_23171 (I396654,I321228);
nor I_23172 (I396671,I396654,I321219);
and I_23173 (I396688,I396671,I321213);
or I_23174 (I396705,I396688,I321237);
DFFARX1 I_23175  ( .D(I396705), .CLK(I2702), .RSTB(I396487), .Q(I396722) );
DFFARX1 I_23176  ( .D(I396722), .CLK(I2702), .RSTB(I396487), .Q(I396455) );
DFFARX1 I_23177  ( .D(I396722), .CLK(I2702), .RSTB(I396487), .Q(I396753) );
DFFARX1 I_23178  ( .D(I396722), .CLK(I2702), .RSTB(I396487), .Q(I396449) );
nand I_23179 (I396784,I396504,I321228);
nand I_23180 (I396801,I396784,I396538);
and I_23181 (I396818,I396620,I396801);
DFFARX1 I_23182  ( .D(I396818), .CLK(I2702), .RSTB(I396487), .Q(I396479) );
and I_23183 (I396452,I396784,I396753);
DFFARX1 I_23184  ( .D(I321234), .CLK(I2702), .RSTB(I396487), .Q(I396863) );
nor I_23185 (I396476,I396863,I396784);
nor I_23186 (I396894,I396863,I396538);
nand I_23187 (I396473,I396572,I396894);
not I_23188 (I396470,I396863);
DFFARX1 I_23189  ( .D(I321216), .CLK(I2702), .RSTB(I396487), .Q(I396939) );
not I_23190 (I396956,I396939);
nor I_23191 (I396973,I396956,I396637);
and I_23192 (I396990,I396863,I396973);
or I_23193 (I397007,I396784,I396990);
DFFARX1 I_23194  ( .D(I397007), .CLK(I2702), .RSTB(I396487), .Q(I396464) );
not I_23195 (I397038,I396956);
nor I_23196 (I397055,I396863,I397038);
nand I_23197 (I396467,I396956,I397055);
nand I_23198 (I396461,I396620,I397038);
not I_23199 (I397133,I2709);
not I_23200 (I397150,I35820);
nor I_23201 (I397167,I35835,I35829);
nand I_23202 (I397184,I397167,I35838);
nor I_23203 (I397201,I397150,I35835);
nand I_23204 (I397218,I397201,I35814);
DFFARX1 I_23205  ( .D(I397218), .CLK(I2702), .RSTB(I397133), .Q(I397235) );
not I_23206 (I397104,I397235);
not I_23207 (I397266,I35835);
not I_23208 (I397283,I397266);
not I_23209 (I397300,I35811);
nor I_23210 (I397317,I397300,I35826);
and I_23211 (I397334,I397317,I35832);
or I_23212 (I397351,I397334,I35841);
DFFARX1 I_23213  ( .D(I397351), .CLK(I2702), .RSTB(I397133), .Q(I397368) );
DFFARX1 I_23214  ( .D(I397368), .CLK(I2702), .RSTB(I397133), .Q(I397101) );
DFFARX1 I_23215  ( .D(I397368), .CLK(I2702), .RSTB(I397133), .Q(I397399) );
DFFARX1 I_23216  ( .D(I397368), .CLK(I2702), .RSTB(I397133), .Q(I397095) );
nand I_23217 (I397430,I397150,I35811);
nand I_23218 (I397447,I397430,I397184);
and I_23219 (I397464,I397266,I397447);
DFFARX1 I_23220  ( .D(I397464), .CLK(I2702), .RSTB(I397133), .Q(I397125) );
and I_23221 (I397098,I397430,I397399);
DFFARX1 I_23222  ( .D(I35823), .CLK(I2702), .RSTB(I397133), .Q(I397509) );
nor I_23223 (I397122,I397509,I397430);
nor I_23224 (I397540,I397509,I397184);
nand I_23225 (I397119,I397218,I397540);
not I_23226 (I397116,I397509);
DFFARX1 I_23227  ( .D(I35817), .CLK(I2702), .RSTB(I397133), .Q(I397585) );
not I_23228 (I397602,I397585);
nor I_23229 (I397619,I397602,I397283);
and I_23230 (I397636,I397509,I397619);
or I_23231 (I397653,I397430,I397636);
DFFARX1 I_23232  ( .D(I397653), .CLK(I2702), .RSTB(I397133), .Q(I397110) );
not I_23233 (I397684,I397602);
nor I_23234 (I397701,I397509,I397684);
nand I_23235 (I397113,I397602,I397701);
nand I_23236 (I397107,I397266,I397684);
not I_23237 (I397779,I2709);
not I_23238 (I397796,I616841);
nor I_23239 (I397813,I616838,I616823);
nand I_23240 (I397830,I397813,I616832);
nor I_23241 (I397847,I397796,I616838);
nand I_23242 (I397864,I397847,I616847);
DFFARX1 I_23243  ( .D(I397864), .CLK(I2702), .RSTB(I397779), .Q(I397881) );
not I_23244 (I397750,I397881);
not I_23245 (I397912,I616838);
not I_23246 (I397929,I397912);
not I_23247 (I397946,I616820);
nor I_23248 (I397963,I397946,I616826);
and I_23249 (I397980,I397963,I616850);
or I_23250 (I397997,I397980,I616844);
DFFARX1 I_23251  ( .D(I397997), .CLK(I2702), .RSTB(I397779), .Q(I398014) );
DFFARX1 I_23252  ( .D(I398014), .CLK(I2702), .RSTB(I397779), .Q(I397747) );
DFFARX1 I_23253  ( .D(I398014), .CLK(I2702), .RSTB(I397779), .Q(I398045) );
DFFARX1 I_23254  ( .D(I398014), .CLK(I2702), .RSTB(I397779), .Q(I397741) );
nand I_23255 (I398076,I397796,I616820);
nand I_23256 (I398093,I398076,I397830);
and I_23257 (I398110,I397912,I398093);
DFFARX1 I_23258  ( .D(I398110), .CLK(I2702), .RSTB(I397779), .Q(I397771) );
and I_23259 (I397744,I398076,I398045);
DFFARX1 I_23260  ( .D(I616829), .CLK(I2702), .RSTB(I397779), .Q(I398155) );
nor I_23261 (I397768,I398155,I398076);
nor I_23262 (I398186,I398155,I397830);
nand I_23263 (I397765,I397864,I398186);
not I_23264 (I397762,I398155);
DFFARX1 I_23265  ( .D(I616835), .CLK(I2702), .RSTB(I397779), .Q(I398231) );
not I_23266 (I398248,I398231);
nor I_23267 (I398265,I398248,I397929);
and I_23268 (I398282,I398155,I398265);
or I_23269 (I398299,I398076,I398282);
DFFARX1 I_23270  ( .D(I398299), .CLK(I2702), .RSTB(I397779), .Q(I397756) );
not I_23271 (I398330,I398248);
nor I_23272 (I398347,I398155,I398330);
nand I_23273 (I397759,I398248,I398347);
nand I_23274 (I397753,I397912,I398330);
not I_23275 (I398425,I2709);
not I_23276 (I398442,I687918);
nor I_23277 (I398459,I687915,I687900);
nand I_23278 (I398476,I398459,I687909);
nor I_23279 (I398493,I398442,I687915);
nand I_23280 (I398510,I398493,I687924);
DFFARX1 I_23281  ( .D(I398510), .CLK(I2702), .RSTB(I398425), .Q(I398527) );
not I_23282 (I398396,I398527);
not I_23283 (I398558,I687915);
not I_23284 (I398575,I398558);
not I_23285 (I398592,I687897);
nor I_23286 (I398609,I398592,I687903);
and I_23287 (I398626,I398609,I687927);
or I_23288 (I398643,I398626,I687921);
DFFARX1 I_23289  ( .D(I398643), .CLK(I2702), .RSTB(I398425), .Q(I398660) );
DFFARX1 I_23290  ( .D(I398660), .CLK(I2702), .RSTB(I398425), .Q(I398393) );
DFFARX1 I_23291  ( .D(I398660), .CLK(I2702), .RSTB(I398425), .Q(I398691) );
DFFARX1 I_23292  ( .D(I398660), .CLK(I2702), .RSTB(I398425), .Q(I398387) );
nand I_23293 (I398722,I398442,I687897);
nand I_23294 (I398739,I398722,I398476);
and I_23295 (I398756,I398558,I398739);
DFFARX1 I_23296  ( .D(I398756), .CLK(I2702), .RSTB(I398425), .Q(I398417) );
and I_23297 (I398390,I398722,I398691);
DFFARX1 I_23298  ( .D(I687906), .CLK(I2702), .RSTB(I398425), .Q(I398801) );
nor I_23299 (I398414,I398801,I398722);
nor I_23300 (I398832,I398801,I398476);
nand I_23301 (I398411,I398510,I398832);
not I_23302 (I398408,I398801);
DFFARX1 I_23303  ( .D(I687912), .CLK(I2702), .RSTB(I398425), .Q(I398877) );
not I_23304 (I398894,I398877);
nor I_23305 (I398911,I398894,I398575);
and I_23306 (I398928,I398801,I398911);
or I_23307 (I398945,I398722,I398928);
DFFARX1 I_23308  ( .D(I398945), .CLK(I2702), .RSTB(I398425), .Q(I398402) );
not I_23309 (I398976,I398894);
nor I_23310 (I398993,I398801,I398976);
nand I_23311 (I398405,I398894,I398993);
nand I_23312 (I398399,I398558,I398976);
not I_23313 (I399071,I2709);
not I_23314 (I399088,I4404);
nor I_23315 (I399105,I4419,I4413);
nand I_23316 (I399122,I399105,I4422);
nor I_23317 (I399139,I399088,I4419);
nand I_23318 (I399156,I399139,I4398);
DFFARX1 I_23319  ( .D(I399156), .CLK(I2702), .RSTB(I399071), .Q(I399173) );
not I_23320 (I399042,I399173);
not I_23321 (I399204,I4419);
not I_23322 (I399221,I399204);
not I_23323 (I399238,I4395);
nor I_23324 (I399255,I399238,I4410);
and I_23325 (I399272,I399255,I4416);
or I_23326 (I399289,I399272,I4425);
DFFARX1 I_23327  ( .D(I399289), .CLK(I2702), .RSTB(I399071), .Q(I399306) );
DFFARX1 I_23328  ( .D(I399306), .CLK(I2702), .RSTB(I399071), .Q(I399039) );
DFFARX1 I_23329  ( .D(I399306), .CLK(I2702), .RSTB(I399071), .Q(I399337) );
DFFARX1 I_23330  ( .D(I399306), .CLK(I2702), .RSTB(I399071), .Q(I399033) );
nand I_23331 (I399368,I399088,I4395);
nand I_23332 (I399385,I399368,I399122);
and I_23333 (I399402,I399204,I399385);
DFFARX1 I_23334  ( .D(I399402), .CLK(I2702), .RSTB(I399071), .Q(I399063) );
and I_23335 (I399036,I399368,I399337);
DFFARX1 I_23336  ( .D(I4407), .CLK(I2702), .RSTB(I399071), .Q(I399447) );
nor I_23337 (I399060,I399447,I399368);
nor I_23338 (I399478,I399447,I399122);
nand I_23339 (I399057,I399156,I399478);
not I_23340 (I399054,I399447);
DFFARX1 I_23341  ( .D(I4401), .CLK(I2702), .RSTB(I399071), .Q(I399523) );
not I_23342 (I399540,I399523);
nor I_23343 (I399557,I399540,I399221);
and I_23344 (I399574,I399447,I399557);
or I_23345 (I399591,I399368,I399574);
DFFARX1 I_23346  ( .D(I399591), .CLK(I2702), .RSTB(I399071), .Q(I399048) );
not I_23347 (I399622,I399540);
nor I_23348 (I399639,I399447,I399622);
nand I_23349 (I399051,I399540,I399639);
nand I_23350 (I399045,I399204,I399622);
not I_23351 (I399717,I2709);
not I_23352 (I399734,I76258);
nor I_23353 (I399751,I76249,I76240);
nand I_23354 (I399768,I399751,I76255);
nor I_23355 (I399785,I399734,I76249);
nand I_23356 (I399802,I399785,I76252);
DFFARX1 I_23357  ( .D(I399802), .CLK(I2702), .RSTB(I399717), .Q(I399819) );
not I_23358 (I399688,I399819);
not I_23359 (I399850,I76249);
not I_23360 (I399867,I399850);
not I_23361 (I399884,I76261);
nor I_23362 (I399901,I399884,I76246);
and I_23363 (I399918,I399901,I76264);
or I_23364 (I399935,I399918,I76237);
DFFARX1 I_23365  ( .D(I399935), .CLK(I2702), .RSTB(I399717), .Q(I399952) );
DFFARX1 I_23366  ( .D(I399952), .CLK(I2702), .RSTB(I399717), .Q(I399685) );
DFFARX1 I_23367  ( .D(I399952), .CLK(I2702), .RSTB(I399717), .Q(I399983) );
DFFARX1 I_23368  ( .D(I399952), .CLK(I2702), .RSTB(I399717), .Q(I399679) );
nand I_23369 (I400014,I399734,I76261);
nand I_23370 (I400031,I400014,I399768);
and I_23371 (I400048,I399850,I400031);
DFFARX1 I_23372  ( .D(I400048), .CLK(I2702), .RSTB(I399717), .Q(I399709) );
and I_23373 (I399682,I400014,I399983);
DFFARX1 I_23374  ( .D(I76267), .CLK(I2702), .RSTB(I399717), .Q(I400093) );
nor I_23375 (I399706,I400093,I400014);
nor I_23376 (I400124,I400093,I399768);
nand I_23377 (I399703,I399802,I400124);
not I_23378 (I399700,I400093);
DFFARX1 I_23379  ( .D(I76243), .CLK(I2702), .RSTB(I399717), .Q(I400169) );
not I_23380 (I400186,I400169);
nor I_23381 (I400203,I400186,I399867);
and I_23382 (I400220,I400093,I400203);
or I_23383 (I400237,I400014,I400220);
DFFARX1 I_23384  ( .D(I400237), .CLK(I2702), .RSTB(I399717), .Q(I399694) );
not I_23385 (I400268,I400186);
nor I_23386 (I400285,I400093,I400268);
nand I_23387 (I399697,I400186,I400285);
nand I_23388 (I399691,I399850,I400268);
not I_23389 (I400363,I2709);
not I_23390 (I400380,I331176);
nor I_23391 (I400397,I331155,I331167);
nand I_23392 (I400414,I400397,I331170);
nor I_23393 (I400431,I400380,I331155);
nand I_23394 (I400448,I400431,I331152);
DFFARX1 I_23395  ( .D(I400448), .CLK(I2702), .RSTB(I400363), .Q(I400465) );
not I_23396 (I400334,I400465);
not I_23397 (I400496,I331155);
not I_23398 (I400513,I400496);
not I_23399 (I400530,I331173);
nor I_23400 (I400547,I400530,I331164);
and I_23401 (I400564,I400547,I331158);
or I_23402 (I400581,I400564,I331182);
DFFARX1 I_23403  ( .D(I400581), .CLK(I2702), .RSTB(I400363), .Q(I400598) );
DFFARX1 I_23404  ( .D(I400598), .CLK(I2702), .RSTB(I400363), .Q(I400331) );
DFFARX1 I_23405  ( .D(I400598), .CLK(I2702), .RSTB(I400363), .Q(I400629) );
DFFARX1 I_23406  ( .D(I400598), .CLK(I2702), .RSTB(I400363), .Q(I400325) );
nand I_23407 (I400660,I400380,I331173);
nand I_23408 (I400677,I400660,I400414);
and I_23409 (I400694,I400496,I400677);
DFFARX1 I_23410  ( .D(I400694), .CLK(I2702), .RSTB(I400363), .Q(I400355) );
and I_23411 (I400328,I400660,I400629);
DFFARX1 I_23412  ( .D(I331179), .CLK(I2702), .RSTB(I400363), .Q(I400739) );
nor I_23413 (I400352,I400739,I400660);
nor I_23414 (I400770,I400739,I400414);
nand I_23415 (I400349,I400448,I400770);
not I_23416 (I400346,I400739);
DFFARX1 I_23417  ( .D(I331161), .CLK(I2702), .RSTB(I400363), .Q(I400815) );
not I_23418 (I400832,I400815);
nor I_23419 (I400849,I400832,I400513);
and I_23420 (I400866,I400739,I400849);
or I_23421 (I400883,I400660,I400866);
DFFARX1 I_23422  ( .D(I400883), .CLK(I2702), .RSTB(I400363), .Q(I400340) );
not I_23423 (I400914,I400832);
nor I_23424 (I400931,I400739,I400914);
nand I_23425 (I400343,I400832,I400931);
nand I_23426 (I400337,I400496,I400914);
not I_23427 (I401009,I2709);
not I_23428 (I401026,I569093);
nor I_23429 (I401043,I569105,I569099);
nand I_23430 (I401060,I401043,I569084);
nor I_23431 (I401077,I401026,I569105);
nand I_23432 (I401094,I401077,I569111);
DFFARX1 I_23433  ( .D(I401094), .CLK(I2702), .RSTB(I401009), .Q(I401111) );
not I_23434 (I400980,I401111);
not I_23435 (I401142,I569105);
not I_23436 (I401159,I401142);
not I_23437 (I401176,I569108);
nor I_23438 (I401193,I401176,I569090);
and I_23439 (I401210,I401193,I569087);
or I_23440 (I401227,I401210,I569114);
DFFARX1 I_23441  ( .D(I401227), .CLK(I2702), .RSTB(I401009), .Q(I401244) );
DFFARX1 I_23442  ( .D(I401244), .CLK(I2702), .RSTB(I401009), .Q(I400977) );
DFFARX1 I_23443  ( .D(I401244), .CLK(I2702), .RSTB(I401009), .Q(I401275) );
DFFARX1 I_23444  ( .D(I401244), .CLK(I2702), .RSTB(I401009), .Q(I400971) );
nand I_23445 (I401306,I401026,I569108);
nand I_23446 (I401323,I401306,I401060);
and I_23447 (I401340,I401142,I401323);
DFFARX1 I_23448  ( .D(I401340), .CLK(I2702), .RSTB(I401009), .Q(I401001) );
and I_23449 (I400974,I401306,I401275);
DFFARX1 I_23450  ( .D(I569102), .CLK(I2702), .RSTB(I401009), .Q(I401385) );
nor I_23451 (I400998,I401385,I401306);
nor I_23452 (I401416,I401385,I401060);
nand I_23453 (I400995,I401094,I401416);
not I_23454 (I400992,I401385);
DFFARX1 I_23455  ( .D(I569096), .CLK(I2702), .RSTB(I401009), .Q(I401461) );
not I_23456 (I401478,I401461);
nor I_23457 (I401495,I401478,I401159);
and I_23458 (I401512,I401385,I401495);
or I_23459 (I401529,I401306,I401512);
DFFARX1 I_23460  ( .D(I401529), .CLK(I2702), .RSTB(I401009), .Q(I400986) );
not I_23461 (I401560,I401478);
nor I_23462 (I401577,I401385,I401560);
nand I_23463 (I400989,I401478,I401577);
nand I_23464 (I400983,I401142,I401560);
not I_23465 (I401655,I2709);
not I_23466 (I401672,I28527);
nor I_23467 (I401689,I28542,I28536);
nand I_23468 (I401706,I401689,I28545);
nor I_23469 (I401723,I401672,I28542);
nand I_23470 (I401740,I401723,I28521);
DFFARX1 I_23471  ( .D(I401740), .CLK(I2702), .RSTB(I401655), .Q(I401757) );
not I_23472 (I401626,I401757);
not I_23473 (I401788,I28542);
not I_23474 (I401805,I401788);
not I_23475 (I401822,I28518);
nor I_23476 (I401839,I401822,I28533);
and I_23477 (I401856,I401839,I28539);
or I_23478 (I401873,I401856,I28548);
DFFARX1 I_23479  ( .D(I401873), .CLK(I2702), .RSTB(I401655), .Q(I401890) );
DFFARX1 I_23480  ( .D(I401890), .CLK(I2702), .RSTB(I401655), .Q(I401623) );
DFFARX1 I_23481  ( .D(I401890), .CLK(I2702), .RSTB(I401655), .Q(I401921) );
DFFARX1 I_23482  ( .D(I401890), .CLK(I2702), .RSTB(I401655), .Q(I401617) );
nand I_23483 (I401952,I401672,I28518);
nand I_23484 (I401969,I401952,I401706);
and I_23485 (I401986,I401788,I401969);
DFFARX1 I_23486  ( .D(I401986), .CLK(I2702), .RSTB(I401655), .Q(I401647) );
and I_23487 (I401620,I401952,I401921);
DFFARX1 I_23488  ( .D(I28530), .CLK(I2702), .RSTB(I401655), .Q(I402031) );
nor I_23489 (I401644,I402031,I401952);
nor I_23490 (I402062,I402031,I401706);
nand I_23491 (I401641,I401740,I402062);
not I_23492 (I401638,I402031);
DFFARX1 I_23493  ( .D(I28524), .CLK(I2702), .RSTB(I401655), .Q(I402107) );
not I_23494 (I402124,I402107);
nor I_23495 (I402141,I402124,I401805);
and I_23496 (I402158,I402031,I402141);
or I_23497 (I402175,I401952,I402158);
DFFARX1 I_23498  ( .D(I402175), .CLK(I2702), .RSTB(I401655), .Q(I401632) );
not I_23499 (I402206,I402124);
nor I_23500 (I402223,I402031,I402206);
nand I_23501 (I401635,I402124,I402223);
nand I_23502 (I401629,I401788,I402206);
not I_23503 (I402301,I2709);
not I_23504 (I402318,I483572);
nor I_23505 (I402335,I483575,I483557);
nand I_23506 (I402352,I402335,I483584);
nor I_23507 (I402369,I402318,I483575);
nand I_23508 (I402386,I402369,I483563);
DFFARX1 I_23509  ( .D(I402386), .CLK(I2702), .RSTB(I402301), .Q(I402403) );
not I_23510 (I402272,I402403);
not I_23511 (I402434,I483575);
not I_23512 (I402451,I402434);
not I_23513 (I402468,I483569);
nor I_23514 (I402485,I402468,I483581);
and I_23515 (I402502,I402485,I483587);
or I_23516 (I402519,I402502,I483566);
DFFARX1 I_23517  ( .D(I402519), .CLK(I2702), .RSTB(I402301), .Q(I402536) );
DFFARX1 I_23518  ( .D(I402536), .CLK(I2702), .RSTB(I402301), .Q(I402269) );
DFFARX1 I_23519  ( .D(I402536), .CLK(I2702), .RSTB(I402301), .Q(I402567) );
DFFARX1 I_23520  ( .D(I402536), .CLK(I2702), .RSTB(I402301), .Q(I402263) );
nand I_23521 (I402598,I402318,I483569);
nand I_23522 (I402615,I402598,I402352);
and I_23523 (I402632,I402434,I402615);
DFFARX1 I_23524  ( .D(I402632), .CLK(I2702), .RSTB(I402301), .Q(I402293) );
and I_23525 (I402266,I402598,I402567);
DFFARX1 I_23526  ( .D(I483578), .CLK(I2702), .RSTB(I402301), .Q(I402677) );
nor I_23527 (I402290,I402677,I402598);
nor I_23528 (I402708,I402677,I402352);
nand I_23529 (I402287,I402386,I402708);
not I_23530 (I402284,I402677);
DFFARX1 I_23531  ( .D(I483560), .CLK(I2702), .RSTB(I402301), .Q(I402753) );
not I_23532 (I402770,I402753);
nor I_23533 (I402787,I402770,I402451);
and I_23534 (I402804,I402677,I402787);
or I_23535 (I402821,I402598,I402804);
DFFARX1 I_23536  ( .D(I402821), .CLK(I2702), .RSTB(I402301), .Q(I402278) );
not I_23537 (I402852,I402770);
nor I_23538 (I402869,I402677,I402852);
nand I_23539 (I402281,I402770,I402869);
nand I_23540 (I402275,I402434,I402852);
not I_23541 (I402947,I2709);
not I_23542 (I402964,I166068);
nor I_23543 (I402981,I166089,I166071);
nand I_23544 (I402998,I402981,I166095);
nor I_23545 (I403015,I402964,I166089);
nand I_23546 (I403032,I403015,I166092);
DFFARX1 I_23547  ( .D(I403032), .CLK(I2702), .RSTB(I402947), .Q(I403049) );
not I_23548 (I402918,I403049);
not I_23549 (I403080,I166089);
not I_23550 (I403097,I403080);
not I_23551 (I403114,I166086);
nor I_23552 (I403131,I403114,I166065);
and I_23553 (I403148,I403131,I166077);
or I_23554 (I403165,I403148,I166074);
DFFARX1 I_23555  ( .D(I403165), .CLK(I2702), .RSTB(I402947), .Q(I403182) );
DFFARX1 I_23556  ( .D(I403182), .CLK(I2702), .RSTB(I402947), .Q(I402915) );
DFFARX1 I_23557  ( .D(I403182), .CLK(I2702), .RSTB(I402947), .Q(I403213) );
DFFARX1 I_23558  ( .D(I403182), .CLK(I2702), .RSTB(I402947), .Q(I402909) );
nand I_23559 (I403244,I402964,I166086);
nand I_23560 (I403261,I403244,I402998);
and I_23561 (I403278,I403080,I403261);
DFFARX1 I_23562  ( .D(I403278), .CLK(I2702), .RSTB(I402947), .Q(I402939) );
and I_23563 (I402912,I403244,I403213);
DFFARX1 I_23564  ( .D(I166080), .CLK(I2702), .RSTB(I402947), .Q(I403323) );
nor I_23565 (I402936,I403323,I403244);
nor I_23566 (I403354,I403323,I402998);
nand I_23567 (I402933,I403032,I403354);
not I_23568 (I402930,I403323);
DFFARX1 I_23569  ( .D(I166083), .CLK(I2702), .RSTB(I402947), .Q(I403399) );
not I_23570 (I403416,I403399);
nor I_23571 (I403433,I403416,I403097);
and I_23572 (I403450,I403323,I403433);
or I_23573 (I403467,I403244,I403450);
DFFARX1 I_23574  ( .D(I403467), .CLK(I2702), .RSTB(I402947), .Q(I402924) );
not I_23575 (I403498,I403416);
nor I_23576 (I403515,I403323,I403498);
nand I_23577 (I402927,I403416,I403515);
nand I_23578 (I402921,I403080,I403498);
not I_23579 (I403593,I2709);
not I_23580 (I403610,I122124);
nor I_23581 (I403627,I122115,I122106);
nand I_23582 (I403644,I403627,I122121);
nor I_23583 (I403661,I403610,I122115);
nand I_23584 (I403678,I403661,I122118);
DFFARX1 I_23585  ( .D(I403678), .CLK(I2702), .RSTB(I403593), .Q(I403695) );
not I_23586 (I403564,I403695);
not I_23587 (I403726,I122115);
not I_23588 (I403743,I403726);
not I_23589 (I403760,I122127);
nor I_23590 (I403777,I403760,I122112);
and I_23591 (I403794,I403777,I122130);
or I_23592 (I403811,I403794,I122103);
DFFARX1 I_23593  ( .D(I403811), .CLK(I2702), .RSTB(I403593), .Q(I403828) );
DFFARX1 I_23594  ( .D(I403828), .CLK(I2702), .RSTB(I403593), .Q(I403561) );
DFFARX1 I_23595  ( .D(I403828), .CLK(I2702), .RSTB(I403593), .Q(I403859) );
DFFARX1 I_23596  ( .D(I403828), .CLK(I2702), .RSTB(I403593), .Q(I403555) );
nand I_23597 (I403890,I403610,I122127);
nand I_23598 (I403907,I403890,I403644);
and I_23599 (I403924,I403726,I403907);
DFFARX1 I_23600  ( .D(I403924), .CLK(I2702), .RSTB(I403593), .Q(I403585) );
and I_23601 (I403558,I403890,I403859);
DFFARX1 I_23602  ( .D(I122133), .CLK(I2702), .RSTB(I403593), .Q(I403969) );
nor I_23603 (I403582,I403969,I403890);
nor I_23604 (I404000,I403969,I403644);
nand I_23605 (I403579,I403678,I404000);
not I_23606 (I403576,I403969);
DFFARX1 I_23607  ( .D(I122109), .CLK(I2702), .RSTB(I403593), .Q(I404045) );
not I_23608 (I404062,I404045);
nor I_23609 (I404079,I404062,I403743);
and I_23610 (I404096,I403969,I404079);
or I_23611 (I404113,I403890,I404096);
DFFARX1 I_23612  ( .D(I404113), .CLK(I2702), .RSTB(I403593), .Q(I403570) );
not I_23613 (I404144,I404062);
nor I_23614 (I404161,I403969,I404144);
nand I_23615 (I403573,I404062,I404161);
nand I_23616 (I403567,I403726,I404144);
not I_23617 (I404239,I2709);
not I_23618 (I404256,I627534);
nor I_23619 (I404273,I627531,I627516);
nand I_23620 (I404290,I404273,I627525);
nor I_23621 (I404307,I404256,I627531);
nand I_23622 (I404324,I404307,I627540);
DFFARX1 I_23623  ( .D(I404324), .CLK(I2702), .RSTB(I404239), .Q(I404341) );
not I_23624 (I404210,I404341);
not I_23625 (I404372,I627531);
not I_23626 (I404389,I404372);
not I_23627 (I404406,I627513);
nor I_23628 (I404423,I404406,I627519);
and I_23629 (I404440,I404423,I627543);
or I_23630 (I404457,I404440,I627537);
DFFARX1 I_23631  ( .D(I404457), .CLK(I2702), .RSTB(I404239), .Q(I404474) );
DFFARX1 I_23632  ( .D(I404474), .CLK(I2702), .RSTB(I404239), .Q(I404207) );
DFFARX1 I_23633  ( .D(I404474), .CLK(I2702), .RSTB(I404239), .Q(I404505) );
DFFARX1 I_23634  ( .D(I404474), .CLK(I2702), .RSTB(I404239), .Q(I404201) );
nand I_23635 (I404536,I404256,I627513);
nand I_23636 (I404553,I404536,I404290);
and I_23637 (I404570,I404372,I404553);
DFFARX1 I_23638  ( .D(I404570), .CLK(I2702), .RSTB(I404239), .Q(I404231) );
and I_23639 (I404204,I404536,I404505);
DFFARX1 I_23640  ( .D(I627522), .CLK(I2702), .RSTB(I404239), .Q(I404615) );
nor I_23641 (I404228,I404615,I404536);
nor I_23642 (I404646,I404615,I404290);
nand I_23643 (I404225,I404324,I404646);
not I_23644 (I404222,I404615);
DFFARX1 I_23645  ( .D(I627528), .CLK(I2702), .RSTB(I404239), .Q(I404691) );
not I_23646 (I404708,I404691);
nor I_23647 (I404725,I404708,I404389);
and I_23648 (I404742,I404615,I404725);
or I_23649 (I404759,I404536,I404742);
DFFARX1 I_23650  ( .D(I404759), .CLK(I2702), .RSTB(I404239), .Q(I404216) );
not I_23651 (I404790,I404708);
nor I_23652 (I404807,I404615,I404790);
nand I_23653 (I404219,I404708,I404807);
nand I_23654 (I404213,I404372,I404790);
not I_23655 (I404885,I2709);
not I_23656 (I404902,I639485);
nor I_23657 (I404919,I639482,I639467);
nand I_23658 (I404936,I404919,I639476);
nor I_23659 (I404953,I404902,I639482);
nand I_23660 (I404970,I404953,I639491);
DFFARX1 I_23661  ( .D(I404970), .CLK(I2702), .RSTB(I404885), .Q(I404987) );
not I_23662 (I404856,I404987);
not I_23663 (I405018,I639482);
not I_23664 (I405035,I405018);
not I_23665 (I405052,I639464);
nor I_23666 (I405069,I405052,I639470);
and I_23667 (I405086,I405069,I639494);
or I_23668 (I405103,I405086,I639488);
DFFARX1 I_23669  ( .D(I405103), .CLK(I2702), .RSTB(I404885), .Q(I405120) );
DFFARX1 I_23670  ( .D(I405120), .CLK(I2702), .RSTB(I404885), .Q(I404853) );
DFFARX1 I_23671  ( .D(I405120), .CLK(I2702), .RSTB(I404885), .Q(I405151) );
DFFARX1 I_23672  ( .D(I405120), .CLK(I2702), .RSTB(I404885), .Q(I404847) );
nand I_23673 (I405182,I404902,I639464);
nand I_23674 (I405199,I405182,I404936);
and I_23675 (I405216,I405018,I405199);
DFFARX1 I_23676  ( .D(I405216), .CLK(I2702), .RSTB(I404885), .Q(I404877) );
and I_23677 (I404850,I405182,I405151);
DFFARX1 I_23678  ( .D(I639473), .CLK(I2702), .RSTB(I404885), .Q(I405261) );
nor I_23679 (I404874,I405261,I405182);
nor I_23680 (I405292,I405261,I404936);
nand I_23681 (I404871,I404970,I405292);
not I_23682 (I404868,I405261);
DFFARX1 I_23683  ( .D(I639479), .CLK(I2702), .RSTB(I404885), .Q(I405337) );
not I_23684 (I405354,I405337);
nor I_23685 (I405371,I405354,I405035);
and I_23686 (I405388,I405261,I405371);
or I_23687 (I405405,I405182,I405388);
DFFARX1 I_23688  ( .D(I405405), .CLK(I2702), .RSTB(I404885), .Q(I404862) );
not I_23689 (I405436,I405354);
nor I_23690 (I405453,I405261,I405436);
nand I_23691 (I404865,I405354,I405453);
nand I_23692 (I404859,I405018,I405436);
not I_23693 (I405531,I2709);
not I_23694 (I405548,I611347);
nor I_23695 (I405565,I611335,I611344);
nand I_23696 (I405582,I405565,I611359);
nor I_23697 (I405599,I405548,I611335);
nand I_23698 (I405616,I405599,I611341);
DFFARX1 I_23699  ( .D(I405616), .CLK(I2702), .RSTB(I405531), .Q(I405633) );
not I_23700 (I405502,I405633);
not I_23701 (I405664,I611335);
not I_23702 (I405681,I405664);
not I_23703 (I405698,I611329);
nor I_23704 (I405715,I405698,I611350);
and I_23705 (I405732,I405715,I611332);
or I_23706 (I405749,I405732,I611338);
DFFARX1 I_23707  ( .D(I405749), .CLK(I2702), .RSTB(I405531), .Q(I405766) );
DFFARX1 I_23708  ( .D(I405766), .CLK(I2702), .RSTB(I405531), .Q(I405499) );
DFFARX1 I_23709  ( .D(I405766), .CLK(I2702), .RSTB(I405531), .Q(I405797) );
DFFARX1 I_23710  ( .D(I405766), .CLK(I2702), .RSTB(I405531), .Q(I405493) );
nand I_23711 (I405828,I405548,I611329);
nand I_23712 (I405845,I405828,I405582);
and I_23713 (I405862,I405664,I405845);
DFFARX1 I_23714  ( .D(I405862), .CLK(I2702), .RSTB(I405531), .Q(I405523) );
and I_23715 (I405496,I405828,I405797);
DFFARX1 I_23716  ( .D(I611356), .CLK(I2702), .RSTB(I405531), .Q(I405907) );
nor I_23717 (I405520,I405907,I405828);
nor I_23718 (I405938,I405907,I405582);
nand I_23719 (I405517,I405616,I405938);
not I_23720 (I405514,I405907);
DFFARX1 I_23721  ( .D(I611353), .CLK(I2702), .RSTB(I405531), .Q(I405983) );
not I_23722 (I406000,I405983);
nor I_23723 (I406017,I406000,I405681);
and I_23724 (I406034,I405907,I406017);
or I_23725 (I406051,I405828,I406034);
DFFARX1 I_23726  ( .D(I406051), .CLK(I2702), .RSTB(I405531), .Q(I405508) );
not I_23727 (I406082,I406000);
nor I_23728 (I406099,I405907,I406082);
nand I_23729 (I405511,I406000,I406099);
nand I_23730 (I405505,I405664,I406082);
not I_23731 (I406177,I2709);
not I_23732 (I406194,I156123);
nor I_23733 (I406211,I156144,I156126);
nand I_23734 (I406228,I406211,I156150);
nor I_23735 (I406245,I406194,I156144);
nand I_23736 (I406262,I406245,I156147);
DFFARX1 I_23737  ( .D(I406262), .CLK(I2702), .RSTB(I406177), .Q(I406279) );
not I_23738 (I406148,I406279);
not I_23739 (I406310,I156144);
not I_23740 (I406327,I406310);
not I_23741 (I406344,I156141);
nor I_23742 (I406361,I406344,I156120);
and I_23743 (I406378,I406361,I156132);
or I_23744 (I406395,I406378,I156129);
DFFARX1 I_23745  ( .D(I406395), .CLK(I2702), .RSTB(I406177), .Q(I406412) );
DFFARX1 I_23746  ( .D(I406412), .CLK(I2702), .RSTB(I406177), .Q(I406145) );
DFFARX1 I_23747  ( .D(I406412), .CLK(I2702), .RSTB(I406177), .Q(I406443) );
DFFARX1 I_23748  ( .D(I406412), .CLK(I2702), .RSTB(I406177), .Q(I406139) );
nand I_23749 (I406474,I406194,I156141);
nand I_23750 (I406491,I406474,I406228);
and I_23751 (I406508,I406310,I406491);
DFFARX1 I_23752  ( .D(I406508), .CLK(I2702), .RSTB(I406177), .Q(I406169) );
and I_23753 (I406142,I406474,I406443);
DFFARX1 I_23754  ( .D(I156135), .CLK(I2702), .RSTB(I406177), .Q(I406553) );
nor I_23755 (I406166,I406553,I406474);
nor I_23756 (I406584,I406553,I406228);
nand I_23757 (I406163,I406262,I406584);
not I_23758 (I406160,I406553);
DFFARX1 I_23759  ( .D(I156138), .CLK(I2702), .RSTB(I406177), .Q(I406629) );
not I_23760 (I406646,I406629);
nor I_23761 (I406663,I406646,I406327);
and I_23762 (I406680,I406553,I406663);
or I_23763 (I406697,I406474,I406680);
DFFARX1 I_23764  ( .D(I406697), .CLK(I2702), .RSTB(I406177), .Q(I406154) );
not I_23765 (I406728,I406646);
nor I_23766 (I406745,I406553,I406728);
nand I_23767 (I406157,I406646,I406745);
nand I_23768 (I406151,I406310,I406728);
not I_23769 (I406823,I2709);
not I_23770 (I406840,I715812);
nor I_23771 (I406857,I715797,I715803);
nand I_23772 (I406874,I406857,I715800);
nor I_23773 (I406891,I406840,I715797);
nand I_23774 (I406908,I406891,I715809);
DFFARX1 I_23775  ( .D(I406908), .CLK(I2702), .RSTB(I406823), .Q(I406925) );
not I_23776 (I406794,I406925);
not I_23777 (I406956,I715797);
not I_23778 (I406973,I406956);
not I_23779 (I406990,I715824);
nor I_23780 (I407007,I406990,I715818);
and I_23781 (I407024,I407007,I715815);
or I_23782 (I407041,I407024,I715794);
DFFARX1 I_23783  ( .D(I407041), .CLK(I2702), .RSTB(I406823), .Q(I407058) );
DFFARX1 I_23784  ( .D(I407058), .CLK(I2702), .RSTB(I406823), .Q(I406791) );
DFFARX1 I_23785  ( .D(I407058), .CLK(I2702), .RSTB(I406823), .Q(I407089) );
DFFARX1 I_23786  ( .D(I407058), .CLK(I2702), .RSTB(I406823), .Q(I406785) );
nand I_23787 (I407120,I406840,I715824);
nand I_23788 (I407137,I407120,I406874);
and I_23789 (I407154,I406956,I407137);
DFFARX1 I_23790  ( .D(I407154), .CLK(I2702), .RSTB(I406823), .Q(I406815) );
and I_23791 (I406788,I407120,I407089);
DFFARX1 I_23792  ( .D(I715821), .CLK(I2702), .RSTB(I406823), .Q(I407199) );
nor I_23793 (I406812,I407199,I407120);
nor I_23794 (I407230,I407199,I406874);
nand I_23795 (I406809,I406908,I407230);
not I_23796 (I406806,I407199);
DFFARX1 I_23797  ( .D(I715806), .CLK(I2702), .RSTB(I406823), .Q(I407275) );
not I_23798 (I407292,I407275);
nor I_23799 (I407309,I407292,I406973);
and I_23800 (I407326,I407199,I407309);
or I_23801 (I407343,I407120,I407326);
DFFARX1 I_23802  ( .D(I407343), .CLK(I2702), .RSTB(I406823), .Q(I406800) );
not I_23803 (I407374,I407292);
nor I_23804 (I407391,I407199,I407374);
nand I_23805 (I406803,I407292,I407391);
nand I_23806 (I406797,I406956,I407374);
not I_23807 (I407469,I2709);
not I_23808 (I407486,I20673);
nor I_23809 (I407503,I20688,I20682);
nand I_23810 (I407520,I407503,I20691);
nor I_23811 (I407537,I407486,I20688);
nand I_23812 (I407554,I407537,I20667);
DFFARX1 I_23813  ( .D(I407554), .CLK(I2702), .RSTB(I407469), .Q(I407571) );
not I_23814 (I407440,I407571);
not I_23815 (I407602,I20688);
not I_23816 (I407619,I407602);
not I_23817 (I407636,I20664);
nor I_23818 (I407653,I407636,I20679);
and I_23819 (I407670,I407653,I20685);
or I_23820 (I407687,I407670,I20694);
DFFARX1 I_23821  ( .D(I407687), .CLK(I2702), .RSTB(I407469), .Q(I407704) );
DFFARX1 I_23822  ( .D(I407704), .CLK(I2702), .RSTB(I407469), .Q(I407437) );
DFFARX1 I_23823  ( .D(I407704), .CLK(I2702), .RSTB(I407469), .Q(I407735) );
DFFARX1 I_23824  ( .D(I407704), .CLK(I2702), .RSTB(I407469), .Q(I407431) );
nand I_23825 (I407766,I407486,I20664);
nand I_23826 (I407783,I407766,I407520);
and I_23827 (I407800,I407602,I407783);
DFFARX1 I_23828  ( .D(I407800), .CLK(I2702), .RSTB(I407469), .Q(I407461) );
and I_23829 (I407434,I407766,I407735);
DFFARX1 I_23830  ( .D(I20676), .CLK(I2702), .RSTB(I407469), .Q(I407845) );
nor I_23831 (I407458,I407845,I407766);
nor I_23832 (I407876,I407845,I407520);
nand I_23833 (I407455,I407554,I407876);
not I_23834 (I407452,I407845);
DFFARX1 I_23835  ( .D(I20670), .CLK(I2702), .RSTB(I407469), .Q(I407921) );
not I_23836 (I407938,I407921);
nor I_23837 (I407955,I407938,I407619);
and I_23838 (I407972,I407845,I407955);
or I_23839 (I407989,I407766,I407972);
DFFARX1 I_23840  ( .D(I407989), .CLK(I2702), .RSTB(I407469), .Q(I407446) );
not I_23841 (I408020,I407938);
nor I_23842 (I408037,I407845,I408020);
nand I_23843 (I407449,I407938,I408037);
nand I_23844 (I407443,I407602,I408020);
not I_23845 (I408115,I2709);
not I_23846 (I408132,I21795);
nor I_23847 (I408149,I21810,I21804);
nand I_23848 (I408166,I408149,I21813);
nor I_23849 (I408183,I408132,I21810);
nand I_23850 (I408200,I408183,I21789);
DFFARX1 I_23851  ( .D(I408200), .CLK(I2702), .RSTB(I408115), .Q(I408217) );
not I_23852 (I408086,I408217);
not I_23853 (I408248,I21810);
not I_23854 (I408265,I408248);
not I_23855 (I408282,I21786);
nor I_23856 (I408299,I408282,I21801);
and I_23857 (I408316,I408299,I21807);
or I_23858 (I408333,I408316,I21816);
DFFARX1 I_23859  ( .D(I408333), .CLK(I2702), .RSTB(I408115), .Q(I408350) );
DFFARX1 I_23860  ( .D(I408350), .CLK(I2702), .RSTB(I408115), .Q(I408083) );
DFFARX1 I_23861  ( .D(I408350), .CLK(I2702), .RSTB(I408115), .Q(I408381) );
DFFARX1 I_23862  ( .D(I408350), .CLK(I2702), .RSTB(I408115), .Q(I408077) );
nand I_23863 (I408412,I408132,I21786);
nand I_23864 (I408429,I408412,I408166);
and I_23865 (I408446,I408248,I408429);
DFFARX1 I_23866  ( .D(I408446), .CLK(I2702), .RSTB(I408115), .Q(I408107) );
and I_23867 (I408080,I408412,I408381);
DFFARX1 I_23868  ( .D(I21798), .CLK(I2702), .RSTB(I408115), .Q(I408491) );
nor I_23869 (I408104,I408491,I408412);
nor I_23870 (I408522,I408491,I408166);
nand I_23871 (I408101,I408200,I408522);
not I_23872 (I408098,I408491);
DFFARX1 I_23873  ( .D(I21792), .CLK(I2702), .RSTB(I408115), .Q(I408567) );
not I_23874 (I408584,I408567);
nor I_23875 (I408601,I408584,I408265);
and I_23876 (I408618,I408491,I408601);
or I_23877 (I408635,I408412,I408618);
DFFARX1 I_23878  ( .D(I408635), .CLK(I2702), .RSTB(I408115), .Q(I408092) );
not I_23879 (I408666,I408584);
nor I_23880 (I408683,I408491,I408666);
nand I_23881 (I408095,I408584,I408683);
nand I_23882 (I408089,I408248,I408666);
not I_23883 (I408761,I2709);
not I_23884 (I408778,I191925);
nor I_23885 (I408795,I191946,I191928);
nand I_23886 (I408812,I408795,I191952);
nor I_23887 (I408829,I408778,I191946);
nand I_23888 (I408846,I408829,I191949);
DFFARX1 I_23889  ( .D(I408846), .CLK(I2702), .RSTB(I408761), .Q(I408863) );
not I_23890 (I408732,I408863);
not I_23891 (I408894,I191946);
not I_23892 (I408911,I408894);
not I_23893 (I408928,I191943);
nor I_23894 (I408945,I408928,I191922);
and I_23895 (I408962,I408945,I191934);
or I_23896 (I408979,I408962,I191931);
DFFARX1 I_23897  ( .D(I408979), .CLK(I2702), .RSTB(I408761), .Q(I408996) );
DFFARX1 I_23898  ( .D(I408996), .CLK(I2702), .RSTB(I408761), .Q(I408729) );
DFFARX1 I_23899  ( .D(I408996), .CLK(I2702), .RSTB(I408761), .Q(I409027) );
DFFARX1 I_23900  ( .D(I408996), .CLK(I2702), .RSTB(I408761), .Q(I408723) );
nand I_23901 (I409058,I408778,I191943);
nand I_23902 (I409075,I409058,I408812);
and I_23903 (I409092,I408894,I409075);
DFFARX1 I_23904  ( .D(I409092), .CLK(I2702), .RSTB(I408761), .Q(I408753) );
and I_23905 (I408726,I409058,I409027);
DFFARX1 I_23906  ( .D(I191937), .CLK(I2702), .RSTB(I408761), .Q(I409137) );
nor I_23907 (I408750,I409137,I409058);
nor I_23908 (I409168,I409137,I408812);
nand I_23909 (I408747,I408846,I409168);
not I_23910 (I408744,I409137);
DFFARX1 I_23911  ( .D(I191940), .CLK(I2702), .RSTB(I408761), .Q(I409213) );
not I_23912 (I409230,I409213);
nor I_23913 (I409247,I409230,I408911);
and I_23914 (I409264,I409137,I409247);
or I_23915 (I409281,I409058,I409264);
DFFARX1 I_23916  ( .D(I409281), .CLK(I2702), .RSTB(I408761), .Q(I408738) );
not I_23917 (I409312,I409230);
nor I_23918 (I409329,I409137,I409312);
nand I_23919 (I408741,I409230,I409329);
nand I_23920 (I408735,I408894,I409312);
not I_23921 (I409407,I2709);
not I_23922 (I409424,I605992);
nor I_23923 (I409441,I605980,I605989);
nand I_23924 (I409458,I409441,I606004);
nor I_23925 (I409475,I409424,I605980);
nand I_23926 (I409492,I409475,I605986);
DFFARX1 I_23927  ( .D(I409492), .CLK(I2702), .RSTB(I409407), .Q(I409509) );
not I_23928 (I409378,I409509);
not I_23929 (I409540,I605980);
not I_23930 (I409557,I409540);
not I_23931 (I409574,I605974);
nor I_23932 (I409591,I409574,I605995);
and I_23933 (I409608,I409591,I605977);
or I_23934 (I409625,I409608,I605983);
DFFARX1 I_23935  ( .D(I409625), .CLK(I2702), .RSTB(I409407), .Q(I409642) );
DFFARX1 I_23936  ( .D(I409642), .CLK(I2702), .RSTB(I409407), .Q(I409375) );
DFFARX1 I_23937  ( .D(I409642), .CLK(I2702), .RSTB(I409407), .Q(I409673) );
DFFARX1 I_23938  ( .D(I409642), .CLK(I2702), .RSTB(I409407), .Q(I409369) );
nand I_23939 (I409704,I409424,I605974);
nand I_23940 (I409721,I409704,I409458);
and I_23941 (I409738,I409540,I409721);
DFFARX1 I_23942  ( .D(I409738), .CLK(I2702), .RSTB(I409407), .Q(I409399) );
and I_23943 (I409372,I409704,I409673);
DFFARX1 I_23944  ( .D(I606001), .CLK(I2702), .RSTB(I409407), .Q(I409783) );
nor I_23945 (I409396,I409783,I409704);
nor I_23946 (I409814,I409783,I409458);
nand I_23947 (I409393,I409492,I409814);
not I_23948 (I409390,I409783);
DFFARX1 I_23949  ( .D(I605998), .CLK(I2702), .RSTB(I409407), .Q(I409859) );
not I_23950 (I409876,I409859);
nor I_23951 (I409893,I409876,I409557);
and I_23952 (I409910,I409783,I409893);
or I_23953 (I409927,I409704,I409910);
DFFARX1 I_23954  ( .D(I409927), .CLK(I2702), .RSTB(I409407), .Q(I409384) );
not I_23955 (I409958,I409876);
nor I_23956 (I409975,I409783,I409958);
nand I_23957 (I409387,I409876,I409975);
nand I_23958 (I409381,I409540,I409958);
not I_23959 (I410053,I2709);
not I_23960 (I410070,I597067);
nor I_23961 (I410087,I597055,I597064);
nand I_23962 (I410104,I410087,I597079);
nor I_23963 (I410121,I410070,I597055);
nand I_23964 (I410138,I410121,I597061);
DFFARX1 I_23965  ( .D(I410138), .CLK(I2702), .RSTB(I410053), .Q(I410155) );
not I_23966 (I410024,I410155);
not I_23967 (I410186,I597055);
not I_23968 (I410203,I410186);
not I_23969 (I410220,I597049);
nor I_23970 (I410237,I410220,I597070);
and I_23971 (I410254,I410237,I597052);
or I_23972 (I410271,I410254,I597058);
DFFARX1 I_23973  ( .D(I410271), .CLK(I2702), .RSTB(I410053), .Q(I410288) );
DFFARX1 I_23974  ( .D(I410288), .CLK(I2702), .RSTB(I410053), .Q(I410021) );
DFFARX1 I_23975  ( .D(I410288), .CLK(I2702), .RSTB(I410053), .Q(I410319) );
DFFARX1 I_23976  ( .D(I410288), .CLK(I2702), .RSTB(I410053), .Q(I410015) );
nand I_23977 (I410350,I410070,I597049);
nand I_23978 (I410367,I410350,I410104);
and I_23979 (I410384,I410186,I410367);
DFFARX1 I_23980  ( .D(I410384), .CLK(I2702), .RSTB(I410053), .Q(I410045) );
and I_23981 (I410018,I410350,I410319);
DFFARX1 I_23982  ( .D(I597076), .CLK(I2702), .RSTB(I410053), .Q(I410429) );
nor I_23983 (I410042,I410429,I410350);
nor I_23984 (I410460,I410429,I410104);
nand I_23985 (I410039,I410138,I410460);
not I_23986 (I410036,I410429);
DFFARX1 I_23987  ( .D(I597073), .CLK(I2702), .RSTB(I410053), .Q(I410505) );
not I_23988 (I410522,I410505);
nor I_23989 (I410539,I410522,I410203);
and I_23990 (I410556,I410429,I410539);
or I_23991 (I410573,I410350,I410556);
DFFARX1 I_23992  ( .D(I410573), .CLK(I2702), .RSTB(I410053), .Q(I410030) );
not I_23993 (I410604,I410522);
nor I_23994 (I410621,I410429,I410604);
nand I_23995 (I410033,I410522,I410621);
nand I_23996 (I410027,I410186,I410604);
not I_23997 (I410699,I2709);
not I_23998 (I410716,I682886);
nor I_23999 (I410733,I682883,I682868);
nand I_24000 (I410750,I410733,I682877);
nor I_24001 (I410767,I410716,I682883);
nand I_24002 (I410784,I410767,I682892);
DFFARX1 I_24003  ( .D(I410784), .CLK(I2702), .RSTB(I410699), .Q(I410801) );
not I_24004 (I410670,I410801);
not I_24005 (I410832,I682883);
not I_24006 (I410849,I410832);
not I_24007 (I410866,I682865);
nor I_24008 (I410883,I410866,I682871);
and I_24009 (I410900,I410883,I682895);
or I_24010 (I410917,I410900,I682889);
DFFARX1 I_24011  ( .D(I410917), .CLK(I2702), .RSTB(I410699), .Q(I410934) );
DFFARX1 I_24012  ( .D(I410934), .CLK(I2702), .RSTB(I410699), .Q(I410667) );
DFFARX1 I_24013  ( .D(I410934), .CLK(I2702), .RSTB(I410699), .Q(I410965) );
DFFARX1 I_24014  ( .D(I410934), .CLK(I2702), .RSTB(I410699), .Q(I410661) );
nand I_24015 (I410996,I410716,I682865);
nand I_24016 (I411013,I410996,I410750);
and I_24017 (I411030,I410832,I411013);
DFFARX1 I_24018  ( .D(I411030), .CLK(I2702), .RSTB(I410699), .Q(I410691) );
and I_24019 (I410664,I410996,I410965);
DFFARX1 I_24020  ( .D(I682874), .CLK(I2702), .RSTB(I410699), .Q(I411075) );
nor I_24021 (I410688,I411075,I410996);
nor I_24022 (I411106,I411075,I410750);
nand I_24023 (I410685,I410784,I411106);
not I_24024 (I410682,I411075);
DFFARX1 I_24025  ( .D(I682880), .CLK(I2702), .RSTB(I410699), .Q(I411151) );
not I_24026 (I411168,I411151);
nor I_24027 (I411185,I411168,I410849);
and I_24028 (I411202,I411075,I411185);
or I_24029 (I411219,I410996,I411202);
DFFARX1 I_24030  ( .D(I411219), .CLK(I2702), .RSTB(I410699), .Q(I410676) );
not I_24031 (I411250,I411168);
nor I_24032 (I411267,I411075,I411250);
nand I_24033 (I410679,I411168,I411267);
nand I_24034 (I410673,I410832,I411250);
not I_24035 (I411345,I2709);
not I_24036 (I411362,I283440);
nor I_24037 (I411379,I283419,I283431);
nand I_24038 (I411396,I411379,I283434);
nor I_24039 (I411413,I411362,I283419);
nand I_24040 (I411430,I411413,I283416);
DFFARX1 I_24041  ( .D(I411430), .CLK(I2702), .RSTB(I411345), .Q(I411447) );
not I_24042 (I411316,I411447);
not I_24043 (I411478,I283419);
not I_24044 (I411495,I411478);
not I_24045 (I411512,I283437);
nor I_24046 (I411529,I411512,I283428);
and I_24047 (I411546,I411529,I283422);
or I_24048 (I411563,I411546,I283446);
DFFARX1 I_24049  ( .D(I411563), .CLK(I2702), .RSTB(I411345), .Q(I411580) );
DFFARX1 I_24050  ( .D(I411580), .CLK(I2702), .RSTB(I411345), .Q(I411313) );
DFFARX1 I_24051  ( .D(I411580), .CLK(I2702), .RSTB(I411345), .Q(I411611) );
DFFARX1 I_24052  ( .D(I411580), .CLK(I2702), .RSTB(I411345), .Q(I411307) );
nand I_24053 (I411642,I411362,I283437);
nand I_24054 (I411659,I411642,I411396);
and I_24055 (I411676,I411478,I411659);
DFFARX1 I_24056  ( .D(I411676), .CLK(I2702), .RSTB(I411345), .Q(I411337) );
and I_24057 (I411310,I411642,I411611);
DFFARX1 I_24058  ( .D(I283443), .CLK(I2702), .RSTB(I411345), .Q(I411721) );
nor I_24059 (I411334,I411721,I411642);
nor I_24060 (I411752,I411721,I411396);
nand I_24061 (I411331,I411430,I411752);
not I_24062 (I411328,I411721);
DFFARX1 I_24063  ( .D(I283425), .CLK(I2702), .RSTB(I411345), .Q(I411797) );
not I_24064 (I411814,I411797);
nor I_24065 (I411831,I411814,I411495);
and I_24066 (I411848,I411721,I411831);
or I_24067 (I411865,I411642,I411848);
DFFARX1 I_24068  ( .D(I411865), .CLK(I2702), .RSTB(I411345), .Q(I411322) );
not I_24069 (I411896,I411814);
nor I_24070 (I411913,I411721,I411896);
nand I_24071 (I411325,I411814,I411913);
nand I_24072 (I411319,I411478,I411896);
not I_24073 (I411991,I2709);
or I_24074 (I412008,I228459,I228468);
or I_24075 (I412025,I228453,I228459);
nor I_24076 (I412042,I228447,I228441);
DFFARX1 I_24077  ( .D(I412042), .CLK(I2702), .RSTB(I411991), .Q(I412059) );
DFFARX1 I_24078  ( .D(I412042), .CLK(I2702), .RSTB(I411991), .Q(I411953) );
not I_24079 (I412090,I228447);
and I_24080 (I412107,I412090,I228438);
nor I_24081 (I412124,I412107,I228468);
nor I_24082 (I412141,I228465,I228462);
DFFARX1 I_24083  ( .D(I412141), .CLK(I2702), .RSTB(I411991), .Q(I412158) );
not I_24084 (I412175,I412158);
DFFARX1 I_24085  ( .D(I412158), .CLK(I2702), .RSTB(I411991), .Q(I411962) );
nor I_24086 (I412206,I228465,I228453);
and I_24087 (I411956,I412206,I412059);
DFFARX1 I_24088  ( .D(I228444), .CLK(I2702), .RSTB(I411991), .Q(I412237) );
and I_24089 (I412254,I412237,I228450);
nand I_24090 (I412271,I412254,I412025);
and I_24091 (I412288,I412158,I412271);
DFFARX1 I_24092  ( .D(I412288), .CLK(I2702), .RSTB(I411991), .Q(I411983) );
nor I_24093 (I411980,I412254,I412124);
not I_24094 (I412333,I412254);
nor I_24095 (I412350,I412008,I412333);
nor I_24096 (I412367,I412254,I412206);
nand I_24097 (I411977,I412025,I412367);
nor I_24098 (I412398,I412254,I412175);
not I_24099 (I411974,I412254);
nand I_24100 (I411965,I412254,I412175);
DFFARX1 I_24101  ( .D(I228456), .CLK(I2702), .RSTB(I411991), .Q(I412443) );
and I_24102 (I412460,I412443,I412350);
or I_24103 (I412477,I412008,I412460);
DFFARX1 I_24104  ( .D(I412477), .CLK(I2702), .RSTB(I411991), .Q(I411968) );
nand I_24105 (I411971,I412443,I412398);
nand I_24106 (I412522,I412443,I412124);
and I_24107 (I412539,I412042,I412522);
DFFARX1 I_24108  ( .D(I412539), .CLK(I2702), .RSTB(I411991), .Q(I411959) );
not I_24109 (I412603,I2709);
or I_24110 (I412620,I721598,I721583);
or I_24111 (I412637,I721580,I721598);
nor I_24112 (I412654,I721574,I721586);
DFFARX1 I_24113  ( .D(I412654), .CLK(I2702), .RSTB(I412603), .Q(I412671) );
DFFARX1 I_24114  ( .D(I412654), .CLK(I2702), .RSTB(I412603), .Q(I412565) );
not I_24115 (I412702,I721574);
and I_24116 (I412719,I412702,I721601);
nor I_24117 (I412736,I412719,I721583);
nor I_24118 (I412753,I721589,I721592);
DFFARX1 I_24119  ( .D(I412753), .CLK(I2702), .RSTB(I412603), .Q(I412770) );
not I_24120 (I412787,I412770);
DFFARX1 I_24121  ( .D(I412770), .CLK(I2702), .RSTB(I412603), .Q(I412574) );
nor I_24122 (I412818,I721589,I721580);
and I_24123 (I412568,I412818,I412671);
DFFARX1 I_24124  ( .D(I721577), .CLK(I2702), .RSTB(I412603), .Q(I412849) );
and I_24125 (I412866,I412849,I721595);
nand I_24126 (I412883,I412866,I412637);
and I_24127 (I412900,I412770,I412883);
DFFARX1 I_24128  ( .D(I412900), .CLK(I2702), .RSTB(I412603), .Q(I412595) );
nor I_24129 (I412592,I412866,I412736);
not I_24130 (I412945,I412866);
nor I_24131 (I412962,I412620,I412945);
nor I_24132 (I412979,I412866,I412818);
nand I_24133 (I412589,I412637,I412979);
nor I_24134 (I413010,I412866,I412787);
not I_24135 (I412586,I412866);
nand I_24136 (I412577,I412866,I412787);
DFFARX1 I_24137  ( .D(I721604), .CLK(I2702), .RSTB(I412603), .Q(I413055) );
and I_24138 (I413072,I413055,I412962);
or I_24139 (I413089,I412620,I413072);
DFFARX1 I_24140  ( .D(I413089), .CLK(I2702), .RSTB(I412603), .Q(I412580) );
nand I_24141 (I412583,I413055,I413010);
nand I_24142 (I413134,I413055,I412736);
and I_24143 (I413151,I412654,I413134);
DFFARX1 I_24144  ( .D(I413151), .CLK(I2702), .RSTB(I412603), .Q(I412571) );
not I_24145 (I413215,I2709);
or I_24146 (I413232,I79467,I79494);
or I_24147 (I413249,I79482,I79467);
nor I_24148 (I413266,I79491,I79470);
DFFARX1 I_24149  ( .D(I413266), .CLK(I2702), .RSTB(I413215), .Q(I413283) );
DFFARX1 I_24150  ( .D(I413266), .CLK(I2702), .RSTB(I413215), .Q(I413177) );
not I_24151 (I413314,I79491);
and I_24152 (I413331,I413314,I79488);
nor I_24153 (I413348,I413331,I79494);
nor I_24154 (I413365,I79485,I79473);
DFFARX1 I_24155  ( .D(I413365), .CLK(I2702), .RSTB(I413215), .Q(I413382) );
not I_24156 (I413399,I413382);
DFFARX1 I_24157  ( .D(I413382), .CLK(I2702), .RSTB(I413215), .Q(I413186) );
nor I_24158 (I413430,I79485,I79482);
and I_24159 (I413180,I413430,I413283);
DFFARX1 I_24160  ( .D(I79497), .CLK(I2702), .RSTB(I413215), .Q(I413461) );
and I_24161 (I413478,I413461,I79479);
nand I_24162 (I413495,I413478,I413249);
and I_24163 (I413512,I413382,I413495);
DFFARX1 I_24164  ( .D(I413512), .CLK(I2702), .RSTB(I413215), .Q(I413207) );
nor I_24165 (I413204,I413478,I413348);
not I_24166 (I413557,I413478);
nor I_24167 (I413574,I413232,I413557);
nor I_24168 (I413591,I413478,I413430);
nand I_24169 (I413201,I413249,I413591);
nor I_24170 (I413622,I413478,I413399);
not I_24171 (I413198,I413478);
nand I_24172 (I413189,I413478,I413399);
DFFARX1 I_24173  ( .D(I79476), .CLK(I2702), .RSTB(I413215), .Q(I413667) );
and I_24174 (I413684,I413667,I413574);
or I_24175 (I413701,I413232,I413684);
DFFARX1 I_24176  ( .D(I413701), .CLK(I2702), .RSTB(I413215), .Q(I413192) );
nand I_24177 (I413195,I413667,I413622);
nand I_24178 (I413746,I413667,I413348);
and I_24179 (I413763,I413266,I413746);
DFFARX1 I_24180  ( .D(I413763), .CLK(I2702), .RSTB(I413215), .Q(I413183) );
not I_24181 (I413827,I2709);
or I_24182 (I413844,I319893,I319881);
or I_24183 (I413861,I319890,I319893);
nor I_24184 (I413878,I319884,I319905);
DFFARX1 I_24185  ( .D(I413878), .CLK(I2702), .RSTB(I413827), .Q(I413895) );
DFFARX1 I_24186  ( .D(I413878), .CLK(I2702), .RSTB(I413827), .Q(I413789) );
not I_24187 (I413926,I319884);
and I_24188 (I413943,I413926,I319899);
nor I_24189 (I413960,I413943,I319881);
nor I_24190 (I413977,I319896,I319911);
DFFARX1 I_24191  ( .D(I413977), .CLK(I2702), .RSTB(I413827), .Q(I413994) );
not I_24192 (I414011,I413994);
DFFARX1 I_24193  ( .D(I413994), .CLK(I2702), .RSTB(I413827), .Q(I413798) );
nor I_24194 (I414042,I319896,I319890);
and I_24195 (I413792,I414042,I413895);
DFFARX1 I_24196  ( .D(I319908), .CLK(I2702), .RSTB(I413827), .Q(I414073) );
and I_24197 (I414090,I414073,I319887);
nand I_24198 (I414107,I414090,I413861);
and I_24199 (I414124,I413994,I414107);
DFFARX1 I_24200  ( .D(I414124), .CLK(I2702), .RSTB(I413827), .Q(I413819) );
nor I_24201 (I413816,I414090,I413960);
not I_24202 (I414169,I414090);
nor I_24203 (I414186,I413844,I414169);
nor I_24204 (I414203,I414090,I414042);
nand I_24205 (I413813,I413861,I414203);
nor I_24206 (I414234,I414090,I414011);
not I_24207 (I413810,I414090);
nand I_24208 (I413801,I414090,I414011);
DFFARX1 I_24209  ( .D(I319902), .CLK(I2702), .RSTB(I413827), .Q(I414279) );
and I_24210 (I414296,I414279,I414186);
or I_24211 (I414313,I413844,I414296);
DFFARX1 I_24212  ( .D(I414313), .CLK(I2702), .RSTB(I413827), .Q(I413804) );
nand I_24213 (I413807,I414279,I414234);
nand I_24214 (I414358,I414279,I413960);
and I_24215 (I414375,I413878,I414358);
DFFARX1 I_24216  ( .D(I414375), .CLK(I2702), .RSTB(I413827), .Q(I413795) );
not I_24217 (I414439,I2709);
or I_24218 (I414456,I469107,I469122);
or I_24219 (I414473,I469137,I469107);
nor I_24220 (I414490,I469119,I469110);
DFFARX1 I_24221  ( .D(I414490), .CLK(I2702), .RSTB(I414439), .Q(I414507) );
DFFARX1 I_24222  ( .D(I414490), .CLK(I2702), .RSTB(I414439), .Q(I414401) );
not I_24223 (I414538,I469119);
and I_24224 (I414555,I414538,I469128);
nor I_24225 (I414572,I414555,I469122);
nor I_24226 (I414589,I469134,I469125);
DFFARX1 I_24227  ( .D(I414589), .CLK(I2702), .RSTB(I414439), .Q(I414606) );
not I_24228 (I414623,I414606);
DFFARX1 I_24229  ( .D(I414606), .CLK(I2702), .RSTB(I414439), .Q(I414410) );
nor I_24230 (I414654,I469134,I469137);
and I_24231 (I414404,I414654,I414507);
DFFARX1 I_24232  ( .D(I469113), .CLK(I2702), .RSTB(I414439), .Q(I414685) );
and I_24233 (I414702,I414685,I469116);
nand I_24234 (I414719,I414702,I414473);
and I_24235 (I414736,I414606,I414719);
DFFARX1 I_24236  ( .D(I414736), .CLK(I2702), .RSTB(I414439), .Q(I414431) );
nor I_24237 (I414428,I414702,I414572);
not I_24238 (I414781,I414702);
nor I_24239 (I414798,I414456,I414781);
nor I_24240 (I414815,I414702,I414654);
nand I_24241 (I414425,I414473,I414815);
nor I_24242 (I414846,I414702,I414623);
not I_24243 (I414422,I414702);
nand I_24244 (I414413,I414702,I414623);
DFFARX1 I_24245  ( .D(I469131), .CLK(I2702), .RSTB(I414439), .Q(I414891) );
and I_24246 (I414908,I414891,I414798);
or I_24247 (I414925,I414456,I414908);
DFFARX1 I_24248  ( .D(I414925), .CLK(I2702), .RSTB(I414439), .Q(I414416) );
nand I_24249 (I414419,I414891,I414846);
nand I_24250 (I414970,I414891,I414572);
and I_24251 (I414987,I414490,I414970);
DFFARX1 I_24252  ( .D(I414987), .CLK(I2702), .RSTB(I414439), .Q(I414407) );
not I_24253 (I415051,I2709);
or I_24254 (I415068,I573258,I573270);
or I_24255 (I415085,I573273,I573258);
nor I_24256 (I415102,I573255,I573249);
DFFARX1 I_24257  ( .D(I415102), .CLK(I2702), .RSTB(I415051), .Q(I415119) );
DFFARX1 I_24258  ( .D(I415102), .CLK(I2702), .RSTB(I415051), .Q(I415013) );
not I_24259 (I415150,I573255);
and I_24260 (I415167,I415150,I573261);
nor I_24261 (I415184,I415167,I573270);
nor I_24262 (I415201,I573264,I573267);
DFFARX1 I_24263  ( .D(I415201), .CLK(I2702), .RSTB(I415051), .Q(I415218) );
not I_24264 (I415235,I415218);
DFFARX1 I_24265  ( .D(I415218), .CLK(I2702), .RSTB(I415051), .Q(I415022) );
nor I_24266 (I415266,I573264,I573273);
and I_24267 (I415016,I415266,I415119);
DFFARX1 I_24268  ( .D(I573279), .CLK(I2702), .RSTB(I415051), .Q(I415297) );
and I_24269 (I415314,I415297,I573252);
nand I_24270 (I415331,I415314,I415085);
and I_24271 (I415348,I415218,I415331);
DFFARX1 I_24272  ( .D(I415348), .CLK(I2702), .RSTB(I415051), .Q(I415043) );
nor I_24273 (I415040,I415314,I415184);
not I_24274 (I415393,I415314);
nor I_24275 (I415410,I415068,I415393);
nor I_24276 (I415427,I415314,I415266);
nand I_24277 (I415037,I415085,I415427);
nor I_24278 (I415458,I415314,I415235);
not I_24279 (I415034,I415314);
nand I_24280 (I415025,I415314,I415235);
DFFARX1 I_24281  ( .D(I573276), .CLK(I2702), .RSTB(I415051), .Q(I415503) );
and I_24282 (I415520,I415503,I415410);
or I_24283 (I415537,I415068,I415520);
DFFARX1 I_24284  ( .D(I415537), .CLK(I2702), .RSTB(I415051), .Q(I415028) );
nand I_24285 (I415031,I415503,I415458);
nand I_24286 (I415582,I415503,I415184);
and I_24287 (I415599,I415102,I415582);
DFFARX1 I_24288  ( .D(I415599), .CLK(I2702), .RSTB(I415051), .Q(I415019) );
not I_24289 (I415663,I2709);
or I_24290 (I415680,I44253,I44238);
or I_24291 (I415697,I44226,I44253);
nor I_24292 (I415714,I44232,I44256);
DFFARX1 I_24293  ( .D(I415714), .CLK(I2702), .RSTB(I415663), .Q(I415731) );
DFFARX1 I_24294  ( .D(I415714), .CLK(I2702), .RSTB(I415663), .Q(I415625) );
not I_24295 (I415762,I44232);
and I_24296 (I415779,I415762,I44229);
nor I_24297 (I415796,I415779,I44238);
nor I_24298 (I415813,I44244,I44241);
DFFARX1 I_24299  ( .D(I415813), .CLK(I2702), .RSTB(I415663), .Q(I415830) );
not I_24300 (I415847,I415830);
DFFARX1 I_24301  ( .D(I415830), .CLK(I2702), .RSTB(I415663), .Q(I415634) );
nor I_24302 (I415878,I44244,I44226);
and I_24303 (I415628,I415878,I415731);
DFFARX1 I_24304  ( .D(I44235), .CLK(I2702), .RSTB(I415663), .Q(I415909) );
and I_24305 (I415926,I415909,I44250);
nand I_24306 (I415943,I415926,I415697);
and I_24307 (I415960,I415830,I415943);
DFFARX1 I_24308  ( .D(I415960), .CLK(I2702), .RSTB(I415663), .Q(I415655) );
nor I_24309 (I415652,I415926,I415796);
not I_24310 (I416005,I415926);
nor I_24311 (I416022,I415680,I416005);
nor I_24312 (I416039,I415926,I415878);
nand I_24313 (I415649,I415697,I416039);
nor I_24314 (I416070,I415926,I415847);
not I_24315 (I415646,I415926);
nand I_24316 (I415637,I415926,I415847);
DFFARX1 I_24317  ( .D(I44247), .CLK(I2702), .RSTB(I415663), .Q(I416115) );
and I_24318 (I416132,I416115,I416022);
or I_24319 (I416149,I415680,I416132);
DFFARX1 I_24320  ( .D(I416149), .CLK(I2702), .RSTB(I415663), .Q(I415640) );
nand I_24321 (I415643,I416115,I416070);
nand I_24322 (I416194,I416115,I415796);
and I_24323 (I416211,I415714,I416194);
DFFARX1 I_24324  ( .D(I416211), .CLK(I2702), .RSTB(I415663), .Q(I415631) );
not I_24325 (I416275,I2709);
or I_24326 (I416292,I488888,I488876);
or I_24327 (I416309,I488891,I488888);
nor I_24328 (I416326,I488873,I488867);
DFFARX1 I_24329  ( .D(I416326), .CLK(I2702), .RSTB(I416275), .Q(I416343) );
DFFARX1 I_24330  ( .D(I416326), .CLK(I2702), .RSTB(I416275), .Q(I416237) );
not I_24331 (I416374,I488873);
and I_24332 (I416391,I416374,I488885);
nor I_24333 (I416408,I416391,I488876);
nor I_24334 (I416425,I488879,I488861);
DFFARX1 I_24335  ( .D(I416425), .CLK(I2702), .RSTB(I416275), .Q(I416442) );
not I_24336 (I416459,I416442);
DFFARX1 I_24337  ( .D(I416442), .CLK(I2702), .RSTB(I416275), .Q(I416246) );
nor I_24338 (I416490,I488879,I488891);
and I_24339 (I416240,I416490,I416343);
DFFARX1 I_24340  ( .D(I488882), .CLK(I2702), .RSTB(I416275), .Q(I416521) );
and I_24341 (I416538,I416521,I488870);
nand I_24342 (I416555,I416538,I416309);
and I_24343 (I416572,I416442,I416555);
DFFARX1 I_24344  ( .D(I416572), .CLK(I2702), .RSTB(I416275), .Q(I416267) );
nor I_24345 (I416264,I416538,I416408);
not I_24346 (I416617,I416538);
nor I_24347 (I416634,I416292,I416617);
nor I_24348 (I416651,I416538,I416490);
nand I_24349 (I416261,I416309,I416651);
nor I_24350 (I416682,I416538,I416459);
not I_24351 (I416258,I416538);
nand I_24352 (I416249,I416538,I416459);
DFFARX1 I_24353  ( .D(I488864), .CLK(I2702), .RSTB(I416275), .Q(I416727) );
and I_24354 (I416744,I416727,I416634);
or I_24355 (I416761,I416292,I416744);
DFFARX1 I_24356  ( .D(I416761), .CLK(I2702), .RSTB(I416275), .Q(I416252) );
nand I_24357 (I416255,I416727,I416682);
nand I_24358 (I416806,I416727,I416408);
and I_24359 (I416823,I416326,I416806);
DFFARX1 I_24360  ( .D(I416823), .CLK(I2702), .RSTB(I416275), .Q(I416243) );
not I_24361 (I416887,I2709);
or I_24362 (I416904,I264864,I264852);
or I_24363 (I416921,I264861,I264864);
nor I_24364 (I416938,I264855,I264876);
DFFARX1 I_24365  ( .D(I416938), .CLK(I2702), .RSTB(I416887), .Q(I416955) );
DFFARX1 I_24366  ( .D(I416938), .CLK(I2702), .RSTB(I416887), .Q(I416849) );
not I_24367 (I416986,I264855);
and I_24368 (I417003,I416986,I264870);
nor I_24369 (I417020,I417003,I264852);
nor I_24370 (I417037,I264867,I264882);
DFFARX1 I_24371  ( .D(I417037), .CLK(I2702), .RSTB(I416887), .Q(I417054) );
not I_24372 (I417071,I417054);
DFFARX1 I_24373  ( .D(I417054), .CLK(I2702), .RSTB(I416887), .Q(I416858) );
nor I_24374 (I417102,I264867,I264861);
and I_24375 (I416852,I417102,I416955);
DFFARX1 I_24376  ( .D(I264879), .CLK(I2702), .RSTB(I416887), .Q(I417133) );
and I_24377 (I417150,I417133,I264858);
nand I_24378 (I417167,I417150,I416921);
and I_24379 (I417184,I417054,I417167);
DFFARX1 I_24380  ( .D(I417184), .CLK(I2702), .RSTB(I416887), .Q(I416879) );
nor I_24381 (I416876,I417150,I417020);
not I_24382 (I417229,I417150);
nor I_24383 (I417246,I416904,I417229);
nor I_24384 (I417263,I417150,I417102);
nand I_24385 (I416873,I416921,I417263);
nor I_24386 (I417294,I417150,I417071);
not I_24387 (I416870,I417150);
nand I_24388 (I416861,I417150,I417071);
DFFARX1 I_24389  ( .D(I264873), .CLK(I2702), .RSTB(I416887), .Q(I417339) );
and I_24390 (I417356,I417339,I417246);
or I_24391 (I417373,I416904,I417356);
DFFARX1 I_24392  ( .D(I417373), .CLK(I2702), .RSTB(I416887), .Q(I416864) );
nand I_24393 (I416867,I417339,I417294);
nand I_24394 (I417418,I417339,I417020);
and I_24395 (I417435,I416938,I417418);
DFFARX1 I_24396  ( .D(I417435), .CLK(I2702), .RSTB(I416887), .Q(I416855) );
not I_24397 (I417499,I2709);
or I_24398 (I417516,I164745,I164766);
or I_24399 (I417533,I164763,I164745);
nor I_24400 (I417550,I164754,I164751);
DFFARX1 I_24401  ( .D(I417550), .CLK(I2702), .RSTB(I417499), .Q(I417567) );
DFFARX1 I_24402  ( .D(I417550), .CLK(I2702), .RSTB(I417499), .Q(I417461) );
not I_24403 (I417598,I164754);
and I_24404 (I417615,I417598,I164760);
nor I_24405 (I417632,I417615,I164766);
nor I_24406 (I417649,I164748,I164739);
DFFARX1 I_24407  ( .D(I417649), .CLK(I2702), .RSTB(I417499), .Q(I417666) );
not I_24408 (I417683,I417666);
DFFARX1 I_24409  ( .D(I417666), .CLK(I2702), .RSTB(I417499), .Q(I417470) );
nor I_24410 (I417714,I164748,I164763);
and I_24411 (I417464,I417714,I417567);
DFFARX1 I_24412  ( .D(I164742), .CLK(I2702), .RSTB(I417499), .Q(I417745) );
and I_24413 (I417762,I417745,I164757);
nand I_24414 (I417779,I417762,I417533);
and I_24415 (I417796,I417666,I417779);
DFFARX1 I_24416  ( .D(I417796), .CLK(I2702), .RSTB(I417499), .Q(I417491) );
nor I_24417 (I417488,I417762,I417632);
not I_24418 (I417841,I417762);
nor I_24419 (I417858,I417516,I417841);
nor I_24420 (I417875,I417762,I417714);
nand I_24421 (I417485,I417533,I417875);
nor I_24422 (I417906,I417762,I417683);
not I_24423 (I417482,I417762);
nand I_24424 (I417473,I417762,I417683);
DFFARX1 I_24425  ( .D(I164769), .CLK(I2702), .RSTB(I417499), .Q(I417951) );
and I_24426 (I417968,I417951,I417858);
or I_24427 (I417985,I417516,I417968);
DFFARX1 I_24428  ( .D(I417985), .CLK(I2702), .RSTB(I417499), .Q(I417476) );
nand I_24429 (I417479,I417951,I417906);
nand I_24430 (I418030,I417951,I417632);
and I_24431 (I418047,I417550,I418030);
DFFARX1 I_24432  ( .D(I418047), .CLK(I2702), .RSTB(I417499), .Q(I417467) );
not I_24433 (I418111,I2709);
or I_24434 (I418128,I128563,I128590);
or I_24435 (I418145,I128578,I128563);
nor I_24436 (I418162,I128587,I128566);
DFFARX1 I_24437  ( .D(I418162), .CLK(I2702), .RSTB(I418111), .Q(I418179) );
DFFARX1 I_24438  ( .D(I418162), .CLK(I2702), .RSTB(I418111), .Q(I418073) );
not I_24439 (I418210,I128587);
and I_24440 (I418227,I418210,I128584);
nor I_24441 (I418244,I418227,I128590);
nor I_24442 (I418261,I128581,I128569);
DFFARX1 I_24443  ( .D(I418261), .CLK(I2702), .RSTB(I418111), .Q(I418278) );
not I_24444 (I418295,I418278);
DFFARX1 I_24445  ( .D(I418278), .CLK(I2702), .RSTB(I418111), .Q(I418082) );
nor I_24446 (I418326,I128581,I128578);
and I_24447 (I418076,I418326,I418179);
DFFARX1 I_24448  ( .D(I128593), .CLK(I2702), .RSTB(I418111), .Q(I418357) );
and I_24449 (I418374,I418357,I128575);
nand I_24450 (I418391,I418374,I418145);
and I_24451 (I418408,I418278,I418391);
DFFARX1 I_24452  ( .D(I418408), .CLK(I2702), .RSTB(I418111), .Q(I418103) );
nor I_24453 (I418100,I418374,I418244);
not I_24454 (I418453,I418374);
nor I_24455 (I418470,I418128,I418453);
nor I_24456 (I418487,I418374,I418326);
nand I_24457 (I418097,I418145,I418487);
nor I_24458 (I418518,I418374,I418295);
not I_24459 (I418094,I418374);
nand I_24460 (I418085,I418374,I418295);
DFFARX1 I_24461  ( .D(I128572), .CLK(I2702), .RSTB(I418111), .Q(I418563) );
and I_24462 (I418580,I418563,I418470);
or I_24463 (I418597,I418128,I418580);
DFFARX1 I_24464  ( .D(I418597), .CLK(I2702), .RSTB(I418111), .Q(I418088) );
nand I_24465 (I418091,I418563,I418518);
nand I_24466 (I418642,I418563,I418244);
and I_24467 (I418659,I418162,I418642);
DFFARX1 I_24468  ( .D(I418659), .CLK(I2702), .RSTB(I418111), .Q(I418079) );
not I_24469 (I418723,I2709);
or I_24470 (I418740,I725066,I725051);
or I_24471 (I418757,I725048,I725066);
nor I_24472 (I418774,I725042,I725054);
DFFARX1 I_24473  ( .D(I418774), .CLK(I2702), .RSTB(I418723), .Q(I418791) );
DFFARX1 I_24474  ( .D(I418774), .CLK(I2702), .RSTB(I418723), .Q(I418685) );
not I_24475 (I418822,I725042);
and I_24476 (I418839,I418822,I725069);
nor I_24477 (I418856,I418839,I725051);
nor I_24478 (I418873,I725057,I725060);
DFFARX1 I_24479  ( .D(I418873), .CLK(I2702), .RSTB(I418723), .Q(I418890) );
not I_24480 (I418907,I418890);
DFFARX1 I_24481  ( .D(I418890), .CLK(I2702), .RSTB(I418723), .Q(I418694) );
nor I_24482 (I418938,I725057,I725048);
and I_24483 (I418688,I418938,I418791);
DFFARX1 I_24484  ( .D(I725045), .CLK(I2702), .RSTB(I418723), .Q(I418969) );
and I_24485 (I418986,I418969,I725063);
nand I_24486 (I419003,I418986,I418757);
and I_24487 (I419020,I418890,I419003);
DFFARX1 I_24488  ( .D(I419020), .CLK(I2702), .RSTB(I418723), .Q(I418715) );
nor I_24489 (I418712,I418986,I418856);
not I_24490 (I419065,I418986);
nor I_24491 (I419082,I418740,I419065);
nor I_24492 (I419099,I418986,I418938);
nand I_24493 (I418709,I418757,I419099);
nor I_24494 (I419130,I418986,I418907);
not I_24495 (I418706,I418986);
nand I_24496 (I418697,I418986,I418907);
DFFARX1 I_24497  ( .D(I725072), .CLK(I2702), .RSTB(I418723), .Q(I419175) );
and I_24498 (I419192,I419175,I419082);
or I_24499 (I419209,I418740,I419192);
DFFARX1 I_24500  ( .D(I419209), .CLK(I2702), .RSTB(I418723), .Q(I418700) );
nand I_24501 (I418703,I419175,I419130);
nand I_24502 (I419254,I419175,I418856);
and I_24503 (I419271,I418774,I419254);
DFFARX1 I_24504  ( .D(I419271), .CLK(I2702), .RSTB(I418723), .Q(I418691) );
not I_24505 (I419335,I2709);
or I_24506 (I419352,I447721,I447736);
or I_24507 (I419369,I447751,I447721);
nor I_24508 (I419386,I447733,I447724);
DFFARX1 I_24509  ( .D(I419386), .CLK(I2702), .RSTB(I419335), .Q(I419403) );
DFFARX1 I_24510  ( .D(I419386), .CLK(I2702), .RSTB(I419335), .Q(I419297) );
not I_24511 (I419434,I447733);
and I_24512 (I419451,I419434,I447742);
nor I_24513 (I419468,I419451,I447736);
nor I_24514 (I419485,I447748,I447739);
DFFARX1 I_24515  ( .D(I419485), .CLK(I2702), .RSTB(I419335), .Q(I419502) );
not I_24516 (I419519,I419502);
DFFARX1 I_24517  ( .D(I419502), .CLK(I2702), .RSTB(I419335), .Q(I419306) );
nor I_24518 (I419550,I447748,I447751);
and I_24519 (I419300,I419550,I419403);
DFFARX1 I_24520  ( .D(I447727), .CLK(I2702), .RSTB(I419335), .Q(I419581) );
and I_24521 (I419598,I419581,I447730);
nand I_24522 (I419615,I419598,I419369);
and I_24523 (I419632,I419502,I419615);
DFFARX1 I_24524  ( .D(I419632), .CLK(I2702), .RSTB(I419335), .Q(I419327) );
nor I_24525 (I419324,I419598,I419468);
not I_24526 (I419677,I419598);
nor I_24527 (I419694,I419352,I419677);
nor I_24528 (I419711,I419598,I419550);
nand I_24529 (I419321,I419369,I419711);
nor I_24530 (I419742,I419598,I419519);
not I_24531 (I419318,I419598);
nand I_24532 (I419309,I419598,I419519);
DFFARX1 I_24533  ( .D(I447745), .CLK(I2702), .RSTB(I419335), .Q(I419787) );
and I_24534 (I419804,I419787,I419694);
or I_24535 (I419821,I419352,I419804);
DFFARX1 I_24536  ( .D(I419821), .CLK(I2702), .RSTB(I419335), .Q(I419312) );
nand I_24537 (I419315,I419787,I419742);
nand I_24538 (I419866,I419787,I419468);
and I_24539 (I419883,I419386,I419866);
DFFARX1 I_24540  ( .D(I419883), .CLK(I2702), .RSTB(I419335), .Q(I419303) );
not I_24541 (I419947,I2709);
or I_24542 (I419964,I392588,I392600);
or I_24543 (I419981,I392582,I392588);
nor I_24544 (I419998,I392603,I392579);
DFFARX1 I_24545  ( .D(I419998), .CLK(I2702), .RSTB(I419947), .Q(I420015) );
DFFARX1 I_24546  ( .D(I419998), .CLK(I2702), .RSTB(I419947), .Q(I419909) );
not I_24547 (I420046,I392603);
and I_24548 (I420063,I420046,I392594);
nor I_24549 (I420080,I420063,I392600);
nor I_24550 (I420097,I392573,I392591);
DFFARX1 I_24551  ( .D(I420097), .CLK(I2702), .RSTB(I419947), .Q(I420114) );
not I_24552 (I420131,I420114);
DFFARX1 I_24553  ( .D(I420114), .CLK(I2702), .RSTB(I419947), .Q(I419918) );
nor I_24554 (I420162,I392573,I392582);
and I_24555 (I419912,I420162,I420015);
DFFARX1 I_24556  ( .D(I392597), .CLK(I2702), .RSTB(I419947), .Q(I420193) );
and I_24557 (I420210,I420193,I392576);
nand I_24558 (I420227,I420210,I419981);
and I_24559 (I420244,I420114,I420227);
DFFARX1 I_24560  ( .D(I420244), .CLK(I2702), .RSTB(I419947), .Q(I419939) );
nor I_24561 (I419936,I420210,I420080);
not I_24562 (I420289,I420210);
nor I_24563 (I420306,I419964,I420289);
nor I_24564 (I420323,I420210,I420162);
nand I_24565 (I419933,I419981,I420323);
nor I_24566 (I420354,I420210,I420131);
not I_24567 (I419930,I420210);
nand I_24568 (I419921,I420210,I420131);
DFFARX1 I_24569  ( .D(I392585), .CLK(I2702), .RSTB(I419947), .Q(I420399) );
and I_24570 (I420416,I420399,I420306);
or I_24571 (I420433,I419964,I420416);
DFFARX1 I_24572  ( .D(I420433), .CLK(I2702), .RSTB(I419947), .Q(I419924) );
nand I_24573 (I419927,I420399,I420354);
nand I_24574 (I420478,I420399,I420080);
and I_24575 (I420495,I419998,I420478);
DFFARX1 I_24576  ( .D(I420495), .CLK(I2702), .RSTB(I419947), .Q(I419915) );
not I_24577 (I420559,I2709);
or I_24578 (I420576,I474309,I474324);
or I_24579 (I420593,I474339,I474309);
nor I_24580 (I420610,I474321,I474312);
DFFARX1 I_24581  ( .D(I420610), .CLK(I2702), .RSTB(I420559), .Q(I420627) );
DFFARX1 I_24582  ( .D(I420610), .CLK(I2702), .RSTB(I420559), .Q(I420521) );
not I_24583 (I420658,I474321);
and I_24584 (I420675,I420658,I474330);
nor I_24585 (I420692,I420675,I474324);
nor I_24586 (I420709,I474336,I474327);
DFFARX1 I_24587  ( .D(I420709), .CLK(I2702), .RSTB(I420559), .Q(I420726) );
not I_24588 (I420743,I420726);
DFFARX1 I_24589  ( .D(I420726), .CLK(I2702), .RSTB(I420559), .Q(I420530) );
nor I_24590 (I420774,I474336,I474339);
and I_24591 (I420524,I420774,I420627);
DFFARX1 I_24592  ( .D(I474315), .CLK(I2702), .RSTB(I420559), .Q(I420805) );
and I_24593 (I420822,I420805,I474318);
nand I_24594 (I420839,I420822,I420593);
and I_24595 (I420856,I420726,I420839);
DFFARX1 I_24596  ( .D(I420856), .CLK(I2702), .RSTB(I420559), .Q(I420551) );
nor I_24597 (I420548,I420822,I420692);
not I_24598 (I420901,I420822);
nor I_24599 (I420918,I420576,I420901);
nor I_24600 (I420935,I420822,I420774);
nand I_24601 (I420545,I420593,I420935);
nor I_24602 (I420966,I420822,I420743);
not I_24603 (I420542,I420822);
nand I_24604 (I420533,I420822,I420743);
DFFARX1 I_24605  ( .D(I474333), .CLK(I2702), .RSTB(I420559), .Q(I421011) );
and I_24606 (I421028,I421011,I420918);
or I_24607 (I421045,I420576,I421028);
DFFARX1 I_24608  ( .D(I421045), .CLK(I2702), .RSTB(I420559), .Q(I420536) );
nand I_24609 (I420539,I421011,I420966);
nand I_24610 (I421090,I421011,I420692);
and I_24611 (I421107,I420610,I421090);
DFFARX1 I_24612  ( .D(I421107), .CLK(I2702), .RSTB(I420559), .Q(I420527) );
not I_24613 (I421171,I2709);
or I_24614 (I421188,I112413,I112440);
or I_24615 (I421205,I112428,I112413);
nor I_24616 (I421222,I112437,I112416);
DFFARX1 I_24617  ( .D(I421222), .CLK(I2702), .RSTB(I421171), .Q(I421239) );
DFFARX1 I_24618  ( .D(I421222), .CLK(I2702), .RSTB(I421171), .Q(I421133) );
not I_24619 (I421270,I112437);
and I_24620 (I421287,I421270,I112434);
nor I_24621 (I421304,I421287,I112440);
nor I_24622 (I421321,I112431,I112419);
DFFARX1 I_24623  ( .D(I421321), .CLK(I2702), .RSTB(I421171), .Q(I421338) );
not I_24624 (I421355,I421338);
DFFARX1 I_24625  ( .D(I421338), .CLK(I2702), .RSTB(I421171), .Q(I421142) );
nor I_24626 (I421386,I112431,I112428);
and I_24627 (I421136,I421386,I421239);
DFFARX1 I_24628  ( .D(I112443), .CLK(I2702), .RSTB(I421171), .Q(I421417) );
and I_24629 (I421434,I421417,I112425);
nand I_24630 (I421451,I421434,I421205);
and I_24631 (I421468,I421338,I421451);
DFFARX1 I_24632  ( .D(I421468), .CLK(I2702), .RSTB(I421171), .Q(I421163) );
nor I_24633 (I421160,I421434,I421304);
not I_24634 (I421513,I421434);
nor I_24635 (I421530,I421188,I421513);
nor I_24636 (I421547,I421434,I421386);
nand I_24637 (I421157,I421205,I421547);
nor I_24638 (I421578,I421434,I421355);
not I_24639 (I421154,I421434);
nand I_24640 (I421145,I421434,I421355);
DFFARX1 I_24641  ( .D(I112422), .CLK(I2702), .RSTB(I421171), .Q(I421623) );
and I_24642 (I421640,I421623,I421530);
or I_24643 (I421657,I421188,I421640);
DFFARX1 I_24644  ( .D(I421657), .CLK(I2702), .RSTB(I421171), .Q(I421148) );
nand I_24645 (I421151,I421623,I421578);
nand I_24646 (I421702,I421623,I421304);
and I_24647 (I421719,I421222,I421702);
DFFARX1 I_24648  ( .D(I421719), .CLK(I2702), .RSTB(I421171), .Q(I421139) );
not I_24649 (I421783,I2709);
or I_24650 (I421800,I473153,I473168);
or I_24651 (I421817,I473183,I473153);
nor I_24652 (I421834,I473165,I473156);
DFFARX1 I_24653  ( .D(I421834), .CLK(I2702), .RSTB(I421783), .Q(I421851) );
DFFARX1 I_24654  ( .D(I421834), .CLK(I2702), .RSTB(I421783), .Q(I421745) );
not I_24655 (I421882,I473165);
and I_24656 (I421899,I421882,I473174);
nor I_24657 (I421916,I421899,I473168);
nor I_24658 (I421933,I473180,I473171);
DFFARX1 I_24659  ( .D(I421933), .CLK(I2702), .RSTB(I421783), .Q(I421950) );
not I_24660 (I421967,I421950);
DFFARX1 I_24661  ( .D(I421950), .CLK(I2702), .RSTB(I421783), .Q(I421754) );
nor I_24662 (I421998,I473180,I473183);
and I_24663 (I421748,I421998,I421851);
DFFARX1 I_24664  ( .D(I473159), .CLK(I2702), .RSTB(I421783), .Q(I422029) );
and I_24665 (I422046,I422029,I473162);
nand I_24666 (I422063,I422046,I421817);
and I_24667 (I422080,I421950,I422063);
DFFARX1 I_24668  ( .D(I422080), .CLK(I2702), .RSTB(I421783), .Q(I421775) );
nor I_24669 (I421772,I422046,I421916);
not I_24670 (I422125,I422046);
nor I_24671 (I422142,I421800,I422125);
nor I_24672 (I422159,I422046,I421998);
nand I_24673 (I421769,I421817,I422159);
nor I_24674 (I422190,I422046,I421967);
not I_24675 (I421766,I422046);
nand I_24676 (I421757,I422046,I421967);
DFFARX1 I_24677  ( .D(I473177), .CLK(I2702), .RSTB(I421783), .Q(I422235) );
and I_24678 (I422252,I422235,I422142);
or I_24679 (I422269,I421800,I422252);
DFFARX1 I_24680  ( .D(I422269), .CLK(I2702), .RSTB(I421783), .Q(I421760) );
nand I_24681 (I421763,I422235,I422190);
nand I_24682 (I422314,I422235,I421916);
and I_24683 (I422331,I421834,I422314);
DFFARX1 I_24684  ( .D(I422331), .CLK(I2702), .RSTB(I421783), .Q(I421751) );
not I_24685 (I422395,I2709);
or I_24686 (I422412,I52981,I53008);
or I_24687 (I422429,I52996,I52981);
nor I_24688 (I422446,I53005,I52984);
DFFARX1 I_24689  ( .D(I422446), .CLK(I2702), .RSTB(I422395), .Q(I422463) );
DFFARX1 I_24690  ( .D(I422446), .CLK(I2702), .RSTB(I422395), .Q(I422357) );
not I_24691 (I422494,I53005);
and I_24692 (I422511,I422494,I53002);
nor I_24693 (I422528,I422511,I53008);
nor I_24694 (I422545,I52999,I52987);
DFFARX1 I_24695  ( .D(I422545), .CLK(I2702), .RSTB(I422395), .Q(I422562) );
not I_24696 (I422579,I422562);
DFFARX1 I_24697  ( .D(I422562), .CLK(I2702), .RSTB(I422395), .Q(I422366) );
nor I_24698 (I422610,I52999,I52996);
and I_24699 (I422360,I422610,I422463);
DFFARX1 I_24700  ( .D(I53011), .CLK(I2702), .RSTB(I422395), .Q(I422641) );
and I_24701 (I422658,I422641,I52993);
nand I_24702 (I422675,I422658,I422429);
and I_24703 (I422692,I422562,I422675);
DFFARX1 I_24704  ( .D(I422692), .CLK(I2702), .RSTB(I422395), .Q(I422387) );
nor I_24705 (I422384,I422658,I422528);
not I_24706 (I422737,I422658);
nor I_24707 (I422754,I422412,I422737);
nor I_24708 (I422771,I422658,I422610);
nand I_24709 (I422381,I422429,I422771);
nor I_24710 (I422802,I422658,I422579);
not I_24711 (I422378,I422658);
nand I_24712 (I422369,I422658,I422579);
DFFARX1 I_24713  ( .D(I52990), .CLK(I2702), .RSTB(I422395), .Q(I422847) );
and I_24714 (I422864,I422847,I422754);
or I_24715 (I422881,I422412,I422864);
DFFARX1 I_24716  ( .D(I422881), .CLK(I2702), .RSTB(I422395), .Q(I422372) );
nand I_24717 (I422375,I422847,I422802);
nand I_24718 (I422926,I422847,I422528);
and I_24719 (I422943,I422446,I422926);
DFFARX1 I_24720  ( .D(I422943), .CLK(I2702), .RSTB(I422395), .Q(I422363) );
not I_24721 (I423007,I2709);
or I_24722 (I423024,I705992,I705977);
or I_24723 (I423041,I705974,I705992);
nor I_24724 (I423058,I705968,I705980);
DFFARX1 I_24725  ( .D(I423058), .CLK(I2702), .RSTB(I423007), .Q(I423075) );
DFFARX1 I_24726  ( .D(I423058), .CLK(I2702), .RSTB(I423007), .Q(I422969) );
not I_24727 (I423106,I705968);
and I_24728 (I423123,I423106,I705995);
nor I_24729 (I423140,I423123,I705977);
nor I_24730 (I423157,I705983,I705986);
DFFARX1 I_24731  ( .D(I423157), .CLK(I2702), .RSTB(I423007), .Q(I423174) );
not I_24732 (I423191,I423174);
DFFARX1 I_24733  ( .D(I423174), .CLK(I2702), .RSTB(I423007), .Q(I422978) );
nor I_24734 (I423222,I705983,I705974);
and I_24735 (I422972,I423222,I423075);
DFFARX1 I_24736  ( .D(I705971), .CLK(I2702), .RSTB(I423007), .Q(I423253) );
and I_24737 (I423270,I423253,I705989);
nand I_24738 (I423287,I423270,I423041);
and I_24739 (I423304,I423174,I423287);
DFFARX1 I_24740  ( .D(I423304), .CLK(I2702), .RSTB(I423007), .Q(I422999) );
nor I_24741 (I422996,I423270,I423140);
not I_24742 (I423349,I423270);
nor I_24743 (I423366,I423024,I423349);
nor I_24744 (I423383,I423270,I423222);
nand I_24745 (I422993,I423041,I423383);
nor I_24746 (I423414,I423270,I423191);
not I_24747 (I422990,I423270);
nand I_24748 (I422981,I423270,I423191);
DFFARX1 I_24749  ( .D(I705998), .CLK(I2702), .RSTB(I423007), .Q(I423459) );
and I_24750 (I423476,I423459,I423366);
or I_24751 (I423493,I423024,I423476);
DFFARX1 I_24752  ( .D(I423493), .CLK(I2702), .RSTB(I423007), .Q(I422984) );
nand I_24753 (I422987,I423459,I423414);
nand I_24754 (I423538,I423459,I423140);
and I_24755 (I423555,I423058,I423538);
DFFARX1 I_24756  ( .D(I423555), .CLK(I2702), .RSTB(I423007), .Q(I422975) );
not I_24757 (I423619,I2709);
or I_24758 (I423636,I490724,I490712);
or I_24759 (I423653,I490727,I490724);
nor I_24760 (I423670,I490709,I490703);
DFFARX1 I_24761  ( .D(I423670), .CLK(I2702), .RSTB(I423619), .Q(I423687) );
DFFARX1 I_24762  ( .D(I423670), .CLK(I2702), .RSTB(I423619), .Q(I423581) );
not I_24763 (I423718,I490709);
and I_24764 (I423735,I423718,I490721);
nor I_24765 (I423752,I423735,I490712);
nor I_24766 (I423769,I490715,I490697);
DFFARX1 I_24767  ( .D(I423769), .CLK(I2702), .RSTB(I423619), .Q(I423786) );
not I_24768 (I423803,I423786);
DFFARX1 I_24769  ( .D(I423786), .CLK(I2702), .RSTB(I423619), .Q(I423590) );
nor I_24770 (I423834,I490715,I490727);
and I_24771 (I423584,I423834,I423687);
DFFARX1 I_24772  ( .D(I490718), .CLK(I2702), .RSTB(I423619), .Q(I423865) );
and I_24773 (I423882,I423865,I490706);
nand I_24774 (I423899,I423882,I423653);
and I_24775 (I423916,I423786,I423899);
DFFARX1 I_24776  ( .D(I423916), .CLK(I2702), .RSTB(I423619), .Q(I423611) );
nor I_24777 (I423608,I423882,I423752);
not I_24778 (I423961,I423882);
nor I_24779 (I423978,I423636,I423961);
nor I_24780 (I423995,I423882,I423834);
nand I_24781 (I423605,I423653,I423995);
nor I_24782 (I424026,I423882,I423803);
not I_24783 (I423602,I423882);
nand I_24784 (I423593,I423882,I423803);
DFFARX1 I_24785  ( .D(I490700), .CLK(I2702), .RSTB(I423619), .Q(I424071) );
and I_24786 (I424088,I424071,I423978);
or I_24787 (I424105,I423636,I424088);
DFFARX1 I_24788  ( .D(I424105), .CLK(I2702), .RSTB(I423619), .Q(I423596) );
nand I_24789 (I423599,I424071,I424026);
nand I_24790 (I424150,I424071,I423752);
and I_24791 (I424167,I423670,I424150);
DFFARX1 I_24792  ( .D(I424167), .CLK(I2702), .RSTB(I423619), .Q(I423587) );
not I_24793 (I424231,I2709);
or I_24794 (I424248,I282765,I282753);
or I_24795 (I424265,I282762,I282765);
nor I_24796 (I424282,I282756,I282777);
DFFARX1 I_24797  ( .D(I424282), .CLK(I2702), .RSTB(I424231), .Q(I424299) );
DFFARX1 I_24798  ( .D(I424282), .CLK(I2702), .RSTB(I424231), .Q(I424193) );
not I_24799 (I424330,I282756);
and I_24800 (I424347,I424330,I282771);
nor I_24801 (I424364,I424347,I282753);
nor I_24802 (I424381,I282768,I282783);
DFFARX1 I_24803  ( .D(I424381), .CLK(I2702), .RSTB(I424231), .Q(I424398) );
not I_24804 (I424415,I424398);
DFFARX1 I_24805  ( .D(I424398), .CLK(I2702), .RSTB(I424231), .Q(I424202) );
nor I_24806 (I424446,I282768,I282762);
and I_24807 (I424196,I424446,I424299);
DFFARX1 I_24808  ( .D(I282780), .CLK(I2702), .RSTB(I424231), .Q(I424477) );
and I_24809 (I424494,I424477,I282759);
nand I_24810 (I424511,I424494,I424265);
and I_24811 (I424528,I424398,I424511);
DFFARX1 I_24812  ( .D(I424528), .CLK(I2702), .RSTB(I424231), .Q(I424223) );
nor I_24813 (I424220,I424494,I424364);
not I_24814 (I424573,I424494);
nor I_24815 (I424590,I424248,I424573);
nor I_24816 (I424607,I424494,I424446);
nand I_24817 (I424217,I424265,I424607);
nor I_24818 (I424638,I424494,I424415);
not I_24819 (I424214,I424494);
nand I_24820 (I424205,I424494,I424415);
DFFARX1 I_24821  ( .D(I282774), .CLK(I2702), .RSTB(I424231), .Q(I424683) );
and I_24822 (I424700,I424683,I424590);
or I_24823 (I424717,I424248,I424700);
DFFARX1 I_24824  ( .D(I424717), .CLK(I2702), .RSTB(I424231), .Q(I424208) );
nand I_24825 (I424211,I424683,I424638);
nand I_24826 (I424762,I424683,I424364);
and I_24827 (I424779,I424282,I424762);
DFFARX1 I_24828  ( .D(I424779), .CLK(I2702), .RSTB(I424231), .Q(I424199) );
not I_24829 (I424843,I2709);
or I_24830 (I424860,I648920,I648923);
or I_24831 (I424877,I648929,I648920);
nor I_24832 (I424894,I648926,I648902);
DFFARX1 I_24833  ( .D(I424894), .CLK(I2702), .RSTB(I424843), .Q(I424911) );
DFFARX1 I_24834  ( .D(I424894), .CLK(I2702), .RSTB(I424843), .Q(I424805) );
not I_24835 (I424942,I648926);
and I_24836 (I424959,I424942,I648905);
nor I_24837 (I424976,I424959,I648923);
nor I_24838 (I424993,I648914,I648899);
DFFARX1 I_24839  ( .D(I424993), .CLK(I2702), .RSTB(I424843), .Q(I425010) );
not I_24840 (I425027,I425010);
DFFARX1 I_24841  ( .D(I425010), .CLK(I2702), .RSTB(I424843), .Q(I424814) );
nor I_24842 (I425058,I648914,I648929);
and I_24843 (I424808,I425058,I424911);
DFFARX1 I_24844  ( .D(I648917), .CLK(I2702), .RSTB(I424843), .Q(I425089) );
and I_24845 (I425106,I425089,I648911);
nand I_24846 (I425123,I425106,I424877);
and I_24847 (I425140,I425010,I425123);
DFFARX1 I_24848  ( .D(I425140), .CLK(I2702), .RSTB(I424843), .Q(I424835) );
nor I_24849 (I424832,I425106,I424976);
not I_24850 (I425185,I425106);
nor I_24851 (I425202,I424860,I425185);
nor I_24852 (I425219,I425106,I425058);
nand I_24853 (I424829,I424877,I425219);
nor I_24854 (I425250,I425106,I425027);
not I_24855 (I424826,I425106);
nand I_24856 (I424817,I425106,I425027);
DFFARX1 I_24857  ( .D(I648908), .CLK(I2702), .RSTB(I424843), .Q(I425295) );
and I_24858 (I425312,I425295,I425202);
or I_24859 (I425329,I424860,I425312);
DFFARX1 I_24860  ( .D(I425329), .CLK(I2702), .RSTB(I424843), .Q(I424820) );
nand I_24861 (I424823,I425295,I425250);
nand I_24862 (I425374,I425295,I424976);
and I_24863 (I425391,I424894,I425374);
DFFARX1 I_24864  ( .D(I425391), .CLK(I2702), .RSTB(I424843), .Q(I424811) );
not I_24865 (I425455,I2709);
or I_24866 (I425472,I490112,I490100);
or I_24867 (I425489,I490115,I490112);
nor I_24868 (I425506,I490097,I490091);
DFFARX1 I_24869  ( .D(I425506), .CLK(I2702), .RSTB(I425455), .Q(I425523) );
DFFARX1 I_24870  ( .D(I425506), .CLK(I2702), .RSTB(I425455), .Q(I425417) );
not I_24871 (I425554,I490097);
and I_24872 (I425571,I425554,I490109);
nor I_24873 (I425588,I425571,I490100);
nor I_24874 (I425605,I490103,I490085);
DFFARX1 I_24875  ( .D(I425605), .CLK(I2702), .RSTB(I425455), .Q(I425622) );
not I_24876 (I425639,I425622);
DFFARX1 I_24877  ( .D(I425622), .CLK(I2702), .RSTB(I425455), .Q(I425426) );
nor I_24878 (I425670,I490103,I490115);
and I_24879 (I425420,I425670,I425523);
DFFARX1 I_24880  ( .D(I490106), .CLK(I2702), .RSTB(I425455), .Q(I425701) );
and I_24881 (I425718,I425701,I490094);
nand I_24882 (I425735,I425718,I425489);
and I_24883 (I425752,I425622,I425735);
DFFARX1 I_24884  ( .D(I425752), .CLK(I2702), .RSTB(I425455), .Q(I425447) );
nor I_24885 (I425444,I425718,I425588);
not I_24886 (I425797,I425718);
nor I_24887 (I425814,I425472,I425797);
nor I_24888 (I425831,I425718,I425670);
nand I_24889 (I425441,I425489,I425831);
nor I_24890 (I425862,I425718,I425639);
not I_24891 (I425438,I425718);
nand I_24892 (I425429,I425718,I425639);
DFFARX1 I_24893  ( .D(I490088), .CLK(I2702), .RSTB(I425455), .Q(I425907) );
and I_24894 (I425924,I425907,I425814);
or I_24895 (I425941,I425472,I425924);
DFFARX1 I_24896  ( .D(I425941), .CLK(I2702), .RSTB(I425455), .Q(I425432) );
nand I_24897 (I425435,I425907,I425862);
nand I_24898 (I425986,I425907,I425588);
and I_24899 (I426003,I425506,I425986);
DFFARX1 I_24900  ( .D(I426003), .CLK(I2702), .RSTB(I425455), .Q(I425423) );
not I_24901 (I426067,I2709);
or I_24902 (I426084,I480089,I480104);
or I_24903 (I426101,I480119,I480089);
nor I_24904 (I426118,I480101,I480092);
DFFARX1 I_24905  ( .D(I426118), .CLK(I2702), .RSTB(I426067), .Q(I426135) );
DFFARX1 I_24906  ( .D(I426118), .CLK(I2702), .RSTB(I426067), .Q(I426029) );
not I_24907 (I426166,I480101);
and I_24908 (I426183,I426166,I480110);
nor I_24909 (I426200,I426183,I480104);
nor I_24910 (I426217,I480116,I480107);
DFFARX1 I_24911  ( .D(I426217), .CLK(I2702), .RSTB(I426067), .Q(I426234) );
not I_24912 (I426251,I426234);
DFFARX1 I_24913  ( .D(I426234), .CLK(I2702), .RSTB(I426067), .Q(I426038) );
nor I_24914 (I426282,I480116,I480119);
and I_24915 (I426032,I426282,I426135);
DFFARX1 I_24916  ( .D(I480095), .CLK(I2702), .RSTB(I426067), .Q(I426313) );
and I_24917 (I426330,I426313,I480098);
nand I_24918 (I426347,I426330,I426101);
and I_24919 (I426364,I426234,I426347);
DFFARX1 I_24920  ( .D(I426364), .CLK(I2702), .RSTB(I426067), .Q(I426059) );
nor I_24921 (I426056,I426330,I426200);
not I_24922 (I426409,I426330);
nor I_24923 (I426426,I426084,I426409);
nor I_24924 (I426443,I426330,I426282);
nand I_24925 (I426053,I426101,I426443);
nor I_24926 (I426474,I426330,I426251);
not I_24927 (I426050,I426330);
nand I_24928 (I426041,I426330,I426251);
DFFARX1 I_24929  ( .D(I480113), .CLK(I2702), .RSTB(I426067), .Q(I426519) );
and I_24930 (I426536,I426519,I426426);
or I_24931 (I426553,I426084,I426536);
DFFARX1 I_24932  ( .D(I426553), .CLK(I2702), .RSTB(I426067), .Q(I426044) );
nand I_24933 (I426047,I426519,I426474);
nand I_24934 (I426598,I426519,I426200);
and I_24935 (I426615,I426118,I426598);
DFFARX1 I_24936  ( .D(I426615), .CLK(I2702), .RSTB(I426067), .Q(I426035) );
not I_24937 (I426679,I2709);
or I_24938 (I426696,I396464,I396476);
or I_24939 (I426713,I396458,I396464);
nor I_24940 (I426730,I396479,I396455);
DFFARX1 I_24941  ( .D(I426730), .CLK(I2702), .RSTB(I426679), .Q(I426747) );
DFFARX1 I_24942  ( .D(I426730), .CLK(I2702), .RSTB(I426679), .Q(I426641) );
not I_24943 (I426778,I396479);
and I_24944 (I426795,I426778,I396470);
nor I_24945 (I426812,I426795,I396476);
nor I_24946 (I426829,I396449,I396467);
DFFARX1 I_24947  ( .D(I426829), .CLK(I2702), .RSTB(I426679), .Q(I426846) );
not I_24948 (I426863,I426846);
DFFARX1 I_24949  ( .D(I426846), .CLK(I2702), .RSTB(I426679), .Q(I426650) );
nor I_24950 (I426894,I396449,I396458);
and I_24951 (I426644,I426894,I426747);
DFFARX1 I_24952  ( .D(I396473), .CLK(I2702), .RSTB(I426679), .Q(I426925) );
and I_24953 (I426942,I426925,I396452);
nand I_24954 (I426959,I426942,I426713);
and I_24955 (I426976,I426846,I426959);
DFFARX1 I_24956  ( .D(I426976), .CLK(I2702), .RSTB(I426679), .Q(I426671) );
nor I_24957 (I426668,I426942,I426812);
not I_24958 (I427021,I426942);
nor I_24959 (I427038,I426696,I427021);
nor I_24960 (I427055,I426942,I426894);
nand I_24961 (I426665,I426713,I427055);
nor I_24962 (I427086,I426942,I426863);
not I_24963 (I426662,I426942);
nand I_24964 (I426653,I426942,I426863);
DFFARX1 I_24965  ( .D(I396461), .CLK(I2702), .RSTB(I426679), .Q(I427131) );
and I_24966 (I427148,I427131,I427038);
or I_24967 (I427165,I426696,I427148);
DFFARX1 I_24968  ( .D(I427165), .CLK(I2702), .RSTB(I426679), .Q(I426656) );
nand I_24969 (I426659,I427131,I427086);
nand I_24970 (I427210,I427131,I426812);
and I_24971 (I427227,I426730,I427210);
DFFARX1 I_24972  ( .D(I427227), .CLK(I2702), .RSTB(I426679), .Q(I426647) );
not I_24973 (I427291,I2709);
or I_24974 (I427308,I610740,I610761);
or I_24975 (I427325,I610746,I610740);
nor I_24976 (I427342,I610749,I610737);
DFFARX1 I_24977  ( .D(I427342), .CLK(I2702), .RSTB(I427291), .Q(I427359) );
DFFARX1 I_24978  ( .D(I427342), .CLK(I2702), .RSTB(I427291), .Q(I427253) );
not I_24979 (I427390,I610749);
and I_24980 (I427407,I427390,I610755);
nor I_24981 (I427424,I427407,I610761);
nor I_24982 (I427441,I610743,I610758);
DFFARX1 I_24983  ( .D(I427441), .CLK(I2702), .RSTB(I427291), .Q(I427458) );
not I_24984 (I427475,I427458);
DFFARX1 I_24985  ( .D(I427458), .CLK(I2702), .RSTB(I427291), .Q(I427262) );
nor I_24986 (I427506,I610743,I610746);
and I_24987 (I427256,I427506,I427359);
DFFARX1 I_24988  ( .D(I610734), .CLK(I2702), .RSTB(I427291), .Q(I427537) );
and I_24989 (I427554,I427537,I610764);
nand I_24990 (I427571,I427554,I427325);
and I_24991 (I427588,I427458,I427571);
DFFARX1 I_24992  ( .D(I427588), .CLK(I2702), .RSTB(I427291), .Q(I427283) );
nor I_24993 (I427280,I427554,I427424);
not I_24994 (I427633,I427554);
nor I_24995 (I427650,I427308,I427633);
nor I_24996 (I427667,I427554,I427506);
nand I_24997 (I427277,I427325,I427667);
nor I_24998 (I427698,I427554,I427475);
not I_24999 (I427274,I427554);
nand I_25000 (I427265,I427554,I427475);
DFFARX1 I_25001  ( .D(I610752), .CLK(I2702), .RSTB(I427291), .Q(I427743) );
and I_25002 (I427760,I427743,I427650);
or I_25003 (I427777,I427308,I427760);
DFFARX1 I_25004  ( .D(I427777), .CLK(I2702), .RSTB(I427291), .Q(I427268) );
nand I_25005 (I427271,I427743,I427698);
nand I_25006 (I427822,I427743,I427424);
and I_25007 (I427839,I427342,I427822);
DFFARX1 I_25008  ( .D(I427839), .CLK(I2702), .RSTB(I427291), .Q(I427259) );
not I_25009 (I427903,I2709);
or I_25010 (I427920,I150159,I150180);
or I_25011 (I427937,I150177,I150159);
nor I_25012 (I427954,I150168,I150165);
DFFARX1 I_25013  ( .D(I427954), .CLK(I2702), .RSTB(I427903), .Q(I427971) );
DFFARX1 I_25014  ( .D(I427954), .CLK(I2702), .RSTB(I427903), .Q(I427865) );
not I_25015 (I428002,I150168);
and I_25016 (I428019,I428002,I150174);
nor I_25017 (I428036,I428019,I150180);
nor I_25018 (I428053,I150162,I150153);
DFFARX1 I_25019  ( .D(I428053), .CLK(I2702), .RSTB(I427903), .Q(I428070) );
not I_25020 (I428087,I428070);
DFFARX1 I_25021  ( .D(I428070), .CLK(I2702), .RSTB(I427903), .Q(I427874) );
nor I_25022 (I428118,I150162,I150177);
and I_25023 (I427868,I428118,I427971);
DFFARX1 I_25024  ( .D(I150156), .CLK(I2702), .RSTB(I427903), .Q(I428149) );
and I_25025 (I428166,I428149,I150171);
nand I_25026 (I428183,I428166,I427937);
and I_25027 (I428200,I428070,I428183);
DFFARX1 I_25028  ( .D(I428200), .CLK(I2702), .RSTB(I427903), .Q(I427895) );
nor I_25029 (I427892,I428166,I428036);
not I_25030 (I428245,I428166);
nor I_25031 (I428262,I427920,I428245);
nor I_25032 (I428279,I428166,I428118);
nand I_25033 (I427889,I427937,I428279);
nor I_25034 (I428310,I428166,I428087);
not I_25035 (I427886,I428166);
nand I_25036 (I427877,I428166,I428087);
DFFARX1 I_25037  ( .D(I150183), .CLK(I2702), .RSTB(I427903), .Q(I428355) );
and I_25038 (I428372,I428355,I428262);
or I_25039 (I428389,I427920,I428372);
DFFARX1 I_25040  ( .D(I428389), .CLK(I2702), .RSTB(I427903), .Q(I427880) );
nand I_25041 (I427883,I428355,I428310);
nand I_25042 (I428434,I428355,I428036);
and I_25043 (I428451,I427954,I428434);
DFFARX1 I_25044  ( .D(I428451), .CLK(I2702), .RSTB(I427903), .Q(I427871) );
not I_25045 (I428515,I2709);
or I_25046 (I428532,I104661,I104688);
or I_25047 (I428549,I104676,I104661);
nor I_25048 (I428566,I104685,I104664);
DFFARX1 I_25049  ( .D(I428566), .CLK(I2702), .RSTB(I428515), .Q(I428583) );
DFFARX1 I_25050  ( .D(I428566), .CLK(I2702), .RSTB(I428515), .Q(I428477) );
not I_25051 (I428614,I104685);
and I_25052 (I428631,I428614,I104682);
nor I_25053 (I428648,I428631,I104688);
nor I_25054 (I428665,I104679,I104667);
DFFARX1 I_25055  ( .D(I428665), .CLK(I2702), .RSTB(I428515), .Q(I428682) );
not I_25056 (I428699,I428682);
DFFARX1 I_25057  ( .D(I428682), .CLK(I2702), .RSTB(I428515), .Q(I428486) );
nor I_25058 (I428730,I104679,I104676);
and I_25059 (I428480,I428730,I428583);
DFFARX1 I_25060  ( .D(I104691), .CLK(I2702), .RSTB(I428515), .Q(I428761) );
and I_25061 (I428778,I428761,I104673);
nand I_25062 (I428795,I428778,I428549);
and I_25063 (I428812,I428682,I428795);
DFFARX1 I_25064  ( .D(I428812), .CLK(I2702), .RSTB(I428515), .Q(I428507) );
nor I_25065 (I428504,I428778,I428648);
not I_25066 (I428857,I428778);
nor I_25067 (I428874,I428532,I428857);
nor I_25068 (I428891,I428778,I428730);
nand I_25069 (I428501,I428549,I428891);
nor I_25070 (I428922,I428778,I428699);
not I_25071 (I428498,I428778);
nand I_25072 (I428489,I428778,I428699);
DFFARX1 I_25073  ( .D(I104670), .CLK(I2702), .RSTB(I428515), .Q(I428967) );
and I_25074 (I428984,I428967,I428874);
or I_25075 (I429001,I428532,I428984);
DFFARX1 I_25076  ( .D(I429001), .CLK(I2702), .RSTB(I428515), .Q(I428492) );
nand I_25077 (I428495,I428967,I428922);
nand I_25078 (I429046,I428967,I428648);
and I_25079 (I429063,I428566,I429046);
DFFARX1 I_25080  ( .D(I429063), .CLK(I2702), .RSTB(I428515), .Q(I428483) );
not I_25081 (I429127,I2709);
or I_25082 (I429144,I708304,I708289);
or I_25083 (I429161,I708286,I708304);
nor I_25084 (I429178,I708280,I708292);
DFFARX1 I_25085  ( .D(I429178), .CLK(I2702), .RSTB(I429127), .Q(I429195) );
DFFARX1 I_25086  ( .D(I429178), .CLK(I2702), .RSTB(I429127), .Q(I429089) );
not I_25087 (I429226,I708280);
and I_25088 (I429243,I429226,I708307);
nor I_25089 (I429260,I429243,I708289);
nor I_25090 (I429277,I708295,I708298);
DFFARX1 I_25091  ( .D(I429277), .CLK(I2702), .RSTB(I429127), .Q(I429294) );
not I_25092 (I429311,I429294);
DFFARX1 I_25093  ( .D(I429294), .CLK(I2702), .RSTB(I429127), .Q(I429098) );
nor I_25094 (I429342,I708295,I708286);
and I_25095 (I429092,I429342,I429195);
DFFARX1 I_25096  ( .D(I708283), .CLK(I2702), .RSTB(I429127), .Q(I429373) );
and I_25097 (I429390,I429373,I708301);
nand I_25098 (I429407,I429390,I429161);
and I_25099 (I429424,I429294,I429407);
DFFARX1 I_25100  ( .D(I429424), .CLK(I2702), .RSTB(I429127), .Q(I429119) );
nor I_25101 (I429116,I429390,I429260);
not I_25102 (I429469,I429390);
nor I_25103 (I429486,I429144,I429469);
nor I_25104 (I429503,I429390,I429342);
nand I_25105 (I429113,I429161,I429503);
nor I_25106 (I429534,I429390,I429311);
not I_25107 (I429110,I429390);
nand I_25108 (I429101,I429390,I429311);
DFFARX1 I_25109  ( .D(I708310), .CLK(I2702), .RSTB(I429127), .Q(I429579) );
and I_25110 (I429596,I429579,I429486);
or I_25111 (I429613,I429144,I429596);
DFFARX1 I_25112  ( .D(I429613), .CLK(I2702), .RSTB(I429127), .Q(I429104) );
nand I_25113 (I429107,I429579,I429534);
nand I_25114 (I429658,I429579,I429260);
and I_25115 (I429675,I429178,I429658);
DFFARX1 I_25116  ( .D(I429675), .CLK(I2702), .RSTB(I429127), .Q(I429095) );
not I_25117 (I429739,I2709);
or I_25118 (I429756,I705414,I705399);
or I_25119 (I429773,I705396,I705414);
nor I_25120 (I429790,I705390,I705402);
DFFARX1 I_25121  ( .D(I429790), .CLK(I2702), .RSTB(I429739), .Q(I429807) );
DFFARX1 I_25122  ( .D(I429790), .CLK(I2702), .RSTB(I429739), .Q(I429701) );
not I_25123 (I429838,I705390);
and I_25124 (I429855,I429838,I705417);
nor I_25125 (I429872,I429855,I705399);
nor I_25126 (I429889,I705405,I705408);
DFFARX1 I_25127  ( .D(I429889), .CLK(I2702), .RSTB(I429739), .Q(I429906) );
not I_25128 (I429923,I429906);
DFFARX1 I_25129  ( .D(I429906), .CLK(I2702), .RSTB(I429739), .Q(I429710) );
nor I_25130 (I429954,I705405,I705396);
and I_25131 (I429704,I429954,I429807);
DFFARX1 I_25132  ( .D(I705393), .CLK(I2702), .RSTB(I429739), .Q(I429985) );
and I_25133 (I430002,I429985,I705411);
nand I_25134 (I430019,I430002,I429773);
and I_25135 (I430036,I429906,I430019);
DFFARX1 I_25136  ( .D(I430036), .CLK(I2702), .RSTB(I429739), .Q(I429731) );
nor I_25137 (I429728,I430002,I429872);
not I_25138 (I430081,I430002);
nor I_25139 (I430098,I429756,I430081);
nor I_25140 (I430115,I430002,I429954);
nand I_25141 (I429725,I429773,I430115);
nor I_25142 (I430146,I430002,I429923);
not I_25143 (I429722,I430002);
nand I_25144 (I429713,I430002,I429923);
DFFARX1 I_25145  ( .D(I705420), .CLK(I2702), .RSTB(I429739), .Q(I430191) );
and I_25146 (I430208,I430191,I430098);
or I_25147 (I430225,I429756,I430208);
DFFARX1 I_25148  ( .D(I430225), .CLK(I2702), .RSTB(I429739), .Q(I429716) );
nand I_25149 (I429719,I430191,I430146);
nand I_25150 (I430270,I430191,I429872);
and I_25151 (I430287,I429790,I430270);
DFFARX1 I_25152  ( .D(I430287), .CLK(I2702), .RSTB(I429739), .Q(I429707) );
not I_25153 (I430351,I2709);
or I_25154 (I430368,I595865,I595886);
or I_25155 (I430385,I595871,I595865);
nor I_25156 (I430402,I595874,I595862);
DFFARX1 I_25157  ( .D(I430402), .CLK(I2702), .RSTB(I430351), .Q(I430419) );
DFFARX1 I_25158  ( .D(I430402), .CLK(I2702), .RSTB(I430351), .Q(I430313) );
not I_25159 (I430450,I595874);
and I_25160 (I430467,I430450,I595880);
nor I_25161 (I430484,I430467,I595886);
nor I_25162 (I430501,I595868,I595883);
DFFARX1 I_25163  ( .D(I430501), .CLK(I2702), .RSTB(I430351), .Q(I430518) );
not I_25164 (I430535,I430518);
DFFARX1 I_25165  ( .D(I430518), .CLK(I2702), .RSTB(I430351), .Q(I430322) );
nor I_25166 (I430566,I595868,I595871);
and I_25167 (I430316,I430566,I430419);
DFFARX1 I_25168  ( .D(I595859), .CLK(I2702), .RSTB(I430351), .Q(I430597) );
and I_25169 (I430614,I430597,I595889);
nand I_25170 (I430631,I430614,I430385);
and I_25171 (I430648,I430518,I430631);
DFFARX1 I_25172  ( .D(I430648), .CLK(I2702), .RSTB(I430351), .Q(I430343) );
nor I_25173 (I430340,I430614,I430484);
not I_25174 (I430693,I430614);
nor I_25175 (I430710,I430368,I430693);
nor I_25176 (I430727,I430614,I430566);
nand I_25177 (I430337,I430385,I430727);
nor I_25178 (I430758,I430614,I430535);
not I_25179 (I430334,I430614);
nand I_25180 (I430325,I430614,I430535);
DFFARX1 I_25181  ( .D(I595877), .CLK(I2702), .RSTB(I430351), .Q(I430803) );
and I_25182 (I430820,I430803,I430710);
or I_25183 (I430837,I430368,I430820);
DFFARX1 I_25184  ( .D(I430837), .CLK(I2702), .RSTB(I430351), .Q(I430328) );
nand I_25185 (I430331,I430803,I430758);
nand I_25186 (I430882,I430803,I430484);
and I_25187 (I430899,I430402,I430882);
DFFARX1 I_25188  ( .D(I430899), .CLK(I2702), .RSTB(I430351), .Q(I430319) );
not I_25189 (I430963,I2709);
or I_25190 (I430980,I70423,I70450);
or I_25191 (I430997,I70438,I70423);
nor I_25192 (I431014,I70447,I70426);
DFFARX1 I_25193  ( .D(I431014), .CLK(I2702), .RSTB(I430963), .Q(I431031) );
DFFARX1 I_25194  ( .D(I431014), .CLK(I2702), .RSTB(I430963), .Q(I430925) );
not I_25195 (I431062,I70447);
and I_25196 (I431079,I431062,I70444);
nor I_25197 (I431096,I431079,I70450);
nor I_25198 (I431113,I70441,I70429);
DFFARX1 I_25199  ( .D(I431113), .CLK(I2702), .RSTB(I430963), .Q(I431130) );
not I_25200 (I431147,I431130);
DFFARX1 I_25201  ( .D(I431130), .CLK(I2702), .RSTB(I430963), .Q(I430934) );
nor I_25202 (I431178,I70441,I70438);
and I_25203 (I430928,I431178,I431031);
DFFARX1 I_25204  ( .D(I70453), .CLK(I2702), .RSTB(I430963), .Q(I431209) );
and I_25205 (I431226,I431209,I70435);
nand I_25206 (I431243,I431226,I430997);
and I_25207 (I431260,I431130,I431243);
DFFARX1 I_25208  ( .D(I431260), .CLK(I2702), .RSTB(I430963), .Q(I430955) );
nor I_25209 (I430952,I431226,I431096);
not I_25210 (I431305,I431226);
nor I_25211 (I431322,I430980,I431305);
nor I_25212 (I431339,I431226,I431178);
nand I_25213 (I430949,I430997,I431339);
nor I_25214 (I431370,I431226,I431147);
not I_25215 (I430946,I431226);
nand I_25216 (I430937,I431226,I431147);
DFFARX1 I_25217  ( .D(I70432), .CLK(I2702), .RSTB(I430963), .Q(I431415) );
and I_25218 (I431432,I431415,I431322);
or I_25219 (I431449,I430980,I431432);
DFFARX1 I_25220  ( .D(I431449), .CLK(I2702), .RSTB(I430963), .Q(I430940) );
nand I_25221 (I430943,I431415,I431370);
nand I_25222 (I431494,I431415,I431096);
and I_25223 (I431511,I431014,I431494);
DFFARX1 I_25224  ( .D(I431511), .CLK(I2702), .RSTB(I430963), .Q(I430931) );
not I_25225 (I431575,I2709);
nand I_25226 (I431592,I726213,I726225);
and I_25227 (I431609,I431592,I726198);
DFFARX1 I_25228  ( .D(I431609), .CLK(I2702), .RSTB(I431575), .Q(I431626) );
not I_25229 (I431643,I431626);
DFFARX1 I_25230  ( .D(I431626), .CLK(I2702), .RSTB(I431575), .Q(I431543) );
nor I_25231 (I431674,I726216,I726225);
DFFARX1 I_25232  ( .D(I726207), .CLK(I2702), .RSTB(I431575), .Q(I431691) );
DFFARX1 I_25233  ( .D(I431691), .CLK(I2702), .RSTB(I431575), .Q(I431708) );
not I_25234 (I431546,I431708);
DFFARX1 I_25235  ( .D(I431691), .CLK(I2702), .RSTB(I431575), .Q(I431739) );
and I_25236 (I431540,I431626,I431739);
nand I_25237 (I431770,I726204,I726210);
and I_25238 (I431787,I431770,I726222);
DFFARX1 I_25239  ( .D(I431787), .CLK(I2702), .RSTB(I431575), .Q(I431804) );
nor I_25240 (I431821,I431804,I431643);
not I_25241 (I431838,I431804);
nand I_25242 (I431549,I431626,I431838);
DFFARX1 I_25243  ( .D(I726228), .CLK(I2702), .RSTB(I431575), .Q(I431869) );
and I_25244 (I431886,I431869,I726219);
nor I_25245 (I431903,I431886,I431804);
nor I_25246 (I431920,I431886,I431838);
nand I_25247 (I431555,I431674,I431920);
not I_25248 (I431558,I431886);
DFFARX1 I_25249  ( .D(I431886), .CLK(I2702), .RSTB(I431575), .Q(I431537) );
DFFARX1 I_25250  ( .D(I726201), .CLK(I2702), .RSTB(I431575), .Q(I431979) );
nand I_25251 (I431996,I431979,I431691);
and I_25252 (I432013,I431674,I431996);
DFFARX1 I_25253  ( .D(I432013), .CLK(I2702), .RSTB(I431575), .Q(I431567) );
nor I_25254 (I431564,I431979,I431886);
and I_25255 (I432058,I431979,I431821);
or I_25256 (I432075,I431674,I432058);
DFFARX1 I_25257  ( .D(I432075), .CLK(I2702), .RSTB(I431575), .Q(I431552) );
nand I_25258 (I431561,I431979,I431903);
not I_25259 (I432153,I2709);
nand I_25260 (I432170,I43119,I43134);
and I_25261 (I432187,I432170,I43122);
DFFARX1 I_25262  ( .D(I432187), .CLK(I2702), .RSTB(I432153), .Q(I432204) );
not I_25263 (I432221,I432204);
DFFARX1 I_25264  ( .D(I432204), .CLK(I2702), .RSTB(I432153), .Q(I432121) );
nor I_25265 (I432252,I43131,I43134);
DFFARX1 I_25266  ( .D(I43116), .CLK(I2702), .RSTB(I432153), .Q(I432269) );
DFFARX1 I_25267  ( .D(I432269), .CLK(I2702), .RSTB(I432153), .Q(I432286) );
not I_25268 (I432124,I432286);
DFFARX1 I_25269  ( .D(I432269), .CLK(I2702), .RSTB(I432153), .Q(I432317) );
and I_25270 (I432118,I432204,I432317);
nand I_25271 (I432348,I43107,I43104);
and I_25272 (I432365,I432348,I43110);
DFFARX1 I_25273  ( .D(I432365), .CLK(I2702), .RSTB(I432153), .Q(I432382) );
nor I_25274 (I432399,I432382,I432221);
not I_25275 (I432416,I432382);
nand I_25276 (I432127,I432204,I432416);
DFFARX1 I_25277  ( .D(I43113), .CLK(I2702), .RSTB(I432153), .Q(I432447) );
and I_25278 (I432464,I432447,I43125);
nor I_25279 (I432481,I432464,I432382);
nor I_25280 (I432498,I432464,I432416);
nand I_25281 (I432133,I432252,I432498);
not I_25282 (I432136,I432464);
DFFARX1 I_25283  ( .D(I432464), .CLK(I2702), .RSTB(I432153), .Q(I432115) );
DFFARX1 I_25284  ( .D(I43128), .CLK(I2702), .RSTB(I432153), .Q(I432557) );
nand I_25285 (I432574,I432557,I432269);
and I_25286 (I432591,I432252,I432574);
DFFARX1 I_25287  ( .D(I432591), .CLK(I2702), .RSTB(I432153), .Q(I432145) );
nor I_25288 (I432142,I432557,I432464);
and I_25289 (I432636,I432557,I432399);
or I_25290 (I432653,I432252,I432636);
DFFARX1 I_25291  ( .D(I432653), .CLK(I2702), .RSTB(I432153), .Q(I432130) );
nand I_25292 (I432139,I432557,I432481);
not I_25293 (I432731,I2709);
nand I_25294 (I432748,I2319,I2431);
and I_25295 (I432765,I432748,I1751);
DFFARX1 I_25296  ( .D(I432765), .CLK(I2702), .RSTB(I432731), .Q(I432782) );
not I_25297 (I432799,I432782);
DFFARX1 I_25298  ( .D(I432782), .CLK(I2702), .RSTB(I432731), .Q(I432699) );
nor I_25299 (I432830,I1791,I2431);
DFFARX1 I_25300  ( .D(I1223), .CLK(I2702), .RSTB(I432731), .Q(I432847) );
DFFARX1 I_25301  ( .D(I432847), .CLK(I2702), .RSTB(I432731), .Q(I432864) );
not I_25302 (I432702,I432864);
DFFARX1 I_25303  ( .D(I432847), .CLK(I2702), .RSTB(I432731), .Q(I432895) );
and I_25304 (I432696,I432782,I432895);
nand I_25305 (I432926,I2119,I2623);
and I_25306 (I432943,I432926,I1591);
DFFARX1 I_25307  ( .D(I432943), .CLK(I2702), .RSTB(I432731), .Q(I432960) );
nor I_25308 (I432977,I432960,I432799);
not I_25309 (I432994,I432960);
nand I_25310 (I432705,I432782,I432994);
DFFARX1 I_25311  ( .D(I2599), .CLK(I2702), .RSTB(I432731), .Q(I433025) );
and I_25312 (I433042,I433025,I1983);
nor I_25313 (I433059,I433042,I432960);
nor I_25314 (I433076,I433042,I432994);
nand I_25315 (I432711,I432830,I433076);
not I_25316 (I432714,I433042);
DFFARX1 I_25317  ( .D(I433042), .CLK(I2702), .RSTB(I432731), .Q(I432693) );
DFFARX1 I_25318  ( .D(I1559), .CLK(I2702), .RSTB(I432731), .Q(I433135) );
nand I_25319 (I433152,I433135,I432847);
and I_25320 (I433169,I432830,I433152);
DFFARX1 I_25321  ( .D(I433169), .CLK(I2702), .RSTB(I432731), .Q(I432723) );
nor I_25322 (I432720,I433135,I433042);
and I_25323 (I433214,I433135,I432977);
or I_25324 (I433231,I432830,I433214);
DFFARX1 I_25325  ( .D(I433231), .CLK(I2702), .RSTB(I432731), .Q(I432708) );
nand I_25326 (I432717,I433135,I433059);
not I_25327 (I433309,I2709);
nand I_25328 (I433326,I2183,I1951);
and I_25329 (I433343,I433326,I1775);
DFFARX1 I_25330  ( .D(I433343), .CLK(I2702), .RSTB(I433309), .Q(I433360) );
not I_25331 (I433377,I433360);
DFFARX1 I_25332  ( .D(I433360), .CLK(I2702), .RSTB(I433309), .Q(I433277) );
nor I_25333 (I433408,I1903,I1951);
DFFARX1 I_25334  ( .D(I1583), .CLK(I2702), .RSTB(I433309), .Q(I433425) );
DFFARX1 I_25335  ( .D(I433425), .CLK(I2702), .RSTB(I433309), .Q(I433442) );
not I_25336 (I433280,I433442);
DFFARX1 I_25337  ( .D(I433425), .CLK(I2702), .RSTB(I433309), .Q(I433473) );
and I_25338 (I433274,I433360,I433473);
nand I_25339 (I433504,I1471,I1391);
and I_25340 (I433521,I433504,I1735);
DFFARX1 I_25341  ( .D(I433521), .CLK(I2702), .RSTB(I433309), .Q(I433538) );
nor I_25342 (I433555,I433538,I433377);
not I_25343 (I433572,I433538);
nand I_25344 (I433283,I433360,I433572);
DFFARX1 I_25345  ( .D(I2471), .CLK(I2702), .RSTB(I433309), .Q(I433603) );
and I_25346 (I433620,I433603,I1327);
nor I_25347 (I433637,I433620,I433538);
nor I_25348 (I433654,I433620,I433572);
nand I_25349 (I433289,I433408,I433654);
not I_25350 (I433292,I433620);
DFFARX1 I_25351  ( .D(I433620), .CLK(I2702), .RSTB(I433309), .Q(I433271) );
DFFARX1 I_25352  ( .D(I2375), .CLK(I2702), .RSTB(I433309), .Q(I433713) );
nand I_25353 (I433730,I433713,I433425);
and I_25354 (I433747,I433408,I433730);
DFFARX1 I_25355  ( .D(I433747), .CLK(I2702), .RSTB(I433309), .Q(I433301) );
nor I_25356 (I433298,I433713,I433620);
and I_25357 (I433792,I433713,I433555);
or I_25358 (I433809,I433408,I433792);
DFFARX1 I_25359  ( .D(I433809), .CLK(I2702), .RSTB(I433309), .Q(I433286) );
nand I_25360 (I433295,I433713,I433637);
not I_25361 (I433887,I2709);
nand I_25362 (I433904,I372562,I372559);
and I_25363 (I433921,I433904,I372571);
DFFARX1 I_25364  ( .D(I433921), .CLK(I2702), .RSTB(I433887), .Q(I433938) );
not I_25365 (I433955,I433938);
DFFARX1 I_25366  ( .D(I433938), .CLK(I2702), .RSTB(I433887), .Q(I433855) );
nor I_25367 (I433986,I372568,I372559);
DFFARX1 I_25368  ( .D(I372574), .CLK(I2702), .RSTB(I433887), .Q(I434003) );
DFFARX1 I_25369  ( .D(I434003), .CLK(I2702), .RSTB(I433887), .Q(I434020) );
not I_25370 (I433858,I434020);
DFFARX1 I_25371  ( .D(I434003), .CLK(I2702), .RSTB(I433887), .Q(I434051) );
and I_25372 (I433852,I433938,I434051);
nand I_25373 (I434082,I372550,I372553);
and I_25374 (I434099,I434082,I372577);
DFFARX1 I_25375  ( .D(I434099), .CLK(I2702), .RSTB(I433887), .Q(I434116) );
nor I_25376 (I434133,I434116,I433955);
not I_25377 (I434150,I434116);
nand I_25378 (I433861,I433938,I434150);
DFFARX1 I_25379  ( .D(I372556), .CLK(I2702), .RSTB(I433887), .Q(I434181) );
and I_25380 (I434198,I434181,I372547);
nor I_25381 (I434215,I434198,I434116);
nor I_25382 (I434232,I434198,I434150);
nand I_25383 (I433867,I433986,I434232);
not I_25384 (I433870,I434198);
DFFARX1 I_25385  ( .D(I434198), .CLK(I2702), .RSTB(I433887), .Q(I433849) );
DFFARX1 I_25386  ( .D(I372565), .CLK(I2702), .RSTB(I433887), .Q(I434291) );
nand I_25387 (I434308,I434291,I434003);
and I_25388 (I434325,I433986,I434308);
DFFARX1 I_25389  ( .D(I434325), .CLK(I2702), .RSTB(I433887), .Q(I433879) );
nor I_25390 (I433876,I434291,I434198);
and I_25391 (I434370,I434291,I434133);
or I_25392 (I434387,I433986,I434370);
DFFARX1 I_25393  ( .D(I434387), .CLK(I2702), .RSTB(I433887), .Q(I433864) );
nand I_25394 (I433873,I434291,I434215);
not I_25395 (I434465,I2709);
nand I_25396 (I434482,I643256,I643259);
and I_25397 (I434499,I434482,I643265);
DFFARX1 I_25398  ( .D(I434499), .CLK(I2702), .RSTB(I434465), .Q(I434516) );
not I_25399 (I434533,I434516);
DFFARX1 I_25400  ( .D(I434516), .CLK(I2702), .RSTB(I434465), .Q(I434433) );
nor I_25401 (I434564,I643262,I643259);
DFFARX1 I_25402  ( .D(I643241), .CLK(I2702), .RSTB(I434465), .Q(I434581) );
DFFARX1 I_25403  ( .D(I434581), .CLK(I2702), .RSTB(I434465), .Q(I434598) );
not I_25404 (I434436,I434598);
DFFARX1 I_25405  ( .D(I434581), .CLK(I2702), .RSTB(I434465), .Q(I434629) );
and I_25406 (I434430,I434516,I434629);
nand I_25407 (I434660,I643238,I643253);
and I_25408 (I434677,I434660,I643250);
DFFARX1 I_25409  ( .D(I434677), .CLK(I2702), .RSTB(I434465), .Q(I434694) );
nor I_25410 (I434711,I434694,I434533);
not I_25411 (I434728,I434694);
nand I_25412 (I434439,I434516,I434728);
DFFARX1 I_25413  ( .D(I643268), .CLK(I2702), .RSTB(I434465), .Q(I434759) );
and I_25414 (I434776,I434759,I643247);
nor I_25415 (I434793,I434776,I434694);
nor I_25416 (I434810,I434776,I434728);
nand I_25417 (I434445,I434564,I434810);
not I_25418 (I434448,I434776);
DFFARX1 I_25419  ( .D(I434776), .CLK(I2702), .RSTB(I434465), .Q(I434427) );
DFFARX1 I_25420  ( .D(I643244), .CLK(I2702), .RSTB(I434465), .Q(I434869) );
nand I_25421 (I434886,I434869,I434581);
and I_25422 (I434903,I434564,I434886);
DFFARX1 I_25423  ( .D(I434903), .CLK(I2702), .RSTB(I434465), .Q(I434457) );
nor I_25424 (I434454,I434869,I434776);
and I_25425 (I434948,I434869,I434711);
or I_25426 (I434965,I434564,I434948);
DFFARX1 I_25427  ( .D(I434965), .CLK(I2702), .RSTB(I434465), .Q(I434442) );
nand I_25428 (I434451,I434869,I434793);
not I_25429 (I435043,I2709);
nand I_25430 (I435060,I600628,I600625);
and I_25431 (I435077,I435060,I600619);
DFFARX1 I_25432  ( .D(I435077), .CLK(I2702), .RSTB(I435043), .Q(I435094) );
not I_25433 (I435111,I435094);
DFFARX1 I_25434  ( .D(I435094), .CLK(I2702), .RSTB(I435043), .Q(I435011) );
nor I_25435 (I435142,I600640,I600625);
DFFARX1 I_25436  ( .D(I600643), .CLK(I2702), .RSTB(I435043), .Q(I435159) );
DFFARX1 I_25437  ( .D(I435159), .CLK(I2702), .RSTB(I435043), .Q(I435176) );
not I_25438 (I435014,I435176);
DFFARX1 I_25439  ( .D(I435159), .CLK(I2702), .RSTB(I435043), .Q(I435207) );
and I_25440 (I435008,I435094,I435207);
nand I_25441 (I435238,I600646,I600637);
and I_25442 (I435255,I435238,I600649);
DFFARX1 I_25443  ( .D(I435255), .CLK(I2702), .RSTB(I435043), .Q(I435272) );
nor I_25444 (I435289,I435272,I435111);
not I_25445 (I435306,I435272);
nand I_25446 (I435017,I435094,I435306);
DFFARX1 I_25447  ( .D(I600622), .CLK(I2702), .RSTB(I435043), .Q(I435337) );
and I_25448 (I435354,I435337,I600631);
nor I_25449 (I435371,I435354,I435272);
nor I_25450 (I435388,I435354,I435306);
nand I_25451 (I435023,I435142,I435388);
not I_25452 (I435026,I435354);
DFFARX1 I_25453  ( .D(I435354), .CLK(I2702), .RSTB(I435043), .Q(I435005) );
DFFARX1 I_25454  ( .D(I600634), .CLK(I2702), .RSTB(I435043), .Q(I435447) );
nand I_25455 (I435464,I435447,I435159);
and I_25456 (I435481,I435142,I435464);
DFFARX1 I_25457  ( .D(I435481), .CLK(I2702), .RSTB(I435043), .Q(I435035) );
nor I_25458 (I435032,I435447,I435354);
and I_25459 (I435526,I435447,I435289);
or I_25460 (I435543,I435142,I435526);
DFFARX1 I_25461  ( .D(I435543), .CLK(I2702), .RSTB(I435043), .Q(I435020) );
nand I_25462 (I435029,I435447,I435371);
not I_25463 (I435621,I2709);
nand I_25464 (I435638,I542931,I542919);
and I_25465 (I435655,I435638,I542913);
DFFARX1 I_25466  ( .D(I435655), .CLK(I2702), .RSTB(I435621), .Q(I435672) );
not I_25467 (I435689,I435672);
DFFARX1 I_25468  ( .D(I435672), .CLK(I2702), .RSTB(I435621), .Q(I435589) );
nor I_25469 (I435720,I542910,I542919);
DFFARX1 I_25470  ( .D(I542904), .CLK(I2702), .RSTB(I435621), .Q(I435737) );
DFFARX1 I_25471  ( .D(I435737), .CLK(I2702), .RSTB(I435621), .Q(I435754) );
not I_25472 (I435592,I435754);
DFFARX1 I_25473  ( .D(I435737), .CLK(I2702), .RSTB(I435621), .Q(I435785) );
and I_25474 (I435586,I435672,I435785);
nand I_25475 (I435816,I542907,I542922);
and I_25476 (I435833,I435816,I542934);
DFFARX1 I_25477  ( .D(I435833), .CLK(I2702), .RSTB(I435621), .Q(I435850) );
nor I_25478 (I435867,I435850,I435689);
not I_25479 (I435884,I435850);
nand I_25480 (I435595,I435672,I435884);
DFFARX1 I_25481  ( .D(I542925), .CLK(I2702), .RSTB(I435621), .Q(I435915) );
and I_25482 (I435932,I435915,I542916);
nor I_25483 (I435949,I435932,I435850);
nor I_25484 (I435966,I435932,I435884);
nand I_25485 (I435601,I435720,I435966);
not I_25486 (I435604,I435932);
DFFARX1 I_25487  ( .D(I435932), .CLK(I2702), .RSTB(I435621), .Q(I435583) );
DFFARX1 I_25488  ( .D(I542928), .CLK(I2702), .RSTB(I435621), .Q(I436025) );
nand I_25489 (I436042,I436025,I435737);
and I_25490 (I436059,I435720,I436042);
DFFARX1 I_25491  ( .D(I436059), .CLK(I2702), .RSTB(I435621), .Q(I435613) );
nor I_25492 (I435610,I436025,I435932);
and I_25493 (I436104,I436025,I435867);
or I_25494 (I436121,I435720,I436104);
DFFARX1 I_25495  ( .D(I436121), .CLK(I2702), .RSTB(I435621), .Q(I435598) );
nand I_25496 (I435607,I436025,I435949);
not I_25497 (I436199,I2709);
nand I_25498 (I436216,I56878,I56860);
and I_25499 (I436233,I436216,I56872);
DFFARX1 I_25500  ( .D(I436233), .CLK(I2702), .RSTB(I436199), .Q(I436250) );
not I_25501 (I436267,I436250);
DFFARX1 I_25502  ( .D(I436250), .CLK(I2702), .RSTB(I436199), .Q(I436167) );
nor I_25503 (I436298,I56875,I56860);
DFFARX1 I_25504  ( .D(I56884), .CLK(I2702), .RSTB(I436199), .Q(I436315) );
DFFARX1 I_25505  ( .D(I436315), .CLK(I2702), .RSTB(I436199), .Q(I436332) );
not I_25506 (I436170,I436332);
DFFARX1 I_25507  ( .D(I436315), .CLK(I2702), .RSTB(I436199), .Q(I436363) );
and I_25508 (I436164,I436250,I436363);
nand I_25509 (I436394,I56863,I56887);
and I_25510 (I436411,I436394,I56866);
DFFARX1 I_25511  ( .D(I436411), .CLK(I2702), .RSTB(I436199), .Q(I436428) );
nor I_25512 (I436445,I436428,I436267);
not I_25513 (I436462,I436428);
nand I_25514 (I436173,I436250,I436462);
DFFARX1 I_25515  ( .D(I56869), .CLK(I2702), .RSTB(I436199), .Q(I436493) );
and I_25516 (I436510,I436493,I56881);
nor I_25517 (I436527,I436510,I436428);
nor I_25518 (I436544,I436510,I436462);
nand I_25519 (I436179,I436298,I436544);
not I_25520 (I436182,I436510);
DFFARX1 I_25521  ( .D(I436510), .CLK(I2702), .RSTB(I436199), .Q(I436161) );
DFFARX1 I_25522  ( .D(I56857), .CLK(I2702), .RSTB(I436199), .Q(I436603) );
nand I_25523 (I436620,I436603,I436315);
and I_25524 (I436637,I436298,I436620);
DFFARX1 I_25525  ( .D(I436637), .CLK(I2702), .RSTB(I436199), .Q(I436191) );
nor I_25526 (I436188,I436603,I436510);
and I_25527 (I436682,I436603,I436445);
or I_25528 (I436699,I436298,I436682);
DFFARX1 I_25529  ( .D(I436699), .CLK(I2702), .RSTB(I436199), .Q(I436176) );
nand I_25530 (I436185,I436603,I436527);
not I_25531 (I436777,I2709);
nand I_25532 (I436794,I336386,I336383);
and I_25533 (I436811,I436794,I336395);
DFFARX1 I_25534  ( .D(I436811), .CLK(I2702), .RSTB(I436777), .Q(I436828) );
not I_25535 (I436845,I436828);
DFFARX1 I_25536  ( .D(I436828), .CLK(I2702), .RSTB(I436777), .Q(I436745) );
nor I_25537 (I436876,I336392,I336383);
DFFARX1 I_25538  ( .D(I336398), .CLK(I2702), .RSTB(I436777), .Q(I436893) );
DFFARX1 I_25539  ( .D(I436893), .CLK(I2702), .RSTB(I436777), .Q(I436910) );
not I_25540 (I436748,I436910);
DFFARX1 I_25541  ( .D(I436893), .CLK(I2702), .RSTB(I436777), .Q(I436941) );
and I_25542 (I436742,I436828,I436941);
nand I_25543 (I436972,I336374,I336377);
and I_25544 (I436989,I436972,I336401);
DFFARX1 I_25545  ( .D(I436989), .CLK(I2702), .RSTB(I436777), .Q(I437006) );
nor I_25546 (I437023,I437006,I436845);
not I_25547 (I437040,I437006);
nand I_25548 (I436751,I436828,I437040);
DFFARX1 I_25549  ( .D(I336380), .CLK(I2702), .RSTB(I436777), .Q(I437071) );
and I_25550 (I437088,I437071,I336371);
nor I_25551 (I437105,I437088,I437006);
nor I_25552 (I437122,I437088,I437040);
nand I_25553 (I436757,I436876,I437122);
not I_25554 (I436760,I437088);
DFFARX1 I_25555  ( .D(I437088), .CLK(I2702), .RSTB(I436777), .Q(I436739) );
DFFARX1 I_25556  ( .D(I336389), .CLK(I2702), .RSTB(I436777), .Q(I437181) );
nand I_25557 (I437198,I437181,I436893);
and I_25558 (I437215,I436876,I437198);
DFFARX1 I_25559  ( .D(I437215), .CLK(I2702), .RSTB(I436777), .Q(I436769) );
nor I_25560 (I436766,I437181,I437088);
and I_25561 (I437260,I437181,I437023);
or I_25562 (I437277,I436876,I437260);
DFFARX1 I_25563  ( .D(I437277), .CLK(I2702), .RSTB(I436777), .Q(I436754) );
nand I_25564 (I436763,I437181,I437105);
not I_25565 (I437355,I2709);
nand I_25566 (I437372,I301983,I302010);
and I_25567 (I437389,I437372,I301998);
DFFARX1 I_25568  ( .D(I437389), .CLK(I2702), .RSTB(I437355), .Q(I437406) );
not I_25569 (I437423,I437406);
DFFARX1 I_25570  ( .D(I437406), .CLK(I2702), .RSTB(I437355), .Q(I437323) );
nor I_25571 (I437454,I301986,I302010);
DFFARX1 I_25572  ( .D(I302001), .CLK(I2702), .RSTB(I437355), .Q(I437471) );
DFFARX1 I_25573  ( .D(I437471), .CLK(I2702), .RSTB(I437355), .Q(I437488) );
not I_25574 (I437326,I437488);
DFFARX1 I_25575  ( .D(I437471), .CLK(I2702), .RSTB(I437355), .Q(I437519) );
and I_25576 (I437320,I437406,I437519);
nand I_25577 (I437550,I301995,I301992);
and I_25578 (I437567,I437550,I301989);
DFFARX1 I_25579  ( .D(I437567), .CLK(I2702), .RSTB(I437355), .Q(I437584) );
nor I_25580 (I437601,I437584,I437423);
not I_25581 (I437618,I437584);
nand I_25582 (I437329,I437406,I437618);
DFFARX1 I_25583  ( .D(I302004), .CLK(I2702), .RSTB(I437355), .Q(I437649) );
and I_25584 (I437666,I437649,I301980);
nor I_25585 (I437683,I437666,I437584);
nor I_25586 (I437700,I437666,I437618);
nand I_25587 (I437335,I437454,I437700);
not I_25588 (I437338,I437666);
DFFARX1 I_25589  ( .D(I437666), .CLK(I2702), .RSTB(I437355), .Q(I437317) );
DFFARX1 I_25590  ( .D(I302007), .CLK(I2702), .RSTB(I437355), .Q(I437759) );
nand I_25591 (I437776,I437759,I437471);
and I_25592 (I437793,I437454,I437776);
DFFARX1 I_25593  ( .D(I437793), .CLK(I2702), .RSTB(I437355), .Q(I437347) );
nor I_25594 (I437344,I437759,I437666);
and I_25595 (I437838,I437759,I437601);
or I_25596 (I437855,I437454,I437838);
DFFARX1 I_25597  ( .D(I437855), .CLK(I2702), .RSTB(I437355), .Q(I437332) );
nand I_25598 (I437341,I437759,I437683);
not I_25599 (I437933,I2709);
nand I_25600 (I437950,I541146,I541134);
and I_25601 (I437967,I437950,I541128);
DFFARX1 I_25602  ( .D(I437967), .CLK(I2702), .RSTB(I437933), .Q(I437984) );
not I_25603 (I438001,I437984);
DFFARX1 I_25604  ( .D(I437984), .CLK(I2702), .RSTB(I437933), .Q(I437901) );
nor I_25605 (I438032,I541125,I541134);
DFFARX1 I_25606  ( .D(I541119), .CLK(I2702), .RSTB(I437933), .Q(I438049) );
DFFARX1 I_25607  ( .D(I438049), .CLK(I2702), .RSTB(I437933), .Q(I438066) );
not I_25608 (I437904,I438066);
DFFARX1 I_25609  ( .D(I438049), .CLK(I2702), .RSTB(I437933), .Q(I438097) );
and I_25610 (I437898,I437984,I438097);
nand I_25611 (I438128,I541122,I541137);
and I_25612 (I438145,I438128,I541149);
DFFARX1 I_25613  ( .D(I438145), .CLK(I2702), .RSTB(I437933), .Q(I438162) );
nor I_25614 (I438179,I438162,I438001);
not I_25615 (I438196,I438162);
nand I_25616 (I437907,I437984,I438196);
DFFARX1 I_25617  ( .D(I541140), .CLK(I2702), .RSTB(I437933), .Q(I438227) );
and I_25618 (I438244,I438227,I541131);
nor I_25619 (I438261,I438244,I438162);
nor I_25620 (I438278,I438244,I438196);
nand I_25621 (I437913,I438032,I438278);
not I_25622 (I437916,I438244);
DFFARX1 I_25623  ( .D(I438244), .CLK(I2702), .RSTB(I437933), .Q(I437895) );
DFFARX1 I_25624  ( .D(I541143), .CLK(I2702), .RSTB(I437933), .Q(I438337) );
nand I_25625 (I438354,I438337,I438049);
and I_25626 (I438371,I438032,I438354);
DFFARX1 I_25627  ( .D(I438371), .CLK(I2702), .RSTB(I437933), .Q(I437925) );
nor I_25628 (I437922,I438337,I438244);
and I_25629 (I438416,I438337,I438179);
or I_25630 (I438433,I438032,I438416);
DFFARX1 I_25631  ( .D(I438433), .CLK(I2702), .RSTB(I437933), .Q(I437910) );
nand I_25632 (I437919,I438337,I438261);
not I_25633 (I438511,I2709);
nand I_25634 (I438528,I660239,I660242);
and I_25635 (I438545,I438528,I660248);
DFFARX1 I_25636  ( .D(I438545), .CLK(I2702), .RSTB(I438511), .Q(I438562) );
not I_25637 (I438579,I438562);
DFFARX1 I_25638  ( .D(I438562), .CLK(I2702), .RSTB(I438511), .Q(I438479) );
nor I_25639 (I438610,I660245,I660242);
DFFARX1 I_25640  ( .D(I660224), .CLK(I2702), .RSTB(I438511), .Q(I438627) );
DFFARX1 I_25641  ( .D(I438627), .CLK(I2702), .RSTB(I438511), .Q(I438644) );
not I_25642 (I438482,I438644);
DFFARX1 I_25643  ( .D(I438627), .CLK(I2702), .RSTB(I438511), .Q(I438675) );
and I_25644 (I438476,I438562,I438675);
nand I_25645 (I438706,I660221,I660236);
and I_25646 (I438723,I438706,I660233);
DFFARX1 I_25647  ( .D(I438723), .CLK(I2702), .RSTB(I438511), .Q(I438740) );
nor I_25648 (I438757,I438740,I438579);
not I_25649 (I438774,I438740);
nand I_25650 (I438485,I438562,I438774);
DFFARX1 I_25651  ( .D(I660251), .CLK(I2702), .RSTB(I438511), .Q(I438805) );
and I_25652 (I438822,I438805,I660230);
nor I_25653 (I438839,I438822,I438740);
nor I_25654 (I438856,I438822,I438774);
nand I_25655 (I438491,I438610,I438856);
not I_25656 (I438494,I438822);
DFFARX1 I_25657  ( .D(I438822), .CLK(I2702), .RSTB(I438511), .Q(I438473) );
DFFARX1 I_25658  ( .D(I660227), .CLK(I2702), .RSTB(I438511), .Q(I438915) );
nand I_25659 (I438932,I438915,I438627);
and I_25660 (I438949,I438610,I438932);
DFFARX1 I_25661  ( .D(I438949), .CLK(I2702), .RSTB(I438511), .Q(I438503) );
nor I_25662 (I438500,I438915,I438822);
and I_25663 (I438994,I438915,I438757);
or I_25664 (I439011,I438610,I438994);
DFFARX1 I_25665  ( .D(I439011), .CLK(I2702), .RSTB(I438511), .Q(I438488) );
nand I_25666 (I438497,I438915,I438839);
not I_25667 (I439089,I2709);
nand I_25668 (I439106,I215967,I215952);
and I_25669 (I439123,I439106,I215961);
DFFARX1 I_25670  ( .D(I439123), .CLK(I2702), .RSTB(I439089), .Q(I439140) );
not I_25671 (I439157,I439140);
DFFARX1 I_25672  ( .D(I439140), .CLK(I2702), .RSTB(I439089), .Q(I439057) );
nor I_25673 (I439188,I215970,I215952);
DFFARX1 I_25674  ( .D(I215949), .CLK(I2702), .RSTB(I439089), .Q(I439205) );
DFFARX1 I_25675  ( .D(I439205), .CLK(I2702), .RSTB(I439089), .Q(I439222) );
not I_25676 (I439060,I439222);
DFFARX1 I_25677  ( .D(I439205), .CLK(I2702), .RSTB(I439089), .Q(I439253) );
and I_25678 (I439054,I439140,I439253);
nand I_25679 (I439284,I215973,I215946);
and I_25680 (I439301,I439284,I215964);
DFFARX1 I_25681  ( .D(I439301), .CLK(I2702), .RSTB(I439089), .Q(I439318) );
nor I_25682 (I439335,I439318,I439157);
not I_25683 (I439352,I439318);
nand I_25684 (I439063,I439140,I439352);
DFFARX1 I_25685  ( .D(I215958), .CLK(I2702), .RSTB(I439089), .Q(I439383) );
and I_25686 (I439400,I439383,I215943);
nor I_25687 (I439417,I439400,I439318);
nor I_25688 (I439434,I439400,I439352);
nand I_25689 (I439069,I439188,I439434);
not I_25690 (I439072,I439400);
DFFARX1 I_25691  ( .D(I439400), .CLK(I2702), .RSTB(I439089), .Q(I439051) );
DFFARX1 I_25692  ( .D(I215955), .CLK(I2702), .RSTB(I439089), .Q(I439493) );
nand I_25693 (I439510,I439493,I439205);
and I_25694 (I439527,I439188,I439510);
DFFARX1 I_25695  ( .D(I439527), .CLK(I2702), .RSTB(I439089), .Q(I439081) );
nor I_25696 (I439078,I439493,I439400);
and I_25697 (I439572,I439493,I439335);
or I_25698 (I439589,I439188,I439572);
DFFARX1 I_25699  ( .D(I439589), .CLK(I2702), .RSTB(I439089), .Q(I439066) );
nand I_25700 (I439075,I439493,I439417);
not I_25701 (I439667,I2709);
nand I_25702 (I439684,I535791,I535779);
and I_25703 (I439701,I439684,I535773);
DFFARX1 I_25704  ( .D(I439701), .CLK(I2702), .RSTB(I439667), .Q(I439718) );
not I_25705 (I439735,I439718);
DFFARX1 I_25706  ( .D(I439718), .CLK(I2702), .RSTB(I439667), .Q(I439635) );
nor I_25707 (I439766,I535770,I535779);
DFFARX1 I_25708  ( .D(I535764), .CLK(I2702), .RSTB(I439667), .Q(I439783) );
DFFARX1 I_25709  ( .D(I439783), .CLK(I2702), .RSTB(I439667), .Q(I439800) );
not I_25710 (I439638,I439800);
DFFARX1 I_25711  ( .D(I439783), .CLK(I2702), .RSTB(I439667), .Q(I439831) );
and I_25712 (I439632,I439718,I439831);
nand I_25713 (I439862,I535767,I535782);
and I_25714 (I439879,I439862,I535794);
DFFARX1 I_25715  ( .D(I439879), .CLK(I2702), .RSTB(I439667), .Q(I439896) );
nor I_25716 (I439913,I439896,I439735);
not I_25717 (I439930,I439896);
nand I_25718 (I439641,I439718,I439930);
DFFARX1 I_25719  ( .D(I535785), .CLK(I2702), .RSTB(I439667), .Q(I439961) );
and I_25720 (I439978,I439961,I535776);
nor I_25721 (I439995,I439978,I439896);
nor I_25722 (I440012,I439978,I439930);
nand I_25723 (I439647,I439766,I440012);
not I_25724 (I439650,I439978);
DFFARX1 I_25725  ( .D(I439978), .CLK(I2702), .RSTB(I439667), .Q(I439629) );
DFFARX1 I_25726  ( .D(I535788), .CLK(I2702), .RSTB(I439667), .Q(I440071) );
nand I_25727 (I440088,I440071,I439783);
and I_25728 (I440105,I439766,I440088);
DFFARX1 I_25729  ( .D(I440105), .CLK(I2702), .RSTB(I439667), .Q(I439659) );
nor I_25730 (I439656,I440071,I439978);
and I_25731 (I440150,I440071,I439913);
or I_25732 (I440167,I439766,I440150);
DFFARX1 I_25733  ( .D(I440167), .CLK(I2702), .RSTB(I439667), .Q(I439644) );
nand I_25734 (I439653,I440071,I439995);
not I_25735 (I440245,I2709);
nand I_25736 (I440262,I595273,I595270);
and I_25737 (I440279,I440262,I595264);
DFFARX1 I_25738  ( .D(I440279), .CLK(I2702), .RSTB(I440245), .Q(I440296) );
not I_25739 (I440313,I440296);
DFFARX1 I_25740  ( .D(I440296), .CLK(I2702), .RSTB(I440245), .Q(I440213) );
nor I_25741 (I440344,I595285,I595270);
DFFARX1 I_25742  ( .D(I595288), .CLK(I2702), .RSTB(I440245), .Q(I440361) );
DFFARX1 I_25743  ( .D(I440361), .CLK(I2702), .RSTB(I440245), .Q(I440378) );
not I_25744 (I440216,I440378);
DFFARX1 I_25745  ( .D(I440361), .CLK(I2702), .RSTB(I440245), .Q(I440409) );
and I_25746 (I440210,I440296,I440409);
nand I_25747 (I440440,I595291,I595282);
and I_25748 (I440457,I440440,I595294);
DFFARX1 I_25749  ( .D(I440457), .CLK(I2702), .RSTB(I440245), .Q(I440474) );
nor I_25750 (I440491,I440474,I440313);
not I_25751 (I440508,I440474);
nand I_25752 (I440219,I440296,I440508);
DFFARX1 I_25753  ( .D(I595267), .CLK(I2702), .RSTB(I440245), .Q(I440539) );
and I_25754 (I440556,I440539,I595276);
nor I_25755 (I440573,I440556,I440474);
nor I_25756 (I440590,I440556,I440508);
nand I_25757 (I440225,I440344,I440590);
not I_25758 (I440228,I440556);
DFFARX1 I_25759  ( .D(I440556), .CLK(I2702), .RSTB(I440245), .Q(I440207) );
DFFARX1 I_25760  ( .D(I595279), .CLK(I2702), .RSTB(I440245), .Q(I440649) );
nand I_25761 (I440666,I440649,I440361);
and I_25762 (I440683,I440344,I440666);
DFFARX1 I_25763  ( .D(I440683), .CLK(I2702), .RSTB(I440245), .Q(I440237) );
nor I_25764 (I440234,I440649,I440556);
and I_25765 (I440728,I440649,I440491);
or I_25766 (I440745,I440344,I440728);
DFFARX1 I_25767  ( .D(I440745), .CLK(I2702), .RSTB(I440245), .Q(I440222) );
nand I_25768 (I440231,I440649,I440573);
not I_25769 (I440823,I2709);
nand I_25770 (I440840,I681625,I681628);
and I_25771 (I440857,I440840,I681634);
DFFARX1 I_25772  ( .D(I440857), .CLK(I2702), .RSTB(I440823), .Q(I440874) );
not I_25773 (I440891,I440874);
DFFARX1 I_25774  ( .D(I440874), .CLK(I2702), .RSTB(I440823), .Q(I440791) );
nor I_25775 (I440922,I681631,I681628);
DFFARX1 I_25776  ( .D(I681610), .CLK(I2702), .RSTB(I440823), .Q(I440939) );
DFFARX1 I_25777  ( .D(I440939), .CLK(I2702), .RSTB(I440823), .Q(I440956) );
not I_25778 (I440794,I440956);
DFFARX1 I_25779  ( .D(I440939), .CLK(I2702), .RSTB(I440823), .Q(I440987) );
and I_25780 (I440788,I440874,I440987);
nand I_25781 (I441018,I681607,I681622);
and I_25782 (I441035,I441018,I681619);
DFFARX1 I_25783  ( .D(I441035), .CLK(I2702), .RSTB(I440823), .Q(I441052) );
nor I_25784 (I441069,I441052,I440891);
not I_25785 (I441086,I441052);
nand I_25786 (I440797,I440874,I441086);
DFFARX1 I_25787  ( .D(I681637), .CLK(I2702), .RSTB(I440823), .Q(I441117) );
and I_25788 (I441134,I441117,I681616);
nor I_25789 (I441151,I441134,I441052);
nor I_25790 (I441168,I441134,I441086);
nand I_25791 (I440803,I440922,I441168);
not I_25792 (I440806,I441134);
DFFARX1 I_25793  ( .D(I441134), .CLK(I2702), .RSTB(I440823), .Q(I440785) );
DFFARX1 I_25794  ( .D(I681613), .CLK(I2702), .RSTB(I440823), .Q(I441227) );
nand I_25795 (I441244,I441227,I440939);
and I_25796 (I441261,I440922,I441244);
DFFARX1 I_25797  ( .D(I441261), .CLK(I2702), .RSTB(I440823), .Q(I440815) );
nor I_25798 (I440812,I441227,I441134);
and I_25799 (I441306,I441227,I441069);
or I_25800 (I441323,I440922,I441306);
DFFARX1 I_25801  ( .D(I441323), .CLK(I2702), .RSTB(I440823), .Q(I440800) );
nand I_25802 (I440809,I441227,I441151);
not I_25803 (I441401,I2709);
nand I_25804 (I441418,I318558,I318585);
and I_25805 (I441435,I441418,I318573);
DFFARX1 I_25806  ( .D(I441435), .CLK(I2702), .RSTB(I441401), .Q(I441452) );
not I_25807 (I441469,I441452);
DFFARX1 I_25808  ( .D(I441452), .CLK(I2702), .RSTB(I441401), .Q(I441369) );
nor I_25809 (I441500,I318561,I318585);
DFFARX1 I_25810  ( .D(I318576), .CLK(I2702), .RSTB(I441401), .Q(I441517) );
DFFARX1 I_25811  ( .D(I441517), .CLK(I2702), .RSTB(I441401), .Q(I441534) );
not I_25812 (I441372,I441534);
DFFARX1 I_25813  ( .D(I441517), .CLK(I2702), .RSTB(I441401), .Q(I441565) );
and I_25814 (I441366,I441452,I441565);
nand I_25815 (I441596,I318570,I318567);
and I_25816 (I441613,I441596,I318564);
DFFARX1 I_25817  ( .D(I441613), .CLK(I2702), .RSTB(I441401), .Q(I441630) );
nor I_25818 (I441647,I441630,I441469);
not I_25819 (I441664,I441630);
nand I_25820 (I441375,I441452,I441664);
DFFARX1 I_25821  ( .D(I318579), .CLK(I2702), .RSTB(I441401), .Q(I441695) );
and I_25822 (I441712,I441695,I318555);
nor I_25823 (I441729,I441712,I441630);
nor I_25824 (I441746,I441712,I441664);
nand I_25825 (I441381,I441500,I441746);
not I_25826 (I441384,I441712);
DFFARX1 I_25827  ( .D(I441712), .CLK(I2702), .RSTB(I441401), .Q(I441363) );
DFFARX1 I_25828  ( .D(I318582), .CLK(I2702), .RSTB(I441401), .Q(I441805) );
nand I_25829 (I441822,I441805,I441517);
and I_25830 (I441839,I441500,I441822);
DFFARX1 I_25831  ( .D(I441839), .CLK(I2702), .RSTB(I441401), .Q(I441393) );
nor I_25832 (I441390,I441805,I441712);
and I_25833 (I441884,I441805,I441647);
or I_25834 (I441901,I441500,I441884);
DFFARX1 I_25835  ( .D(I441901), .CLK(I2702), .RSTB(I441401), .Q(I441378) );
nand I_25836 (I441387,I441805,I441729);
not I_25837 (I441979,I2709);
nand I_25838 (I441996,I72382,I72364);
and I_25839 (I442013,I441996,I72376);
DFFARX1 I_25840  ( .D(I442013), .CLK(I2702), .RSTB(I441979), .Q(I442030) );
not I_25841 (I442047,I442030);
DFFARX1 I_25842  ( .D(I442030), .CLK(I2702), .RSTB(I441979), .Q(I441947) );
nor I_25843 (I442078,I72379,I72364);
DFFARX1 I_25844  ( .D(I72388), .CLK(I2702), .RSTB(I441979), .Q(I442095) );
DFFARX1 I_25845  ( .D(I442095), .CLK(I2702), .RSTB(I441979), .Q(I442112) );
not I_25846 (I441950,I442112);
DFFARX1 I_25847  ( .D(I442095), .CLK(I2702), .RSTB(I441979), .Q(I442143) );
and I_25848 (I441944,I442030,I442143);
nand I_25849 (I442174,I72367,I72391);
and I_25850 (I442191,I442174,I72370);
DFFARX1 I_25851  ( .D(I442191), .CLK(I2702), .RSTB(I441979), .Q(I442208) );
nor I_25852 (I442225,I442208,I442047);
not I_25853 (I442242,I442208);
nand I_25854 (I441953,I442030,I442242);
DFFARX1 I_25855  ( .D(I72373), .CLK(I2702), .RSTB(I441979), .Q(I442273) );
and I_25856 (I442290,I442273,I72385);
nor I_25857 (I442307,I442290,I442208);
nor I_25858 (I442324,I442290,I442242);
nand I_25859 (I441959,I442078,I442324);
not I_25860 (I441962,I442290);
DFFARX1 I_25861  ( .D(I442290), .CLK(I2702), .RSTB(I441979), .Q(I441941) );
DFFARX1 I_25862  ( .D(I72361), .CLK(I2702), .RSTB(I441979), .Q(I442383) );
nand I_25863 (I442400,I442383,I442095);
and I_25864 (I442417,I442078,I442400);
DFFARX1 I_25865  ( .D(I442417), .CLK(I2702), .RSTB(I441979), .Q(I441971) );
nor I_25866 (I441968,I442383,I442290);
and I_25867 (I442462,I442383,I442225);
or I_25868 (I442479,I442078,I442462);
DFFARX1 I_25869  ( .D(I442479), .CLK(I2702), .RSTB(I441979), .Q(I441956) );
nand I_25870 (I441965,I442383,I442307);
not I_25871 (I442557,I2709);
nand I_25872 (I442574,I10581,I10596);
and I_25873 (I442591,I442574,I10584);
DFFARX1 I_25874  ( .D(I442591), .CLK(I2702), .RSTB(I442557), .Q(I442608) );
not I_25875 (I442625,I442608);
DFFARX1 I_25876  ( .D(I442608), .CLK(I2702), .RSTB(I442557), .Q(I442525) );
nor I_25877 (I442656,I10593,I10596);
DFFARX1 I_25878  ( .D(I10578), .CLK(I2702), .RSTB(I442557), .Q(I442673) );
DFFARX1 I_25879  ( .D(I442673), .CLK(I2702), .RSTB(I442557), .Q(I442690) );
not I_25880 (I442528,I442690);
DFFARX1 I_25881  ( .D(I442673), .CLK(I2702), .RSTB(I442557), .Q(I442721) );
and I_25882 (I442522,I442608,I442721);
nand I_25883 (I442752,I10569,I10566);
and I_25884 (I442769,I442752,I10572);
DFFARX1 I_25885  ( .D(I442769), .CLK(I2702), .RSTB(I442557), .Q(I442786) );
nor I_25886 (I442803,I442786,I442625);
not I_25887 (I442820,I442786);
nand I_25888 (I442531,I442608,I442820);
DFFARX1 I_25889  ( .D(I10575), .CLK(I2702), .RSTB(I442557), .Q(I442851) );
and I_25890 (I442868,I442851,I10587);
nor I_25891 (I442885,I442868,I442786);
nor I_25892 (I442902,I442868,I442820);
nand I_25893 (I442537,I442656,I442902);
not I_25894 (I442540,I442868);
DFFARX1 I_25895  ( .D(I442868), .CLK(I2702), .RSTB(I442557), .Q(I442519) );
DFFARX1 I_25896  ( .D(I10590), .CLK(I2702), .RSTB(I442557), .Q(I442961) );
nand I_25897 (I442978,I442961,I442673);
and I_25898 (I442995,I442656,I442978);
DFFARX1 I_25899  ( .D(I442995), .CLK(I2702), .RSTB(I442557), .Q(I442549) );
nor I_25900 (I442546,I442961,I442868);
and I_25901 (I443040,I442961,I442803);
or I_25902 (I443057,I442656,I443040);
DFFARX1 I_25903  ( .D(I443057), .CLK(I2702), .RSTB(I442557), .Q(I442534) );
nand I_25904 (I442543,I442961,I442885);
not I_25905 (I443135,I2709);
nand I_25906 (I443152,I630676,I630679);
and I_25907 (I443169,I443152,I630685);
DFFARX1 I_25908  ( .D(I443169), .CLK(I2702), .RSTB(I443135), .Q(I443186) );
not I_25909 (I443203,I443186);
DFFARX1 I_25910  ( .D(I443186), .CLK(I2702), .RSTB(I443135), .Q(I443103) );
nor I_25911 (I443234,I630682,I630679);
DFFARX1 I_25912  ( .D(I630661), .CLK(I2702), .RSTB(I443135), .Q(I443251) );
DFFARX1 I_25913  ( .D(I443251), .CLK(I2702), .RSTB(I443135), .Q(I443268) );
not I_25914 (I443106,I443268);
DFFARX1 I_25915  ( .D(I443251), .CLK(I2702), .RSTB(I443135), .Q(I443299) );
and I_25916 (I443100,I443186,I443299);
nand I_25917 (I443330,I630658,I630673);
and I_25918 (I443347,I443330,I630670);
DFFARX1 I_25919  ( .D(I443347), .CLK(I2702), .RSTB(I443135), .Q(I443364) );
nor I_25920 (I443381,I443364,I443203);
not I_25921 (I443398,I443364);
nand I_25922 (I443109,I443186,I443398);
DFFARX1 I_25923  ( .D(I630688), .CLK(I2702), .RSTB(I443135), .Q(I443429) );
and I_25924 (I443446,I443429,I630667);
nor I_25925 (I443463,I443446,I443364);
nor I_25926 (I443480,I443446,I443398);
nand I_25927 (I443115,I443234,I443480);
not I_25928 (I443118,I443446);
DFFARX1 I_25929  ( .D(I443446), .CLK(I2702), .RSTB(I443135), .Q(I443097) );
DFFARX1 I_25930  ( .D(I630664), .CLK(I2702), .RSTB(I443135), .Q(I443539) );
nand I_25931 (I443556,I443539,I443251);
and I_25932 (I443573,I443234,I443556);
DFFARX1 I_25933  ( .D(I443573), .CLK(I2702), .RSTB(I443135), .Q(I443127) );
nor I_25934 (I443124,I443539,I443446);
and I_25935 (I443618,I443539,I443381);
or I_25936 (I443635,I443234,I443618);
DFFARX1 I_25937  ( .D(I443635), .CLK(I2702), .RSTB(I443135), .Q(I443112) );
nand I_25938 (I443121,I443539,I443463);
not I_25939 (I443713,I2709);
nand I_25940 (I443730,I305961,I305988);
and I_25941 (I443747,I443730,I305976);
DFFARX1 I_25942  ( .D(I443747), .CLK(I2702), .RSTB(I443713), .Q(I443764) );
not I_25943 (I443781,I443764);
DFFARX1 I_25944  ( .D(I443764), .CLK(I2702), .RSTB(I443713), .Q(I443681) );
nor I_25945 (I443812,I305964,I305988);
DFFARX1 I_25946  ( .D(I305979), .CLK(I2702), .RSTB(I443713), .Q(I443829) );
DFFARX1 I_25947  ( .D(I443829), .CLK(I2702), .RSTB(I443713), .Q(I443846) );
not I_25948 (I443684,I443846);
DFFARX1 I_25949  ( .D(I443829), .CLK(I2702), .RSTB(I443713), .Q(I443877) );
and I_25950 (I443678,I443764,I443877);
nand I_25951 (I443908,I305973,I305970);
and I_25952 (I443925,I443908,I305967);
DFFARX1 I_25953  ( .D(I443925), .CLK(I2702), .RSTB(I443713), .Q(I443942) );
nor I_25954 (I443959,I443942,I443781);
not I_25955 (I443976,I443942);
nand I_25956 (I443687,I443764,I443976);
DFFARX1 I_25957  ( .D(I305982), .CLK(I2702), .RSTB(I443713), .Q(I444007) );
and I_25958 (I444024,I444007,I305958);
nor I_25959 (I444041,I444024,I443942);
nor I_25960 (I444058,I444024,I443976);
nand I_25961 (I443693,I443812,I444058);
not I_25962 (I443696,I444024);
DFFARX1 I_25963  ( .D(I444024), .CLK(I2702), .RSTB(I443713), .Q(I443675) );
DFFARX1 I_25964  ( .D(I305985), .CLK(I2702), .RSTB(I443713), .Q(I444117) );
nand I_25965 (I444134,I444117,I443829);
and I_25966 (I444151,I443812,I444134);
DFFARX1 I_25967  ( .D(I444151), .CLK(I2702), .RSTB(I443713), .Q(I443705) );
nor I_25968 (I443702,I444117,I444024);
and I_25969 (I444196,I444117,I443959);
or I_25970 (I444213,I443812,I444196);
DFFARX1 I_25971  ( .D(I444213), .CLK(I2702), .RSTB(I443713), .Q(I443690) );
nand I_25972 (I443699,I444117,I444041);
not I_25973 (I444291,I2709);
nand I_25974 (I444308,I563161,I563149);
and I_25975 (I444325,I444308,I563143);
DFFARX1 I_25976  ( .D(I444325), .CLK(I2702), .RSTB(I444291), .Q(I444342) );
not I_25977 (I444359,I444342);
DFFARX1 I_25978  ( .D(I444342), .CLK(I2702), .RSTB(I444291), .Q(I444259) );
nor I_25979 (I444390,I563140,I563149);
DFFARX1 I_25980  ( .D(I563134), .CLK(I2702), .RSTB(I444291), .Q(I444407) );
DFFARX1 I_25981  ( .D(I444407), .CLK(I2702), .RSTB(I444291), .Q(I444424) );
not I_25982 (I444262,I444424);
DFFARX1 I_25983  ( .D(I444407), .CLK(I2702), .RSTB(I444291), .Q(I444455) );
and I_25984 (I444256,I444342,I444455);
nand I_25985 (I444486,I563137,I563152);
and I_25986 (I444503,I444486,I563164);
DFFARX1 I_25987  ( .D(I444503), .CLK(I2702), .RSTB(I444291), .Q(I444520) );
nor I_25988 (I444537,I444520,I444359);
not I_25989 (I444554,I444520);
nand I_25990 (I444265,I444342,I444554);
DFFARX1 I_25991  ( .D(I563155), .CLK(I2702), .RSTB(I444291), .Q(I444585) );
and I_25992 (I444602,I444585,I563146);
nor I_25993 (I444619,I444602,I444520);
nor I_25994 (I444636,I444602,I444554);
nand I_25995 (I444271,I444390,I444636);
not I_25996 (I444274,I444602);
DFFARX1 I_25997  ( .D(I444602), .CLK(I2702), .RSTB(I444291), .Q(I444253) );
DFFARX1 I_25998  ( .D(I563158), .CLK(I2702), .RSTB(I444291), .Q(I444695) );
nand I_25999 (I444712,I444695,I444407);
and I_26000 (I444729,I444390,I444712);
DFFARX1 I_26001  ( .D(I444729), .CLK(I2702), .RSTB(I444291), .Q(I444283) );
nor I_26002 (I444280,I444695,I444602);
and I_26003 (I444774,I444695,I444537);
or I_26004 (I444791,I444390,I444774);
DFFARX1 I_26005  ( .D(I444791), .CLK(I2702), .RSTB(I444291), .Q(I444268) );
nand I_26006 (I444277,I444695,I444619);
not I_26007 (I444869,I2709);
nand I_26008 (I444886,I407446,I407443);
and I_26009 (I444903,I444886,I407455);
DFFARX1 I_26010  ( .D(I444903), .CLK(I2702), .RSTB(I444869), .Q(I444920) );
not I_26011 (I444937,I444920);
DFFARX1 I_26012  ( .D(I444920), .CLK(I2702), .RSTB(I444869), .Q(I444837) );
nor I_26013 (I444968,I407452,I407443);
DFFARX1 I_26014  ( .D(I407458), .CLK(I2702), .RSTB(I444869), .Q(I444985) );
DFFARX1 I_26015  ( .D(I444985), .CLK(I2702), .RSTB(I444869), .Q(I445002) );
not I_26016 (I444840,I445002);
DFFARX1 I_26017  ( .D(I444985), .CLK(I2702), .RSTB(I444869), .Q(I445033) );
and I_26018 (I444834,I444920,I445033);
nand I_26019 (I445064,I407434,I407437);
and I_26020 (I445081,I445064,I407461);
DFFARX1 I_26021  ( .D(I445081), .CLK(I2702), .RSTB(I444869), .Q(I445098) );
nor I_26022 (I445115,I445098,I444937);
not I_26023 (I445132,I445098);
nand I_26024 (I444843,I444920,I445132);
DFFARX1 I_26025  ( .D(I407440), .CLK(I2702), .RSTB(I444869), .Q(I445163) );
and I_26026 (I445180,I445163,I407431);
nor I_26027 (I445197,I445180,I445098);
nor I_26028 (I445214,I445180,I445132);
nand I_26029 (I444849,I444968,I445214);
not I_26030 (I444852,I445180);
DFFARX1 I_26031  ( .D(I445180), .CLK(I2702), .RSTB(I444869), .Q(I444831) );
DFFARX1 I_26032  ( .D(I407449), .CLK(I2702), .RSTB(I444869), .Q(I445273) );
nand I_26033 (I445290,I445273,I444985);
and I_26034 (I445307,I444968,I445290);
DFFARX1 I_26035  ( .D(I445307), .CLK(I2702), .RSTB(I444869), .Q(I444861) );
nor I_26036 (I444858,I445273,I445180);
and I_26037 (I445352,I445273,I445115);
or I_26038 (I445369,I444968,I445352);
DFFARX1 I_26039  ( .D(I445369), .CLK(I2702), .RSTB(I444869), .Q(I444846) );
nand I_26040 (I444855,I445273,I445197);
not I_26041 (I445447,I2709);
nand I_26042 (I445464,I250932,I250959);
and I_26043 (I445481,I445464,I250947);
DFFARX1 I_26044  ( .D(I445481), .CLK(I2702), .RSTB(I445447), .Q(I445498) );
not I_26045 (I445515,I445498);
DFFARX1 I_26046  ( .D(I445498), .CLK(I2702), .RSTB(I445447), .Q(I445415) );
nor I_26047 (I445546,I250935,I250959);
DFFARX1 I_26048  ( .D(I250950), .CLK(I2702), .RSTB(I445447), .Q(I445563) );
DFFARX1 I_26049  ( .D(I445563), .CLK(I2702), .RSTB(I445447), .Q(I445580) );
not I_26050 (I445418,I445580);
DFFARX1 I_26051  ( .D(I445563), .CLK(I2702), .RSTB(I445447), .Q(I445611) );
and I_26052 (I445412,I445498,I445611);
nand I_26053 (I445642,I250944,I250941);
and I_26054 (I445659,I445642,I250938);
DFFARX1 I_26055  ( .D(I445659), .CLK(I2702), .RSTB(I445447), .Q(I445676) );
nor I_26056 (I445693,I445676,I445515);
not I_26057 (I445710,I445676);
nand I_26058 (I445421,I445498,I445710);
DFFARX1 I_26059  ( .D(I250953), .CLK(I2702), .RSTB(I445447), .Q(I445741) );
and I_26060 (I445758,I445741,I250929);
nor I_26061 (I445775,I445758,I445676);
nor I_26062 (I445792,I445758,I445710);
nand I_26063 (I445427,I445546,I445792);
not I_26064 (I445430,I445758);
DFFARX1 I_26065  ( .D(I445758), .CLK(I2702), .RSTB(I445447), .Q(I445409) );
DFFARX1 I_26066  ( .D(I250956), .CLK(I2702), .RSTB(I445447), .Q(I445851) );
nand I_26067 (I445868,I445851,I445563);
and I_26068 (I445885,I445546,I445868);
DFFARX1 I_26069  ( .D(I445885), .CLK(I2702), .RSTB(I445447), .Q(I445439) );
nor I_26070 (I445436,I445851,I445758);
and I_26071 (I445930,I445851,I445693);
or I_26072 (I445947,I445546,I445930);
DFFARX1 I_26073  ( .D(I445947), .CLK(I2702), .RSTB(I445447), .Q(I445424) );
nand I_26074 (I445433,I445851,I445775);
not I_26075 (I446025,I2709);
nand I_26076 (I446042,I617467,I617470);
and I_26077 (I446059,I446042,I617476);
DFFARX1 I_26078  ( .D(I446059), .CLK(I2702), .RSTB(I446025), .Q(I446076) );
not I_26079 (I446093,I446076);
DFFARX1 I_26080  ( .D(I446076), .CLK(I2702), .RSTB(I446025), .Q(I445993) );
nor I_26081 (I446124,I617473,I617470);
DFFARX1 I_26082  ( .D(I617452), .CLK(I2702), .RSTB(I446025), .Q(I446141) );
DFFARX1 I_26083  ( .D(I446141), .CLK(I2702), .RSTB(I446025), .Q(I446158) );
not I_26084 (I445996,I446158);
DFFARX1 I_26085  ( .D(I446141), .CLK(I2702), .RSTB(I446025), .Q(I446189) );
and I_26086 (I445990,I446076,I446189);
nand I_26087 (I446220,I617449,I617464);
and I_26088 (I446237,I446220,I617461);
DFFARX1 I_26089  ( .D(I446237), .CLK(I2702), .RSTB(I446025), .Q(I446254) );
nor I_26090 (I446271,I446254,I446093);
not I_26091 (I446288,I446254);
nand I_26092 (I445999,I446076,I446288);
DFFARX1 I_26093  ( .D(I617479), .CLK(I2702), .RSTB(I446025), .Q(I446319) );
and I_26094 (I446336,I446319,I617458);
nor I_26095 (I446353,I446336,I446254);
nor I_26096 (I446370,I446336,I446288);
nand I_26097 (I446005,I446124,I446370);
not I_26098 (I446008,I446336);
DFFARX1 I_26099  ( .D(I446336), .CLK(I2702), .RSTB(I446025), .Q(I445987) );
DFFARX1 I_26100  ( .D(I617455), .CLK(I2702), .RSTB(I446025), .Q(I446429) );
nand I_26101 (I446446,I446429,I446141);
and I_26102 (I446463,I446124,I446446);
DFFARX1 I_26103  ( .D(I446463), .CLK(I2702), .RSTB(I446025), .Q(I446017) );
nor I_26104 (I446014,I446429,I446336);
and I_26105 (I446508,I446429,I446271);
or I_26106 (I446525,I446124,I446508);
DFFARX1 I_26107  ( .D(I446525), .CLK(I2702), .RSTB(I446025), .Q(I446002) );
nand I_26108 (I446011,I446429,I446353);
not I_26109 (I446603,I2709);
nand I_26110 (I446620,I107266,I107248);
and I_26111 (I446637,I446620,I107260);
DFFARX1 I_26112  ( .D(I446637), .CLK(I2702), .RSTB(I446603), .Q(I446654) );
not I_26113 (I446671,I446654);
DFFARX1 I_26114  ( .D(I446654), .CLK(I2702), .RSTB(I446603), .Q(I446571) );
nor I_26115 (I446702,I107263,I107248);
DFFARX1 I_26116  ( .D(I107272), .CLK(I2702), .RSTB(I446603), .Q(I446719) );
DFFARX1 I_26117  ( .D(I446719), .CLK(I2702), .RSTB(I446603), .Q(I446736) );
not I_26118 (I446574,I446736);
DFFARX1 I_26119  ( .D(I446719), .CLK(I2702), .RSTB(I446603), .Q(I446767) );
and I_26120 (I446568,I446654,I446767);
nand I_26121 (I446798,I107251,I107275);
and I_26122 (I446815,I446798,I107254);
DFFARX1 I_26123  ( .D(I446815), .CLK(I2702), .RSTB(I446603), .Q(I446832) );
nor I_26124 (I446849,I446832,I446671);
not I_26125 (I446866,I446832);
nand I_26126 (I446577,I446654,I446866);
DFFARX1 I_26127  ( .D(I107257), .CLK(I2702), .RSTB(I446603), .Q(I446897) );
and I_26128 (I446914,I446897,I107269);
nor I_26129 (I446931,I446914,I446832);
nor I_26130 (I446948,I446914,I446866);
nand I_26131 (I446583,I446702,I446948);
not I_26132 (I446586,I446914);
DFFARX1 I_26133  ( .D(I446914), .CLK(I2702), .RSTB(I446603), .Q(I446565) );
DFFARX1 I_26134  ( .D(I107245), .CLK(I2702), .RSTB(I446603), .Q(I447007) );
nand I_26135 (I447024,I447007,I446719);
and I_26136 (I447041,I446702,I447024);
DFFARX1 I_26137  ( .D(I447041), .CLK(I2702), .RSTB(I446603), .Q(I446595) );
nor I_26138 (I446592,I447007,I446914);
and I_26139 (I447086,I447007,I446849);
or I_26140 (I447103,I446702,I447086);
DFFARX1 I_26141  ( .D(I447103), .CLK(I2702), .RSTB(I446603), .Q(I446580) );
nand I_26142 (I446589,I447007,I446931);
not I_26143 (I447181,I2709);
nand I_26144 (I447198,I530436,I530424);
and I_26145 (I447215,I447198,I530418);
DFFARX1 I_26146  ( .D(I447215), .CLK(I2702), .RSTB(I447181), .Q(I447232) );
not I_26147 (I447249,I447232);
DFFARX1 I_26148  ( .D(I447232), .CLK(I2702), .RSTB(I447181), .Q(I447149) );
nor I_26149 (I447280,I530415,I530424);
DFFARX1 I_26150  ( .D(I530409), .CLK(I2702), .RSTB(I447181), .Q(I447297) );
DFFARX1 I_26151  ( .D(I447297), .CLK(I2702), .RSTB(I447181), .Q(I447314) );
not I_26152 (I447152,I447314);
DFFARX1 I_26153  ( .D(I447297), .CLK(I2702), .RSTB(I447181), .Q(I447345) );
and I_26154 (I447146,I447232,I447345);
nand I_26155 (I447376,I530412,I530427);
and I_26156 (I447393,I447376,I530439);
DFFARX1 I_26157  ( .D(I447393), .CLK(I2702), .RSTB(I447181), .Q(I447410) );
nor I_26158 (I447427,I447410,I447249);
not I_26159 (I447444,I447410);
nand I_26160 (I447155,I447232,I447444);
DFFARX1 I_26161  ( .D(I530430), .CLK(I2702), .RSTB(I447181), .Q(I447475) );
and I_26162 (I447492,I447475,I530421);
nor I_26163 (I447509,I447492,I447410);
nor I_26164 (I447526,I447492,I447444);
nand I_26165 (I447161,I447280,I447526);
not I_26166 (I447164,I447492);
DFFARX1 I_26167  ( .D(I447492), .CLK(I2702), .RSTB(I447181), .Q(I447143) );
DFFARX1 I_26168  ( .D(I530433), .CLK(I2702), .RSTB(I447181), .Q(I447585) );
nand I_26169 (I447602,I447585,I447297);
and I_26170 (I447619,I447280,I447602);
DFFARX1 I_26171  ( .D(I447619), .CLK(I2702), .RSTB(I447181), .Q(I447173) );
nor I_26172 (I447170,I447585,I447492);
and I_26173 (I447664,I447585,I447427);
or I_26174 (I447681,I447280,I447664);
DFFARX1 I_26175  ( .D(I447681), .CLK(I2702), .RSTB(I447181), .Q(I447158) );
nand I_26176 (I447167,I447585,I447509);
not I_26177 (I447759,I2709);
nand I_26178 (I447776,I585158,I585155);
and I_26179 (I447793,I447776,I585149);
DFFARX1 I_26180  ( .D(I447793), .CLK(I2702), .RSTB(I447759), .Q(I447810) );
not I_26181 (I447827,I447810);
DFFARX1 I_26182  ( .D(I447810), .CLK(I2702), .RSTB(I447759), .Q(I447727) );
nor I_26183 (I447858,I585170,I585155);
DFFARX1 I_26184  ( .D(I585173), .CLK(I2702), .RSTB(I447759), .Q(I447875) );
DFFARX1 I_26185  ( .D(I447875), .CLK(I2702), .RSTB(I447759), .Q(I447892) );
not I_26186 (I447730,I447892);
DFFARX1 I_26187  ( .D(I447875), .CLK(I2702), .RSTB(I447759), .Q(I447923) );
and I_26188 (I447724,I447810,I447923);
nand I_26189 (I447954,I585176,I585167);
and I_26190 (I447971,I447954,I585179);
DFFARX1 I_26191  ( .D(I447971), .CLK(I2702), .RSTB(I447759), .Q(I447988) );
nor I_26192 (I448005,I447988,I447827);
not I_26193 (I448022,I447988);
nand I_26194 (I447733,I447810,I448022);
DFFARX1 I_26195  ( .D(I585152), .CLK(I2702), .RSTB(I447759), .Q(I448053) );
and I_26196 (I448070,I448053,I585161);
nor I_26197 (I448087,I448070,I447988);
nor I_26198 (I448104,I448070,I448022);
nand I_26199 (I447739,I447858,I448104);
not I_26200 (I447742,I448070);
DFFARX1 I_26201  ( .D(I448070), .CLK(I2702), .RSTB(I447759), .Q(I447721) );
DFFARX1 I_26202  ( .D(I585164), .CLK(I2702), .RSTB(I447759), .Q(I448163) );
nand I_26203 (I448180,I448163,I447875);
and I_26204 (I448197,I447858,I448180);
DFFARX1 I_26205  ( .D(I448197), .CLK(I2702), .RSTB(I447759), .Q(I447751) );
nor I_26206 (I447748,I448163,I448070);
and I_26207 (I448242,I448163,I448005);
or I_26208 (I448259,I447858,I448242);
DFFARX1 I_26209  ( .D(I448259), .CLK(I2702), .RSTB(I447759), .Q(I447736) );
nand I_26210 (I447745,I448163,I448087);
not I_26211 (I448337,I2709);
nand I_26212 (I448354,I521511,I521499);
and I_26213 (I448371,I448354,I521493);
DFFARX1 I_26214  ( .D(I448371), .CLK(I2702), .RSTB(I448337), .Q(I448388) );
not I_26215 (I448405,I448388);
DFFARX1 I_26216  ( .D(I448388), .CLK(I2702), .RSTB(I448337), .Q(I448305) );
nor I_26217 (I448436,I521490,I521499);
DFFARX1 I_26218  ( .D(I521484), .CLK(I2702), .RSTB(I448337), .Q(I448453) );
DFFARX1 I_26219  ( .D(I448453), .CLK(I2702), .RSTB(I448337), .Q(I448470) );
not I_26220 (I448308,I448470);
DFFARX1 I_26221  ( .D(I448453), .CLK(I2702), .RSTB(I448337), .Q(I448501) );
and I_26222 (I448302,I448388,I448501);
nand I_26223 (I448532,I521487,I521502);
and I_26224 (I448549,I448532,I521514);
DFFARX1 I_26225  ( .D(I448549), .CLK(I2702), .RSTB(I448337), .Q(I448566) );
nor I_26226 (I448583,I448566,I448405);
not I_26227 (I448600,I448566);
nand I_26228 (I448311,I448388,I448600);
DFFARX1 I_26229  ( .D(I521505), .CLK(I2702), .RSTB(I448337), .Q(I448631) );
and I_26230 (I448648,I448631,I521496);
nor I_26231 (I448665,I448648,I448566);
nor I_26232 (I448682,I448648,I448600);
nand I_26233 (I448317,I448436,I448682);
not I_26234 (I448320,I448648);
DFFARX1 I_26235  ( .D(I448648), .CLK(I2702), .RSTB(I448337), .Q(I448299) );
DFFARX1 I_26236  ( .D(I521508), .CLK(I2702), .RSTB(I448337), .Q(I448741) );
nand I_26237 (I448758,I448741,I448453);
and I_26238 (I448775,I448436,I448758);
DFFARX1 I_26239  ( .D(I448775), .CLK(I2702), .RSTB(I448337), .Q(I448329) );
nor I_26240 (I448326,I448741,I448648);
and I_26241 (I448820,I448741,I448583);
or I_26242 (I448837,I448436,I448820);
DFFARX1 I_26243  ( .D(I448837), .CLK(I2702), .RSTB(I448337), .Q(I448314) );
nand I_26244 (I448323,I448741,I448665);
not I_26245 (I448915,I2709);
nand I_26246 (I448932,I116956,I116938);
and I_26247 (I448949,I448932,I116950);
DFFARX1 I_26248  ( .D(I448949), .CLK(I2702), .RSTB(I448915), .Q(I448966) );
not I_26249 (I448983,I448966);
DFFARX1 I_26250  ( .D(I448966), .CLK(I2702), .RSTB(I448915), .Q(I448883) );
nor I_26251 (I449014,I116953,I116938);
DFFARX1 I_26252  ( .D(I116962), .CLK(I2702), .RSTB(I448915), .Q(I449031) );
DFFARX1 I_26253  ( .D(I449031), .CLK(I2702), .RSTB(I448915), .Q(I449048) );
not I_26254 (I448886,I449048);
DFFARX1 I_26255  ( .D(I449031), .CLK(I2702), .RSTB(I448915), .Q(I449079) );
and I_26256 (I448880,I448966,I449079);
nand I_26257 (I449110,I116941,I116965);
and I_26258 (I449127,I449110,I116944);
DFFARX1 I_26259  ( .D(I449127), .CLK(I2702), .RSTB(I448915), .Q(I449144) );
nor I_26260 (I449161,I449144,I448983);
not I_26261 (I449178,I449144);
nand I_26262 (I448889,I448966,I449178);
DFFARX1 I_26263  ( .D(I116947), .CLK(I2702), .RSTB(I448915), .Q(I449209) );
and I_26264 (I449226,I449209,I116959);
nor I_26265 (I449243,I449226,I449144);
nor I_26266 (I449260,I449226,I449178);
nand I_26267 (I448895,I449014,I449260);
not I_26268 (I448898,I449226);
DFFARX1 I_26269  ( .D(I449226), .CLK(I2702), .RSTB(I448915), .Q(I448877) );
DFFARX1 I_26270  ( .D(I116935), .CLK(I2702), .RSTB(I448915), .Q(I449319) );
nand I_26271 (I449336,I449319,I449031);
and I_26272 (I449353,I449014,I449336);
DFFARX1 I_26273  ( .D(I449353), .CLK(I2702), .RSTB(I448915), .Q(I448907) );
nor I_26274 (I448904,I449319,I449226);
and I_26275 (I449398,I449319,I449161);
or I_26276 (I449415,I449014,I449398);
DFFARX1 I_26277  ( .D(I449415), .CLK(I2702), .RSTB(I448915), .Q(I448892) );
nand I_26278 (I448901,I449319,I449243);
not I_26279 (I449493,I2709);
nand I_26280 (I449510,I137628,I137610);
and I_26281 (I449527,I449510,I137622);
DFFARX1 I_26282  ( .D(I449527), .CLK(I2702), .RSTB(I449493), .Q(I449544) );
not I_26283 (I449561,I449544);
DFFARX1 I_26284  ( .D(I449544), .CLK(I2702), .RSTB(I449493), .Q(I449461) );
nor I_26285 (I449592,I137625,I137610);
DFFARX1 I_26286  ( .D(I137634), .CLK(I2702), .RSTB(I449493), .Q(I449609) );
DFFARX1 I_26287  ( .D(I449609), .CLK(I2702), .RSTB(I449493), .Q(I449626) );
not I_26288 (I449464,I449626);
DFFARX1 I_26289  ( .D(I449609), .CLK(I2702), .RSTB(I449493), .Q(I449657) );
and I_26290 (I449458,I449544,I449657);
nand I_26291 (I449688,I137613,I137637);
and I_26292 (I449705,I449688,I137616);
DFFARX1 I_26293  ( .D(I449705), .CLK(I2702), .RSTB(I449493), .Q(I449722) );
nor I_26294 (I449739,I449722,I449561);
not I_26295 (I449756,I449722);
nand I_26296 (I449467,I449544,I449756);
DFFARX1 I_26297  ( .D(I137619), .CLK(I2702), .RSTB(I449493), .Q(I449787) );
and I_26298 (I449804,I449787,I137631);
nor I_26299 (I449821,I449804,I449722);
nor I_26300 (I449838,I449804,I449756);
nand I_26301 (I449473,I449592,I449838);
not I_26302 (I449476,I449804);
DFFARX1 I_26303  ( .D(I449804), .CLK(I2702), .RSTB(I449493), .Q(I449455) );
DFFARX1 I_26304  ( .D(I137607), .CLK(I2702), .RSTB(I449493), .Q(I449897) );
nand I_26305 (I449914,I449897,I449609);
and I_26306 (I449931,I449592,I449914);
DFFARX1 I_26307  ( .D(I449931), .CLK(I2702), .RSTB(I449493), .Q(I449485) );
nor I_26308 (I449482,I449897,I449804);
and I_26309 (I449976,I449897,I449739);
or I_26310 (I449993,I449592,I449976);
DFFARX1 I_26311  ( .D(I449993), .CLK(I2702), .RSTB(I449493), .Q(I449470) );
nand I_26312 (I449479,I449897,I449821);
not I_26313 (I450071,I2709);
nand I_26314 (I450088,I4971,I4986);
and I_26315 (I450105,I450088,I4974);
DFFARX1 I_26316  ( .D(I450105), .CLK(I2702), .RSTB(I450071), .Q(I450122) );
not I_26317 (I450139,I450122);
DFFARX1 I_26318  ( .D(I450122), .CLK(I2702), .RSTB(I450071), .Q(I450039) );
nor I_26319 (I450170,I4983,I4986);
DFFARX1 I_26320  ( .D(I4968), .CLK(I2702), .RSTB(I450071), .Q(I450187) );
DFFARX1 I_26321  ( .D(I450187), .CLK(I2702), .RSTB(I450071), .Q(I450204) );
not I_26322 (I450042,I450204);
DFFARX1 I_26323  ( .D(I450187), .CLK(I2702), .RSTB(I450071), .Q(I450235) );
and I_26324 (I450036,I450122,I450235);
nand I_26325 (I450266,I4959,I4956);
and I_26326 (I450283,I450266,I4962);
DFFARX1 I_26327  ( .D(I450283), .CLK(I2702), .RSTB(I450071), .Q(I450300) );
nor I_26328 (I450317,I450300,I450139);
not I_26329 (I450334,I450300);
nand I_26330 (I450045,I450122,I450334);
DFFARX1 I_26331  ( .D(I4965), .CLK(I2702), .RSTB(I450071), .Q(I450365) );
and I_26332 (I450382,I450365,I4977);
nor I_26333 (I450399,I450382,I450300);
nor I_26334 (I450416,I450382,I450334);
nand I_26335 (I450051,I450170,I450416);
not I_26336 (I450054,I450382);
DFFARX1 I_26337  ( .D(I450382), .CLK(I2702), .RSTB(I450071), .Q(I450033) );
DFFARX1 I_26338  ( .D(I4980), .CLK(I2702), .RSTB(I450071), .Q(I450475) );
nand I_26339 (I450492,I450475,I450187);
and I_26340 (I450509,I450170,I450492);
DFFARX1 I_26341  ( .D(I450509), .CLK(I2702), .RSTB(I450071), .Q(I450063) );
nor I_26342 (I450060,I450475,I450382);
and I_26343 (I450554,I450475,I450317);
or I_26344 (I450571,I450170,I450554);
DFFARX1 I_26345  ( .D(I450571), .CLK(I2702), .RSTB(I450071), .Q(I450048) );
nand I_26346 (I450057,I450475,I450399);
not I_26347 (I450649,I2709);
nand I_26348 (I450666,I496171,I496198);
and I_26349 (I450683,I450666,I496186);
DFFARX1 I_26350  ( .D(I450683), .CLK(I2702), .RSTB(I450649), .Q(I450700) );
not I_26351 (I450717,I450700);
DFFARX1 I_26352  ( .D(I450700), .CLK(I2702), .RSTB(I450649), .Q(I450617) );
nor I_26353 (I450748,I496177,I496198);
DFFARX1 I_26354  ( .D(I496174), .CLK(I2702), .RSTB(I450649), .Q(I450765) );
DFFARX1 I_26355  ( .D(I450765), .CLK(I2702), .RSTB(I450649), .Q(I450782) );
not I_26356 (I450620,I450782);
DFFARX1 I_26357  ( .D(I450765), .CLK(I2702), .RSTB(I450649), .Q(I450813) );
and I_26358 (I450614,I450700,I450813);
nand I_26359 (I450844,I496192,I496195);
and I_26360 (I450861,I450844,I496183);
DFFARX1 I_26361  ( .D(I450861), .CLK(I2702), .RSTB(I450649), .Q(I450878) );
nor I_26362 (I450895,I450878,I450717);
not I_26363 (I450912,I450878);
nand I_26364 (I450623,I450700,I450912);
DFFARX1 I_26365  ( .D(I496180), .CLK(I2702), .RSTB(I450649), .Q(I450943) );
and I_26366 (I450960,I450943,I496201);
nor I_26367 (I450977,I450960,I450878);
nor I_26368 (I450994,I450960,I450912);
nand I_26369 (I450629,I450748,I450994);
not I_26370 (I450632,I450960);
DFFARX1 I_26371  ( .D(I450960), .CLK(I2702), .RSTB(I450649), .Q(I450611) );
DFFARX1 I_26372  ( .D(I496189), .CLK(I2702), .RSTB(I450649), .Q(I451053) );
nand I_26373 (I451070,I451053,I450765);
and I_26374 (I451087,I450748,I451070);
DFFARX1 I_26375  ( .D(I451087), .CLK(I2702), .RSTB(I450649), .Q(I450641) );
nor I_26376 (I450638,I451053,I450960);
and I_26377 (I451132,I451053,I450895);
or I_26378 (I451149,I450748,I451132);
DFFARX1 I_26379  ( .D(I451149), .CLK(I2702), .RSTB(I450649), .Q(I450626) );
nand I_26380 (I450635,I451053,I450977);
not I_26381 (I451227,I2709);
nand I_26382 (I451244,I661497,I661500);
and I_26383 (I451261,I451244,I661506);
DFFARX1 I_26384  ( .D(I451261), .CLK(I2702), .RSTB(I451227), .Q(I451278) );
not I_26385 (I451295,I451278);
DFFARX1 I_26386  ( .D(I451278), .CLK(I2702), .RSTB(I451227), .Q(I451195) );
nor I_26387 (I451326,I661503,I661500);
DFFARX1 I_26388  ( .D(I661482), .CLK(I2702), .RSTB(I451227), .Q(I451343) );
DFFARX1 I_26389  ( .D(I451343), .CLK(I2702), .RSTB(I451227), .Q(I451360) );
not I_26390 (I451198,I451360);
DFFARX1 I_26391  ( .D(I451343), .CLK(I2702), .RSTB(I451227), .Q(I451391) );
and I_26392 (I451192,I451278,I451391);
nand I_26393 (I451422,I661479,I661494);
and I_26394 (I451439,I451422,I661491);
DFFARX1 I_26395  ( .D(I451439), .CLK(I2702), .RSTB(I451227), .Q(I451456) );
nor I_26396 (I451473,I451456,I451295);
not I_26397 (I451490,I451456);
nand I_26398 (I451201,I451278,I451490);
DFFARX1 I_26399  ( .D(I661509), .CLK(I2702), .RSTB(I451227), .Q(I451521) );
and I_26400 (I451538,I451521,I661488);
nor I_26401 (I451555,I451538,I451456);
nor I_26402 (I451572,I451538,I451490);
nand I_26403 (I451207,I451326,I451572);
not I_26404 (I451210,I451538);
DFFARX1 I_26405  ( .D(I451538), .CLK(I2702), .RSTB(I451227), .Q(I451189) );
DFFARX1 I_26406  ( .D(I661485), .CLK(I2702), .RSTB(I451227), .Q(I451631) );
nand I_26407 (I451648,I451631,I451343);
and I_26408 (I451665,I451326,I451648);
DFFARX1 I_26409  ( .D(I451665), .CLK(I2702), .RSTB(I451227), .Q(I451219) );
nor I_26410 (I451216,I451631,I451538);
and I_26411 (I451710,I451631,I451473);
or I_26412 (I451727,I451326,I451710);
DFFARX1 I_26413  ( .D(I451727), .CLK(I2702), .RSTB(I451227), .Q(I451204) );
nand I_26414 (I451213,I451631,I451555);
not I_26415 (I451805,I2709);
nand I_26416 (I451822,I198579,I198558);
and I_26417 (I451839,I451822,I198555);
DFFARX1 I_26418  ( .D(I451839), .CLK(I2702), .RSTB(I451805), .Q(I451856) );
not I_26419 (I451873,I451856);
DFFARX1 I_26420  ( .D(I451856), .CLK(I2702), .RSTB(I451805), .Q(I451773) );
nor I_26421 (I451904,I198564,I198558);
DFFARX1 I_26422  ( .D(I198552), .CLK(I2702), .RSTB(I451805), .Q(I451921) );
DFFARX1 I_26423  ( .D(I451921), .CLK(I2702), .RSTB(I451805), .Q(I451938) );
not I_26424 (I451776,I451938);
DFFARX1 I_26425  ( .D(I451921), .CLK(I2702), .RSTB(I451805), .Q(I451969) );
and I_26426 (I451770,I451856,I451969);
nand I_26427 (I452000,I198582,I198573);
and I_26428 (I452017,I452000,I198570);
DFFARX1 I_26429  ( .D(I452017), .CLK(I2702), .RSTB(I451805), .Q(I452034) );
nor I_26430 (I452051,I452034,I451873);
not I_26431 (I452068,I452034);
nand I_26432 (I451779,I451856,I452068);
DFFARX1 I_26433  ( .D(I198567), .CLK(I2702), .RSTB(I451805), .Q(I452099) );
and I_26434 (I452116,I452099,I198576);
nor I_26435 (I452133,I452116,I452034);
nor I_26436 (I452150,I452116,I452068);
nand I_26437 (I451785,I451904,I452150);
not I_26438 (I451788,I452116);
DFFARX1 I_26439  ( .D(I452116), .CLK(I2702), .RSTB(I451805), .Q(I451767) );
DFFARX1 I_26440  ( .D(I198561), .CLK(I2702), .RSTB(I451805), .Q(I452209) );
nand I_26441 (I452226,I452209,I451921);
and I_26442 (I452243,I451904,I452226);
DFFARX1 I_26443  ( .D(I452243), .CLK(I2702), .RSTB(I451805), .Q(I451797) );
nor I_26444 (I451794,I452209,I452116);
and I_26445 (I452288,I452209,I452051);
or I_26446 (I452305,I451904,I452288);
DFFARX1 I_26447  ( .D(I452305), .CLK(I2702), .RSTB(I451805), .Q(I451782) );
nand I_26448 (I451791,I452209,I452133);
not I_26449 (I452383,I2709);
nand I_26450 (I452400,I390004,I390001);
and I_26451 (I452417,I452400,I390013);
DFFARX1 I_26452  ( .D(I452417), .CLK(I2702), .RSTB(I452383), .Q(I452434) );
not I_26453 (I452451,I452434);
DFFARX1 I_26454  ( .D(I452434), .CLK(I2702), .RSTB(I452383), .Q(I452351) );
nor I_26455 (I452482,I390010,I390001);
DFFARX1 I_26456  ( .D(I390016), .CLK(I2702), .RSTB(I452383), .Q(I452499) );
DFFARX1 I_26457  ( .D(I452499), .CLK(I2702), .RSTB(I452383), .Q(I452516) );
not I_26458 (I452354,I452516);
DFFARX1 I_26459  ( .D(I452499), .CLK(I2702), .RSTB(I452383), .Q(I452547) );
and I_26460 (I452348,I452434,I452547);
nand I_26461 (I452578,I389992,I389995);
and I_26462 (I452595,I452578,I390019);
DFFARX1 I_26463  ( .D(I452595), .CLK(I2702), .RSTB(I452383), .Q(I452612) );
nor I_26464 (I452629,I452612,I452451);
not I_26465 (I452646,I452612);
nand I_26466 (I452357,I452434,I452646);
DFFARX1 I_26467  ( .D(I389998), .CLK(I2702), .RSTB(I452383), .Q(I452677) );
and I_26468 (I452694,I452677,I389989);
nor I_26469 (I452711,I452694,I452612);
nor I_26470 (I452728,I452694,I452646);
nand I_26471 (I452363,I452482,I452728);
not I_26472 (I452366,I452694);
DFFARX1 I_26473  ( .D(I452694), .CLK(I2702), .RSTB(I452383), .Q(I452345) );
DFFARX1 I_26474  ( .D(I390007), .CLK(I2702), .RSTB(I452383), .Q(I452787) );
nand I_26475 (I452804,I452787,I452499);
and I_26476 (I452821,I452482,I452804);
DFFARX1 I_26477  ( .D(I452821), .CLK(I2702), .RSTB(I452383), .Q(I452375) );
nor I_26478 (I452372,I452787,I452694);
and I_26479 (I452866,I452787,I452629);
or I_26480 (I452883,I452482,I452866);
DFFARX1 I_26481  ( .D(I452883), .CLK(I2702), .RSTB(I452383), .Q(I452360) );
nand I_26482 (I452369,I452787,I452711);
not I_26483 (I452961,I2709);
nand I_26484 (I452978,I118894,I118876);
and I_26485 (I452995,I452978,I118888);
DFFARX1 I_26486  ( .D(I452995), .CLK(I2702), .RSTB(I452961), .Q(I453012) );
not I_26487 (I453029,I453012);
DFFARX1 I_26488  ( .D(I453012), .CLK(I2702), .RSTB(I452961), .Q(I452929) );
nor I_26489 (I453060,I118891,I118876);
DFFARX1 I_26490  ( .D(I118900), .CLK(I2702), .RSTB(I452961), .Q(I453077) );
DFFARX1 I_26491  ( .D(I453077), .CLK(I2702), .RSTB(I452961), .Q(I453094) );
not I_26492 (I452932,I453094);
DFFARX1 I_26493  ( .D(I453077), .CLK(I2702), .RSTB(I452961), .Q(I453125) );
and I_26494 (I452926,I453012,I453125);
nand I_26495 (I453156,I118879,I118903);
and I_26496 (I453173,I453156,I118882);
DFFARX1 I_26497  ( .D(I453173), .CLK(I2702), .RSTB(I452961), .Q(I453190) );
nor I_26498 (I453207,I453190,I453029);
not I_26499 (I453224,I453190);
nand I_26500 (I452935,I453012,I453224);
DFFARX1 I_26501  ( .D(I118885), .CLK(I2702), .RSTB(I452961), .Q(I453255) );
and I_26502 (I453272,I453255,I118897);
nor I_26503 (I453289,I453272,I453190);
nor I_26504 (I453306,I453272,I453224);
nand I_26505 (I452941,I453060,I453306);
not I_26506 (I452944,I453272);
DFFARX1 I_26507  ( .D(I453272), .CLK(I2702), .RSTB(I452961), .Q(I452923) );
DFFARX1 I_26508  ( .D(I118873), .CLK(I2702), .RSTB(I452961), .Q(I453365) );
nand I_26509 (I453382,I453365,I453077);
and I_26510 (I453399,I453060,I453382);
DFFARX1 I_26511  ( .D(I453399), .CLK(I2702), .RSTB(I452961), .Q(I452953) );
nor I_26512 (I452950,I453365,I453272);
and I_26513 (I453444,I453365,I453207);
or I_26514 (I453461,I453060,I453444);
DFFARX1 I_26515  ( .D(I453461), .CLK(I2702), .RSTB(I452961), .Q(I452938) );
nand I_26516 (I452947,I453365,I453289);
not I_26517 (I453539,I2709);
nand I_26518 (I453556,I26850,I26865);
and I_26519 (I453573,I453556,I26853);
DFFARX1 I_26520  ( .D(I453573), .CLK(I2702), .RSTB(I453539), .Q(I453590) );
not I_26521 (I453607,I453590);
DFFARX1 I_26522  ( .D(I453590), .CLK(I2702), .RSTB(I453539), .Q(I453507) );
nor I_26523 (I453638,I26862,I26865);
DFFARX1 I_26524  ( .D(I26847), .CLK(I2702), .RSTB(I453539), .Q(I453655) );
DFFARX1 I_26525  ( .D(I453655), .CLK(I2702), .RSTB(I453539), .Q(I453672) );
not I_26526 (I453510,I453672);
DFFARX1 I_26527  ( .D(I453655), .CLK(I2702), .RSTB(I453539), .Q(I453703) );
and I_26528 (I453504,I453590,I453703);
nand I_26529 (I453734,I26838,I26835);
and I_26530 (I453751,I453734,I26841);
DFFARX1 I_26531  ( .D(I453751), .CLK(I2702), .RSTB(I453539), .Q(I453768) );
nor I_26532 (I453785,I453768,I453607);
not I_26533 (I453802,I453768);
nand I_26534 (I453513,I453590,I453802);
DFFARX1 I_26535  ( .D(I26844), .CLK(I2702), .RSTB(I453539), .Q(I453833) );
and I_26536 (I453850,I453833,I26856);
nor I_26537 (I453867,I453850,I453768);
nor I_26538 (I453884,I453850,I453802);
nand I_26539 (I453519,I453638,I453884);
not I_26540 (I453522,I453850);
DFFARX1 I_26541  ( .D(I453850), .CLK(I2702), .RSTB(I453539), .Q(I453501) );
DFFARX1 I_26542  ( .D(I26859), .CLK(I2702), .RSTB(I453539), .Q(I453943) );
nand I_26543 (I453960,I453943,I453655);
and I_26544 (I453977,I453638,I453960);
DFFARX1 I_26545  ( .D(I453977), .CLK(I2702), .RSTB(I453539), .Q(I453531) );
nor I_26546 (I453528,I453943,I453850);
and I_26547 (I454022,I453943,I453785);
or I_26548 (I454039,I453638,I454022);
DFFARX1 I_26549  ( .D(I454039), .CLK(I2702), .RSTB(I453539), .Q(I453516) );
nand I_26550 (I453525,I453943,I453867);
not I_26551 (I454117,I2709);
nand I_26552 (I454134,I628160,I628163);
and I_26553 (I454151,I454134,I628169);
DFFARX1 I_26554  ( .D(I454151), .CLK(I2702), .RSTB(I454117), .Q(I454168) );
not I_26555 (I454185,I454168);
DFFARX1 I_26556  ( .D(I454168), .CLK(I2702), .RSTB(I454117), .Q(I454085) );
nor I_26557 (I454216,I628166,I628163);
DFFARX1 I_26558  ( .D(I628145), .CLK(I2702), .RSTB(I454117), .Q(I454233) );
DFFARX1 I_26559  ( .D(I454233), .CLK(I2702), .RSTB(I454117), .Q(I454250) );
not I_26560 (I454088,I454250);
DFFARX1 I_26561  ( .D(I454233), .CLK(I2702), .RSTB(I454117), .Q(I454281) );
and I_26562 (I454082,I454168,I454281);
nand I_26563 (I454312,I628142,I628157);
and I_26564 (I454329,I454312,I628154);
DFFARX1 I_26565  ( .D(I454329), .CLK(I2702), .RSTB(I454117), .Q(I454346) );
nor I_26566 (I454363,I454346,I454185);
not I_26567 (I454380,I454346);
nand I_26568 (I454091,I454168,I454380);
DFFARX1 I_26569  ( .D(I628172), .CLK(I2702), .RSTB(I454117), .Q(I454411) );
and I_26570 (I454428,I454411,I628151);
nor I_26571 (I454445,I454428,I454346);
nor I_26572 (I454462,I454428,I454380);
nand I_26573 (I454097,I454216,I454462);
not I_26574 (I454100,I454428);
DFFARX1 I_26575  ( .D(I454428), .CLK(I2702), .RSTB(I454117), .Q(I454079) );
DFFARX1 I_26576  ( .D(I628148), .CLK(I2702), .RSTB(I454117), .Q(I454521) );
nand I_26577 (I454538,I454521,I454233);
and I_26578 (I454555,I454216,I454538);
DFFARX1 I_26579  ( .D(I454555), .CLK(I2702), .RSTB(I454117), .Q(I454109) );
nor I_26580 (I454106,I454521,I454428);
and I_26581 (I454600,I454521,I454363);
or I_26582 (I454617,I454216,I454600);
DFFARX1 I_26583  ( .D(I454617), .CLK(I2702), .RSTB(I454117), .Q(I454094) );
nand I_26584 (I454103,I454521,I454445);
not I_26585 (I454695,I2709);
nand I_26586 (I454712,I611933,I611930);
and I_26587 (I454729,I454712,I611924);
DFFARX1 I_26588  ( .D(I454729), .CLK(I2702), .RSTB(I454695), .Q(I454746) );
not I_26589 (I454763,I454746);
DFFARX1 I_26590  ( .D(I454746), .CLK(I2702), .RSTB(I454695), .Q(I454663) );
nor I_26591 (I454794,I611945,I611930);
DFFARX1 I_26592  ( .D(I611948), .CLK(I2702), .RSTB(I454695), .Q(I454811) );
DFFARX1 I_26593  ( .D(I454811), .CLK(I2702), .RSTB(I454695), .Q(I454828) );
not I_26594 (I454666,I454828);
DFFARX1 I_26595  ( .D(I454811), .CLK(I2702), .RSTB(I454695), .Q(I454859) );
and I_26596 (I454660,I454746,I454859);
nand I_26597 (I454890,I611951,I611942);
and I_26598 (I454907,I454890,I611954);
DFFARX1 I_26599  ( .D(I454907), .CLK(I2702), .RSTB(I454695), .Q(I454924) );
nor I_26600 (I454941,I454924,I454763);
not I_26601 (I454958,I454924);
nand I_26602 (I454669,I454746,I454958);
DFFARX1 I_26603  ( .D(I611927), .CLK(I2702), .RSTB(I454695), .Q(I454989) );
and I_26604 (I455006,I454989,I611936);
nor I_26605 (I455023,I455006,I454924);
nor I_26606 (I455040,I455006,I454958);
nand I_26607 (I454675,I454794,I455040);
not I_26608 (I454678,I455006);
DFFARX1 I_26609  ( .D(I455006), .CLK(I2702), .RSTB(I454695), .Q(I454657) );
DFFARX1 I_26610  ( .D(I611939), .CLK(I2702), .RSTB(I454695), .Q(I455099) );
nand I_26611 (I455116,I455099,I454811);
and I_26612 (I455133,I454794,I455116);
DFFARX1 I_26613  ( .D(I455133), .CLK(I2702), .RSTB(I454695), .Q(I454687) );
nor I_26614 (I454684,I455099,I455006);
and I_26615 (I455178,I455099,I454941);
or I_26616 (I455195,I454794,I455178);
DFFARX1 I_26617  ( .D(I455195), .CLK(I2702), .RSTB(I454695), .Q(I454672) );
nand I_26618 (I454681,I455099,I455023);
not I_26619 (I455273,I2709);
nand I_26620 (I455290,I580993,I580990);
and I_26621 (I455307,I455290,I580984);
DFFARX1 I_26622  ( .D(I455307), .CLK(I2702), .RSTB(I455273), .Q(I455324) );
not I_26623 (I455341,I455324);
DFFARX1 I_26624  ( .D(I455324), .CLK(I2702), .RSTB(I455273), .Q(I455241) );
nor I_26625 (I455372,I581005,I580990);
DFFARX1 I_26626  ( .D(I581008), .CLK(I2702), .RSTB(I455273), .Q(I455389) );
DFFARX1 I_26627  ( .D(I455389), .CLK(I2702), .RSTB(I455273), .Q(I455406) );
not I_26628 (I455244,I455406);
DFFARX1 I_26629  ( .D(I455389), .CLK(I2702), .RSTB(I455273), .Q(I455437) );
and I_26630 (I455238,I455324,I455437);
nand I_26631 (I455468,I581011,I581002);
and I_26632 (I455485,I455468,I581014);
DFFARX1 I_26633  ( .D(I455485), .CLK(I2702), .RSTB(I455273), .Q(I455502) );
nor I_26634 (I455519,I455502,I455341);
not I_26635 (I455536,I455502);
nand I_26636 (I455247,I455324,I455536);
DFFARX1 I_26637  ( .D(I580987), .CLK(I2702), .RSTB(I455273), .Q(I455567) );
and I_26638 (I455584,I455567,I580996);
nor I_26639 (I455601,I455584,I455502);
nor I_26640 (I455618,I455584,I455536);
nand I_26641 (I455253,I455372,I455618);
not I_26642 (I455256,I455584);
DFFARX1 I_26643  ( .D(I455584), .CLK(I2702), .RSTB(I455273), .Q(I455235) );
DFFARX1 I_26644  ( .D(I580999), .CLK(I2702), .RSTB(I455273), .Q(I455677) );
nand I_26645 (I455694,I455677,I455389);
and I_26646 (I455711,I455372,I455694);
DFFARX1 I_26647  ( .D(I455711), .CLK(I2702), .RSTB(I455273), .Q(I455265) );
nor I_26648 (I455262,I455677,I455584);
and I_26649 (I455756,I455677,I455519);
or I_26650 (I455773,I455372,I455756);
DFFARX1 I_26651  ( .D(I455773), .CLK(I2702), .RSTB(I455273), .Q(I455250) );
nand I_26652 (I455259,I455677,I455601);
not I_26653 (I455851,I2709);
nand I_26654 (I455868,I712919,I712931);
and I_26655 (I455885,I455868,I712904);
DFFARX1 I_26656  ( .D(I455885), .CLK(I2702), .RSTB(I455851), .Q(I455902) );
not I_26657 (I455919,I455902);
DFFARX1 I_26658  ( .D(I455902), .CLK(I2702), .RSTB(I455851), .Q(I455819) );
nor I_26659 (I455950,I712922,I712931);
DFFARX1 I_26660  ( .D(I712913), .CLK(I2702), .RSTB(I455851), .Q(I455967) );
DFFARX1 I_26661  ( .D(I455967), .CLK(I2702), .RSTB(I455851), .Q(I455984) );
not I_26662 (I455822,I455984);
DFFARX1 I_26663  ( .D(I455967), .CLK(I2702), .RSTB(I455851), .Q(I456015) );
and I_26664 (I455816,I455902,I456015);
nand I_26665 (I456046,I712910,I712916);
and I_26666 (I456063,I456046,I712928);
DFFARX1 I_26667  ( .D(I456063), .CLK(I2702), .RSTB(I455851), .Q(I456080) );
nor I_26668 (I456097,I456080,I455919);
not I_26669 (I456114,I456080);
nand I_26670 (I455825,I455902,I456114);
DFFARX1 I_26671  ( .D(I712934), .CLK(I2702), .RSTB(I455851), .Q(I456145) );
and I_26672 (I456162,I456145,I712925);
nor I_26673 (I456179,I456162,I456080);
nor I_26674 (I456196,I456162,I456114);
nand I_26675 (I455831,I455950,I456196);
not I_26676 (I455834,I456162);
DFFARX1 I_26677  ( .D(I456162), .CLK(I2702), .RSTB(I455851), .Q(I455813) );
DFFARX1 I_26678  ( .D(I712907), .CLK(I2702), .RSTB(I455851), .Q(I456255) );
nand I_26679 (I456272,I456255,I455967);
and I_26680 (I456289,I455950,I456272);
DFFARX1 I_26681  ( .D(I456289), .CLK(I2702), .RSTB(I455851), .Q(I455843) );
nor I_26682 (I455840,I456255,I456162);
and I_26683 (I456334,I456255,I456097);
or I_26684 (I456351,I455950,I456334);
DFFARX1 I_26685  ( .D(I456351), .CLK(I2702), .RSTB(I455851), .Q(I455828) );
nand I_26686 (I455837,I456255,I456179);
not I_26687 (I456429,I2709);
nand I_26688 (I456446,I534601,I534589);
and I_26689 (I456463,I456446,I534583);
DFFARX1 I_26690  ( .D(I456463), .CLK(I2702), .RSTB(I456429), .Q(I456480) );
not I_26691 (I456497,I456480);
DFFARX1 I_26692  ( .D(I456480), .CLK(I2702), .RSTB(I456429), .Q(I456397) );
nor I_26693 (I456528,I534580,I534589);
DFFARX1 I_26694  ( .D(I534574), .CLK(I2702), .RSTB(I456429), .Q(I456545) );
DFFARX1 I_26695  ( .D(I456545), .CLK(I2702), .RSTB(I456429), .Q(I456562) );
not I_26696 (I456400,I456562);
DFFARX1 I_26697  ( .D(I456545), .CLK(I2702), .RSTB(I456429), .Q(I456593) );
and I_26698 (I456394,I456480,I456593);
nand I_26699 (I456624,I534577,I534592);
and I_26700 (I456641,I456624,I534604);
DFFARX1 I_26701  ( .D(I456641), .CLK(I2702), .RSTB(I456429), .Q(I456658) );
nor I_26702 (I456675,I456658,I456497);
not I_26703 (I456692,I456658);
nand I_26704 (I456403,I456480,I456692);
DFFARX1 I_26705  ( .D(I534595), .CLK(I2702), .RSTB(I456429), .Q(I456723) );
and I_26706 (I456740,I456723,I534586);
nor I_26707 (I456757,I456740,I456658);
nor I_26708 (I456774,I456740,I456692);
nand I_26709 (I456409,I456528,I456774);
not I_26710 (I456412,I456740);
DFFARX1 I_26711  ( .D(I456740), .CLK(I2702), .RSTB(I456429), .Q(I456391) );
DFFARX1 I_26712  ( .D(I534598), .CLK(I2702), .RSTB(I456429), .Q(I456833) );
nand I_26713 (I456850,I456833,I456545);
and I_26714 (I456867,I456528,I456850);
DFFARX1 I_26715  ( .D(I456867), .CLK(I2702), .RSTB(I456429), .Q(I456421) );
nor I_26716 (I456418,I456833,I456740);
and I_26717 (I456912,I456833,I456675);
or I_26718 (I456929,I456528,I456912);
DFFARX1 I_26719  ( .D(I456929), .CLK(I2702), .RSTB(I456429), .Q(I456406) );
nand I_26720 (I456415,I456833,I456757);
not I_26721 (I457007,I2709);
nand I_26722 (I457024,I511396,I511384);
and I_26723 (I457041,I457024,I511378);
DFFARX1 I_26724  ( .D(I457041), .CLK(I2702), .RSTB(I457007), .Q(I457058) );
not I_26725 (I457075,I457058);
DFFARX1 I_26726  ( .D(I457058), .CLK(I2702), .RSTB(I457007), .Q(I456975) );
nor I_26727 (I457106,I511375,I511384);
DFFARX1 I_26728  ( .D(I511369), .CLK(I2702), .RSTB(I457007), .Q(I457123) );
DFFARX1 I_26729  ( .D(I457123), .CLK(I2702), .RSTB(I457007), .Q(I457140) );
not I_26730 (I456978,I457140);
DFFARX1 I_26731  ( .D(I457123), .CLK(I2702), .RSTB(I457007), .Q(I457171) );
and I_26732 (I456972,I457058,I457171);
nand I_26733 (I457202,I511372,I511387);
and I_26734 (I457219,I457202,I511399);
DFFARX1 I_26735  ( .D(I457219), .CLK(I2702), .RSTB(I457007), .Q(I457236) );
nor I_26736 (I457253,I457236,I457075);
not I_26737 (I457270,I457236);
nand I_26738 (I456981,I457058,I457270);
DFFARX1 I_26739  ( .D(I511390), .CLK(I2702), .RSTB(I457007), .Q(I457301) );
and I_26740 (I457318,I457301,I511381);
nor I_26741 (I457335,I457318,I457236);
nor I_26742 (I457352,I457318,I457270);
nand I_26743 (I456987,I457106,I457352);
not I_26744 (I456990,I457318);
DFFARX1 I_26745  ( .D(I457318), .CLK(I2702), .RSTB(I457007), .Q(I456969) );
DFFARX1 I_26746  ( .D(I511393), .CLK(I2702), .RSTB(I457007), .Q(I457411) );
nand I_26747 (I457428,I457411,I457123);
and I_26748 (I457445,I457106,I457428);
DFFARX1 I_26749  ( .D(I457445), .CLK(I2702), .RSTB(I457007), .Q(I456999) );
nor I_26750 (I456996,I457411,I457318);
and I_26751 (I457490,I457411,I457253);
or I_26752 (I457507,I457106,I457490);
DFFARX1 I_26753  ( .D(I457507), .CLK(I2702), .RSTB(I457007), .Q(I456984) );
nand I_26754 (I456993,I457411,I457335);
not I_26755 (I457585,I2709);
nand I_26756 (I457602,I684770,I684773);
and I_26757 (I457619,I457602,I684779);
DFFARX1 I_26758  ( .D(I457619), .CLK(I2702), .RSTB(I457585), .Q(I457636) );
not I_26759 (I457653,I457636);
DFFARX1 I_26760  ( .D(I457636), .CLK(I2702), .RSTB(I457585), .Q(I457553) );
nor I_26761 (I457684,I684776,I684773);
DFFARX1 I_26762  ( .D(I684755), .CLK(I2702), .RSTB(I457585), .Q(I457701) );
DFFARX1 I_26763  ( .D(I457701), .CLK(I2702), .RSTB(I457585), .Q(I457718) );
not I_26764 (I457556,I457718);
DFFARX1 I_26765  ( .D(I457701), .CLK(I2702), .RSTB(I457585), .Q(I457749) );
and I_26766 (I457550,I457636,I457749);
nand I_26767 (I457780,I684752,I684767);
and I_26768 (I457797,I457780,I684764);
DFFARX1 I_26769  ( .D(I457797), .CLK(I2702), .RSTB(I457585), .Q(I457814) );
nor I_26770 (I457831,I457814,I457653);
not I_26771 (I457848,I457814);
nand I_26772 (I457559,I457636,I457848);
DFFARX1 I_26773  ( .D(I684782), .CLK(I2702), .RSTB(I457585), .Q(I457879) );
and I_26774 (I457896,I457879,I684761);
nor I_26775 (I457913,I457896,I457814);
nor I_26776 (I457930,I457896,I457848);
nand I_26777 (I457565,I457684,I457930);
not I_26778 (I457568,I457896);
DFFARX1 I_26779  ( .D(I457896), .CLK(I2702), .RSTB(I457585), .Q(I457547) );
DFFARX1 I_26780  ( .D(I684758), .CLK(I2702), .RSTB(I457585), .Q(I457989) );
nand I_26781 (I458006,I457989,I457701);
and I_26782 (I458023,I457684,I458006);
DFFARX1 I_26783  ( .D(I458023), .CLK(I2702), .RSTB(I457585), .Q(I457577) );
nor I_26784 (I457574,I457989,I457896);
and I_26785 (I458068,I457989,I457831);
or I_26786 (I458085,I457684,I458068);
DFFARX1 I_26787  ( .D(I458085), .CLK(I2702), .RSTB(I457585), .Q(I457562) );
nand I_26788 (I457571,I457989,I457913);
not I_26789 (I458163,I2709);
nand I_26790 (I458180,I679738,I679741);
and I_26791 (I458197,I458180,I679747);
DFFARX1 I_26792  ( .D(I458197), .CLK(I2702), .RSTB(I458163), .Q(I458214) );
not I_26793 (I458231,I458214);
DFFARX1 I_26794  ( .D(I458214), .CLK(I2702), .RSTB(I458163), .Q(I458131) );
nor I_26795 (I458262,I679744,I679741);
DFFARX1 I_26796  ( .D(I679723), .CLK(I2702), .RSTB(I458163), .Q(I458279) );
DFFARX1 I_26797  ( .D(I458279), .CLK(I2702), .RSTB(I458163), .Q(I458296) );
not I_26798 (I458134,I458296);
DFFARX1 I_26799  ( .D(I458279), .CLK(I2702), .RSTB(I458163), .Q(I458327) );
and I_26800 (I458128,I458214,I458327);
nand I_26801 (I458358,I679720,I679735);
and I_26802 (I458375,I458358,I679732);
DFFARX1 I_26803  ( .D(I458375), .CLK(I2702), .RSTB(I458163), .Q(I458392) );
nor I_26804 (I458409,I458392,I458231);
not I_26805 (I458426,I458392);
nand I_26806 (I458137,I458214,I458426);
DFFARX1 I_26807  ( .D(I679750), .CLK(I2702), .RSTB(I458163), .Q(I458457) );
and I_26808 (I458474,I458457,I679729);
nor I_26809 (I458491,I458474,I458392);
nor I_26810 (I458508,I458474,I458426);
nand I_26811 (I458143,I458262,I458508);
not I_26812 (I458146,I458474);
DFFARX1 I_26813  ( .D(I458474), .CLK(I2702), .RSTB(I458163), .Q(I458125) );
DFFARX1 I_26814  ( .D(I679726), .CLK(I2702), .RSTB(I458163), .Q(I458567) );
nand I_26815 (I458584,I458567,I458279);
and I_26816 (I458601,I458262,I458584);
DFFARX1 I_26817  ( .D(I458601), .CLK(I2702), .RSTB(I458163), .Q(I458155) );
nor I_26818 (I458152,I458567,I458474);
and I_26819 (I458646,I458567,I458409);
or I_26820 (I458663,I458262,I458646);
DFFARX1 I_26821  ( .D(I458663), .CLK(I2702), .RSTB(I458163), .Q(I458140) );
nand I_26822 (I458149,I458567,I458491);
not I_26823 (I458741,I2709);
nand I_26824 (I458758,I221322,I221307);
and I_26825 (I458775,I458758,I221316);
DFFARX1 I_26826  ( .D(I458775), .CLK(I2702), .RSTB(I458741), .Q(I458792) );
not I_26827 (I458809,I458792);
DFFARX1 I_26828  ( .D(I458792), .CLK(I2702), .RSTB(I458741), .Q(I458709) );
nor I_26829 (I458840,I221325,I221307);
DFFARX1 I_26830  ( .D(I221304), .CLK(I2702), .RSTB(I458741), .Q(I458857) );
DFFARX1 I_26831  ( .D(I458857), .CLK(I2702), .RSTB(I458741), .Q(I458874) );
not I_26832 (I458712,I458874);
DFFARX1 I_26833  ( .D(I458857), .CLK(I2702), .RSTB(I458741), .Q(I458905) );
and I_26834 (I458706,I458792,I458905);
nand I_26835 (I458936,I221328,I221301);
and I_26836 (I458953,I458936,I221319);
DFFARX1 I_26837  ( .D(I458953), .CLK(I2702), .RSTB(I458741), .Q(I458970) );
nor I_26838 (I458987,I458970,I458809);
not I_26839 (I459004,I458970);
nand I_26840 (I458715,I458792,I459004);
DFFARX1 I_26841  ( .D(I221313), .CLK(I2702), .RSTB(I458741), .Q(I459035) );
and I_26842 (I459052,I459035,I221298);
nor I_26843 (I459069,I459052,I458970);
nor I_26844 (I459086,I459052,I459004);
nand I_26845 (I458721,I458840,I459086);
not I_26846 (I458724,I459052);
DFFARX1 I_26847  ( .D(I459052), .CLK(I2702), .RSTB(I458741), .Q(I458703) );
DFFARX1 I_26848  ( .D(I221310), .CLK(I2702), .RSTB(I458741), .Q(I459145) );
nand I_26849 (I459162,I459145,I458857);
and I_26850 (I459179,I458840,I459162);
DFFARX1 I_26851  ( .D(I459179), .CLK(I2702), .RSTB(I458741), .Q(I458733) );
nor I_26852 (I458730,I459145,I459052);
and I_26853 (I459224,I459145,I458987);
or I_26854 (I459241,I458840,I459224);
DFFARX1 I_26855  ( .D(I459241), .CLK(I2702), .RSTB(I458741), .Q(I458718) );
nand I_26856 (I458727,I459145,I459069);
not I_26857 (I459319,I2709);
nand I_26858 (I459336,I69798,I69780);
and I_26859 (I459353,I459336,I69792);
DFFARX1 I_26860  ( .D(I459353), .CLK(I2702), .RSTB(I459319), .Q(I459370) );
not I_26861 (I459387,I459370);
DFFARX1 I_26862  ( .D(I459370), .CLK(I2702), .RSTB(I459319), .Q(I459287) );
nor I_26863 (I459418,I69795,I69780);
DFFARX1 I_26864  ( .D(I69804), .CLK(I2702), .RSTB(I459319), .Q(I459435) );
DFFARX1 I_26865  ( .D(I459435), .CLK(I2702), .RSTB(I459319), .Q(I459452) );
not I_26866 (I459290,I459452);
DFFARX1 I_26867  ( .D(I459435), .CLK(I2702), .RSTB(I459319), .Q(I459483) );
and I_26868 (I459284,I459370,I459483);
nand I_26869 (I459514,I69783,I69807);
and I_26870 (I459531,I459514,I69786);
DFFARX1 I_26871  ( .D(I459531), .CLK(I2702), .RSTB(I459319), .Q(I459548) );
nor I_26872 (I459565,I459548,I459387);
not I_26873 (I459582,I459548);
nand I_26874 (I459293,I459370,I459582);
DFFARX1 I_26875  ( .D(I69789), .CLK(I2702), .RSTB(I459319), .Q(I459613) );
and I_26876 (I459630,I459613,I69801);
nor I_26877 (I459647,I459630,I459548);
nor I_26878 (I459664,I459630,I459582);
nand I_26879 (I459299,I459418,I459664);
not I_26880 (I459302,I459630);
DFFARX1 I_26881  ( .D(I459630), .CLK(I2702), .RSTB(I459319), .Q(I459281) );
DFFARX1 I_26882  ( .D(I69777), .CLK(I2702), .RSTB(I459319), .Q(I459723) );
nand I_26883 (I459740,I459723,I459435);
and I_26884 (I459757,I459418,I459740);
DFFARX1 I_26885  ( .D(I459757), .CLK(I2702), .RSTB(I459319), .Q(I459311) );
nor I_26886 (I459308,I459723,I459630);
and I_26887 (I459802,I459723,I459565);
or I_26888 (I459819,I459418,I459802);
DFFARX1 I_26889  ( .D(I459819), .CLK(I2702), .RSTB(I459319), .Q(I459296) );
nand I_26890 (I459305,I459723,I459647);
not I_26891 (I459897,I2709);
nand I_26892 (I459914,I323199,I323226);
and I_26893 (I459931,I459914,I323214);
DFFARX1 I_26894  ( .D(I459931), .CLK(I2702), .RSTB(I459897), .Q(I459948) );
not I_26895 (I459965,I459948);
DFFARX1 I_26896  ( .D(I459948), .CLK(I2702), .RSTB(I459897), .Q(I459865) );
nor I_26897 (I459996,I323202,I323226);
DFFARX1 I_26898  ( .D(I323217), .CLK(I2702), .RSTB(I459897), .Q(I460013) );
DFFARX1 I_26899  ( .D(I460013), .CLK(I2702), .RSTB(I459897), .Q(I460030) );
not I_26900 (I459868,I460030);
DFFARX1 I_26901  ( .D(I460013), .CLK(I2702), .RSTB(I459897), .Q(I460061) );
and I_26902 (I459862,I459948,I460061);
nand I_26903 (I460092,I323211,I323208);
and I_26904 (I460109,I460092,I323205);
DFFARX1 I_26905  ( .D(I460109), .CLK(I2702), .RSTB(I459897), .Q(I460126) );
nor I_26906 (I460143,I460126,I459965);
not I_26907 (I460160,I460126);
nand I_26908 (I459871,I459948,I460160);
DFFARX1 I_26909  ( .D(I323220), .CLK(I2702), .RSTB(I459897), .Q(I460191) );
and I_26910 (I460208,I460191,I323196);
nor I_26911 (I460225,I460208,I460126);
nor I_26912 (I460242,I460208,I460160);
nand I_26913 (I459877,I459996,I460242);
not I_26914 (I459880,I460208);
DFFARX1 I_26915  ( .D(I460208), .CLK(I2702), .RSTB(I459897), .Q(I459859) );
DFFARX1 I_26916  ( .D(I323223), .CLK(I2702), .RSTB(I459897), .Q(I460301) );
nand I_26917 (I460318,I460301,I460013);
and I_26918 (I460335,I459996,I460318);
DFFARX1 I_26919  ( .D(I460335), .CLK(I2702), .RSTB(I459897), .Q(I459889) );
nor I_26920 (I459886,I460301,I460208);
and I_26921 (I460380,I460301,I460143);
or I_26922 (I460397,I459996,I460380);
DFFARX1 I_26923  ( .D(I460397), .CLK(I2702), .RSTB(I459897), .Q(I459874) );
nand I_26924 (I459883,I460301,I460225);
not I_26925 (I460475,I2709);
nand I_26926 (I460492,I240338,I240341);
and I_26927 (I460509,I460492,I240347);
DFFARX1 I_26928  ( .D(I460509), .CLK(I2702), .RSTB(I460475), .Q(I460526) );
not I_26929 (I460543,I460526);
DFFARX1 I_26930  ( .D(I460526), .CLK(I2702), .RSTB(I460475), .Q(I460443) );
nor I_26931 (I460574,I240359,I240341);
DFFARX1 I_26932  ( .D(I240350), .CLK(I2702), .RSTB(I460475), .Q(I460591) );
DFFARX1 I_26933  ( .D(I460591), .CLK(I2702), .RSTB(I460475), .Q(I460608) );
not I_26934 (I460446,I460608);
DFFARX1 I_26935  ( .D(I460591), .CLK(I2702), .RSTB(I460475), .Q(I460639) );
and I_26936 (I460440,I460526,I460639);
nand I_26937 (I460670,I240356,I240353);
and I_26938 (I460687,I460670,I240365);
DFFARX1 I_26939  ( .D(I460687), .CLK(I2702), .RSTB(I460475), .Q(I460704) );
nor I_26940 (I460721,I460704,I460543);
not I_26941 (I460738,I460704);
nand I_26942 (I460449,I460526,I460738);
DFFARX1 I_26943  ( .D(I240362), .CLK(I2702), .RSTB(I460475), .Q(I460769) );
and I_26944 (I460786,I460769,I240368);
nor I_26945 (I460803,I460786,I460704);
nor I_26946 (I460820,I460786,I460738);
nand I_26947 (I460455,I460574,I460820);
not I_26948 (I460458,I460786);
DFFARX1 I_26949  ( .D(I460786), .CLK(I2702), .RSTB(I460475), .Q(I460437) );
DFFARX1 I_26950  ( .D(I240344), .CLK(I2702), .RSTB(I460475), .Q(I460879) );
nand I_26951 (I460896,I460879,I460591);
and I_26952 (I460913,I460574,I460896);
DFFARX1 I_26953  ( .D(I460913), .CLK(I2702), .RSTB(I460475), .Q(I460467) );
nor I_26954 (I460464,I460879,I460786);
and I_26955 (I460958,I460879,I460721);
or I_26956 (I460975,I460574,I460958);
DFFARX1 I_26957  ( .D(I460975), .CLK(I2702), .RSTB(I460475), .Q(I460452) );
nand I_26958 (I460461,I460879,I460803);
not I_26959 (I461053,I2709);
nand I_26960 (I461070,I44802,I44817);
and I_26961 (I461087,I461070,I44805);
DFFARX1 I_26962  ( .D(I461087), .CLK(I2702), .RSTB(I461053), .Q(I461104) );
not I_26963 (I461121,I461104);
DFFARX1 I_26964  ( .D(I461104), .CLK(I2702), .RSTB(I461053), .Q(I461021) );
nor I_26965 (I461152,I44814,I44817);
DFFARX1 I_26966  ( .D(I44799), .CLK(I2702), .RSTB(I461053), .Q(I461169) );
DFFARX1 I_26967  ( .D(I461169), .CLK(I2702), .RSTB(I461053), .Q(I461186) );
not I_26968 (I461024,I461186);
DFFARX1 I_26969  ( .D(I461169), .CLK(I2702), .RSTB(I461053), .Q(I461217) );
and I_26970 (I461018,I461104,I461217);
nand I_26971 (I461248,I44790,I44787);
and I_26972 (I461265,I461248,I44793);
DFFARX1 I_26973  ( .D(I461265), .CLK(I2702), .RSTB(I461053), .Q(I461282) );
nor I_26974 (I461299,I461282,I461121);
not I_26975 (I461316,I461282);
nand I_26976 (I461027,I461104,I461316);
DFFARX1 I_26977  ( .D(I44796), .CLK(I2702), .RSTB(I461053), .Q(I461347) );
and I_26978 (I461364,I461347,I44808);
nor I_26979 (I461381,I461364,I461282);
nor I_26980 (I461398,I461364,I461316);
nand I_26981 (I461033,I461152,I461398);
not I_26982 (I461036,I461364);
DFFARX1 I_26983  ( .D(I461364), .CLK(I2702), .RSTB(I461053), .Q(I461015) );
DFFARX1 I_26984  ( .D(I44811), .CLK(I2702), .RSTB(I461053), .Q(I461457) );
nand I_26985 (I461474,I461457,I461169);
and I_26986 (I461491,I461152,I461474);
DFFARX1 I_26987  ( .D(I461491), .CLK(I2702), .RSTB(I461053), .Q(I461045) );
nor I_26988 (I461042,I461457,I461364);
and I_26989 (I461536,I461457,I461299);
or I_26990 (I461553,I461152,I461536);
DFFARX1 I_26991  ( .D(I461553), .CLK(I2702), .RSTB(I461053), .Q(I461030) );
nand I_26992 (I461039,I461457,I461381);
not I_26993 (I461631,I2709);
nand I_26994 (I461648,I544716,I544704);
and I_26995 (I461665,I461648,I544698);
DFFARX1 I_26996  ( .D(I461665), .CLK(I2702), .RSTB(I461631), .Q(I461682) );
not I_26997 (I461699,I461682);
DFFARX1 I_26998  ( .D(I461682), .CLK(I2702), .RSTB(I461631), .Q(I461599) );
nor I_26999 (I461730,I544695,I544704);
DFFARX1 I_27000  ( .D(I544689), .CLK(I2702), .RSTB(I461631), .Q(I461747) );
DFFARX1 I_27001  ( .D(I461747), .CLK(I2702), .RSTB(I461631), .Q(I461764) );
not I_27002 (I461602,I461764);
DFFARX1 I_27003  ( .D(I461747), .CLK(I2702), .RSTB(I461631), .Q(I461795) );
and I_27004 (I461596,I461682,I461795);
nand I_27005 (I461826,I544692,I544707);
and I_27006 (I461843,I461826,I544719);
DFFARX1 I_27007  ( .D(I461843), .CLK(I2702), .RSTB(I461631), .Q(I461860) );
nor I_27008 (I461877,I461860,I461699);
not I_27009 (I461894,I461860);
nand I_27010 (I461605,I461682,I461894);
DFFARX1 I_27011  ( .D(I544710), .CLK(I2702), .RSTB(I461631), .Q(I461925) );
and I_27012 (I461942,I461925,I544701);
nor I_27013 (I461959,I461942,I461860);
nor I_27014 (I461976,I461942,I461894);
nand I_27015 (I461611,I461730,I461976);
not I_27016 (I461614,I461942);
DFFARX1 I_27017  ( .D(I461942), .CLK(I2702), .RSTB(I461631), .Q(I461593) );
DFFARX1 I_27018  ( .D(I544713), .CLK(I2702), .RSTB(I461631), .Q(I462035) );
nand I_27019 (I462052,I462035,I461747);
and I_27020 (I462069,I461730,I462052);
DFFARX1 I_27021  ( .D(I462069), .CLK(I2702), .RSTB(I461631), .Q(I461623) );
nor I_27022 (I461620,I462035,I461942);
and I_27023 (I462114,I462035,I461877);
or I_27024 (I462131,I461730,I462114);
DFFARX1 I_27025  ( .D(I462131), .CLK(I2702), .RSTB(I461631), .Q(I461608) );
nand I_27026 (I461617,I462035,I461959);
not I_27027 (I462209,I2709);
nand I_27028 (I462226,I292038,I292065);
and I_27029 (I462243,I462226,I292053);
DFFARX1 I_27030  ( .D(I462243), .CLK(I2702), .RSTB(I462209), .Q(I462260) );
not I_27031 (I462277,I462260);
DFFARX1 I_27032  ( .D(I462260), .CLK(I2702), .RSTB(I462209), .Q(I462177) );
nor I_27033 (I462308,I292041,I292065);
DFFARX1 I_27034  ( .D(I292056), .CLK(I2702), .RSTB(I462209), .Q(I462325) );
DFFARX1 I_27035  ( .D(I462325), .CLK(I2702), .RSTB(I462209), .Q(I462342) );
not I_27036 (I462180,I462342);
DFFARX1 I_27037  ( .D(I462325), .CLK(I2702), .RSTB(I462209), .Q(I462373) );
and I_27038 (I462174,I462260,I462373);
nand I_27039 (I462404,I292050,I292047);
and I_27040 (I462421,I462404,I292044);
DFFARX1 I_27041  ( .D(I462421), .CLK(I2702), .RSTB(I462209), .Q(I462438) );
nor I_27042 (I462455,I462438,I462277);
not I_27043 (I462472,I462438);
nand I_27044 (I462183,I462260,I462472);
DFFARX1 I_27045  ( .D(I292059), .CLK(I2702), .RSTB(I462209), .Q(I462503) );
and I_27046 (I462520,I462503,I292035);
nor I_27047 (I462537,I462520,I462438);
nor I_27048 (I462554,I462520,I462472);
nand I_27049 (I462189,I462308,I462554);
not I_27050 (I462192,I462520);
DFFARX1 I_27051  ( .D(I462520), .CLK(I2702), .RSTB(I462209), .Q(I462171) );
DFFARX1 I_27052  ( .D(I292062), .CLK(I2702), .RSTB(I462209), .Q(I462613) );
nand I_27053 (I462630,I462613,I462325);
and I_27054 (I462647,I462308,I462630);
DFFARX1 I_27055  ( .D(I462647), .CLK(I2702), .RSTB(I462209), .Q(I462201) );
nor I_27056 (I462198,I462613,I462520);
and I_27057 (I462692,I462613,I462455);
or I_27058 (I462709,I462308,I462692);
DFFARX1 I_27059  ( .D(I462709), .CLK(I2702), .RSTB(I462209), .Q(I462186) );
nand I_27060 (I462195,I462613,I462537);
not I_27061 (I462787,I2709);
nand I_27062 (I462804,I370624,I370621);
and I_27063 (I462821,I462804,I370633);
DFFARX1 I_27064  ( .D(I462821), .CLK(I2702), .RSTB(I462787), .Q(I462838) );
not I_27065 (I462855,I462838);
DFFARX1 I_27066  ( .D(I462838), .CLK(I2702), .RSTB(I462787), .Q(I462755) );
nor I_27067 (I462886,I370630,I370621);
DFFARX1 I_27068  ( .D(I370636), .CLK(I2702), .RSTB(I462787), .Q(I462903) );
DFFARX1 I_27069  ( .D(I462903), .CLK(I2702), .RSTB(I462787), .Q(I462920) );
not I_27070 (I462758,I462920);
DFFARX1 I_27071  ( .D(I462903), .CLK(I2702), .RSTB(I462787), .Q(I462951) );
and I_27072 (I462752,I462838,I462951);
nand I_27073 (I462982,I370612,I370615);
and I_27074 (I462999,I462982,I370639);
DFFARX1 I_27075  ( .D(I462999), .CLK(I2702), .RSTB(I462787), .Q(I463016) );
nor I_27076 (I463033,I463016,I462855);
not I_27077 (I463050,I463016);
nand I_27078 (I462761,I462838,I463050);
DFFARX1 I_27079  ( .D(I370618), .CLK(I2702), .RSTB(I462787), .Q(I463081) );
and I_27080 (I463098,I463081,I370609);
nor I_27081 (I463115,I463098,I463016);
nor I_27082 (I463132,I463098,I463050);
nand I_27083 (I462767,I462886,I463132);
not I_27084 (I462770,I463098);
DFFARX1 I_27085  ( .D(I463098), .CLK(I2702), .RSTB(I462787), .Q(I462749) );
DFFARX1 I_27086  ( .D(I370627), .CLK(I2702), .RSTB(I462787), .Q(I463191) );
nand I_27087 (I463208,I463191,I462903);
and I_27088 (I463225,I462886,I463208);
DFFARX1 I_27089  ( .D(I463225), .CLK(I2702), .RSTB(I462787), .Q(I462779) );
nor I_27090 (I462776,I463191,I463098);
and I_27091 (I463270,I463191,I463033);
or I_27092 (I463287,I462886,I463270);
DFFARX1 I_27093  ( .D(I463287), .CLK(I2702), .RSTB(I462787), .Q(I462764) );
nand I_27094 (I462773,I463191,I463115);
not I_27095 (I463365,I2709);
nand I_27096 (I463382,I118248,I118230);
and I_27097 (I463399,I463382,I118242);
DFFARX1 I_27098  ( .D(I463399), .CLK(I2702), .RSTB(I463365), .Q(I463416) );
not I_27099 (I463433,I463416);
DFFARX1 I_27100  ( .D(I463416), .CLK(I2702), .RSTB(I463365), .Q(I463333) );
nor I_27101 (I463464,I118245,I118230);
DFFARX1 I_27102  ( .D(I118254), .CLK(I2702), .RSTB(I463365), .Q(I463481) );
DFFARX1 I_27103  ( .D(I463481), .CLK(I2702), .RSTB(I463365), .Q(I463498) );
not I_27104 (I463336,I463498);
DFFARX1 I_27105  ( .D(I463481), .CLK(I2702), .RSTB(I463365), .Q(I463529) );
and I_27106 (I463330,I463416,I463529);
nand I_27107 (I463560,I118233,I118257);
and I_27108 (I463577,I463560,I118236);
DFFARX1 I_27109  ( .D(I463577), .CLK(I2702), .RSTB(I463365), .Q(I463594) );
nor I_27110 (I463611,I463594,I463433);
not I_27111 (I463628,I463594);
nand I_27112 (I463339,I463416,I463628);
DFFARX1 I_27113  ( .D(I118239), .CLK(I2702), .RSTB(I463365), .Q(I463659) );
and I_27114 (I463676,I463659,I118251);
nor I_27115 (I463693,I463676,I463594);
nor I_27116 (I463710,I463676,I463628);
nand I_27117 (I463345,I463464,I463710);
not I_27118 (I463348,I463676);
DFFARX1 I_27119  ( .D(I463676), .CLK(I2702), .RSTB(I463365), .Q(I463327) );
DFFARX1 I_27120  ( .D(I118227), .CLK(I2702), .RSTB(I463365), .Q(I463769) );
nand I_27121 (I463786,I463769,I463481);
and I_27122 (I463803,I463464,I463786);
DFFARX1 I_27123  ( .D(I463803), .CLK(I2702), .RSTB(I463365), .Q(I463357) );
nor I_27124 (I463354,I463769,I463676);
and I_27125 (I463848,I463769,I463611);
or I_27126 (I463865,I463464,I463848);
DFFARX1 I_27127  ( .D(I463865), .CLK(I2702), .RSTB(I463365), .Q(I463342) );
nand I_27128 (I463351,I463769,I463693);
not I_27129 (I463943,I2709);
nand I_27130 (I463960,I271485,I271512);
and I_27131 (I463977,I463960,I271500);
DFFARX1 I_27132  ( .D(I463977), .CLK(I2702), .RSTB(I463943), .Q(I463994) );
not I_27133 (I464011,I463994);
DFFARX1 I_27134  ( .D(I463994), .CLK(I2702), .RSTB(I463943), .Q(I463911) );
nor I_27135 (I464042,I271488,I271512);
DFFARX1 I_27136  ( .D(I271503), .CLK(I2702), .RSTB(I463943), .Q(I464059) );
DFFARX1 I_27137  ( .D(I464059), .CLK(I2702), .RSTB(I463943), .Q(I464076) );
not I_27138 (I463914,I464076);
DFFARX1 I_27139  ( .D(I464059), .CLK(I2702), .RSTB(I463943), .Q(I464107) );
and I_27140 (I463908,I463994,I464107);
nand I_27141 (I464138,I271497,I271494);
and I_27142 (I464155,I464138,I271491);
DFFARX1 I_27143  ( .D(I464155), .CLK(I2702), .RSTB(I463943), .Q(I464172) );
nor I_27144 (I464189,I464172,I464011);
not I_27145 (I464206,I464172);
nand I_27146 (I463917,I463994,I464206);
DFFARX1 I_27147  ( .D(I271506), .CLK(I2702), .RSTB(I463943), .Q(I464237) );
and I_27148 (I464254,I464237,I271482);
nor I_27149 (I464271,I464254,I464172);
nor I_27150 (I464288,I464254,I464206);
nand I_27151 (I463923,I464042,I464288);
not I_27152 (I463926,I464254);
DFFARX1 I_27153  ( .D(I464254), .CLK(I2702), .RSTB(I463943), .Q(I463905) );
DFFARX1 I_27154  ( .D(I271509), .CLK(I2702), .RSTB(I463943), .Q(I464347) );
nand I_27155 (I464364,I464347,I464059);
and I_27156 (I464381,I464042,I464364);
DFFARX1 I_27157  ( .D(I464381), .CLK(I2702), .RSTB(I463943), .Q(I463935) );
nor I_27158 (I463932,I464347,I464254);
and I_27159 (I464426,I464347,I464189);
or I_27160 (I464443,I464042,I464426);
DFFARX1 I_27161  ( .D(I464443), .CLK(I2702), .RSTB(I463943), .Q(I463920) );
nand I_27162 (I463929,I464347,I464271);
not I_27163 (I464521,I2709);
nand I_27164 (I464538,I340908,I340905);
and I_27165 (I464555,I464538,I340917);
DFFARX1 I_27166  ( .D(I464555), .CLK(I2702), .RSTB(I464521), .Q(I464572) );
not I_27167 (I464589,I464572);
DFFARX1 I_27168  ( .D(I464572), .CLK(I2702), .RSTB(I464521), .Q(I464489) );
nor I_27169 (I464620,I340914,I340905);
DFFARX1 I_27170  ( .D(I340920), .CLK(I2702), .RSTB(I464521), .Q(I464637) );
DFFARX1 I_27171  ( .D(I464637), .CLK(I2702), .RSTB(I464521), .Q(I464654) );
not I_27172 (I464492,I464654);
DFFARX1 I_27173  ( .D(I464637), .CLK(I2702), .RSTB(I464521), .Q(I464685) );
and I_27174 (I464486,I464572,I464685);
nand I_27175 (I464716,I340896,I340899);
and I_27176 (I464733,I464716,I340923);
DFFARX1 I_27177  ( .D(I464733), .CLK(I2702), .RSTB(I464521), .Q(I464750) );
nor I_27178 (I464767,I464750,I464589);
not I_27179 (I464784,I464750);
nand I_27180 (I464495,I464572,I464784);
DFFARX1 I_27181  ( .D(I340902), .CLK(I2702), .RSTB(I464521), .Q(I464815) );
and I_27182 (I464832,I464815,I340893);
nor I_27183 (I464849,I464832,I464750);
nor I_27184 (I464866,I464832,I464784);
nand I_27185 (I464501,I464620,I464866);
not I_27186 (I464504,I464832);
DFFARX1 I_27187  ( .D(I464832), .CLK(I2702), .RSTB(I464521), .Q(I464483) );
DFFARX1 I_27188  ( .D(I340911), .CLK(I2702), .RSTB(I464521), .Q(I464925) );
nand I_27189 (I464942,I464925,I464637);
and I_27190 (I464959,I464620,I464942);
DFFARX1 I_27191  ( .D(I464959), .CLK(I2702), .RSTB(I464521), .Q(I464513) );
nor I_27192 (I464510,I464925,I464832);
and I_27193 (I465004,I464925,I464767);
or I_27194 (I465021,I464620,I465004);
DFFARX1 I_27195  ( .D(I465021), .CLK(I2702), .RSTB(I464521), .Q(I464498) );
nand I_27196 (I464507,I464925,I464849);
not I_27197 (I465099,I2709);
nand I_27198 (I465116,I626902,I626905);
and I_27199 (I465133,I465116,I626911);
DFFARX1 I_27200  ( .D(I465133), .CLK(I2702), .RSTB(I465099), .Q(I465150) );
not I_27201 (I465167,I465150);
DFFARX1 I_27202  ( .D(I465150), .CLK(I2702), .RSTB(I465099), .Q(I465067) );
nor I_27203 (I465198,I626908,I626905);
DFFARX1 I_27204  ( .D(I626887), .CLK(I2702), .RSTB(I465099), .Q(I465215) );
DFFARX1 I_27205  ( .D(I465215), .CLK(I2702), .RSTB(I465099), .Q(I465232) );
not I_27206 (I465070,I465232);
DFFARX1 I_27207  ( .D(I465215), .CLK(I2702), .RSTB(I465099), .Q(I465263) );
and I_27208 (I465064,I465150,I465263);
nand I_27209 (I465294,I626884,I626899);
and I_27210 (I465311,I465294,I626896);
DFFARX1 I_27211  ( .D(I465311), .CLK(I2702), .RSTB(I465099), .Q(I465328) );
nor I_27212 (I465345,I465328,I465167);
not I_27213 (I465362,I465328);
nand I_27214 (I465073,I465150,I465362);
DFFARX1 I_27215  ( .D(I626914), .CLK(I2702), .RSTB(I465099), .Q(I465393) );
and I_27216 (I465410,I465393,I626893);
nor I_27217 (I465427,I465410,I465328);
nor I_27218 (I465444,I465410,I465362);
nand I_27219 (I465079,I465198,I465444);
not I_27220 (I465082,I465410);
DFFARX1 I_27221  ( .D(I465410), .CLK(I2702), .RSTB(I465099), .Q(I465061) );
DFFARX1 I_27222  ( .D(I626890), .CLK(I2702), .RSTB(I465099), .Q(I465503) );
nand I_27223 (I465520,I465503,I465215);
and I_27224 (I465537,I465198,I465520);
DFFARX1 I_27225  ( .D(I465537), .CLK(I2702), .RSTB(I465099), .Q(I465091) );
nor I_27226 (I465088,I465503,I465410);
and I_27227 (I465582,I465503,I465345);
or I_27228 (I465599,I465198,I465582);
DFFARX1 I_27229  ( .D(I465599), .CLK(I2702), .RSTB(I465099), .Q(I465076) );
nand I_27230 (I465085,I465503,I465427);
not I_27231 (I465677,I2709);
nand I_27232 (I465694,I51064,I51046);
and I_27233 (I465711,I465694,I51058);
DFFARX1 I_27234  ( .D(I465711), .CLK(I2702), .RSTB(I465677), .Q(I465728) );
not I_27235 (I465745,I465728);
DFFARX1 I_27236  ( .D(I465728), .CLK(I2702), .RSTB(I465677), .Q(I465645) );
nor I_27237 (I465776,I51061,I51046);
DFFARX1 I_27238  ( .D(I51070), .CLK(I2702), .RSTB(I465677), .Q(I465793) );
DFFARX1 I_27239  ( .D(I465793), .CLK(I2702), .RSTB(I465677), .Q(I465810) );
not I_27240 (I465648,I465810);
DFFARX1 I_27241  ( .D(I465793), .CLK(I2702), .RSTB(I465677), .Q(I465841) );
and I_27242 (I465642,I465728,I465841);
nand I_27243 (I465872,I51049,I51073);
and I_27244 (I465889,I465872,I51052);
DFFARX1 I_27245  ( .D(I465889), .CLK(I2702), .RSTB(I465677), .Q(I465906) );
nor I_27246 (I465923,I465906,I465745);
not I_27247 (I465940,I465906);
nand I_27248 (I465651,I465728,I465940);
DFFARX1 I_27249  ( .D(I51055), .CLK(I2702), .RSTB(I465677), .Q(I465971) );
and I_27250 (I465988,I465971,I51067);
nor I_27251 (I466005,I465988,I465906);
nor I_27252 (I466022,I465988,I465940);
nand I_27253 (I465657,I465776,I466022);
not I_27254 (I465660,I465988);
DFFARX1 I_27255  ( .D(I465988), .CLK(I2702), .RSTB(I465677), .Q(I465639) );
DFFARX1 I_27256  ( .D(I51043), .CLK(I2702), .RSTB(I465677), .Q(I466081) );
nand I_27257 (I466098,I466081,I465793);
and I_27258 (I466115,I465776,I466098);
DFFARX1 I_27259  ( .D(I466115), .CLK(I2702), .RSTB(I465677), .Q(I465669) );
nor I_27260 (I465666,I466081,I465988);
and I_27261 (I466160,I466081,I465923);
or I_27262 (I466177,I465776,I466160);
DFFARX1 I_27263  ( .D(I466177), .CLK(I2702), .RSTB(I465677), .Q(I465654) );
nand I_27264 (I465663,I466081,I466005);
not I_27265 (I466255,I2709);
nand I_27266 (I466272,I393234,I393231);
and I_27267 (I466289,I466272,I393243);
DFFARX1 I_27268  ( .D(I466289), .CLK(I2702), .RSTB(I466255), .Q(I466306) );
not I_27269 (I466323,I466306);
DFFARX1 I_27270  ( .D(I466306), .CLK(I2702), .RSTB(I466255), .Q(I466223) );
nor I_27271 (I466354,I393240,I393231);
DFFARX1 I_27272  ( .D(I393246), .CLK(I2702), .RSTB(I466255), .Q(I466371) );
DFFARX1 I_27273  ( .D(I466371), .CLK(I2702), .RSTB(I466255), .Q(I466388) );
not I_27274 (I466226,I466388);
DFFARX1 I_27275  ( .D(I466371), .CLK(I2702), .RSTB(I466255), .Q(I466419) );
and I_27276 (I466220,I466306,I466419);
nand I_27277 (I466450,I393222,I393225);
and I_27278 (I466467,I466450,I393249);
DFFARX1 I_27279  ( .D(I466467), .CLK(I2702), .RSTB(I466255), .Q(I466484) );
nor I_27280 (I466501,I466484,I466323);
not I_27281 (I466518,I466484);
nand I_27282 (I466229,I466306,I466518);
DFFARX1 I_27283  ( .D(I393228), .CLK(I2702), .RSTB(I466255), .Q(I466549) );
and I_27284 (I466566,I466549,I393219);
nor I_27285 (I466583,I466566,I466484);
nor I_27286 (I466600,I466566,I466518);
nand I_27287 (I466235,I466354,I466600);
not I_27288 (I466238,I466566);
DFFARX1 I_27289  ( .D(I466566), .CLK(I2702), .RSTB(I466255), .Q(I466217) );
DFFARX1 I_27290  ( .D(I393237), .CLK(I2702), .RSTB(I466255), .Q(I466659) );
nand I_27291 (I466676,I466659,I466371);
and I_27292 (I466693,I466354,I466676);
DFFARX1 I_27293  ( .D(I466693), .CLK(I2702), .RSTB(I466255), .Q(I466247) );
nor I_27294 (I466244,I466659,I466566);
and I_27295 (I466738,I466659,I466501);
or I_27296 (I466755,I466354,I466738);
DFFARX1 I_27297  ( .D(I466755), .CLK(I2702), .RSTB(I466255), .Q(I466232) );
nand I_27298 (I466241,I466659,I466583);
not I_27299 (I466833,I2709);
nand I_27300 (I466850,I534006,I533994);
and I_27301 (I466867,I466850,I533988);
DFFARX1 I_27302  ( .D(I466867), .CLK(I2702), .RSTB(I466833), .Q(I466884) );
not I_27303 (I466901,I466884);
DFFARX1 I_27304  ( .D(I466884), .CLK(I2702), .RSTB(I466833), .Q(I466801) );
nor I_27305 (I466932,I533985,I533994);
DFFARX1 I_27306  ( .D(I533979), .CLK(I2702), .RSTB(I466833), .Q(I466949) );
DFFARX1 I_27307  ( .D(I466949), .CLK(I2702), .RSTB(I466833), .Q(I466966) );
not I_27308 (I466804,I466966);
DFFARX1 I_27309  ( .D(I466949), .CLK(I2702), .RSTB(I466833), .Q(I466997) );
and I_27310 (I466798,I466884,I466997);
nand I_27311 (I467028,I533982,I533997);
and I_27312 (I467045,I467028,I534009);
DFFARX1 I_27313  ( .D(I467045), .CLK(I2702), .RSTB(I466833), .Q(I467062) );
nor I_27314 (I467079,I467062,I466901);
not I_27315 (I467096,I467062);
nand I_27316 (I466807,I466884,I467096);
DFFARX1 I_27317  ( .D(I534000), .CLK(I2702), .RSTB(I466833), .Q(I467127) );
and I_27318 (I467144,I467127,I533991);
nor I_27319 (I467161,I467144,I467062);
nor I_27320 (I467178,I467144,I467096);
nand I_27321 (I466813,I466932,I467178);
not I_27322 (I466816,I467144);
DFFARX1 I_27323  ( .D(I467144), .CLK(I2702), .RSTB(I466833), .Q(I466795) );
DFFARX1 I_27324  ( .D(I534003), .CLK(I2702), .RSTB(I466833), .Q(I467237) );
nand I_27325 (I467254,I467237,I466949);
and I_27326 (I467271,I466932,I467254);
DFFARX1 I_27327  ( .D(I467271), .CLK(I2702), .RSTB(I466833), .Q(I466825) );
nor I_27328 (I466822,I467237,I467144);
and I_27329 (I467316,I467237,I467079);
or I_27330 (I467333,I466932,I467316);
DFFARX1 I_27331  ( .D(I467333), .CLK(I2702), .RSTB(I466833), .Q(I466810) );
nand I_27332 (I466819,I467237,I467161);
not I_27333 (I467411,I2709);
nand I_27334 (I467428,I343492,I343489);
and I_27335 (I467445,I467428,I343501);
DFFARX1 I_27336  ( .D(I467445), .CLK(I2702), .RSTB(I467411), .Q(I467462) );
not I_27337 (I467479,I467462);
DFFARX1 I_27338  ( .D(I467462), .CLK(I2702), .RSTB(I467411), .Q(I467379) );
nor I_27339 (I467510,I343498,I343489);
DFFARX1 I_27340  ( .D(I343504), .CLK(I2702), .RSTB(I467411), .Q(I467527) );
DFFARX1 I_27341  ( .D(I467527), .CLK(I2702), .RSTB(I467411), .Q(I467544) );
not I_27342 (I467382,I467544);
DFFARX1 I_27343  ( .D(I467527), .CLK(I2702), .RSTB(I467411), .Q(I467575) );
and I_27344 (I467376,I467462,I467575);
nand I_27345 (I467606,I343480,I343483);
and I_27346 (I467623,I467606,I343507);
DFFARX1 I_27347  ( .D(I467623), .CLK(I2702), .RSTB(I467411), .Q(I467640) );
nor I_27348 (I467657,I467640,I467479);
not I_27349 (I467674,I467640);
nand I_27350 (I467385,I467462,I467674);
DFFARX1 I_27351  ( .D(I343486), .CLK(I2702), .RSTB(I467411), .Q(I467705) );
and I_27352 (I467722,I467705,I343477);
nor I_27353 (I467739,I467722,I467640);
nor I_27354 (I467756,I467722,I467674);
nand I_27355 (I467391,I467510,I467756);
not I_27356 (I467394,I467722);
DFFARX1 I_27357  ( .D(I467722), .CLK(I2702), .RSTB(I467411), .Q(I467373) );
DFFARX1 I_27358  ( .D(I343495), .CLK(I2702), .RSTB(I467411), .Q(I467815) );
nand I_27359 (I467832,I467815,I467527);
and I_27360 (I467849,I467510,I467832);
DFFARX1 I_27361  ( .D(I467849), .CLK(I2702), .RSTB(I467411), .Q(I467403) );
nor I_27362 (I467400,I467815,I467722);
and I_27363 (I467894,I467815,I467657);
or I_27364 (I467911,I467510,I467894);
DFFARX1 I_27365  ( .D(I467911), .CLK(I2702), .RSTB(I467411), .Q(I467388) );
nand I_27366 (I467397,I467815,I467739);
not I_27367 (I467989,I2709);
nand I_27368 (I468006,I492539,I492563);
and I_27369 (I468023,I468006,I492545);
DFFARX1 I_27370  ( .D(I468023), .CLK(I2702), .RSTB(I467989), .Q(I468040) );
not I_27371 (I468057,I468040);
DFFARX1 I_27372  ( .D(I468040), .CLK(I2702), .RSTB(I467989), .Q(I467957) );
nor I_27373 (I468088,I492533,I492563);
DFFARX1 I_27374  ( .D(I492548), .CLK(I2702), .RSTB(I467989), .Q(I468105) );
DFFARX1 I_27375  ( .D(I468105), .CLK(I2702), .RSTB(I467989), .Q(I468122) );
not I_27376 (I467960,I468122);
DFFARX1 I_27377  ( .D(I468105), .CLK(I2702), .RSTB(I467989), .Q(I468153) );
and I_27378 (I467954,I468040,I468153);
nand I_27379 (I468184,I492554,I492536);
and I_27380 (I468201,I468184,I492557);
DFFARX1 I_27381  ( .D(I468201), .CLK(I2702), .RSTB(I467989), .Q(I468218) );
nor I_27382 (I468235,I468218,I468057);
not I_27383 (I468252,I468218);
nand I_27384 (I467963,I468040,I468252);
DFFARX1 I_27385  ( .D(I492542), .CLK(I2702), .RSTB(I467989), .Q(I468283) );
and I_27386 (I468300,I468283,I492551);
nor I_27387 (I468317,I468300,I468218);
nor I_27388 (I468334,I468300,I468252);
nand I_27389 (I467969,I468088,I468334);
not I_27390 (I467972,I468300);
DFFARX1 I_27391  ( .D(I468300), .CLK(I2702), .RSTB(I467989), .Q(I467951) );
DFFARX1 I_27392  ( .D(I492560), .CLK(I2702), .RSTB(I467989), .Q(I468393) );
nand I_27393 (I468410,I468393,I468105);
and I_27394 (I468427,I468088,I468410);
DFFARX1 I_27395  ( .D(I468427), .CLK(I2702), .RSTB(I467989), .Q(I467981) );
nor I_27396 (I467978,I468393,I468300);
and I_27397 (I468472,I468393,I468235);
or I_27398 (I468489,I468088,I468472);
DFFARX1 I_27399  ( .D(I468489), .CLK(I2702), .RSTB(I467989), .Q(I467966) );
nand I_27400 (I467975,I468393,I468317);
not I_27401 (I468567,I2709);
nand I_27402 (I468584,I196590,I196569);
and I_27403 (I468601,I468584,I196566);
DFFARX1 I_27404  ( .D(I468601), .CLK(I2702), .RSTB(I468567), .Q(I468618) );
not I_27405 (I468635,I468618);
DFFARX1 I_27406  ( .D(I468618), .CLK(I2702), .RSTB(I468567), .Q(I468535) );
nor I_27407 (I468666,I196575,I196569);
DFFARX1 I_27408  ( .D(I196563), .CLK(I2702), .RSTB(I468567), .Q(I468683) );
DFFARX1 I_27409  ( .D(I468683), .CLK(I2702), .RSTB(I468567), .Q(I468700) );
not I_27410 (I468538,I468700);
DFFARX1 I_27411  ( .D(I468683), .CLK(I2702), .RSTB(I468567), .Q(I468731) );
and I_27412 (I468532,I468618,I468731);
nand I_27413 (I468762,I196593,I196584);
and I_27414 (I468779,I468762,I196581);
DFFARX1 I_27415  ( .D(I468779), .CLK(I2702), .RSTB(I468567), .Q(I468796) );
nor I_27416 (I468813,I468796,I468635);
not I_27417 (I468830,I468796);
nand I_27418 (I468541,I468618,I468830);
DFFARX1 I_27419  ( .D(I196578), .CLK(I2702), .RSTB(I468567), .Q(I468861) );
and I_27420 (I468878,I468861,I196587);
nor I_27421 (I468895,I468878,I468796);
nor I_27422 (I468912,I468878,I468830);
nand I_27423 (I468547,I468666,I468912);
not I_27424 (I468550,I468878);
DFFARX1 I_27425  ( .D(I468878), .CLK(I2702), .RSTB(I468567), .Q(I468529) );
DFFARX1 I_27426  ( .D(I196572), .CLK(I2702), .RSTB(I468567), .Q(I468971) );
nand I_27427 (I468988,I468971,I468683);
and I_27428 (I469005,I468666,I468988);
DFFARX1 I_27429  ( .D(I469005), .CLK(I2702), .RSTB(I468567), .Q(I468559) );
nor I_27430 (I468556,I468971,I468878);
and I_27431 (I469050,I468971,I468813);
or I_27432 (I469067,I468666,I469050);
DFFARX1 I_27433  ( .D(I469067), .CLK(I2702), .RSTB(I468567), .Q(I468544) );
nand I_27434 (I468553,I468971,I468895);
not I_27435 (I469145,I2709);
nand I_27436 (I469162,I55586,I55568);
and I_27437 (I469179,I469162,I55580);
DFFARX1 I_27438  ( .D(I469179), .CLK(I2702), .RSTB(I469145), .Q(I469196) );
not I_27439 (I469213,I469196);
DFFARX1 I_27440  ( .D(I469196), .CLK(I2702), .RSTB(I469145), .Q(I469113) );
nor I_27441 (I469244,I55583,I55568);
DFFARX1 I_27442  ( .D(I55592), .CLK(I2702), .RSTB(I469145), .Q(I469261) );
DFFARX1 I_27443  ( .D(I469261), .CLK(I2702), .RSTB(I469145), .Q(I469278) );
not I_27444 (I469116,I469278);
DFFARX1 I_27445  ( .D(I469261), .CLK(I2702), .RSTB(I469145), .Q(I469309) );
and I_27446 (I469110,I469196,I469309);
nand I_27447 (I469340,I55571,I55595);
and I_27448 (I469357,I469340,I55574);
DFFARX1 I_27449  ( .D(I469357), .CLK(I2702), .RSTB(I469145), .Q(I469374) );
nor I_27450 (I469391,I469374,I469213);
not I_27451 (I469408,I469374);
nand I_27452 (I469119,I469196,I469408);
DFFARX1 I_27453  ( .D(I55577), .CLK(I2702), .RSTB(I469145), .Q(I469439) );
and I_27454 (I469456,I469439,I55589);
nor I_27455 (I469473,I469456,I469374);
nor I_27456 (I469490,I469456,I469408);
nand I_27457 (I469125,I469244,I469490);
not I_27458 (I469128,I469456);
DFFARX1 I_27459  ( .D(I469456), .CLK(I2702), .RSTB(I469145), .Q(I469107) );
DFFARX1 I_27460  ( .D(I55565), .CLK(I2702), .RSTB(I469145), .Q(I469549) );
nand I_27461 (I469566,I469549,I469261);
and I_27462 (I469583,I469244,I469566);
DFFARX1 I_27463  ( .D(I469583), .CLK(I2702), .RSTB(I469145), .Q(I469137) );
nor I_27464 (I469134,I469549,I469456);
and I_27465 (I469628,I469549,I469391);
or I_27466 (I469645,I469244,I469628);
DFFARX1 I_27467  ( .D(I469645), .CLK(I2702), .RSTB(I469145), .Q(I469122) );
nand I_27468 (I469131,I469549,I469473);
not I_27469 (I469723,I2709);
nand I_27470 (I469740,I142887,I142866);
and I_27471 (I469757,I469740,I142863);
DFFARX1 I_27472  ( .D(I469757), .CLK(I2702), .RSTB(I469723), .Q(I469774) );
not I_27473 (I469791,I469774);
DFFARX1 I_27474  ( .D(I469774), .CLK(I2702), .RSTB(I469723), .Q(I469691) );
nor I_27475 (I469822,I142872,I142866);
DFFARX1 I_27476  ( .D(I142860), .CLK(I2702), .RSTB(I469723), .Q(I469839) );
DFFARX1 I_27477  ( .D(I469839), .CLK(I2702), .RSTB(I469723), .Q(I469856) );
not I_27478 (I469694,I469856);
DFFARX1 I_27479  ( .D(I469839), .CLK(I2702), .RSTB(I469723), .Q(I469887) );
and I_27480 (I469688,I469774,I469887);
nand I_27481 (I469918,I142890,I142881);
and I_27482 (I469935,I469918,I142878);
DFFARX1 I_27483  ( .D(I469935), .CLK(I2702), .RSTB(I469723), .Q(I469952) );
nor I_27484 (I469969,I469952,I469791);
not I_27485 (I469986,I469952);
nand I_27486 (I469697,I469774,I469986);
DFFARX1 I_27487  ( .D(I142875), .CLK(I2702), .RSTB(I469723), .Q(I470017) );
and I_27488 (I470034,I470017,I142884);
nor I_27489 (I470051,I470034,I469952);
nor I_27490 (I470068,I470034,I469986);
nand I_27491 (I469703,I469822,I470068);
not I_27492 (I469706,I470034);
DFFARX1 I_27493  ( .D(I470034), .CLK(I2702), .RSTB(I469723), .Q(I469685) );
DFFARX1 I_27494  ( .D(I142869), .CLK(I2702), .RSTB(I469723), .Q(I470127) );
nand I_27495 (I470144,I470127,I469839);
and I_27496 (I470161,I469822,I470144);
DFFARX1 I_27497  ( .D(I470161), .CLK(I2702), .RSTB(I469723), .Q(I469715) );
nor I_27498 (I469712,I470127,I470034);
and I_27499 (I470206,I470127,I469969);
or I_27500 (I470223,I469822,I470206);
DFFARX1 I_27501  ( .D(I470223), .CLK(I2702), .RSTB(I469723), .Q(I469700) );
nand I_27502 (I469709,I470127,I470051);
not I_27503 (I470301,I2709);
nand I_27504 (I470318,I96930,I96912);
and I_27505 (I470335,I470318,I96924);
DFFARX1 I_27506  ( .D(I470335), .CLK(I2702), .RSTB(I470301), .Q(I470352) );
not I_27507 (I470369,I470352);
DFFARX1 I_27508  ( .D(I470352), .CLK(I2702), .RSTB(I470301), .Q(I470269) );
nor I_27509 (I470400,I96927,I96912);
DFFARX1 I_27510  ( .D(I96936), .CLK(I2702), .RSTB(I470301), .Q(I470417) );
DFFARX1 I_27511  ( .D(I470417), .CLK(I2702), .RSTB(I470301), .Q(I470434) );
not I_27512 (I470272,I470434);
DFFARX1 I_27513  ( .D(I470417), .CLK(I2702), .RSTB(I470301), .Q(I470465) );
and I_27514 (I470266,I470352,I470465);
nand I_27515 (I470496,I96915,I96939);
and I_27516 (I470513,I470496,I96918);
DFFARX1 I_27517  ( .D(I470513), .CLK(I2702), .RSTB(I470301), .Q(I470530) );
nor I_27518 (I470547,I470530,I470369);
not I_27519 (I470564,I470530);
nand I_27520 (I470275,I470352,I470564);
DFFARX1 I_27521  ( .D(I96921), .CLK(I2702), .RSTB(I470301), .Q(I470595) );
and I_27522 (I470612,I470595,I96933);
nor I_27523 (I470629,I470612,I470530);
nor I_27524 (I470646,I470612,I470564);
nand I_27525 (I470281,I470400,I470646);
not I_27526 (I470284,I470612);
DFFARX1 I_27527  ( .D(I470612), .CLK(I2702), .RSTB(I470301), .Q(I470263) );
DFFARX1 I_27528  ( .D(I96909), .CLK(I2702), .RSTB(I470301), .Q(I470705) );
nand I_27529 (I470722,I470705,I470417);
and I_27530 (I470739,I470400,I470722);
DFFARX1 I_27531  ( .D(I470739), .CLK(I2702), .RSTB(I470301), .Q(I470293) );
nor I_27532 (I470290,I470705,I470612);
and I_27533 (I470784,I470705,I470547);
or I_27534 (I470801,I470400,I470784);
DFFARX1 I_27535  ( .D(I470801), .CLK(I2702), .RSTB(I470301), .Q(I470278) );
nand I_27536 (I470287,I470705,I470629);
not I_27537 (I470879,I2709);
nand I_27538 (I470896,I568516,I568504);
and I_27539 (I470913,I470896,I568498);
DFFARX1 I_27540  ( .D(I470913), .CLK(I2702), .RSTB(I470879), .Q(I470930) );
not I_27541 (I470947,I470930);
DFFARX1 I_27542  ( .D(I470930), .CLK(I2702), .RSTB(I470879), .Q(I470847) );
nor I_27543 (I470978,I568495,I568504);
DFFARX1 I_27544  ( .D(I568489), .CLK(I2702), .RSTB(I470879), .Q(I470995) );
DFFARX1 I_27545  ( .D(I470995), .CLK(I2702), .RSTB(I470879), .Q(I471012) );
not I_27546 (I470850,I471012);
DFFARX1 I_27547  ( .D(I470995), .CLK(I2702), .RSTB(I470879), .Q(I471043) );
and I_27548 (I470844,I470930,I471043);
nand I_27549 (I471074,I568492,I568507);
and I_27550 (I471091,I471074,I568519);
DFFARX1 I_27551  ( .D(I471091), .CLK(I2702), .RSTB(I470879), .Q(I471108) );
nor I_27552 (I471125,I471108,I470947);
not I_27553 (I471142,I471108);
nand I_27554 (I470853,I470930,I471142);
DFFARX1 I_27555  ( .D(I568510), .CLK(I2702), .RSTB(I470879), .Q(I471173) );
and I_27556 (I471190,I471173,I568501);
nor I_27557 (I471207,I471190,I471108);
nor I_27558 (I471224,I471190,I471142);
nand I_27559 (I470859,I470978,I471224);
not I_27560 (I470862,I471190);
DFFARX1 I_27561  ( .D(I471190), .CLK(I2702), .RSTB(I470879), .Q(I470841) );
DFFARX1 I_27562  ( .D(I568513), .CLK(I2702), .RSTB(I470879), .Q(I471283) );
nand I_27563 (I471300,I471283,I470995);
and I_27564 (I471317,I470978,I471300);
DFFARX1 I_27565  ( .D(I471317), .CLK(I2702), .RSTB(I470879), .Q(I470871) );
nor I_27566 (I470868,I471283,I471190);
and I_27567 (I471362,I471283,I471125);
or I_27568 (I471379,I470978,I471362);
DFFARX1 I_27569  ( .D(I471379), .CLK(I2702), .RSTB(I470879), .Q(I470856) );
nand I_27570 (I470865,I471283,I471207);
not I_27571 (I471457,I2709);
nand I_27572 (I471474,I47607,I47622);
and I_27573 (I471491,I471474,I47610);
DFFARX1 I_27574  ( .D(I471491), .CLK(I2702), .RSTB(I471457), .Q(I471508) );
not I_27575 (I471525,I471508);
DFFARX1 I_27576  ( .D(I471508), .CLK(I2702), .RSTB(I471457), .Q(I471425) );
nor I_27577 (I471556,I47619,I47622);
DFFARX1 I_27578  ( .D(I47604), .CLK(I2702), .RSTB(I471457), .Q(I471573) );
DFFARX1 I_27579  ( .D(I471573), .CLK(I2702), .RSTB(I471457), .Q(I471590) );
not I_27580 (I471428,I471590);
DFFARX1 I_27581  ( .D(I471573), .CLK(I2702), .RSTB(I471457), .Q(I471621) );
and I_27582 (I471422,I471508,I471621);
nand I_27583 (I471652,I47595,I47592);
and I_27584 (I471669,I471652,I47598);
DFFARX1 I_27585  ( .D(I471669), .CLK(I2702), .RSTB(I471457), .Q(I471686) );
nor I_27586 (I471703,I471686,I471525);
not I_27587 (I471720,I471686);
nand I_27588 (I471431,I471508,I471720);
DFFARX1 I_27589  ( .D(I47601), .CLK(I2702), .RSTB(I471457), .Q(I471751) );
and I_27590 (I471768,I471751,I47613);
nor I_27591 (I471785,I471768,I471686);
nor I_27592 (I471802,I471768,I471720);
nand I_27593 (I471437,I471556,I471802);
not I_27594 (I471440,I471768);
DFFARX1 I_27595  ( .D(I471768), .CLK(I2702), .RSTB(I471457), .Q(I471419) );
DFFARX1 I_27596  ( .D(I47616), .CLK(I2702), .RSTB(I471457), .Q(I471861) );
nand I_27597 (I471878,I471861,I471573);
and I_27598 (I471895,I471556,I471878);
DFFARX1 I_27599  ( .D(I471895), .CLK(I2702), .RSTB(I471457), .Q(I471449) );
nor I_27600 (I471446,I471861,I471768);
and I_27601 (I471940,I471861,I471703);
or I_27602 (I471957,I471556,I471940);
DFFARX1 I_27603  ( .D(I471957), .CLK(I2702), .RSTB(I471457), .Q(I471434) );
nand I_27604 (I471443,I471861,I471785);
not I_27605 (I472035,I2709);
nand I_27606 (I472052,I346076,I346073);
and I_27607 (I472069,I472052,I346085);
DFFARX1 I_27608  ( .D(I472069), .CLK(I2702), .RSTB(I472035), .Q(I472086) );
not I_27609 (I472103,I472086);
DFFARX1 I_27610  ( .D(I472086), .CLK(I2702), .RSTB(I472035), .Q(I472003) );
nor I_27611 (I472134,I346082,I346073);
DFFARX1 I_27612  ( .D(I346088), .CLK(I2702), .RSTB(I472035), .Q(I472151) );
DFFARX1 I_27613  ( .D(I472151), .CLK(I2702), .RSTB(I472035), .Q(I472168) );
not I_27614 (I472006,I472168);
DFFARX1 I_27615  ( .D(I472151), .CLK(I2702), .RSTB(I472035), .Q(I472199) );
and I_27616 (I472000,I472086,I472199);
nand I_27617 (I472230,I346064,I346067);
and I_27618 (I472247,I472230,I346091);
DFFARX1 I_27619  ( .D(I472247), .CLK(I2702), .RSTB(I472035), .Q(I472264) );
nor I_27620 (I472281,I472264,I472103);
not I_27621 (I472298,I472264);
nand I_27622 (I472009,I472086,I472298);
DFFARX1 I_27623  ( .D(I346070), .CLK(I2702), .RSTB(I472035), .Q(I472329) );
and I_27624 (I472346,I472329,I346061);
nor I_27625 (I472363,I472346,I472264);
nor I_27626 (I472380,I472346,I472298);
nand I_27627 (I472015,I472134,I472380);
not I_27628 (I472018,I472346);
DFFARX1 I_27629  ( .D(I472346), .CLK(I2702), .RSTB(I472035), .Q(I471997) );
DFFARX1 I_27630  ( .D(I346079), .CLK(I2702), .RSTB(I472035), .Q(I472439) );
nand I_27631 (I472456,I472439,I472151);
and I_27632 (I472473,I472134,I472456);
DFFARX1 I_27633  ( .D(I472473), .CLK(I2702), .RSTB(I472035), .Q(I472027) );
nor I_27634 (I472024,I472439,I472346);
and I_27635 (I472518,I472439,I472281);
or I_27636 (I472535,I472134,I472518);
DFFARX1 I_27637  ( .D(I472535), .CLK(I2702), .RSTB(I472035), .Q(I472012) );
nand I_27638 (I472021,I472439,I472363);
not I_27639 (I472613,I2709);
nand I_27640 (I472630,I677222,I677225);
and I_27641 (I472647,I472630,I677231);
DFFARX1 I_27642  ( .D(I472647), .CLK(I2702), .RSTB(I472613), .Q(I472664) );
not I_27643 (I472681,I472664);
DFFARX1 I_27644  ( .D(I472664), .CLK(I2702), .RSTB(I472613), .Q(I472581) );
nor I_27645 (I472712,I677228,I677225);
DFFARX1 I_27646  ( .D(I677207), .CLK(I2702), .RSTB(I472613), .Q(I472729) );
DFFARX1 I_27647  ( .D(I472729), .CLK(I2702), .RSTB(I472613), .Q(I472746) );
not I_27648 (I472584,I472746);
DFFARX1 I_27649  ( .D(I472729), .CLK(I2702), .RSTB(I472613), .Q(I472777) );
and I_27650 (I472578,I472664,I472777);
nand I_27651 (I472808,I677204,I677219);
and I_27652 (I472825,I472808,I677216);
DFFARX1 I_27653  ( .D(I472825), .CLK(I2702), .RSTB(I472613), .Q(I472842) );
nor I_27654 (I472859,I472842,I472681);
not I_27655 (I472876,I472842);
nand I_27656 (I472587,I472664,I472876);
DFFARX1 I_27657  ( .D(I677234), .CLK(I2702), .RSTB(I472613), .Q(I472907) );
and I_27658 (I472924,I472907,I677213);
nor I_27659 (I472941,I472924,I472842);
nor I_27660 (I472958,I472924,I472876);
nand I_27661 (I472593,I472712,I472958);
not I_27662 (I472596,I472924);
DFFARX1 I_27663  ( .D(I472924), .CLK(I2702), .RSTB(I472613), .Q(I472575) );
DFFARX1 I_27664  ( .D(I677210), .CLK(I2702), .RSTB(I472613), .Q(I473017) );
nand I_27665 (I473034,I473017,I472729);
and I_27666 (I473051,I472712,I473034);
DFFARX1 I_27667  ( .D(I473051), .CLK(I2702), .RSTB(I472613), .Q(I472605) );
nor I_27668 (I472602,I473017,I472924);
and I_27669 (I473096,I473017,I472859);
or I_27670 (I473113,I472712,I473096);
DFFARX1 I_27671  ( .D(I473113), .CLK(I2702), .RSTB(I472613), .Q(I472590) );
nand I_27672 (I472599,I473017,I472941);
not I_27673 (I473191,I2709);
nand I_27674 (I473208,I202877,I202862);
and I_27675 (I473225,I473208,I202871);
DFFARX1 I_27676  ( .D(I473225), .CLK(I2702), .RSTB(I473191), .Q(I473242) );
not I_27677 (I473259,I473242);
DFFARX1 I_27678  ( .D(I473242), .CLK(I2702), .RSTB(I473191), .Q(I473159) );
nor I_27679 (I473290,I202880,I202862);
DFFARX1 I_27680  ( .D(I202859), .CLK(I2702), .RSTB(I473191), .Q(I473307) );
DFFARX1 I_27681  ( .D(I473307), .CLK(I2702), .RSTB(I473191), .Q(I473324) );
not I_27682 (I473162,I473324);
DFFARX1 I_27683  ( .D(I473307), .CLK(I2702), .RSTB(I473191), .Q(I473355) );
and I_27684 (I473156,I473242,I473355);
nand I_27685 (I473386,I202883,I202856);
and I_27686 (I473403,I473386,I202874);
DFFARX1 I_27687  ( .D(I473403), .CLK(I2702), .RSTB(I473191), .Q(I473420) );
nor I_27688 (I473437,I473420,I473259);
not I_27689 (I473454,I473420);
nand I_27690 (I473165,I473242,I473454);
DFFARX1 I_27691  ( .D(I202868), .CLK(I2702), .RSTB(I473191), .Q(I473485) );
and I_27692 (I473502,I473485,I202853);
nor I_27693 (I473519,I473502,I473420);
nor I_27694 (I473536,I473502,I473454);
nand I_27695 (I473171,I473290,I473536);
not I_27696 (I473174,I473502);
DFFARX1 I_27697  ( .D(I473502), .CLK(I2702), .RSTB(I473191), .Q(I473153) );
DFFARX1 I_27698  ( .D(I202865), .CLK(I2702), .RSTB(I473191), .Q(I473595) );
nand I_27699 (I473612,I473595,I473307);
and I_27700 (I473629,I473290,I473612);
DFFARX1 I_27701  ( .D(I473629), .CLK(I2702), .RSTB(I473191), .Q(I473183) );
nor I_27702 (I473180,I473595,I473502);
and I_27703 (I473674,I473595,I473437);
or I_27704 (I473691,I473290,I473674);
DFFARX1 I_27705  ( .D(I473691), .CLK(I2702), .RSTB(I473191), .Q(I473168) );
nand I_27706 (I473177,I473595,I473519);
not I_27707 (I473769,I2709);
nand I_27708 (I473786,I551261,I551249);
and I_27709 (I473803,I473786,I551243);
DFFARX1 I_27710  ( .D(I473803), .CLK(I2702), .RSTB(I473769), .Q(I473820) );
not I_27711 (I473837,I473820);
DFFARX1 I_27712  ( .D(I473820), .CLK(I2702), .RSTB(I473769), .Q(I473737) );
nor I_27713 (I473868,I551240,I551249);
DFFARX1 I_27714  ( .D(I551234), .CLK(I2702), .RSTB(I473769), .Q(I473885) );
DFFARX1 I_27715  ( .D(I473885), .CLK(I2702), .RSTB(I473769), .Q(I473902) );
not I_27716 (I473740,I473902);
DFFARX1 I_27717  ( .D(I473885), .CLK(I2702), .RSTB(I473769), .Q(I473933) );
and I_27718 (I473734,I473820,I473933);
nand I_27719 (I473964,I551237,I551252);
and I_27720 (I473981,I473964,I551264);
DFFARX1 I_27721  ( .D(I473981), .CLK(I2702), .RSTB(I473769), .Q(I473998) );
nor I_27722 (I474015,I473998,I473837);
not I_27723 (I474032,I473998);
nand I_27724 (I473743,I473820,I474032);
DFFARX1 I_27725  ( .D(I551255), .CLK(I2702), .RSTB(I473769), .Q(I474063) );
and I_27726 (I474080,I474063,I551246);
nor I_27727 (I474097,I474080,I473998);
nor I_27728 (I474114,I474080,I474032);
nand I_27729 (I473749,I473868,I474114);
not I_27730 (I473752,I474080);
DFFARX1 I_27731  ( .D(I474080), .CLK(I2702), .RSTB(I473769), .Q(I473731) );
DFFARX1 I_27732  ( .D(I551258), .CLK(I2702), .RSTB(I473769), .Q(I474173) );
nand I_27733 (I474190,I474173,I473885);
and I_27734 (I474207,I473868,I474190);
DFFARX1 I_27735  ( .D(I474207), .CLK(I2702), .RSTB(I473769), .Q(I473761) );
nor I_27736 (I473758,I474173,I474080);
and I_27737 (I474252,I474173,I474015);
or I_27738 (I474269,I473868,I474252);
DFFARX1 I_27739  ( .D(I474269), .CLK(I2702), .RSTB(I473769), .Q(I473746) );
nand I_27740 (I473755,I474173,I474097);
not I_27741 (I474347,I2709);
nand I_27742 (I474364,I80780,I80762);
and I_27743 (I474381,I474364,I80774);
DFFARX1 I_27744  ( .D(I474381), .CLK(I2702), .RSTB(I474347), .Q(I474398) );
not I_27745 (I474415,I474398);
DFFARX1 I_27746  ( .D(I474398), .CLK(I2702), .RSTB(I474347), .Q(I474315) );
nor I_27747 (I474446,I80777,I80762);
DFFARX1 I_27748  ( .D(I80786), .CLK(I2702), .RSTB(I474347), .Q(I474463) );
DFFARX1 I_27749  ( .D(I474463), .CLK(I2702), .RSTB(I474347), .Q(I474480) );
not I_27750 (I474318,I474480);
DFFARX1 I_27751  ( .D(I474463), .CLK(I2702), .RSTB(I474347), .Q(I474511) );
and I_27752 (I474312,I474398,I474511);
nand I_27753 (I474542,I80765,I80789);
and I_27754 (I474559,I474542,I80768);
DFFARX1 I_27755  ( .D(I474559), .CLK(I2702), .RSTB(I474347), .Q(I474576) );
nor I_27756 (I474593,I474576,I474415);
not I_27757 (I474610,I474576);
nand I_27758 (I474321,I474398,I474610);
DFFARX1 I_27759  ( .D(I80771), .CLK(I2702), .RSTB(I474347), .Q(I474641) );
and I_27760 (I474658,I474641,I80783);
nor I_27761 (I474675,I474658,I474576);
nor I_27762 (I474692,I474658,I474610);
nand I_27763 (I474327,I474446,I474692);
not I_27764 (I474330,I474658);
DFFARX1 I_27765  ( .D(I474658), .CLK(I2702), .RSTB(I474347), .Q(I474309) );
DFFARX1 I_27766  ( .D(I80759), .CLK(I2702), .RSTB(I474347), .Q(I474751) );
nand I_27767 (I474768,I474751,I474463);
and I_27768 (I474785,I474446,I474768);
DFFARX1 I_27769  ( .D(I474785), .CLK(I2702), .RSTB(I474347), .Q(I474339) );
nor I_27770 (I474336,I474751,I474658);
and I_27771 (I474830,I474751,I474593);
or I_27772 (I474847,I474446,I474830);
DFFARX1 I_27773  ( .D(I474847), .CLK(I2702), .RSTB(I474347), .Q(I474324) );
nand I_27774 (I474333,I474751,I474675);
not I_27775 (I474925,I2709);
nand I_27776 (I474942,I678480,I678483);
and I_27777 (I474959,I474942,I678489);
DFFARX1 I_27778  ( .D(I474959), .CLK(I2702), .RSTB(I474925), .Q(I474976) );
not I_27779 (I474993,I474976);
DFFARX1 I_27780  ( .D(I474976), .CLK(I2702), .RSTB(I474925), .Q(I474893) );
nor I_27781 (I475024,I678486,I678483);
DFFARX1 I_27782  ( .D(I678465), .CLK(I2702), .RSTB(I474925), .Q(I475041) );
DFFARX1 I_27783  ( .D(I475041), .CLK(I2702), .RSTB(I474925), .Q(I475058) );
not I_27784 (I474896,I475058);
DFFARX1 I_27785  ( .D(I475041), .CLK(I2702), .RSTB(I474925), .Q(I475089) );
and I_27786 (I474890,I474976,I475089);
nand I_27787 (I475120,I678462,I678477);
and I_27788 (I475137,I475120,I678474);
DFFARX1 I_27789  ( .D(I475137), .CLK(I2702), .RSTB(I474925), .Q(I475154) );
nor I_27790 (I475171,I475154,I474993);
not I_27791 (I475188,I475154);
nand I_27792 (I474899,I474976,I475188);
DFFARX1 I_27793  ( .D(I678492), .CLK(I2702), .RSTB(I474925), .Q(I475219) );
and I_27794 (I475236,I475219,I678471);
nor I_27795 (I475253,I475236,I475154);
nor I_27796 (I475270,I475236,I475188);
nand I_27797 (I474905,I475024,I475270);
not I_27798 (I474908,I475236);
DFFARX1 I_27799  ( .D(I475236), .CLK(I2702), .RSTB(I474925), .Q(I474887) );
DFFARX1 I_27800  ( .D(I678468), .CLK(I2702), .RSTB(I474925), .Q(I475329) );
nand I_27801 (I475346,I475329,I475041);
and I_27802 (I475363,I475024,I475346);
DFFARX1 I_27803  ( .D(I475363), .CLK(I2702), .RSTB(I474925), .Q(I474917) );
nor I_27804 (I474914,I475329,I475236);
and I_27805 (I475408,I475329,I475171);
or I_27806 (I475425,I475024,I475408);
DFFARX1 I_27807  ( .D(I475425), .CLK(I2702), .RSTB(I474925), .Q(I474902) );
nand I_27808 (I474911,I475329,I475253);
not I_27809 (I475503,I2709);
nand I_27810 (I475520,I606578,I606575);
and I_27811 (I475537,I475520,I606569);
DFFARX1 I_27812  ( .D(I475537), .CLK(I2702), .RSTB(I475503), .Q(I475554) );
not I_27813 (I475571,I475554);
DFFARX1 I_27814  ( .D(I475554), .CLK(I2702), .RSTB(I475503), .Q(I475471) );
nor I_27815 (I475602,I606590,I606575);
DFFARX1 I_27816  ( .D(I606593), .CLK(I2702), .RSTB(I475503), .Q(I475619) );
DFFARX1 I_27817  ( .D(I475619), .CLK(I2702), .RSTB(I475503), .Q(I475636) );
not I_27818 (I475474,I475636);
DFFARX1 I_27819  ( .D(I475619), .CLK(I2702), .RSTB(I475503), .Q(I475667) );
and I_27820 (I475468,I475554,I475667);
nand I_27821 (I475698,I606596,I606587);
and I_27822 (I475715,I475698,I606599);
DFFARX1 I_27823  ( .D(I475715), .CLK(I2702), .RSTB(I475503), .Q(I475732) );
nor I_27824 (I475749,I475732,I475571);
not I_27825 (I475766,I475732);
nand I_27826 (I475477,I475554,I475766);
DFFARX1 I_27827  ( .D(I606572), .CLK(I2702), .RSTB(I475503), .Q(I475797) );
and I_27828 (I475814,I475797,I606581);
nor I_27829 (I475831,I475814,I475732);
nor I_27830 (I475848,I475814,I475766);
nand I_27831 (I475483,I475602,I475848);
not I_27832 (I475486,I475814);
DFFARX1 I_27833  ( .D(I475814), .CLK(I2702), .RSTB(I475503), .Q(I475465) );
DFFARX1 I_27834  ( .D(I606584), .CLK(I2702), .RSTB(I475503), .Q(I475907) );
nand I_27835 (I475924,I475907,I475619);
and I_27836 (I475941,I475602,I475924);
DFFARX1 I_27837  ( .D(I475941), .CLK(I2702), .RSTB(I475503), .Q(I475495) );
nor I_27838 (I475492,I475907,I475814);
and I_27839 (I475986,I475907,I475749);
or I_27840 (I476003,I475602,I475986);
DFFARX1 I_27841  ( .D(I476003), .CLK(I2702), .RSTB(I475503), .Q(I475480) );
nand I_27842 (I475489,I475907,I475831);
not I_27843 (I476081,I2709);
nand I_27844 (I476098,I618725,I618728);
and I_27845 (I476115,I476098,I618734);
DFFARX1 I_27846  ( .D(I476115), .CLK(I2702), .RSTB(I476081), .Q(I476132) );
not I_27847 (I476149,I476132);
DFFARX1 I_27848  ( .D(I476132), .CLK(I2702), .RSTB(I476081), .Q(I476049) );
nor I_27849 (I476180,I618731,I618728);
DFFARX1 I_27850  ( .D(I618710), .CLK(I2702), .RSTB(I476081), .Q(I476197) );
DFFARX1 I_27851  ( .D(I476197), .CLK(I2702), .RSTB(I476081), .Q(I476214) );
not I_27852 (I476052,I476214);
DFFARX1 I_27853  ( .D(I476197), .CLK(I2702), .RSTB(I476081), .Q(I476245) );
and I_27854 (I476046,I476132,I476245);
nand I_27855 (I476276,I618707,I618722);
and I_27856 (I476293,I476276,I618719);
DFFARX1 I_27857  ( .D(I476293), .CLK(I2702), .RSTB(I476081), .Q(I476310) );
nor I_27858 (I476327,I476310,I476149);
not I_27859 (I476344,I476310);
nand I_27860 (I476055,I476132,I476344);
DFFARX1 I_27861  ( .D(I618737), .CLK(I2702), .RSTB(I476081), .Q(I476375) );
and I_27862 (I476392,I476375,I618716);
nor I_27863 (I476409,I476392,I476310);
nor I_27864 (I476426,I476392,I476344);
nand I_27865 (I476061,I476180,I476426);
not I_27866 (I476064,I476392);
DFFARX1 I_27867  ( .D(I476392), .CLK(I2702), .RSTB(I476081), .Q(I476043) );
DFFARX1 I_27868  ( .D(I618713), .CLK(I2702), .RSTB(I476081), .Q(I476485) );
nand I_27869 (I476502,I476485,I476197);
and I_27870 (I476519,I476180,I476502);
DFFARX1 I_27871  ( .D(I476519), .CLK(I2702), .RSTB(I476081), .Q(I476073) );
nor I_27872 (I476070,I476485,I476392);
and I_27873 (I476564,I476485,I476327);
or I_27874 (I476581,I476180,I476564);
DFFARX1 I_27875  ( .D(I476581), .CLK(I2702), .RSTB(I476081), .Q(I476058) );
nand I_27876 (I476067,I476485,I476409);
not I_27877 (I476659,I2709);
nand I_27878 (I476676,I15630,I15645);
and I_27879 (I476693,I476676,I15633);
DFFARX1 I_27880  ( .D(I476693), .CLK(I2702), .RSTB(I476659), .Q(I476710) );
not I_27881 (I476727,I476710);
DFFARX1 I_27882  ( .D(I476710), .CLK(I2702), .RSTB(I476659), .Q(I476627) );
nor I_27883 (I476758,I15642,I15645);
DFFARX1 I_27884  ( .D(I15627), .CLK(I2702), .RSTB(I476659), .Q(I476775) );
DFFARX1 I_27885  ( .D(I476775), .CLK(I2702), .RSTB(I476659), .Q(I476792) );
not I_27886 (I476630,I476792);
DFFARX1 I_27887  ( .D(I476775), .CLK(I2702), .RSTB(I476659), .Q(I476823) );
and I_27888 (I476624,I476710,I476823);
nand I_27889 (I476854,I15618,I15615);
and I_27890 (I476871,I476854,I15621);
DFFARX1 I_27891  ( .D(I476871), .CLK(I2702), .RSTB(I476659), .Q(I476888) );
nor I_27892 (I476905,I476888,I476727);
not I_27893 (I476922,I476888);
nand I_27894 (I476633,I476710,I476922);
DFFARX1 I_27895  ( .D(I15624), .CLK(I2702), .RSTB(I476659), .Q(I476953) );
and I_27896 (I476970,I476953,I15636);
nor I_27897 (I476987,I476970,I476888);
nor I_27898 (I477004,I476970,I476922);
nand I_27899 (I476639,I476758,I477004);
not I_27900 (I476642,I476970);
DFFARX1 I_27901  ( .D(I476970), .CLK(I2702), .RSTB(I476659), .Q(I476621) );
DFFARX1 I_27902  ( .D(I15639), .CLK(I2702), .RSTB(I476659), .Q(I477063) );
nand I_27903 (I477080,I477063,I476775);
and I_27904 (I477097,I476758,I477080);
DFFARX1 I_27905  ( .D(I477097), .CLK(I2702), .RSTB(I476659), .Q(I476651) );
nor I_27906 (I476648,I477063,I476970);
and I_27907 (I477142,I477063,I476905);
or I_27908 (I477159,I476758,I477142);
DFFARX1 I_27909  ( .D(I477159), .CLK(I2702), .RSTB(I476659), .Q(I476636) );
nand I_27910 (I476645,I477063,I476987);
not I_27911 (I477237,I2709);
nand I_27912 (I477254,I84010,I83992);
and I_27913 (I477271,I477254,I84004);
DFFARX1 I_27914  ( .D(I477271), .CLK(I2702), .RSTB(I477237), .Q(I477288) );
not I_27915 (I477305,I477288);
DFFARX1 I_27916  ( .D(I477288), .CLK(I2702), .RSTB(I477237), .Q(I477205) );
nor I_27917 (I477336,I84007,I83992);
DFFARX1 I_27918  ( .D(I84016), .CLK(I2702), .RSTB(I477237), .Q(I477353) );
DFFARX1 I_27919  ( .D(I477353), .CLK(I2702), .RSTB(I477237), .Q(I477370) );
not I_27920 (I477208,I477370);
DFFARX1 I_27921  ( .D(I477353), .CLK(I2702), .RSTB(I477237), .Q(I477401) );
and I_27922 (I477202,I477288,I477401);
nand I_27923 (I477432,I83995,I84019);
and I_27924 (I477449,I477432,I83998);
DFFARX1 I_27925  ( .D(I477449), .CLK(I2702), .RSTB(I477237), .Q(I477466) );
nor I_27926 (I477483,I477466,I477305);
not I_27927 (I477500,I477466);
nand I_27928 (I477211,I477288,I477500);
DFFARX1 I_27929  ( .D(I84001), .CLK(I2702), .RSTB(I477237), .Q(I477531) );
and I_27930 (I477548,I477531,I84013);
nor I_27931 (I477565,I477548,I477466);
nor I_27932 (I477582,I477548,I477500);
nand I_27933 (I477217,I477336,I477582);
not I_27934 (I477220,I477548);
DFFARX1 I_27935  ( .D(I477548), .CLK(I2702), .RSTB(I477237), .Q(I477199) );
DFFARX1 I_27936  ( .D(I83989), .CLK(I2702), .RSTB(I477237), .Q(I477641) );
nand I_27937 (I477658,I477641,I477353);
and I_27938 (I477675,I477336,I477658);
DFFARX1 I_27939  ( .D(I477675), .CLK(I2702), .RSTB(I477237), .Q(I477229) );
nor I_27940 (I477226,I477641,I477548);
and I_27941 (I477720,I477641,I477483);
or I_27942 (I477737,I477336,I477720);
DFFARX1 I_27943  ( .D(I477737), .CLK(I2702), .RSTB(I477237), .Q(I477214) );
nand I_27944 (I477223,I477641,I477565);
not I_27945 (I477815,I2709);
nand I_27946 (I477832,I538766,I538754);
and I_27947 (I477849,I477832,I538748);
DFFARX1 I_27948  ( .D(I477849), .CLK(I2702), .RSTB(I477815), .Q(I477866) );
not I_27949 (I477883,I477866);
DFFARX1 I_27950  ( .D(I477866), .CLK(I2702), .RSTB(I477815), .Q(I477783) );
nor I_27951 (I477914,I538745,I538754);
DFFARX1 I_27952  ( .D(I538739), .CLK(I2702), .RSTB(I477815), .Q(I477931) );
DFFARX1 I_27953  ( .D(I477931), .CLK(I2702), .RSTB(I477815), .Q(I477948) );
not I_27954 (I477786,I477948);
DFFARX1 I_27955  ( .D(I477931), .CLK(I2702), .RSTB(I477815), .Q(I477979) );
and I_27956 (I477780,I477866,I477979);
nand I_27957 (I478010,I538742,I538757);
and I_27958 (I478027,I478010,I538769);
DFFARX1 I_27959  ( .D(I478027), .CLK(I2702), .RSTB(I477815), .Q(I478044) );
nor I_27960 (I478061,I478044,I477883);
not I_27961 (I478078,I478044);
nand I_27962 (I477789,I477866,I478078);
DFFARX1 I_27963  ( .D(I538760), .CLK(I2702), .RSTB(I477815), .Q(I478109) );
and I_27964 (I478126,I478109,I538751);
nor I_27965 (I478143,I478126,I478044);
nor I_27966 (I478160,I478126,I478078);
nand I_27967 (I477795,I477914,I478160);
not I_27968 (I477798,I478126);
DFFARX1 I_27969  ( .D(I478126), .CLK(I2702), .RSTB(I477815), .Q(I477777) );
DFFARX1 I_27970  ( .D(I538763), .CLK(I2702), .RSTB(I477815), .Q(I478219) );
nand I_27971 (I478236,I478219,I477931);
and I_27972 (I478253,I477914,I478236);
DFFARX1 I_27973  ( .D(I478253), .CLK(I2702), .RSTB(I477815), .Q(I477807) );
nor I_27974 (I477804,I478219,I478126);
and I_27975 (I478298,I478219,I478061);
or I_27976 (I478315,I477914,I478298);
DFFARX1 I_27977  ( .D(I478315), .CLK(I2702), .RSTB(I477815), .Q(I477792) );
nand I_27978 (I477801,I478219,I478143);
not I_27979 (I478393,I2709);
nand I_27980 (I478410,I628789,I628792);
and I_27981 (I478427,I478410,I628798);
DFFARX1 I_27982  ( .D(I478427), .CLK(I2702), .RSTB(I478393), .Q(I478444) );
not I_27983 (I478461,I478444);
DFFARX1 I_27984  ( .D(I478444), .CLK(I2702), .RSTB(I478393), .Q(I478361) );
nor I_27985 (I478492,I628795,I628792);
DFFARX1 I_27986  ( .D(I628774), .CLK(I2702), .RSTB(I478393), .Q(I478509) );
DFFARX1 I_27987  ( .D(I478509), .CLK(I2702), .RSTB(I478393), .Q(I478526) );
not I_27988 (I478364,I478526);
DFFARX1 I_27989  ( .D(I478509), .CLK(I2702), .RSTB(I478393), .Q(I478557) );
and I_27990 (I478358,I478444,I478557);
nand I_27991 (I478588,I628771,I628786);
and I_27992 (I478605,I478588,I628783);
DFFARX1 I_27993  ( .D(I478605), .CLK(I2702), .RSTB(I478393), .Q(I478622) );
nor I_27994 (I478639,I478622,I478461);
not I_27995 (I478656,I478622);
nand I_27996 (I478367,I478444,I478656);
DFFARX1 I_27997  ( .D(I628801), .CLK(I2702), .RSTB(I478393), .Q(I478687) );
and I_27998 (I478704,I478687,I628780);
nor I_27999 (I478721,I478704,I478622);
nor I_28000 (I478738,I478704,I478656);
nand I_28001 (I478373,I478492,I478738);
not I_28002 (I478376,I478704);
DFFARX1 I_28003  ( .D(I478704), .CLK(I2702), .RSTB(I478393), .Q(I478355) );
DFFARX1 I_28004  ( .D(I628777), .CLK(I2702), .RSTB(I478393), .Q(I478797) );
nand I_28005 (I478814,I478797,I478509);
and I_28006 (I478831,I478492,I478814);
DFFARX1 I_28007  ( .D(I478831), .CLK(I2702), .RSTB(I478393), .Q(I478385) );
nor I_28008 (I478382,I478797,I478704);
and I_28009 (I478876,I478797,I478639);
or I_28010 (I478893,I478492,I478876);
DFFARX1 I_28011  ( .D(I478893), .CLK(I2702), .RSTB(I478393), .Q(I478370) );
nand I_28012 (I478379,I478797,I478721);
not I_28013 (I478971,I2709);
nand I_28014 (I478988,I413177,I413207);
and I_28015 (I479005,I478988,I413204);
DFFARX1 I_28016  ( .D(I479005), .CLK(I2702), .RSTB(I478971), .Q(I479022) );
not I_28017 (I479039,I479022);
DFFARX1 I_28018  ( .D(I479022), .CLK(I2702), .RSTB(I478971), .Q(I478939) );
nor I_28019 (I479070,I413195,I413207);
DFFARX1 I_28020  ( .D(I413183), .CLK(I2702), .RSTB(I478971), .Q(I479087) );
DFFARX1 I_28021  ( .D(I479087), .CLK(I2702), .RSTB(I478971), .Q(I479104) );
not I_28022 (I478942,I479104);
DFFARX1 I_28023  ( .D(I479087), .CLK(I2702), .RSTB(I478971), .Q(I479135) );
and I_28024 (I478936,I479022,I479135);
nand I_28025 (I479166,I413186,I413192);
and I_28026 (I479183,I479166,I413198);
DFFARX1 I_28027  ( .D(I479183), .CLK(I2702), .RSTB(I478971), .Q(I479200) );
nor I_28028 (I479217,I479200,I479039);
not I_28029 (I479234,I479200);
nand I_28030 (I478945,I479022,I479234);
DFFARX1 I_28031  ( .D(I413189), .CLK(I2702), .RSTB(I478971), .Q(I479265) );
and I_28032 (I479282,I479265,I413180);
nor I_28033 (I479299,I479282,I479200);
nor I_28034 (I479316,I479282,I479234);
nand I_28035 (I478951,I479070,I479316);
not I_28036 (I478954,I479282);
DFFARX1 I_28037  ( .D(I479282), .CLK(I2702), .RSTB(I478971), .Q(I478933) );
DFFARX1 I_28038  ( .D(I413201), .CLK(I2702), .RSTB(I478971), .Q(I479375) );
nand I_28039 (I479392,I479375,I479087);
and I_28040 (I479409,I479070,I479392);
DFFARX1 I_28041  ( .D(I479409), .CLK(I2702), .RSTB(I478971), .Q(I478963) );
nor I_28042 (I478960,I479375,I479282);
and I_28043 (I479454,I479375,I479217);
or I_28044 (I479471,I479070,I479454);
DFFARX1 I_28045  ( .D(I479471), .CLK(I2702), .RSTB(I478971), .Q(I478948) );
nand I_28046 (I478957,I479375,I479299);
not I_28047 (I479549,I2709);
nand I_28048 (I479566,I184656,I184635);
and I_28049 (I479583,I479566,I184632);
DFFARX1 I_28050  ( .D(I479583), .CLK(I2702), .RSTB(I479549), .Q(I479600) );
not I_28051 (I479617,I479600);
DFFARX1 I_28052  ( .D(I479600), .CLK(I2702), .RSTB(I479549), .Q(I479517) );
nor I_28053 (I479648,I184641,I184635);
DFFARX1 I_28054  ( .D(I184629), .CLK(I2702), .RSTB(I479549), .Q(I479665) );
DFFARX1 I_28055  ( .D(I479665), .CLK(I2702), .RSTB(I479549), .Q(I479682) );
not I_28056 (I479520,I479682);
DFFARX1 I_28057  ( .D(I479665), .CLK(I2702), .RSTB(I479549), .Q(I479713) );
and I_28058 (I479514,I479600,I479713);
nand I_28059 (I479744,I184659,I184650);
and I_28060 (I479761,I479744,I184647);
DFFARX1 I_28061  ( .D(I479761), .CLK(I2702), .RSTB(I479549), .Q(I479778) );
nor I_28062 (I479795,I479778,I479617);
not I_28063 (I479812,I479778);
nand I_28064 (I479523,I479600,I479812);
DFFARX1 I_28065  ( .D(I184644), .CLK(I2702), .RSTB(I479549), .Q(I479843) );
and I_28066 (I479860,I479843,I184653);
nor I_28067 (I479877,I479860,I479778);
nor I_28068 (I479894,I479860,I479812);
nand I_28069 (I479529,I479648,I479894);
not I_28070 (I479532,I479860);
DFFARX1 I_28071  ( .D(I479860), .CLK(I2702), .RSTB(I479549), .Q(I479511) );
DFFARX1 I_28072  ( .D(I184638), .CLK(I2702), .RSTB(I479549), .Q(I479953) );
nand I_28073 (I479970,I479953,I479665);
and I_28074 (I479987,I479648,I479970);
DFFARX1 I_28075  ( .D(I479987), .CLK(I2702), .RSTB(I479549), .Q(I479541) );
nor I_28076 (I479538,I479953,I479860);
and I_28077 (I480032,I479953,I479795);
or I_28078 (I480049,I479648,I480032);
DFFARX1 I_28079  ( .D(I480049), .CLK(I2702), .RSTB(I479549), .Q(I479526) );
nand I_28080 (I479535,I479953,I479877);
not I_28081 (I480127,I2709);
nand I_28082 (I480144,I201687,I201672);
and I_28083 (I480161,I480144,I201681);
DFFARX1 I_28084  ( .D(I480161), .CLK(I2702), .RSTB(I480127), .Q(I480178) );
not I_28085 (I480195,I480178);
DFFARX1 I_28086  ( .D(I480178), .CLK(I2702), .RSTB(I480127), .Q(I480095) );
nor I_28087 (I480226,I201690,I201672);
DFFARX1 I_28088  ( .D(I201669), .CLK(I2702), .RSTB(I480127), .Q(I480243) );
DFFARX1 I_28089  ( .D(I480243), .CLK(I2702), .RSTB(I480127), .Q(I480260) );
not I_28090 (I480098,I480260);
DFFARX1 I_28091  ( .D(I480243), .CLK(I2702), .RSTB(I480127), .Q(I480291) );
and I_28092 (I480092,I480178,I480291);
nand I_28093 (I480322,I201693,I201666);
and I_28094 (I480339,I480322,I201684);
DFFARX1 I_28095  ( .D(I480339), .CLK(I2702), .RSTB(I480127), .Q(I480356) );
nor I_28096 (I480373,I480356,I480195);
not I_28097 (I480390,I480356);
nand I_28098 (I480101,I480178,I480390);
DFFARX1 I_28099  ( .D(I201678), .CLK(I2702), .RSTB(I480127), .Q(I480421) );
and I_28100 (I480438,I480421,I201663);
nor I_28101 (I480455,I480438,I480356);
nor I_28102 (I480472,I480438,I480390);
nand I_28103 (I480107,I480226,I480472);
not I_28104 (I480110,I480438);
DFFARX1 I_28105  ( .D(I480438), .CLK(I2702), .RSTB(I480127), .Q(I480089) );
DFFARX1 I_28106  ( .D(I201675), .CLK(I2702), .RSTB(I480127), .Q(I480531) );
nand I_28107 (I480548,I480531,I480243);
and I_28108 (I480565,I480226,I480548);
DFFARX1 I_28109  ( .D(I480565), .CLK(I2702), .RSTB(I480127), .Q(I480119) );
nor I_28110 (I480116,I480531,I480438);
and I_28111 (I480610,I480531,I480373);
or I_28112 (I480627,I480226,I480610);
DFFARX1 I_28113  ( .D(I480627), .CLK(I2702), .RSTB(I480127), .Q(I480104) );
nand I_28114 (I480113,I480531,I480455);
not I_28115 (I480705,I2709);
nand I_28116 (I480722,I658352,I658355);
and I_28117 (I480739,I480722,I658361);
DFFARX1 I_28118  ( .D(I480739), .CLK(I2702), .RSTB(I480705), .Q(I480756) );
not I_28119 (I480773,I480756);
DFFARX1 I_28120  ( .D(I480756), .CLK(I2702), .RSTB(I480705), .Q(I480673) );
nor I_28121 (I480804,I658358,I658355);
DFFARX1 I_28122  ( .D(I658337), .CLK(I2702), .RSTB(I480705), .Q(I480821) );
DFFARX1 I_28123  ( .D(I480821), .CLK(I2702), .RSTB(I480705), .Q(I480838) );
not I_28124 (I480676,I480838);
DFFARX1 I_28125  ( .D(I480821), .CLK(I2702), .RSTB(I480705), .Q(I480869) );
and I_28126 (I480670,I480756,I480869);
nand I_28127 (I480900,I658334,I658349);
and I_28128 (I480917,I480900,I658346);
DFFARX1 I_28129  ( .D(I480917), .CLK(I2702), .RSTB(I480705), .Q(I480934) );
nor I_28130 (I480951,I480934,I480773);
not I_28131 (I480968,I480934);
nand I_28132 (I480679,I480756,I480968);
DFFARX1 I_28133  ( .D(I658364), .CLK(I2702), .RSTB(I480705), .Q(I480999) );
and I_28134 (I481016,I480999,I658343);
nor I_28135 (I481033,I481016,I480934);
nor I_28136 (I481050,I481016,I480968);
nand I_28137 (I480685,I480804,I481050);
not I_28138 (I480688,I481016);
DFFARX1 I_28139  ( .D(I481016), .CLK(I2702), .RSTB(I480705), .Q(I480667) );
DFFARX1 I_28140  ( .D(I658340), .CLK(I2702), .RSTB(I480705), .Q(I481109) );
nand I_28141 (I481126,I481109,I480821);
and I_28142 (I481143,I480804,I481126);
DFFARX1 I_28143  ( .D(I481143), .CLK(I2702), .RSTB(I480705), .Q(I480697) );
nor I_28144 (I480694,I481109,I481016);
and I_28145 (I481188,I481109,I480951);
or I_28146 (I481205,I480804,I481188);
DFFARX1 I_28147  ( .D(I481205), .CLK(I2702), .RSTB(I480705), .Q(I480682) );
nand I_28148 (I480691,I481109,I481033);
not I_28149 (I481283,I2709);
nand I_28150 (I481300,I609553,I609550);
and I_28151 (I481317,I481300,I609544);
DFFARX1 I_28152  ( .D(I481317), .CLK(I2702), .RSTB(I481283), .Q(I481334) );
not I_28153 (I481351,I481334);
DFFARX1 I_28154  ( .D(I481334), .CLK(I2702), .RSTB(I481283), .Q(I481251) );
nor I_28155 (I481382,I609565,I609550);
DFFARX1 I_28156  ( .D(I609568), .CLK(I2702), .RSTB(I481283), .Q(I481399) );
DFFARX1 I_28157  ( .D(I481399), .CLK(I2702), .RSTB(I481283), .Q(I481416) );
not I_28158 (I481254,I481416);
DFFARX1 I_28159  ( .D(I481399), .CLK(I2702), .RSTB(I481283), .Q(I481447) );
and I_28160 (I481248,I481334,I481447);
nand I_28161 (I481478,I609571,I609562);
and I_28162 (I481495,I481478,I609574);
DFFARX1 I_28163  ( .D(I481495), .CLK(I2702), .RSTB(I481283), .Q(I481512) );
nor I_28164 (I481529,I481512,I481351);
not I_28165 (I481546,I481512);
nand I_28166 (I481257,I481334,I481546);
DFFARX1 I_28167  ( .D(I609547), .CLK(I2702), .RSTB(I481283), .Q(I481577) );
and I_28168 (I481594,I481577,I609556);
nor I_28169 (I481611,I481594,I481512);
nor I_28170 (I481628,I481594,I481546);
nand I_28171 (I481263,I481382,I481628);
not I_28172 (I481266,I481594);
DFFARX1 I_28173  ( .D(I481594), .CLK(I2702), .RSTB(I481283), .Q(I481245) );
DFFARX1 I_28174  ( .D(I609559), .CLK(I2702), .RSTB(I481283), .Q(I481687) );
nand I_28175 (I481704,I481687,I481399);
and I_28176 (I481721,I481382,I481704);
DFFARX1 I_28177  ( .D(I481721), .CLK(I2702), .RSTB(I481283), .Q(I481275) );
nor I_28178 (I481272,I481687,I481594);
and I_28179 (I481766,I481687,I481529);
or I_28180 (I481783,I481382,I481766);
DFFARX1 I_28181  ( .D(I481783), .CLK(I2702), .RSTB(I481283), .Q(I481260) );
nand I_28182 (I481269,I481687,I481611);
not I_28183 (I481861,I2709);
nand I_28184 (I481878,I421133,I421163);
and I_28185 (I481895,I481878,I421160);
DFFARX1 I_28186  ( .D(I481895), .CLK(I2702), .RSTB(I481861), .Q(I481912) );
not I_28187 (I481929,I481912);
DFFARX1 I_28188  ( .D(I481912), .CLK(I2702), .RSTB(I481861), .Q(I481829) );
nor I_28189 (I481960,I421151,I421163);
DFFARX1 I_28190  ( .D(I421139), .CLK(I2702), .RSTB(I481861), .Q(I481977) );
DFFARX1 I_28191  ( .D(I481977), .CLK(I2702), .RSTB(I481861), .Q(I481994) );
not I_28192 (I481832,I481994);
DFFARX1 I_28193  ( .D(I481977), .CLK(I2702), .RSTB(I481861), .Q(I482025) );
and I_28194 (I481826,I481912,I482025);
nand I_28195 (I482056,I421142,I421148);
and I_28196 (I482073,I482056,I421154);
DFFARX1 I_28197  ( .D(I482073), .CLK(I2702), .RSTB(I481861), .Q(I482090) );
nor I_28198 (I482107,I482090,I481929);
not I_28199 (I482124,I482090);
nand I_28200 (I481835,I481912,I482124);
DFFARX1 I_28201  ( .D(I421145), .CLK(I2702), .RSTB(I481861), .Q(I482155) );
and I_28202 (I482172,I482155,I421136);
nor I_28203 (I482189,I482172,I482090);
nor I_28204 (I482206,I482172,I482124);
nand I_28205 (I481841,I481960,I482206);
not I_28206 (I481844,I482172);
DFFARX1 I_28207  ( .D(I482172), .CLK(I2702), .RSTB(I481861), .Q(I481823) );
DFFARX1 I_28208  ( .D(I421157), .CLK(I2702), .RSTB(I481861), .Q(I482265) );
nand I_28209 (I482282,I482265,I481977);
and I_28210 (I482299,I481960,I482282);
DFFARX1 I_28211  ( .D(I482299), .CLK(I2702), .RSTB(I481861), .Q(I481853) );
nor I_28212 (I481850,I482265,I482172);
and I_28213 (I482344,I482265,I482107);
or I_28214 (I482361,I481960,I482344);
DFFARX1 I_28215  ( .D(I482361), .CLK(I2702), .RSTB(I481861), .Q(I481838) );
nand I_28216 (I481847,I482265,I482189);
not I_28217 (I482439,I2709);
nand I_28218 (I482456,I652062,I652065);
and I_28219 (I482473,I482456,I652071);
DFFARX1 I_28220  ( .D(I482473), .CLK(I2702), .RSTB(I482439), .Q(I482490) );
not I_28221 (I482507,I482490);
DFFARX1 I_28222  ( .D(I482490), .CLK(I2702), .RSTB(I482439), .Q(I482407) );
nor I_28223 (I482538,I652068,I652065);
DFFARX1 I_28224  ( .D(I652047), .CLK(I2702), .RSTB(I482439), .Q(I482555) );
DFFARX1 I_28225  ( .D(I482555), .CLK(I2702), .RSTB(I482439), .Q(I482572) );
not I_28226 (I482410,I482572);
DFFARX1 I_28227  ( .D(I482555), .CLK(I2702), .RSTB(I482439), .Q(I482603) );
and I_28228 (I482404,I482490,I482603);
nand I_28229 (I482634,I652044,I652059);
and I_28230 (I482651,I482634,I652056);
DFFARX1 I_28231  ( .D(I482651), .CLK(I2702), .RSTB(I482439), .Q(I482668) );
nor I_28232 (I482685,I482668,I482507);
not I_28233 (I482702,I482668);
nand I_28234 (I482413,I482490,I482702);
DFFARX1 I_28235  ( .D(I652074), .CLK(I2702), .RSTB(I482439), .Q(I482733) );
and I_28236 (I482750,I482733,I652053);
nor I_28237 (I482767,I482750,I482668);
nor I_28238 (I482784,I482750,I482702);
nand I_28239 (I482419,I482538,I482784);
not I_28240 (I482422,I482750);
DFFARX1 I_28241  ( .D(I482750), .CLK(I2702), .RSTB(I482439), .Q(I482401) );
DFFARX1 I_28242  ( .D(I652050), .CLK(I2702), .RSTB(I482439), .Q(I482843) );
nand I_28243 (I482860,I482843,I482555);
and I_28244 (I482877,I482538,I482860);
DFFARX1 I_28245  ( .D(I482877), .CLK(I2702), .RSTB(I482439), .Q(I482431) );
nor I_28246 (I482428,I482843,I482750);
and I_28247 (I482922,I482843,I482685);
or I_28248 (I482939,I482538,I482922);
DFFARX1 I_28249  ( .D(I482939), .CLK(I2702), .RSTB(I482439), .Q(I482416) );
nand I_28250 (I482425,I482843,I482767);
not I_28251 (I483017,I2709);
nand I_28252 (I483034,I513181,I513169);
and I_28253 (I483051,I483034,I513163);
DFFARX1 I_28254  ( .D(I483051), .CLK(I2702), .RSTB(I483017), .Q(I483068) );
not I_28255 (I483085,I483068);
DFFARX1 I_28256  ( .D(I483068), .CLK(I2702), .RSTB(I483017), .Q(I482985) );
nor I_28257 (I483116,I513160,I513169);
DFFARX1 I_28258  ( .D(I513154), .CLK(I2702), .RSTB(I483017), .Q(I483133) );
DFFARX1 I_28259  ( .D(I483133), .CLK(I2702), .RSTB(I483017), .Q(I483150) );
not I_28260 (I482988,I483150);
DFFARX1 I_28261  ( .D(I483133), .CLK(I2702), .RSTB(I483017), .Q(I483181) );
and I_28262 (I482982,I483068,I483181);
nand I_28263 (I483212,I513157,I513172);
and I_28264 (I483229,I483212,I513184);
DFFARX1 I_28265  ( .D(I483229), .CLK(I2702), .RSTB(I483017), .Q(I483246) );
nor I_28266 (I483263,I483246,I483085);
not I_28267 (I483280,I483246);
nand I_28268 (I482991,I483068,I483280);
DFFARX1 I_28269  ( .D(I513175), .CLK(I2702), .RSTB(I483017), .Q(I483311) );
and I_28270 (I483328,I483311,I513166);
nor I_28271 (I483345,I483328,I483246);
nor I_28272 (I483362,I483328,I483280);
nand I_28273 (I482997,I483116,I483362);
not I_28274 (I483000,I483328);
DFFARX1 I_28275  ( .D(I483328), .CLK(I2702), .RSTB(I483017), .Q(I482979) );
DFFARX1 I_28276  ( .D(I513178), .CLK(I2702), .RSTB(I483017), .Q(I483421) );
nand I_28277 (I483438,I483421,I483133);
and I_28278 (I483455,I483116,I483438);
DFFARX1 I_28279  ( .D(I483455), .CLK(I2702), .RSTB(I483017), .Q(I483009) );
nor I_28280 (I483006,I483421,I483328);
and I_28281 (I483500,I483421,I483263);
or I_28282 (I483517,I483116,I483500);
DFFARX1 I_28283  ( .D(I483517), .CLK(I2702), .RSTB(I483017), .Q(I482994) );
nand I_28284 (I483003,I483421,I483345);
not I_28285 (I483595,I2709);
nand I_28286 (I483612,I124062,I124044);
and I_28287 (I483629,I483612,I124056);
DFFARX1 I_28288  ( .D(I483629), .CLK(I2702), .RSTB(I483595), .Q(I483646) );
not I_28289 (I483663,I483646);
DFFARX1 I_28290  ( .D(I483646), .CLK(I2702), .RSTB(I483595), .Q(I483563) );
nor I_28291 (I483694,I124059,I124044);
DFFARX1 I_28292  ( .D(I124068), .CLK(I2702), .RSTB(I483595), .Q(I483711) );
DFFARX1 I_28293  ( .D(I483711), .CLK(I2702), .RSTB(I483595), .Q(I483728) );
not I_28294 (I483566,I483728);
DFFARX1 I_28295  ( .D(I483711), .CLK(I2702), .RSTB(I483595), .Q(I483759) );
and I_28296 (I483560,I483646,I483759);
nand I_28297 (I483790,I124047,I124071);
and I_28298 (I483807,I483790,I124050);
DFFARX1 I_28299  ( .D(I483807), .CLK(I2702), .RSTB(I483595), .Q(I483824) );
nor I_28300 (I483841,I483824,I483663);
not I_28301 (I483858,I483824);
nand I_28302 (I483569,I483646,I483858);
DFFARX1 I_28303  ( .D(I124053), .CLK(I2702), .RSTB(I483595), .Q(I483889) );
and I_28304 (I483906,I483889,I124065);
nor I_28305 (I483923,I483906,I483824);
nor I_28306 (I483940,I483906,I483858);
nand I_28307 (I483575,I483694,I483940);
not I_28308 (I483578,I483906);
DFFARX1 I_28309  ( .D(I483906), .CLK(I2702), .RSTB(I483595), .Q(I483557) );
DFFARX1 I_28310  ( .D(I124041), .CLK(I2702), .RSTB(I483595), .Q(I483999) );
nand I_28311 (I484016,I483999,I483711);
and I_28312 (I484033,I483694,I484016);
DFFARX1 I_28313  ( .D(I484033), .CLK(I2702), .RSTB(I483595), .Q(I483587) );
nor I_28314 (I483584,I483999,I483906);
and I_28315 (I484078,I483999,I483841);
or I_28316 (I484095,I483694,I484078);
DFFARX1 I_28317  ( .D(I484095), .CLK(I2702), .RSTB(I483595), .Q(I483572) );
nand I_28318 (I483581,I483999,I483923);
not I_28319 (I484173,I2709);
nand I_28320 (I484190,I286071,I286098);
and I_28321 (I484207,I484190,I286086);
DFFARX1 I_28322  ( .D(I484207), .CLK(I2702), .RSTB(I484173), .Q(I484224) );
not I_28323 (I484241,I484224);
DFFARX1 I_28324  ( .D(I484224), .CLK(I2702), .RSTB(I484173), .Q(I484141) );
nor I_28325 (I484272,I286074,I286098);
DFFARX1 I_28326  ( .D(I286089), .CLK(I2702), .RSTB(I484173), .Q(I484289) );
DFFARX1 I_28327  ( .D(I484289), .CLK(I2702), .RSTB(I484173), .Q(I484306) );
not I_28328 (I484144,I484306);
DFFARX1 I_28329  ( .D(I484289), .CLK(I2702), .RSTB(I484173), .Q(I484337) );
and I_28330 (I484138,I484224,I484337);
nand I_28331 (I484368,I286083,I286080);
and I_28332 (I484385,I484368,I286077);
DFFARX1 I_28333  ( .D(I484385), .CLK(I2702), .RSTB(I484173), .Q(I484402) );
nor I_28334 (I484419,I484402,I484241);
not I_28335 (I484436,I484402);
nand I_28336 (I484147,I484224,I484436);
DFFARX1 I_28337  ( .D(I286092), .CLK(I2702), .RSTB(I484173), .Q(I484467) );
and I_28338 (I484484,I484467,I286068);
nor I_28339 (I484501,I484484,I484402);
nor I_28340 (I484518,I484484,I484436);
nand I_28341 (I484153,I484272,I484518);
not I_28342 (I484156,I484484);
DFFARX1 I_28343  ( .D(I484484), .CLK(I2702), .RSTB(I484173), .Q(I484135) );
DFFARX1 I_28344  ( .D(I286095), .CLK(I2702), .RSTB(I484173), .Q(I484577) );
nand I_28345 (I484594,I484577,I484289);
and I_28346 (I484611,I484272,I484594);
DFFARX1 I_28347  ( .D(I484611), .CLK(I2702), .RSTB(I484173), .Q(I484165) );
nor I_28348 (I484162,I484577,I484484);
and I_28349 (I484656,I484577,I484419);
or I_28350 (I484673,I484272,I484656);
DFFARX1 I_28351  ( .D(I484673), .CLK(I2702), .RSTB(I484173), .Q(I484150) );
nand I_28352 (I484159,I484577,I484501);
not I_28353 (I484751,I2709);
nand I_28354 (I484768,I402924,I402921);
and I_28355 (I484785,I484768,I402933);
DFFARX1 I_28356  ( .D(I484785), .CLK(I2702), .RSTB(I484751), .Q(I484802) );
not I_28357 (I484819,I484802);
DFFARX1 I_28358  ( .D(I484802), .CLK(I2702), .RSTB(I484751), .Q(I484719) );
nor I_28359 (I484850,I402930,I402921);
DFFARX1 I_28360  ( .D(I402936), .CLK(I2702), .RSTB(I484751), .Q(I484867) );
DFFARX1 I_28361  ( .D(I484867), .CLK(I2702), .RSTB(I484751), .Q(I484884) );
not I_28362 (I484722,I484884);
DFFARX1 I_28363  ( .D(I484867), .CLK(I2702), .RSTB(I484751), .Q(I484915) );
and I_28364 (I484716,I484802,I484915);
nand I_28365 (I484946,I402912,I402915);
and I_28366 (I484963,I484946,I402939);
DFFARX1 I_28367  ( .D(I484963), .CLK(I2702), .RSTB(I484751), .Q(I484980) );
nor I_28368 (I484997,I484980,I484819);
not I_28369 (I485014,I484980);
nand I_28370 (I484725,I484802,I485014);
DFFARX1 I_28371  ( .D(I402918), .CLK(I2702), .RSTB(I484751), .Q(I485045) );
and I_28372 (I485062,I485045,I402909);
nor I_28373 (I485079,I485062,I484980);
nor I_28374 (I485096,I485062,I485014);
nand I_28375 (I484731,I484850,I485096);
not I_28376 (I484734,I485062);
DFFARX1 I_28377  ( .D(I485062), .CLK(I2702), .RSTB(I484751), .Q(I484713) );
DFFARX1 I_28378  ( .D(I402927), .CLK(I2702), .RSTB(I484751), .Q(I485155) );
nand I_28379 (I485172,I485155,I484867);
and I_28380 (I485189,I484850,I485172);
DFFARX1 I_28381  ( .D(I485189), .CLK(I2702), .RSTB(I484751), .Q(I484743) );
nor I_28382 (I484740,I485155,I485062);
and I_28383 (I485234,I485155,I484997);
or I_28384 (I485251,I484850,I485234);
DFFARX1 I_28385  ( .D(I485251), .CLK(I2702), .RSTB(I484751), .Q(I484728) );
nand I_28386 (I484737,I485155,I485079);
not I_28387 (I485329,I2709);
nand I_28388 (I485346,I413789,I413819);
and I_28389 (I485363,I485346,I413816);
DFFARX1 I_28390  ( .D(I485363), .CLK(I2702), .RSTB(I485329), .Q(I485380) );
not I_28391 (I485397,I485380);
DFFARX1 I_28392  ( .D(I485380), .CLK(I2702), .RSTB(I485329), .Q(I485297) );
nor I_28393 (I485428,I413807,I413819);
DFFARX1 I_28394  ( .D(I413795), .CLK(I2702), .RSTB(I485329), .Q(I485445) );
DFFARX1 I_28395  ( .D(I485445), .CLK(I2702), .RSTB(I485329), .Q(I485462) );
not I_28396 (I485300,I485462);
DFFARX1 I_28397  ( .D(I485445), .CLK(I2702), .RSTB(I485329), .Q(I485493) );
and I_28398 (I485294,I485380,I485493);
nand I_28399 (I485524,I413798,I413804);
and I_28400 (I485541,I485524,I413810);
DFFARX1 I_28401  ( .D(I485541), .CLK(I2702), .RSTB(I485329), .Q(I485558) );
nor I_28402 (I485575,I485558,I485397);
not I_28403 (I485592,I485558);
nand I_28404 (I485303,I485380,I485592);
DFFARX1 I_28405  ( .D(I413801), .CLK(I2702), .RSTB(I485329), .Q(I485623) );
and I_28406 (I485640,I485623,I413792);
nor I_28407 (I485657,I485640,I485558);
nor I_28408 (I485674,I485640,I485592);
nand I_28409 (I485309,I485428,I485674);
not I_28410 (I485312,I485640);
DFFARX1 I_28411  ( .D(I485640), .CLK(I2702), .RSTB(I485329), .Q(I485291) );
DFFARX1 I_28412  ( .D(I413813), .CLK(I2702), .RSTB(I485329), .Q(I485733) );
nand I_28413 (I485750,I485733,I485445);
and I_28414 (I485767,I485428,I485750);
DFFARX1 I_28415  ( .D(I485767), .CLK(I2702), .RSTB(I485329), .Q(I485321) );
nor I_28416 (I485318,I485733,I485640);
and I_28417 (I485812,I485733,I485575);
or I_28418 (I485829,I485428,I485812);
DFFARX1 I_28419  ( .D(I485829), .CLK(I2702), .RSTB(I485329), .Q(I485306) );
nand I_28420 (I485315,I485733,I485657);
not I_28421 (I485907,I2709);
nand I_28422 (I485924,I702515,I702527);
and I_28423 (I485941,I485924,I702500);
DFFARX1 I_28424  ( .D(I485941), .CLK(I2702), .RSTB(I485907), .Q(I485958) );
not I_28425 (I485975,I485958);
DFFARX1 I_28426  ( .D(I485958), .CLK(I2702), .RSTB(I485907), .Q(I485875) );
nor I_28427 (I486006,I702518,I702527);
DFFARX1 I_28428  ( .D(I702509), .CLK(I2702), .RSTB(I485907), .Q(I486023) );
DFFARX1 I_28429  ( .D(I486023), .CLK(I2702), .RSTB(I485907), .Q(I486040) );
not I_28430 (I485878,I486040);
DFFARX1 I_28431  ( .D(I486023), .CLK(I2702), .RSTB(I485907), .Q(I486071) );
and I_28432 (I485872,I485958,I486071);
nand I_28433 (I486102,I702506,I702512);
and I_28434 (I486119,I486102,I702524);
DFFARX1 I_28435  ( .D(I486119), .CLK(I2702), .RSTB(I485907), .Q(I486136) );
nor I_28436 (I486153,I486136,I485975);
not I_28437 (I486170,I486136);
nand I_28438 (I485881,I485958,I486170);
DFFARX1 I_28439  ( .D(I702530), .CLK(I2702), .RSTB(I485907), .Q(I486201) );
and I_28440 (I486218,I486201,I702521);
nor I_28441 (I486235,I486218,I486136);
nor I_28442 (I486252,I486218,I486170);
nand I_28443 (I485887,I486006,I486252);
not I_28444 (I485890,I486218);
DFFARX1 I_28445  ( .D(I486218), .CLK(I2702), .RSTB(I485907), .Q(I485869) );
DFFARX1 I_28446  ( .D(I702503), .CLK(I2702), .RSTB(I485907), .Q(I486311) );
nand I_28447 (I486328,I486311,I486023);
and I_28448 (I486345,I486006,I486328);
DFFARX1 I_28449  ( .D(I486345), .CLK(I2702), .RSTB(I485907), .Q(I485899) );
nor I_28450 (I485896,I486311,I486218);
and I_28451 (I486390,I486311,I486153);
or I_28452 (I486407,I486006,I486390);
DFFARX1 I_28453  ( .D(I486407), .CLK(I2702), .RSTB(I485907), .Q(I485884) );
nand I_28454 (I485893,I486311,I486235);
not I_28455 (I486485,I2709);
nand I_28456 (I486502,I416237,I416267);
and I_28457 (I486519,I486502,I416264);
DFFARX1 I_28458  ( .D(I486519), .CLK(I2702), .RSTB(I486485), .Q(I486536) );
not I_28459 (I486553,I486536);
DFFARX1 I_28460  ( .D(I486536), .CLK(I2702), .RSTB(I486485), .Q(I486453) );
nor I_28461 (I486584,I416255,I416267);
DFFARX1 I_28462  ( .D(I416243), .CLK(I2702), .RSTB(I486485), .Q(I486601) );
DFFARX1 I_28463  ( .D(I486601), .CLK(I2702), .RSTB(I486485), .Q(I486618) );
not I_28464 (I486456,I486618);
DFFARX1 I_28465  ( .D(I486601), .CLK(I2702), .RSTB(I486485), .Q(I486649) );
and I_28466 (I486450,I486536,I486649);
nand I_28467 (I486680,I416246,I416252);
and I_28468 (I486697,I486680,I416258);
DFFARX1 I_28469  ( .D(I486697), .CLK(I2702), .RSTB(I486485), .Q(I486714) );
nor I_28470 (I486731,I486714,I486553);
not I_28471 (I486748,I486714);
nand I_28472 (I486459,I486536,I486748);
DFFARX1 I_28473  ( .D(I416249), .CLK(I2702), .RSTB(I486485), .Q(I486779) );
and I_28474 (I486796,I486779,I416240);
nor I_28475 (I486813,I486796,I486714);
nor I_28476 (I486830,I486796,I486748);
nand I_28477 (I486465,I486584,I486830);
not I_28478 (I486468,I486796);
DFFARX1 I_28479  ( .D(I486796), .CLK(I2702), .RSTB(I486485), .Q(I486447) );
DFFARX1 I_28480  ( .D(I416261), .CLK(I2702), .RSTB(I486485), .Q(I486889) );
nand I_28481 (I486906,I486889,I486601);
and I_28482 (I486923,I486584,I486906);
DFFARX1 I_28483  ( .D(I486923), .CLK(I2702), .RSTB(I486485), .Q(I486477) );
nor I_28484 (I486474,I486889,I486796);
and I_28485 (I486968,I486889,I486731);
or I_28486 (I486985,I486584,I486968);
DFFARX1 I_28487  ( .D(I486985), .CLK(I2702), .RSTB(I486485), .Q(I486462) );
nand I_28488 (I486471,I486889,I486813);
not I_28489 (I487063,I2709);
or I_28490 (I487080,I311265,I311262);
or I_28491 (I487097,I311277,I311265);
nor I_28492 (I487114,I311292,I311268);
not I_28493 (I487131,I487114);
DFFARX1 I_28494  ( .D(I487114), .CLK(I2702), .RSTB(I487063), .Q(I487031) );
nand I_28495 (I487162,I487114,I487080);
not I_28496 (I487179,I311292);
and I_28497 (I487196,I487179,I311286);
nor I_28498 (I487213,I487196,I311262);
nor I_28499 (I487230,I311280,I311289);
DFFARX1 I_28500  ( .D(I487230), .CLK(I2702), .RSTB(I487063), .Q(I487247) );
nor I_28501 (I487264,I487247,I487131);
not I_28502 (I487281,I487247);
nand I_28503 (I487037,I487114,I487281);
DFFARX1 I_28504  ( .D(I487247), .CLK(I2702), .RSTB(I487063), .Q(I487028) );
nor I_28505 (I487326,I311280,I311277);
nand I_28506 (I487343,I487097,I487326);
nor I_28507 (I487052,I487080,I487326);
and I_28508 (I487374,I487326,I487264);
or I_28509 (I487391,I487213,I487374);
DFFARX1 I_28510  ( .D(I487391), .CLK(I2702), .RSTB(I487063), .Q(I487040) );
DFFARX1 I_28511  ( .D(I311274), .CLK(I2702), .RSTB(I487063), .Q(I487422) );
and I_28512 (I487439,I487422,I311271);
not I_28513 (I487046,I487439);
DFFARX1 I_28514  ( .D(I487439), .CLK(I2702), .RSTB(I487063), .Q(I487470) );
not I_28515 (I487034,I487470);
and I_28516 (I487501,I487439,I487162);
DFFARX1 I_28517  ( .D(I487501), .CLK(I2702), .RSTB(I487063), .Q(I487025) );
DFFARX1 I_28518  ( .D(I311283), .CLK(I2702), .RSTB(I487063), .Q(I487532) );
and I_28519 (I487549,I487532,I487343);
DFFARX1 I_28520  ( .D(I487549), .CLK(I2702), .RSTB(I487063), .Q(I487055) );
nor I_28521 (I487580,I487532,I487439);
nand I_28522 (I487049,I487213,I487580);
nor I_28523 (I487611,I487532,I487281);
nand I_28524 (I487043,I487097,I487611);
not I_28525 (I487675,I2709);
or I_28526 (I487692,I625653,I625647);
or I_28527 (I487709,I625656,I625653);
nor I_28528 (I487726,I625650,I625632);
not I_28529 (I487743,I487726);
DFFARX1 I_28530  ( .D(I487726), .CLK(I2702), .RSTB(I487675), .Q(I487643) );
nand I_28531 (I487774,I487726,I487692);
not I_28532 (I487791,I625650);
and I_28533 (I487808,I487791,I625629);
nor I_28534 (I487825,I487808,I625647);
nor I_28535 (I487842,I625644,I625626);
DFFARX1 I_28536  ( .D(I487842), .CLK(I2702), .RSTB(I487675), .Q(I487859) );
nor I_28537 (I487876,I487859,I487743);
not I_28538 (I487893,I487859);
nand I_28539 (I487649,I487726,I487893);
DFFARX1 I_28540  ( .D(I487859), .CLK(I2702), .RSTB(I487675), .Q(I487640) );
nor I_28541 (I487938,I625644,I625656);
nand I_28542 (I487955,I487709,I487938);
nor I_28543 (I487664,I487692,I487938);
and I_28544 (I487986,I487938,I487876);
or I_28545 (I488003,I487825,I487986);
DFFARX1 I_28546  ( .D(I488003), .CLK(I2702), .RSTB(I487675), .Q(I487652) );
DFFARX1 I_28547  ( .D(I625638), .CLK(I2702), .RSTB(I487675), .Q(I488034) );
and I_28548 (I488051,I488034,I625641);
not I_28549 (I487658,I488051);
DFFARX1 I_28550  ( .D(I488051), .CLK(I2702), .RSTB(I487675), .Q(I488082) );
not I_28551 (I487646,I488082);
and I_28552 (I488113,I488051,I487774);
DFFARX1 I_28553  ( .D(I488113), .CLK(I2702), .RSTB(I487675), .Q(I487637) );
DFFARX1 I_28554  ( .D(I625635), .CLK(I2702), .RSTB(I487675), .Q(I488144) );
and I_28555 (I488161,I488144,I487955);
DFFARX1 I_28556  ( .D(I488161), .CLK(I2702), .RSTB(I487675), .Q(I487667) );
nor I_28557 (I488192,I488144,I488051);
nand I_28558 (I487661,I487825,I488192);
nor I_28559 (I488223,I488144,I487893);
nand I_28560 (I487655,I487709,I488223);
not I_28561 (I488287,I2709);
or I_28562 (I488304,I312591,I312588);
or I_28563 (I488321,I312603,I312591);
nor I_28564 (I488338,I312618,I312594);
not I_28565 (I488355,I488338);
DFFARX1 I_28566  ( .D(I488338), .CLK(I2702), .RSTB(I488287), .Q(I488255) );
nand I_28567 (I488386,I488338,I488304);
not I_28568 (I488403,I312618);
and I_28569 (I488420,I488403,I312612);
nor I_28570 (I488437,I488420,I312588);
nor I_28571 (I488454,I312606,I312615);
DFFARX1 I_28572  ( .D(I488454), .CLK(I2702), .RSTB(I488287), .Q(I488471) );
nor I_28573 (I488488,I488471,I488355);
not I_28574 (I488505,I488471);
nand I_28575 (I488261,I488338,I488505);
DFFARX1 I_28576  ( .D(I488471), .CLK(I2702), .RSTB(I488287), .Q(I488252) );
nor I_28577 (I488550,I312606,I312603);
nand I_28578 (I488567,I488321,I488550);
nor I_28579 (I488276,I488304,I488550);
and I_28580 (I488598,I488550,I488488);
or I_28581 (I488615,I488437,I488598);
DFFARX1 I_28582  ( .D(I488615), .CLK(I2702), .RSTB(I488287), .Q(I488264) );
DFFARX1 I_28583  ( .D(I312600), .CLK(I2702), .RSTB(I488287), .Q(I488646) );
and I_28584 (I488663,I488646,I312597);
not I_28585 (I488270,I488663);
DFFARX1 I_28586  ( .D(I488663), .CLK(I2702), .RSTB(I488287), .Q(I488694) );
not I_28587 (I488258,I488694);
and I_28588 (I488725,I488663,I488386);
DFFARX1 I_28589  ( .D(I488725), .CLK(I2702), .RSTB(I488287), .Q(I488249) );
DFFARX1 I_28590  ( .D(I312609), .CLK(I2702), .RSTB(I488287), .Q(I488756) );
and I_28591 (I488773,I488756,I488567);
DFFARX1 I_28592  ( .D(I488773), .CLK(I2702), .RSTB(I488287), .Q(I488279) );
nor I_28593 (I488804,I488756,I488663);
nand I_28594 (I488273,I488437,I488804);
nor I_28595 (I488835,I488756,I488505);
nand I_28596 (I488267,I488321,I488835);
not I_28597 (I488899,I2709);
or I_28598 (I488916,I426050,I426035);
or I_28599 (I488933,I426047,I426050);
nor I_28600 (I488950,I426032,I426059);
not I_28601 (I488967,I488950);
DFFARX1 I_28602  ( .D(I488950), .CLK(I2702), .RSTB(I488899), .Q(I488867) );
nand I_28603 (I488998,I488950,I488916);
not I_28604 (I489015,I426032);
and I_28605 (I489032,I489015,I426053);
nor I_28606 (I489049,I489032,I426035);
nor I_28607 (I489066,I426056,I426029);
DFFARX1 I_28608  ( .D(I489066), .CLK(I2702), .RSTB(I488899), .Q(I489083) );
nor I_28609 (I489100,I489083,I488967);
not I_28610 (I489117,I489083);
nand I_28611 (I488873,I488950,I489117);
DFFARX1 I_28612  ( .D(I489083), .CLK(I2702), .RSTB(I488899), .Q(I488864) );
nor I_28613 (I489162,I426056,I426047);
nand I_28614 (I489179,I488933,I489162);
nor I_28615 (I488888,I488916,I489162);
and I_28616 (I489210,I489162,I489100);
or I_28617 (I489227,I489049,I489210);
DFFARX1 I_28618  ( .D(I489227), .CLK(I2702), .RSTB(I488899), .Q(I488876) );
DFFARX1 I_28619  ( .D(I426041), .CLK(I2702), .RSTB(I488899), .Q(I489258) );
and I_28620 (I489275,I489258,I426044);
not I_28621 (I488882,I489275);
DFFARX1 I_28622  ( .D(I489275), .CLK(I2702), .RSTB(I488899), .Q(I489306) );
not I_28623 (I488870,I489306);
and I_28624 (I489337,I489275,I488998);
DFFARX1 I_28625  ( .D(I489337), .CLK(I2702), .RSTB(I488899), .Q(I488861) );
DFFARX1 I_28626  ( .D(I426038), .CLK(I2702), .RSTB(I488899), .Q(I489368) );
and I_28627 (I489385,I489368,I489179);
DFFARX1 I_28628  ( .D(I489385), .CLK(I2702), .RSTB(I488899), .Q(I488891) );
nor I_28629 (I489416,I489368,I489275);
nand I_28630 (I488885,I489049,I489416);
nor I_28631 (I489447,I489368,I489117);
nand I_28632 (I488879,I488933,I489447);
not I_28633 (I489511,I2709);
or I_28634 (I489528,I560778,I560784);
or I_28635 (I489545,I560781,I560778);
nor I_28636 (I489562,I560754,I560772);
not I_28637 (I489579,I489562);
DFFARX1 I_28638  ( .D(I489562), .CLK(I2702), .RSTB(I489511), .Q(I489479) );
nand I_28639 (I489610,I489562,I489528);
not I_28640 (I489627,I560754);
and I_28641 (I489644,I489627,I560766);
nor I_28642 (I489661,I489644,I560784);
nor I_28643 (I489678,I560769,I560757);
DFFARX1 I_28644  ( .D(I489678), .CLK(I2702), .RSTB(I489511), .Q(I489695) );
nor I_28645 (I489712,I489695,I489579);
not I_28646 (I489729,I489695);
nand I_28647 (I489485,I489562,I489729);
DFFARX1 I_28648  ( .D(I489695), .CLK(I2702), .RSTB(I489511), .Q(I489476) );
nor I_28649 (I489774,I560769,I560781);
nand I_28650 (I489791,I489545,I489774);
nor I_28651 (I489500,I489528,I489774);
and I_28652 (I489822,I489774,I489712);
or I_28653 (I489839,I489661,I489822);
DFFARX1 I_28654  ( .D(I489839), .CLK(I2702), .RSTB(I489511), .Q(I489488) );
DFFARX1 I_28655  ( .D(I560760), .CLK(I2702), .RSTB(I489511), .Q(I489870) );
and I_28656 (I489887,I489870,I560775);
not I_28657 (I489494,I489887);
DFFARX1 I_28658  ( .D(I489887), .CLK(I2702), .RSTB(I489511), .Q(I489918) );
not I_28659 (I489482,I489918);
and I_28660 (I489949,I489887,I489610);
DFFARX1 I_28661  ( .D(I489949), .CLK(I2702), .RSTB(I489511), .Q(I489473) );
DFFARX1 I_28662  ( .D(I560763), .CLK(I2702), .RSTB(I489511), .Q(I489980) );
and I_28663 (I489997,I489980,I489791);
DFFARX1 I_28664  ( .D(I489997), .CLK(I2702), .RSTB(I489511), .Q(I489503) );
nor I_28665 (I490028,I489980,I489887);
nand I_28666 (I489497,I489661,I490028);
nor I_28667 (I490059,I489980,I489729);
nand I_28668 (I489491,I489545,I490059);
not I_28669 (I490123,I2709);
or I_28670 (I490140,I131817,I131808);
or I_28671 (I490157,I131805,I131817);
nor I_28672 (I490174,I131802,I131820);
not I_28673 (I490191,I490174);
DFFARX1 I_28674  ( .D(I490174), .CLK(I2702), .RSTB(I490123), .Q(I490091) );
nand I_28675 (I490222,I490174,I490140);
not I_28676 (I490239,I131802);
and I_28677 (I490256,I490239,I131793);
nor I_28678 (I490273,I490256,I131808);
nor I_28679 (I490290,I131796,I131799);
DFFARX1 I_28680  ( .D(I490290), .CLK(I2702), .RSTB(I490123), .Q(I490307) );
nor I_28681 (I490324,I490307,I490191);
not I_28682 (I490341,I490307);
nand I_28683 (I490097,I490174,I490341);
DFFARX1 I_28684  ( .D(I490307), .CLK(I2702), .RSTB(I490123), .Q(I490088) );
nor I_28685 (I490386,I131796,I131805);
nand I_28686 (I490403,I490157,I490386);
nor I_28687 (I490112,I490140,I490386);
and I_28688 (I490434,I490386,I490324);
or I_28689 (I490451,I490273,I490434);
DFFARX1 I_28690  ( .D(I490451), .CLK(I2702), .RSTB(I490123), .Q(I490100) );
DFFARX1 I_28691  ( .D(I131811), .CLK(I2702), .RSTB(I490123), .Q(I490482) );
and I_28692 (I490499,I490482,I131823);
not I_28693 (I490106,I490499);
DFFARX1 I_28694  ( .D(I490499), .CLK(I2702), .RSTB(I490123), .Q(I490530) );
not I_28695 (I490094,I490530);
and I_28696 (I490561,I490499,I490222);
DFFARX1 I_28697  ( .D(I490561), .CLK(I2702), .RSTB(I490123), .Q(I490085) );
DFFARX1 I_28698  ( .D(I131814), .CLK(I2702), .RSTB(I490123), .Q(I490592) );
and I_28699 (I490609,I490592,I490403);
DFFARX1 I_28700  ( .D(I490609), .CLK(I2702), .RSTB(I490123), .Q(I490115) );
nor I_28701 (I490640,I490592,I490499);
nand I_28702 (I490109,I490273,I490640);
nor I_28703 (I490671,I490592,I490341);
nand I_28704 (I490103,I490157,I490671);
not I_28705 (I490735,I2709);
or I_28706 (I490752,I704234,I704249);
or I_28707 (I490769,I704243,I704234);
nor I_28708 (I490786,I704240,I704237);
not I_28709 (I490803,I490786);
DFFARX1 I_28710  ( .D(I490786), .CLK(I2702), .RSTB(I490735), .Q(I490703) );
nand I_28711 (I490834,I490786,I490752);
not I_28712 (I490851,I704240);
and I_28713 (I490868,I490851,I704255);
nor I_28714 (I490885,I490868,I704249);
nor I_28715 (I490902,I704246,I704252);
DFFARX1 I_28716  ( .D(I490902), .CLK(I2702), .RSTB(I490735), .Q(I490919) );
nor I_28717 (I490936,I490919,I490803);
not I_28718 (I490953,I490919);
nand I_28719 (I490709,I490786,I490953);
DFFARX1 I_28720  ( .D(I490919), .CLK(I2702), .RSTB(I490735), .Q(I490700) );
nor I_28721 (I490998,I704246,I704243);
nand I_28722 (I491015,I490769,I490998);
nor I_28723 (I490724,I490752,I490998);
and I_28724 (I491046,I490998,I490936);
or I_28725 (I491063,I490885,I491046);
DFFARX1 I_28726  ( .D(I491063), .CLK(I2702), .RSTB(I490735), .Q(I490712) );
DFFARX1 I_28727  ( .D(I704264), .CLK(I2702), .RSTB(I490735), .Q(I491094) );
and I_28728 (I491111,I491094,I704261);
not I_28729 (I490718,I491111);
DFFARX1 I_28730  ( .D(I491111), .CLK(I2702), .RSTB(I490735), .Q(I491142) );
not I_28731 (I490706,I491142);
and I_28732 (I491173,I491111,I490834);
DFFARX1 I_28733  ( .D(I491173), .CLK(I2702), .RSTB(I490735), .Q(I490697) );
DFFARX1 I_28734  ( .D(I704258), .CLK(I2702), .RSTB(I490735), .Q(I491204) );
and I_28735 (I491221,I491204,I491015);
DFFARX1 I_28736  ( .D(I491221), .CLK(I2702), .RSTB(I490735), .Q(I490727) );
nor I_28737 (I491252,I491204,I491111);
nand I_28738 (I490721,I490885,I491252);
nor I_28739 (I491283,I491204,I490953);
nand I_28740 (I490715,I490769,I491283);
not I_28741 (I491347,I2709);
or I_28742 (I491364,I536383,I536389);
or I_28743 (I491381,I536386,I536383);
nor I_28744 (I491398,I536359,I536377);
not I_28745 (I491415,I491398);
DFFARX1 I_28746  ( .D(I491398), .CLK(I2702), .RSTB(I491347), .Q(I491315) );
nand I_28747 (I491446,I491398,I491364);
not I_28748 (I491463,I536359);
and I_28749 (I491480,I491463,I536371);
nor I_28750 (I491497,I491480,I536389);
nor I_28751 (I491514,I536374,I536362);
DFFARX1 I_28752  ( .D(I491514), .CLK(I2702), .RSTB(I491347), .Q(I491531) );
nor I_28753 (I491548,I491531,I491415);
not I_28754 (I491565,I491531);
nand I_28755 (I491321,I491398,I491565);
DFFARX1 I_28756  ( .D(I491531), .CLK(I2702), .RSTB(I491347), .Q(I491312) );
nor I_28757 (I491610,I536374,I536386);
nand I_28758 (I491627,I491381,I491610);
nor I_28759 (I491336,I491364,I491610);
and I_28760 (I491658,I491610,I491548);
or I_28761 (I491675,I491497,I491658);
DFFARX1 I_28762  ( .D(I491675), .CLK(I2702), .RSTB(I491347), .Q(I491324) );
DFFARX1 I_28763  ( .D(I536365), .CLK(I2702), .RSTB(I491347), .Q(I491706) );
and I_28764 (I491723,I491706,I536380);
not I_28765 (I491330,I491723);
DFFARX1 I_28766  ( .D(I491723), .CLK(I2702), .RSTB(I491347), .Q(I491754) );
not I_28767 (I491318,I491754);
and I_28768 (I491785,I491723,I491446);
DFFARX1 I_28769  ( .D(I491785), .CLK(I2702), .RSTB(I491347), .Q(I491309) );
DFFARX1 I_28770  ( .D(I536368), .CLK(I2702), .RSTB(I491347), .Q(I491816) );
and I_28771 (I491833,I491816,I491627);
DFFARX1 I_28772  ( .D(I491833), .CLK(I2702), .RSTB(I491347), .Q(I491339) );
nor I_28773 (I491864,I491816,I491723);
nand I_28774 (I491333,I491497,I491864);
nor I_28775 (I491895,I491816,I491565);
nand I_28776 (I491327,I491381,I491895);
not I_28777 (I491959,I2709);
or I_28778 (I491976,I714060,I714075);
or I_28779 (I491993,I714069,I714060);
nor I_28780 (I492010,I714066,I714063);
not I_28781 (I492027,I492010);
DFFARX1 I_28782  ( .D(I492010), .CLK(I2702), .RSTB(I491959), .Q(I491927) );
nand I_28783 (I492058,I492010,I491976);
not I_28784 (I492075,I714066);
and I_28785 (I492092,I492075,I714081);
nor I_28786 (I492109,I492092,I714075);
nor I_28787 (I492126,I714072,I714078);
DFFARX1 I_28788  ( .D(I492126), .CLK(I2702), .RSTB(I491959), .Q(I492143) );
nor I_28789 (I492160,I492143,I492027);
not I_28790 (I492177,I492143);
nand I_28791 (I491933,I492010,I492177);
DFFARX1 I_28792  ( .D(I492143), .CLK(I2702), .RSTB(I491959), .Q(I491924) );
nor I_28793 (I492222,I714072,I714069);
nand I_28794 (I492239,I491993,I492222);
nor I_28795 (I491948,I491976,I492222);
and I_28796 (I492270,I492222,I492160);
or I_28797 (I492287,I492109,I492270);
DFFARX1 I_28798  ( .D(I492287), .CLK(I2702), .RSTB(I491959), .Q(I491936) );
DFFARX1 I_28799  ( .D(I714090), .CLK(I2702), .RSTB(I491959), .Q(I492318) );
and I_28800 (I492335,I492318,I714087);
not I_28801 (I491942,I492335);
DFFARX1 I_28802  ( .D(I492335), .CLK(I2702), .RSTB(I491959), .Q(I492366) );
not I_28803 (I491930,I492366);
and I_28804 (I492397,I492335,I492058);
DFFARX1 I_28805  ( .D(I492397), .CLK(I2702), .RSTB(I491959), .Q(I491921) );
DFFARX1 I_28806  ( .D(I714084), .CLK(I2702), .RSTB(I491959), .Q(I492428) );
and I_28807 (I492445,I492428,I492239);
DFFARX1 I_28808  ( .D(I492445), .CLK(I2702), .RSTB(I491959), .Q(I491951) );
nor I_28809 (I492476,I492428,I492335);
nand I_28810 (I491945,I492109,I492476);
nor I_28811 (I492507,I492428,I492177);
nand I_28812 (I491939,I491993,I492507);
not I_28813 (I492571,I2709);
or I_28814 (I492588,I498510,I498489);
or I_28815 (I492605,I498492,I498510);
nor I_28816 (I492622,I498486,I498498);
not I_28817 (I492639,I492622);
DFFARX1 I_28818  ( .D(I492622), .CLK(I2702), .RSTB(I492571), .Q(I492539) );
nand I_28819 (I492670,I492622,I492588);
not I_28820 (I492687,I498486);
and I_28821 (I492704,I492687,I498495);
nor I_28822 (I492721,I492704,I498489);
nor I_28823 (I492738,I498507,I498513);
DFFARX1 I_28824  ( .D(I492738), .CLK(I2702), .RSTB(I492571), .Q(I492755) );
nor I_28825 (I492772,I492755,I492639);
not I_28826 (I492789,I492755);
nand I_28827 (I492545,I492622,I492789);
DFFARX1 I_28828  ( .D(I492755), .CLK(I2702), .RSTB(I492571), .Q(I492536) );
nor I_28829 (I492834,I498507,I498492);
nand I_28830 (I492851,I492605,I492834);
nor I_28831 (I492560,I492588,I492834);
and I_28832 (I492882,I492834,I492772);
or I_28833 (I492899,I492721,I492882);
DFFARX1 I_28834  ( .D(I492899), .CLK(I2702), .RSTB(I492571), .Q(I492548) );
DFFARX1 I_28835  ( .D(I498483), .CLK(I2702), .RSTB(I492571), .Q(I492930) );
and I_28836 (I492947,I492930,I498501);
not I_28837 (I492554,I492947);
DFFARX1 I_28838  ( .D(I492947), .CLK(I2702), .RSTB(I492571), .Q(I492978) );
not I_28839 (I492542,I492978);
and I_28840 (I493009,I492947,I492670);
DFFARX1 I_28841  ( .D(I493009), .CLK(I2702), .RSTB(I492571), .Q(I492533) );
DFFARX1 I_28842  ( .D(I498504), .CLK(I2702), .RSTB(I492571), .Q(I493040) );
and I_28843 (I493057,I493040,I492851);
DFFARX1 I_28844  ( .D(I493057), .CLK(I2702), .RSTB(I492571), .Q(I492563) );
nor I_28845 (I493088,I493040,I492947);
nand I_28846 (I492557,I492721,I493088);
nor I_28847 (I493119,I493040,I492789);
nand I_28848 (I492551,I492605,I493119);
not I_28849 (I493183,I2709);
or I_28850 (I493200,I411974,I411959);
or I_28851 (I493217,I411971,I411974);
nor I_28852 (I493234,I411956,I411983);
not I_28853 (I493251,I493234);
DFFARX1 I_28854  ( .D(I493234), .CLK(I2702), .RSTB(I493183), .Q(I493151) );
nand I_28855 (I493282,I493234,I493200);
not I_28856 (I493299,I411956);
and I_28857 (I493316,I493299,I411977);
nor I_28858 (I493333,I493316,I411959);
nor I_28859 (I493350,I411980,I411953);
DFFARX1 I_28860  ( .D(I493350), .CLK(I2702), .RSTB(I493183), .Q(I493367) );
nor I_28861 (I493384,I493367,I493251);
not I_28862 (I493401,I493367);
nand I_28863 (I493157,I493234,I493401);
DFFARX1 I_28864  ( .D(I493367), .CLK(I2702), .RSTB(I493183), .Q(I493148) );
nor I_28865 (I493446,I411980,I411971);
nand I_28866 (I493463,I493217,I493446);
nor I_28867 (I493172,I493200,I493446);
and I_28868 (I493494,I493446,I493384);
or I_28869 (I493511,I493333,I493494);
DFFARX1 I_28870  ( .D(I493511), .CLK(I2702), .RSTB(I493183), .Q(I493160) );
DFFARX1 I_28871  ( .D(I411965), .CLK(I2702), .RSTB(I493183), .Q(I493542) );
and I_28872 (I493559,I493542,I411968);
not I_28873 (I493166,I493559);
DFFARX1 I_28874  ( .D(I493559), .CLK(I2702), .RSTB(I493183), .Q(I493590) );
not I_28875 (I493154,I493590);
and I_28876 (I493621,I493559,I493282);
DFFARX1 I_28877  ( .D(I493621), .CLK(I2702), .RSTB(I493183), .Q(I493145) );
DFFARX1 I_28878  ( .D(I411962), .CLK(I2702), .RSTB(I493183), .Q(I493652) );
and I_28879 (I493669,I493652,I493463);
DFFARX1 I_28880  ( .D(I493669), .CLK(I2702), .RSTB(I493183), .Q(I493175) );
nor I_28881 (I493700,I493652,I493559);
nand I_28882 (I493169,I493333,I493700);
nor I_28883 (I493731,I493652,I493401);
nand I_28884 (I493163,I493217,I493731);
not I_28885 (I493795,I2709);
or I_28886 (I493812,I258225,I258222);
or I_28887 (I493829,I258237,I258225);
nor I_28888 (I493846,I258252,I258228);
not I_28889 (I493863,I493846);
DFFARX1 I_28890  ( .D(I493846), .CLK(I2702), .RSTB(I493795), .Q(I493763) );
nand I_28891 (I493894,I493846,I493812);
not I_28892 (I493911,I258252);
and I_28893 (I493928,I493911,I258246);
nor I_28894 (I493945,I493928,I258222);
nor I_28895 (I493962,I258240,I258249);
DFFARX1 I_28896  ( .D(I493962), .CLK(I2702), .RSTB(I493795), .Q(I493979) );
nor I_28897 (I493996,I493979,I493863);
not I_28898 (I494013,I493979);
nand I_28899 (I493769,I493846,I494013);
DFFARX1 I_28900  ( .D(I493979), .CLK(I2702), .RSTB(I493795), .Q(I493760) );
nor I_28901 (I494058,I258240,I258237);
nand I_28902 (I494075,I493829,I494058);
nor I_28903 (I493784,I493812,I494058);
and I_28904 (I494106,I494058,I493996);
or I_28905 (I494123,I493945,I494106);
DFFARX1 I_28906  ( .D(I494123), .CLK(I2702), .RSTB(I493795), .Q(I493772) );
DFFARX1 I_28907  ( .D(I258234), .CLK(I2702), .RSTB(I493795), .Q(I494154) );
and I_28908 (I494171,I494154,I258231);
not I_28909 (I493778,I494171);
DFFARX1 I_28910  ( .D(I494171), .CLK(I2702), .RSTB(I493795), .Q(I494202) );
not I_28911 (I493766,I494202);
and I_28912 (I494233,I494171,I493894);
DFFARX1 I_28913  ( .D(I494233), .CLK(I2702), .RSTB(I493795), .Q(I493757) );
DFFARX1 I_28914  ( .D(I258243), .CLK(I2702), .RSTB(I493795), .Q(I494264) );
and I_28915 (I494281,I494264,I494075);
DFFARX1 I_28916  ( .D(I494281), .CLK(I2702), .RSTB(I493795), .Q(I493787) );
nor I_28917 (I494312,I494264,I494171);
nand I_28918 (I493781,I493945,I494312);
nor I_28919 (I494343,I494264,I494013);
nand I_28920 (I493775,I493829,I494343);
not I_28921 (I494407,I2709);
or I_28922 (I494424,I418706,I418691);
or I_28923 (I494441,I418703,I418706);
nor I_28924 (I494458,I418688,I418715);
not I_28925 (I494475,I494458);
DFFARX1 I_28926  ( .D(I494458), .CLK(I2702), .RSTB(I494407), .Q(I494375) );
nand I_28927 (I494506,I494458,I494424);
not I_28928 (I494523,I418688);
and I_28929 (I494540,I494523,I418709);
nor I_28930 (I494557,I494540,I418691);
nor I_28931 (I494574,I418712,I418685);
DFFARX1 I_28932  ( .D(I494574), .CLK(I2702), .RSTB(I494407), .Q(I494591) );
nor I_28933 (I494608,I494591,I494475);
not I_28934 (I494625,I494591);
nand I_28935 (I494381,I494458,I494625);
DFFARX1 I_28936  ( .D(I494591), .CLK(I2702), .RSTB(I494407), .Q(I494372) );
nor I_28937 (I494670,I418712,I418703);
nand I_28938 (I494687,I494441,I494670);
nor I_28939 (I494396,I494424,I494670);
and I_28940 (I494718,I494670,I494608);
or I_28941 (I494735,I494557,I494718);
DFFARX1 I_28942  ( .D(I494735), .CLK(I2702), .RSTB(I494407), .Q(I494384) );
DFFARX1 I_28943  ( .D(I418697), .CLK(I2702), .RSTB(I494407), .Q(I494766) );
and I_28944 (I494783,I494766,I418700);
not I_28945 (I494390,I494783);
DFFARX1 I_28946  ( .D(I494783), .CLK(I2702), .RSTB(I494407), .Q(I494814) );
not I_28947 (I494378,I494814);
and I_28948 (I494845,I494783,I494506);
DFFARX1 I_28949  ( .D(I494845), .CLK(I2702), .RSTB(I494407), .Q(I494369) );
DFFARX1 I_28950  ( .D(I418694), .CLK(I2702), .RSTB(I494407), .Q(I494876) );
and I_28951 (I494893,I494876,I494687);
DFFARX1 I_28952  ( .D(I494893), .CLK(I2702), .RSTB(I494407), .Q(I494399) );
nor I_28953 (I494924,I494876,I494783);
nand I_28954 (I494393,I494557,I494924);
nor I_28955 (I494955,I494876,I494625);
nand I_28956 (I494387,I494441,I494955);
not I_28957 (I495019,I2709);
or I_28958 (I495036,I277452,I277449);
or I_28959 (I495053,I277464,I277452);
nor I_28960 (I495070,I277479,I277455);
not I_28961 (I495087,I495070);
DFFARX1 I_28962  ( .D(I495070), .CLK(I2702), .RSTB(I495019), .Q(I494987) );
nand I_28963 (I495118,I495070,I495036);
not I_28964 (I495135,I277479);
and I_28965 (I495152,I495135,I277473);
nor I_28966 (I495169,I495152,I277449);
nor I_28967 (I495186,I277467,I277476);
DFFARX1 I_28968  ( .D(I495186), .CLK(I2702), .RSTB(I495019), .Q(I495203) );
nor I_28969 (I495220,I495203,I495087);
not I_28970 (I495237,I495203);
nand I_28971 (I494993,I495070,I495237);
DFFARX1 I_28972  ( .D(I495203), .CLK(I2702), .RSTB(I495019), .Q(I494984) );
nor I_28973 (I495282,I277467,I277464);
nand I_28974 (I495299,I495053,I495282);
nor I_28975 (I495008,I495036,I495282);
and I_28976 (I495330,I495282,I495220);
or I_28977 (I495347,I495169,I495330);
DFFARX1 I_28978  ( .D(I495347), .CLK(I2702), .RSTB(I495019), .Q(I494996) );
DFFARX1 I_28979  ( .D(I277461), .CLK(I2702), .RSTB(I495019), .Q(I495378) );
and I_28980 (I495395,I495378,I277458);
not I_28981 (I495002,I495395);
DFFARX1 I_28982  ( .D(I495395), .CLK(I2702), .RSTB(I495019), .Q(I495426) );
not I_28983 (I494990,I495426);
and I_28984 (I495457,I495395,I495118);
DFFARX1 I_28985  ( .D(I495457), .CLK(I2702), .RSTB(I495019), .Q(I494981) );
DFFARX1 I_28986  ( .D(I277470), .CLK(I2702), .RSTB(I495019), .Q(I495488) );
and I_28987 (I495505,I495488,I495299);
DFFARX1 I_28988  ( .D(I495505), .CLK(I2702), .RSTB(I495019), .Q(I495011) );
nor I_28989 (I495536,I495488,I495395);
nand I_28990 (I495005,I495169,I495536);
nor I_28991 (I495567,I495488,I495237);
nand I_28992 (I494999,I495053,I495567);
not I_28993 (I495631,I2709);
or I_28994 (I495648,I36393,I36387);
or I_28995 (I495665,I36375,I36393);
nor I_28996 (I495682,I36402,I36396);
or I_28997 (I495620,I495682,I495648);
not I_28998 (I495713,I36402);
and I_28999 (I495730,I495713,I36378);
nor I_29000 (I495747,I495730,I36387);
not I_29001 (I495764,I495747);
nor I_29002 (I495781,I36372,I36399);
DFFARX1 I_29003  ( .D(I495781), .CLK(I2702), .RSTB(I495631), .Q(I495798) );
nor I_29004 (I495815,I495798,I495747);
nand I_29005 (I495605,I495648,I495815);
nor I_29006 (I495846,I495798,I495764);
not I_29007 (I495602,I495798);
nor I_29008 (I495877,I36372,I36375);
or I_29009 (I495614,I495648,I495877);
DFFARX1 I_29010  ( .D(I36381), .CLK(I2702), .RSTB(I495631), .Q(I495908) );
and I_29011 (I495925,I495908,I36390);
nor I_29012 (I495942,I495925,I495798);
DFFARX1 I_29013  ( .D(I495942), .CLK(I2702), .RSTB(I495631), .Q(I495608) );
nor I_29014 (I495623,I495925,I495877);
not I_29015 (I495987,I495925);
nor I_29016 (I496004,I495665,I495987);
nand I_29017 (I495593,I495925,I495764);
DFFARX1 I_29018  ( .D(I36384), .CLK(I2702), .RSTB(I495631), .Q(I496035) );
nor I_29019 (I495611,I496035,I495665);
not I_29020 (I496066,I496035);
and I_29021 (I496083,I495877,I496066);
nor I_29022 (I495617,I495682,I496083);
and I_29023 (I496114,I496035,I496004);
or I_29024 (I496131,I495682,I496114);
DFFARX1 I_29025  ( .D(I496131), .CLK(I2702), .RSTB(I495631), .Q(I495596) );
nand I_29026 (I495599,I496035,I495846);
not I_29027 (I496209,I2709);
or I_29028 (I496226,I604210,I604207);
or I_29029 (I496243,I604195,I604210);
nor I_29030 (I496260,I604189,I604216);
or I_29031 (I496198,I496260,I496226);
not I_29032 (I496291,I604189);
and I_29033 (I496308,I496291,I604201);
nor I_29034 (I496325,I496308,I604207);
not I_29035 (I496342,I496325);
nor I_29036 (I496359,I604192,I604213);
DFFARX1 I_29037  ( .D(I496359), .CLK(I2702), .RSTB(I496209), .Q(I496376) );
nor I_29038 (I496393,I496376,I496325);
nand I_29039 (I496183,I496226,I496393);
nor I_29040 (I496424,I496376,I496342);
not I_29041 (I496180,I496376);
nor I_29042 (I496455,I604192,I604195);
or I_29043 (I496192,I496226,I496455);
DFFARX1 I_29044  ( .D(I604204), .CLK(I2702), .RSTB(I496209), .Q(I496486) );
and I_29045 (I496503,I496486,I604198);
nor I_29046 (I496520,I496503,I496376);
DFFARX1 I_29047  ( .D(I496520), .CLK(I2702), .RSTB(I496209), .Q(I496186) );
nor I_29048 (I496201,I496503,I496455);
not I_29049 (I496565,I496503);
nor I_29050 (I496582,I496243,I496565);
nand I_29051 (I496171,I496503,I496342);
DFFARX1 I_29052  ( .D(I604219), .CLK(I2702), .RSTB(I496209), .Q(I496613) );
nor I_29053 (I496189,I496613,I496243);
not I_29054 (I496644,I496613);
and I_29055 (I496661,I496455,I496644);
nor I_29056 (I496195,I496260,I496661);
and I_29057 (I496692,I496613,I496582);
or I_29058 (I496709,I496260,I496692);
DFFARX1 I_29059  ( .D(I496709), .CLK(I2702), .RSTB(I496209), .Q(I496174) );
nand I_29060 (I496177,I496613,I496424);
not I_29061 (I496787,I2709);
or I_29062 (I496804,I669659,I669662);
or I_29063 (I496821,I669680,I669659);
nor I_29064 (I496838,I669674,I669683);
or I_29065 (I496776,I496838,I496804);
not I_29066 (I496869,I669674);
and I_29067 (I496886,I496869,I669686);
nor I_29068 (I496903,I496886,I669662);
not I_29069 (I496920,I496903);
nor I_29070 (I496937,I669671,I669656);
DFFARX1 I_29071  ( .D(I496937), .CLK(I2702), .RSTB(I496787), .Q(I496954) );
nor I_29072 (I496971,I496954,I496903);
nand I_29073 (I496761,I496804,I496971);
nor I_29074 (I497002,I496954,I496920);
not I_29075 (I496758,I496954);
nor I_29076 (I497033,I669671,I669680);
or I_29077 (I496770,I496804,I497033);
DFFARX1 I_29078  ( .D(I669668), .CLK(I2702), .RSTB(I496787), .Q(I497064) );
and I_29079 (I497081,I497064,I669677);
nor I_29080 (I497098,I497081,I496954);
DFFARX1 I_29081  ( .D(I497098), .CLK(I2702), .RSTB(I496787), .Q(I496764) );
nor I_29082 (I496779,I497081,I497033);
not I_29083 (I497143,I497081);
nor I_29084 (I497160,I496821,I497143);
nand I_29085 (I496749,I497081,I496920);
DFFARX1 I_29086  ( .D(I669665), .CLK(I2702), .RSTB(I496787), .Q(I497191) );
nor I_29087 (I496767,I497191,I496821);
not I_29088 (I497222,I497191);
and I_29089 (I497239,I497033,I497222);
nor I_29090 (I496773,I496838,I497239);
and I_29091 (I497270,I497191,I497160);
or I_29092 (I497287,I496838,I497270);
DFFARX1 I_29093  ( .D(I497287), .CLK(I2702), .RSTB(I496787), .Q(I496752) );
nand I_29094 (I496755,I497191,I497002);
not I_29095 (I497365,I2709);
or I_29096 (I497382,I349321,I349306);
or I_29097 (I497399,I349315,I349321);
nor I_29098 (I497416,I349309,I349297);
or I_29099 (I497354,I497416,I497382);
not I_29100 (I497447,I349309);
and I_29101 (I497464,I497447,I349318);
nor I_29102 (I497481,I497464,I349306);
not I_29103 (I497498,I497481);
nor I_29104 (I497515,I349303,I349294);
DFFARX1 I_29105  ( .D(I497515), .CLK(I2702), .RSTB(I497365), .Q(I497532) );
nor I_29106 (I497549,I497532,I497481);
nand I_29107 (I497339,I497382,I497549);
nor I_29108 (I497580,I497532,I497498);
not I_29109 (I497336,I497532);
nor I_29110 (I497611,I349303,I349315);
or I_29111 (I497348,I497382,I497611);
DFFARX1 I_29112  ( .D(I349312), .CLK(I2702), .RSTB(I497365), .Q(I497642) );
and I_29113 (I497659,I497642,I349291);
nor I_29114 (I497676,I497659,I497532);
DFFARX1 I_29115  ( .D(I497676), .CLK(I2702), .RSTB(I497365), .Q(I497342) );
nor I_29116 (I497357,I497659,I497611);
not I_29117 (I497721,I497659);
nor I_29118 (I497738,I497399,I497721);
nand I_29119 (I497327,I497659,I497498);
DFFARX1 I_29120  ( .D(I349300), .CLK(I2702), .RSTB(I497365), .Q(I497769) );
nor I_29121 (I497345,I497769,I497399);
not I_29122 (I497800,I497769);
and I_29123 (I497817,I497611,I497800);
nor I_29124 (I497351,I497416,I497817);
and I_29125 (I497848,I497769,I497738);
or I_29126 (I497865,I497416,I497848);
DFFARX1 I_29127  ( .D(I497865), .CLK(I2702), .RSTB(I497365), .Q(I497330) );
nand I_29128 (I497333,I497769,I497580);
not I_29129 (I497943,I2709);
or I_29130 (I497960,I364825,I364810);
or I_29131 (I497977,I364819,I364825);
nor I_29132 (I497994,I364813,I364801);
or I_29133 (I497932,I497994,I497960);
not I_29134 (I498025,I364813);
and I_29135 (I498042,I498025,I364822);
nor I_29136 (I498059,I498042,I364810);
not I_29137 (I498076,I498059);
nor I_29138 (I498093,I364807,I364798);
DFFARX1 I_29139  ( .D(I498093), .CLK(I2702), .RSTB(I497943), .Q(I498110) );
nor I_29140 (I498127,I498110,I498059);
nand I_29141 (I497917,I497960,I498127);
nor I_29142 (I498158,I498110,I498076);
not I_29143 (I497914,I498110);
nor I_29144 (I498189,I364807,I364819);
or I_29145 (I497926,I497960,I498189);
DFFARX1 I_29146  ( .D(I364816), .CLK(I2702), .RSTB(I497943), .Q(I498220) );
and I_29147 (I498237,I498220,I364795);
nor I_29148 (I498254,I498237,I498110);
DFFARX1 I_29149  ( .D(I498254), .CLK(I2702), .RSTB(I497943), .Q(I497920) );
nor I_29150 (I497935,I498237,I498189);
not I_29151 (I498299,I498237);
nor I_29152 (I498316,I497977,I498299);
nand I_29153 (I497905,I498237,I498076);
DFFARX1 I_29154  ( .D(I364804), .CLK(I2702), .RSTB(I497943), .Q(I498347) );
nor I_29155 (I497923,I498347,I497977);
not I_29156 (I498378,I498347);
and I_29157 (I498395,I498189,I498378);
nor I_29158 (I497929,I497994,I498395);
and I_29159 (I498426,I498347,I498316);
or I_29160 (I498443,I497994,I498426);
DFFARX1 I_29161  ( .D(I498443), .CLK(I2702), .RSTB(I497943), .Q(I497908) );
nand I_29162 (I497911,I498347,I498158);
not I_29163 (I498521,I2709);
or I_29164 (I498538,I234992,I235010);
or I_29165 (I498555,I235007,I234992);
nor I_29166 (I498572,I234986,I234983);
or I_29167 (I498510,I498572,I498538);
not I_29168 (I498603,I234986);
and I_29169 (I498620,I498603,I234989);
nor I_29170 (I498637,I498620,I235010);
not I_29171 (I498654,I498637);
nor I_29172 (I498671,I235013,I235001);
DFFARX1 I_29173  ( .D(I498671), .CLK(I2702), .RSTB(I498521), .Q(I498688) );
nor I_29174 (I498705,I498688,I498637);
nand I_29175 (I498495,I498538,I498705);
nor I_29176 (I498736,I498688,I498654);
not I_29177 (I498492,I498688);
nor I_29178 (I498767,I235013,I235007);
or I_29179 (I498504,I498538,I498767);
DFFARX1 I_29180  ( .D(I234998), .CLK(I2702), .RSTB(I498521), .Q(I498798) );
and I_29181 (I498815,I498798,I235004);
nor I_29182 (I498832,I498815,I498688);
DFFARX1 I_29183  ( .D(I498832), .CLK(I2702), .RSTB(I498521), .Q(I498498) );
nor I_29184 (I498513,I498815,I498767);
not I_29185 (I498877,I498815);
nor I_29186 (I498894,I498555,I498877);
nand I_29187 (I498483,I498815,I498654);
DFFARX1 I_29188  ( .D(I234995), .CLK(I2702), .RSTB(I498521), .Q(I498925) );
nor I_29189 (I498501,I498925,I498555);
not I_29190 (I498956,I498925);
and I_29191 (I498973,I498767,I498956);
nor I_29192 (I498507,I498572,I498973);
and I_29193 (I499004,I498925,I498894);
or I_29194 (I499021,I498572,I499004);
DFFARX1 I_29195  ( .D(I499021), .CLK(I2702), .RSTB(I498521), .Q(I498486) );
nand I_29196 (I498489,I498925,I498736);
not I_29197 (I499099,I2709);
or I_29198 (I499116,I549470,I549464);
or I_29199 (I499133,I549458,I549470);
nor I_29200 (I499150,I549479,I549467);
or I_29201 (I499088,I499150,I499116);
not I_29202 (I499181,I549479);
and I_29203 (I499198,I499181,I549452);
nor I_29204 (I499215,I499198,I549464);
not I_29205 (I499232,I499215);
nor I_29206 (I499249,I549455,I549449);
DFFARX1 I_29207  ( .D(I499249), .CLK(I2702), .RSTB(I499099), .Q(I499266) );
nor I_29208 (I499283,I499266,I499215);
nand I_29209 (I499073,I499116,I499283);
nor I_29210 (I499314,I499266,I499232);
not I_29211 (I499070,I499266);
nor I_29212 (I499345,I549455,I549458);
or I_29213 (I499082,I499116,I499345);
DFFARX1 I_29214  ( .D(I549476), .CLK(I2702), .RSTB(I499099), .Q(I499376) );
and I_29215 (I499393,I499376,I549473);
nor I_29216 (I499410,I499393,I499266);
DFFARX1 I_29217  ( .D(I499410), .CLK(I2702), .RSTB(I499099), .Q(I499076) );
nor I_29218 (I499091,I499393,I499345);
not I_29219 (I499455,I499393);
nor I_29220 (I499472,I499133,I499455);
nand I_29221 (I499061,I499393,I499232);
DFFARX1 I_29222  ( .D(I549461), .CLK(I2702), .RSTB(I499099), .Q(I499503) );
nor I_29223 (I499079,I499503,I499133);
not I_29224 (I499534,I499503);
and I_29225 (I499551,I499345,I499534);
nor I_29226 (I499085,I499150,I499551);
and I_29227 (I499582,I499503,I499472);
or I_29228 (I499599,I499150,I499582);
DFFARX1 I_29229  ( .D(I499599), .CLK(I2702), .RSTB(I499099), .Q(I499064) );
nand I_29230 (I499067,I499503,I499314);
not I_29231 (I499677,I2709);
or I_29232 (I499694,I429722,I429713);
or I_29233 (I499711,I429707,I429722);
nor I_29234 (I499728,I429704,I429728);
or I_29235 (I499666,I499728,I499694);
not I_29236 (I499759,I429704);
and I_29237 (I499776,I499759,I429719);
nor I_29238 (I499793,I499776,I429713);
not I_29239 (I499810,I499793);
nor I_29240 (I499827,I429701,I429731);
DFFARX1 I_29241  ( .D(I499827), .CLK(I2702), .RSTB(I499677), .Q(I499844) );
nor I_29242 (I499861,I499844,I499793);
nand I_29243 (I499651,I499694,I499861);
nor I_29244 (I499892,I499844,I499810);
not I_29245 (I499648,I499844);
nor I_29246 (I499923,I429701,I429707);
or I_29247 (I499660,I499694,I499923);
DFFARX1 I_29248  ( .D(I429710), .CLK(I2702), .RSTB(I499677), .Q(I499954) );
and I_29249 (I499971,I499954,I429716);
nor I_29250 (I499988,I499971,I499844);
DFFARX1 I_29251  ( .D(I499988), .CLK(I2702), .RSTB(I499677), .Q(I499654) );
nor I_29252 (I499669,I499971,I499923);
not I_29253 (I500033,I499971);
nor I_29254 (I500050,I499711,I500033);
nand I_29255 (I499639,I499971,I499810);
DFFARX1 I_29256  ( .D(I429725), .CLK(I2702), .RSTB(I499677), .Q(I500081) );
nor I_29257 (I499657,I500081,I499711);
not I_29258 (I500112,I500081);
and I_29259 (I500129,I499923,I500112);
nor I_29260 (I499663,I499728,I500129);
and I_29261 (I500160,I500081,I500050);
or I_29262 (I500177,I499728,I500160);
DFFARX1 I_29263  ( .D(I500177), .CLK(I2702), .RSTB(I499677), .Q(I499642) );
nand I_29264 (I499645,I500081,I499892);
not I_29265 (I500255,I2709);
or I_29266 (I500272,I650160,I650163);
or I_29267 (I500289,I650181,I650160);
nor I_29268 (I500306,I650175,I650184);
or I_29269 (I500244,I500306,I500272);
not I_29270 (I500337,I650175);
and I_29271 (I500354,I500337,I650187);
nor I_29272 (I500371,I500354,I650163);
not I_29273 (I500388,I500371);
nor I_29274 (I500405,I650172,I650157);
DFFARX1 I_29275  ( .D(I500405), .CLK(I2702), .RSTB(I500255), .Q(I500422) );
nor I_29276 (I500439,I500422,I500371);
nand I_29277 (I500229,I500272,I500439);
nor I_29278 (I500470,I500422,I500388);
not I_29279 (I500226,I500422);
nor I_29280 (I500501,I650172,I650181);
or I_29281 (I500238,I500272,I500501);
DFFARX1 I_29282  ( .D(I650169), .CLK(I2702), .RSTB(I500255), .Q(I500532) );
and I_29283 (I500549,I500532,I650178);
nor I_29284 (I500566,I500549,I500422);
DFFARX1 I_29285  ( .D(I500566), .CLK(I2702), .RSTB(I500255), .Q(I500232) );
nor I_29286 (I500247,I500549,I500501);
not I_29287 (I500611,I500549);
nor I_29288 (I500628,I500289,I500611);
nand I_29289 (I500217,I500549,I500388);
DFFARX1 I_29290  ( .D(I650166), .CLK(I2702), .RSTB(I500255), .Q(I500659) );
nor I_29291 (I500235,I500659,I500289);
not I_29292 (I500690,I500659);
and I_29293 (I500707,I500501,I500690);
nor I_29294 (I500241,I500306,I500707);
and I_29295 (I500738,I500659,I500628);
or I_29296 (I500755,I500306,I500738);
DFFARX1 I_29297  ( .D(I500755), .CLK(I2702), .RSTB(I500255), .Q(I500220) );
nand I_29298 (I500223,I500659,I500470);
not I_29299 (I500833,I2709);
or I_29300 (I500850,I342861,I342846);
or I_29301 (I500867,I342855,I342861);
nor I_29302 (I500884,I342849,I342837);
or I_29303 (I500822,I500884,I500850);
not I_29304 (I500915,I342849);
and I_29305 (I500932,I500915,I342858);
nor I_29306 (I500949,I500932,I342846);
not I_29307 (I500966,I500949);
nor I_29308 (I500983,I342843,I342834);
DFFARX1 I_29309  ( .D(I500983), .CLK(I2702), .RSTB(I500833), .Q(I501000) );
nor I_29310 (I501017,I501000,I500949);
nand I_29311 (I500807,I500850,I501017);
nor I_29312 (I501048,I501000,I500966);
not I_29313 (I500804,I501000);
nor I_29314 (I501079,I342843,I342855);
or I_29315 (I500816,I500850,I501079);
DFFARX1 I_29316  ( .D(I342852), .CLK(I2702), .RSTB(I500833), .Q(I501110) );
and I_29317 (I501127,I501110,I342831);
nor I_29318 (I501144,I501127,I501000);
DFFARX1 I_29319  ( .D(I501144), .CLK(I2702), .RSTB(I500833), .Q(I500810) );
nor I_29320 (I500825,I501127,I501079);
not I_29321 (I501189,I501127);
nor I_29322 (I501206,I500867,I501189);
nand I_29323 (I500795,I501127,I500966);
DFFARX1 I_29324  ( .D(I342840), .CLK(I2702), .RSTB(I500833), .Q(I501237) );
nor I_29325 (I500813,I501237,I500867);
not I_29326 (I501268,I501237);
and I_29327 (I501285,I501079,I501268);
nor I_29328 (I500819,I500884,I501285);
and I_29329 (I501316,I501237,I501206);
or I_29330 (I501333,I500884,I501316);
DFFARX1 I_29331  ( .D(I501333), .CLK(I2702), .RSTB(I500833), .Q(I500798) );
nand I_29332 (I500801,I501237,I501048);
not I_29333 (I501411,I2709);
or I_29334 (I501428,I161451,I161439);
or I_29335 (I501445,I161424,I161451);
nor I_29336 (I501462,I161436,I161433);
or I_29337 (I501400,I501462,I501428);
not I_29338 (I501493,I161436);
and I_29339 (I501510,I501493,I161448);
nor I_29340 (I501527,I501510,I161439);
not I_29341 (I501544,I501527);
nor I_29342 (I501561,I161430,I161445);
DFFARX1 I_29343  ( .D(I501561), .CLK(I2702), .RSTB(I501411), .Q(I501578) );
nor I_29344 (I501595,I501578,I501527);
nand I_29345 (I501385,I501428,I501595);
nor I_29346 (I501626,I501578,I501544);
not I_29347 (I501382,I501578);
nor I_29348 (I501657,I161430,I161424);
or I_29349 (I501394,I501428,I501657);
DFFARX1 I_29350  ( .D(I161454), .CLK(I2702), .RSTB(I501411), .Q(I501688) );
and I_29351 (I501705,I501688,I161427);
nor I_29352 (I501722,I501705,I501578);
DFFARX1 I_29353  ( .D(I501722), .CLK(I2702), .RSTB(I501411), .Q(I501388) );
nor I_29354 (I501403,I501705,I501657);
not I_29355 (I501767,I501705);
nor I_29356 (I501784,I501445,I501767);
nand I_29357 (I501373,I501705,I501544);
DFFARX1 I_29358  ( .D(I161442), .CLK(I2702), .RSTB(I501411), .Q(I501815) );
nor I_29359 (I501391,I501815,I501445);
not I_29360 (I501846,I501815);
and I_29361 (I501863,I501657,I501846);
nor I_29362 (I501397,I501462,I501863);
and I_29363 (I501894,I501815,I501784);
or I_29364 (I501911,I501462,I501894);
DFFARX1 I_29365  ( .D(I501911), .CLK(I2702), .RSTB(I501411), .Q(I501376) );
nand I_29366 (I501379,I501815,I501626);
not I_29367 (I501989,I2709);
or I_29368 (I502006,I638209,I638212);
or I_29369 (I502023,I638230,I638209);
nor I_29370 (I502040,I638224,I638233);
or I_29371 (I501978,I502040,I502006);
not I_29372 (I502071,I638224);
and I_29373 (I502088,I502071,I638236);
nor I_29374 (I502105,I502088,I638212);
not I_29375 (I502122,I502105);
nor I_29376 (I502139,I638221,I638206);
DFFARX1 I_29377  ( .D(I502139), .CLK(I2702), .RSTB(I501989), .Q(I502156) );
nor I_29378 (I502173,I502156,I502105);
nand I_29379 (I501963,I502006,I502173);
nor I_29380 (I502204,I502156,I502122);
not I_29381 (I501960,I502156);
nor I_29382 (I502235,I638221,I638230);
or I_29383 (I501972,I502006,I502235);
DFFARX1 I_29384  ( .D(I638218), .CLK(I2702), .RSTB(I501989), .Q(I502266) );
and I_29385 (I502283,I502266,I638227);
nor I_29386 (I502300,I502283,I502156);
DFFARX1 I_29387  ( .D(I502300), .CLK(I2702), .RSTB(I501989), .Q(I501966) );
nor I_29388 (I501981,I502283,I502235);
not I_29389 (I502345,I502283);
nor I_29390 (I502362,I502023,I502345);
nand I_29391 (I501951,I502283,I502122);
DFFARX1 I_29392  ( .D(I638215), .CLK(I2702), .RSTB(I501989), .Q(I502393) );
nor I_29393 (I501969,I502393,I502023);
not I_29394 (I502424,I502393);
and I_29395 (I502441,I502235,I502424);
nor I_29396 (I501975,I502040,I502441);
and I_29397 (I502472,I502393,I502362);
or I_29398 (I502489,I502040,I502472);
DFFARX1 I_29399  ( .D(I502489), .CLK(I2702), .RSTB(I501989), .Q(I501954) );
nand I_29400 (I501957,I502393,I502204);
not I_29401 (I502567,I2709);
or I_29402 (I502584,I287403,I287397);
or I_29403 (I502601,I287415,I287403);
nor I_29404 (I502618,I287394,I287421);
or I_29405 (I502556,I502618,I502584);
not I_29406 (I502649,I287394);
and I_29407 (I502666,I502649,I287418);
nor I_29408 (I502683,I502666,I287397);
not I_29409 (I502700,I502683);
nor I_29410 (I502717,I287409,I287424);
DFFARX1 I_29411  ( .D(I502717), .CLK(I2702), .RSTB(I502567), .Q(I502734) );
nor I_29412 (I502751,I502734,I502683);
nand I_29413 (I502541,I502584,I502751);
nor I_29414 (I502782,I502734,I502700);
not I_29415 (I502538,I502734);
nor I_29416 (I502813,I287409,I287415);
or I_29417 (I502550,I502584,I502813);
DFFARX1 I_29418  ( .D(I287406), .CLK(I2702), .RSTB(I502567), .Q(I502844) );
and I_29419 (I502861,I502844,I287412);
nor I_29420 (I502878,I502861,I502734);
DFFARX1 I_29421  ( .D(I502878), .CLK(I2702), .RSTB(I502567), .Q(I502544) );
nor I_29422 (I502559,I502861,I502813);
not I_29423 (I502923,I502861);
nor I_29424 (I502940,I502601,I502923);
nand I_29425 (I502529,I502861,I502700);
DFFARX1 I_29426  ( .D(I287400), .CLK(I2702), .RSTB(I502567), .Q(I502971) );
nor I_29427 (I502547,I502971,I502601);
not I_29428 (I503002,I502971);
and I_29429 (I503019,I502813,I503002);
nor I_29430 (I502553,I502618,I503019);
and I_29431 (I503050,I502971,I502940);
or I_29432 (I503067,I502618,I503050);
DFFARX1 I_29433  ( .D(I503067), .CLK(I2702), .RSTB(I502567), .Q(I502532) );
nand I_29434 (I502535,I502971,I502782);
not I_29435 (I503145,I2709);
or I_29436 (I503162,I180015,I180003);
or I_29437 (I503179,I179988,I180015);
nor I_29438 (I503196,I180000,I179997);
or I_29439 (I503134,I503196,I503162);
not I_29440 (I503227,I180000);
and I_29441 (I503244,I503227,I180012);
nor I_29442 (I503261,I503244,I180003);
not I_29443 (I503278,I503261);
nor I_29444 (I503295,I179994,I180009);
DFFARX1 I_29445  ( .D(I503295), .CLK(I2702), .RSTB(I503145), .Q(I503312) );
nor I_29446 (I503329,I503312,I503261);
nand I_29447 (I503119,I503162,I503329);
nor I_29448 (I503360,I503312,I503278);
not I_29449 (I503116,I503312);
nor I_29450 (I503391,I179994,I179988);
or I_29451 (I503128,I503162,I503391);
DFFARX1 I_29452  ( .D(I180018), .CLK(I2702), .RSTB(I503145), .Q(I503422) );
and I_29453 (I503439,I503422,I179991);
nor I_29454 (I503456,I503439,I503312);
DFFARX1 I_29455  ( .D(I503456), .CLK(I2702), .RSTB(I503145), .Q(I503122) );
nor I_29456 (I503137,I503439,I503391);
not I_29457 (I503501,I503439);
nor I_29458 (I503518,I503179,I503501);
nand I_29459 (I503107,I503439,I503278);
DFFARX1 I_29460  ( .D(I180006), .CLK(I2702), .RSTB(I503145), .Q(I503549) );
nor I_29461 (I503125,I503549,I503179);
not I_29462 (I503580,I503549);
and I_29463 (I503597,I503391,I503580);
nor I_29464 (I503131,I503196,I503597);
and I_29465 (I503628,I503549,I503518);
or I_29466 (I503645,I503196,I503628);
DFFARX1 I_29467  ( .D(I503645), .CLK(I2702), .RSTB(I503145), .Q(I503110) );
nand I_29468 (I503113,I503549,I503360);
not I_29469 (I503723,I2709);
or I_29470 (I503740,I433879,I433852);
or I_29471 (I503757,I433849,I433879);
nor I_29472 (I503774,I433861,I433873);
or I_29473 (I503712,I503774,I503740);
not I_29474 (I503805,I433861);
and I_29475 (I503822,I503805,I433867);
nor I_29476 (I503839,I503822,I433852);
not I_29477 (I503856,I503839);
nor I_29478 (I503873,I433855,I433876);
DFFARX1 I_29479  ( .D(I503873), .CLK(I2702), .RSTB(I503723), .Q(I503890) );
nor I_29480 (I503907,I503890,I503839);
nand I_29481 (I503697,I503740,I503907);
nor I_29482 (I503938,I503890,I503856);
not I_29483 (I503694,I503890);
nor I_29484 (I503969,I433855,I433849);
or I_29485 (I503706,I503740,I503969);
DFFARX1 I_29486  ( .D(I433870), .CLK(I2702), .RSTB(I503723), .Q(I504000) );
and I_29487 (I504017,I504000,I433858);
nor I_29488 (I504034,I504017,I503890);
DFFARX1 I_29489  ( .D(I504034), .CLK(I2702), .RSTB(I503723), .Q(I503700) );
nor I_29490 (I503715,I504017,I503969);
not I_29491 (I504079,I504017);
nor I_29492 (I504096,I503757,I504079);
nand I_29493 (I503685,I504017,I503856);
DFFARX1 I_29494  ( .D(I433864), .CLK(I2702), .RSTB(I503723), .Q(I504127) );
nor I_29495 (I503703,I504127,I503757);
not I_29496 (I504158,I504127);
and I_29497 (I504175,I503969,I504158);
nor I_29498 (I503709,I503774,I504175);
and I_29499 (I504206,I504127,I504096);
or I_29500 (I504223,I503774,I504206);
DFFARX1 I_29501  ( .D(I504223), .CLK(I2702), .RSTB(I503723), .Q(I503688) );
nand I_29502 (I503691,I504127,I503938);
not I_29503 (I504301,I2709);
or I_29504 (I504318,I249612,I249606);
or I_29505 (I504335,I249624,I249612);
nor I_29506 (I504352,I249603,I249630);
or I_29507 (I504290,I504352,I504318);
not I_29508 (I504383,I249603);
and I_29509 (I504400,I504383,I249627);
nor I_29510 (I504417,I504400,I249606);
not I_29511 (I504434,I504417);
nor I_29512 (I504451,I249618,I249633);
DFFARX1 I_29513  ( .D(I504451), .CLK(I2702), .RSTB(I504301), .Q(I504468) );
nor I_29514 (I504485,I504468,I504417);
nand I_29515 (I504275,I504318,I504485);
nor I_29516 (I504516,I504468,I504434);
not I_29517 (I504272,I504468);
nor I_29518 (I504547,I249618,I249624);
or I_29519 (I504284,I504318,I504547);
DFFARX1 I_29520  ( .D(I249615), .CLK(I2702), .RSTB(I504301), .Q(I504578) );
and I_29521 (I504595,I504578,I249621);
nor I_29522 (I504612,I504595,I504468);
DFFARX1 I_29523  ( .D(I504612), .CLK(I2702), .RSTB(I504301), .Q(I504278) );
nor I_29524 (I504293,I504595,I504547);
not I_29525 (I504657,I504595);
nor I_29526 (I504674,I504335,I504657);
nand I_29527 (I504263,I504595,I504434);
DFFARX1 I_29528  ( .D(I249609), .CLK(I2702), .RSTB(I504301), .Q(I504705) );
nor I_29529 (I504281,I504705,I504335);
not I_29530 (I504736,I504705);
and I_29531 (I504753,I504547,I504736);
nor I_29532 (I504287,I504352,I504753);
and I_29533 (I504784,I504705,I504674);
or I_29534 (I504801,I504352,I504784);
DFFARX1 I_29535  ( .D(I504801), .CLK(I2702), .RSTB(I504301), .Q(I504266) );
nand I_29536 (I504269,I504705,I504516);
not I_29537 (I504879,I2709);
or I_29538 (I504896,I422378,I422369);
or I_29539 (I504913,I422363,I422378);
nor I_29540 (I504930,I422360,I422384);
or I_29541 (I504868,I504930,I504896);
not I_29542 (I504961,I422360);
and I_29543 (I504978,I504961,I422375);
nor I_29544 (I504995,I504978,I422369);
not I_29545 (I505012,I504995);
nor I_29546 (I505029,I422357,I422387);
DFFARX1 I_29547  ( .D(I505029), .CLK(I2702), .RSTB(I504879), .Q(I505046) );
nor I_29548 (I505063,I505046,I504995);
nand I_29549 (I504853,I504896,I505063);
nor I_29550 (I505094,I505046,I505012);
not I_29551 (I504850,I505046);
nor I_29552 (I505125,I422357,I422363);
or I_29553 (I504862,I504896,I505125);
DFFARX1 I_29554  ( .D(I422366), .CLK(I2702), .RSTB(I504879), .Q(I505156) );
and I_29555 (I505173,I505156,I422372);
nor I_29556 (I505190,I505173,I505046);
DFFARX1 I_29557  ( .D(I505190), .CLK(I2702), .RSTB(I504879), .Q(I504856) );
nor I_29558 (I504871,I505173,I505125);
not I_29559 (I505235,I505173);
nor I_29560 (I505252,I504913,I505235);
nand I_29561 (I504841,I505173,I505012);
DFFARX1 I_29562  ( .D(I422381), .CLK(I2702), .RSTB(I504879), .Q(I505283) );
nor I_29563 (I504859,I505283,I504913);
not I_29564 (I505314,I505283);
and I_29565 (I505331,I505125,I505314);
nor I_29566 (I504865,I504930,I505331);
and I_29567 (I505362,I505283,I505252);
or I_29568 (I505379,I504930,I505362);
DFFARX1 I_29569  ( .D(I505379), .CLK(I2702), .RSTB(I504879), .Q(I504844) );
nand I_29570 (I504847,I505283,I505094);
not I_29571 (I505457,I2709);
nand I_29572 (I505474,I6081,I6087);
and I_29573 (I505491,I505474,I6084);
DFFARX1 I_29574  ( .D(I505491), .CLK(I2702), .RSTB(I505457), .Q(I505508) );
nor I_29575 (I505525,I6108,I6087);
nor I_29576 (I505542,I505525,I505508);
not I_29577 (I505440,I505525);
DFFARX1 I_29578  ( .D(I6099), .CLK(I2702), .RSTB(I505457), .Q(I505573) );
not I_29579 (I505590,I505573);
nor I_29580 (I505607,I505525,I505590);
nand I_29581 (I505443,I505573,I505542);
DFFARX1 I_29582  ( .D(I505573), .CLK(I2702), .RSTB(I505457), .Q(I505425) );
nand I_29583 (I505652,I6102,I6105);
and I_29584 (I505669,I505652,I6078);
DFFARX1 I_29585  ( .D(I505669), .CLK(I2702), .RSTB(I505457), .Q(I505686) );
nor I_29586 (I505446,I505686,I505508);
nand I_29587 (I505437,I505686,I505607);
DFFARX1 I_29588  ( .D(I6096), .CLK(I2702), .RSTB(I505457), .Q(I505731) );
and I_29589 (I505748,I505731,I6090);
DFFARX1 I_29590  ( .D(I505748), .CLK(I2702), .RSTB(I505457), .Q(I505765) );
not I_29591 (I505428,I505765);
nand I_29592 (I505796,I505748,I505686);
and I_29593 (I505813,I505508,I505796);
DFFARX1 I_29594  ( .D(I505813), .CLK(I2702), .RSTB(I505457), .Q(I505419) );
DFFARX1 I_29595  ( .D(I6093), .CLK(I2702), .RSTB(I505457), .Q(I505844) );
nand I_29596 (I505861,I505844,I505508);
and I_29597 (I505878,I505686,I505861);
DFFARX1 I_29598  ( .D(I505878), .CLK(I2702), .RSTB(I505457), .Q(I505449) );
not I_29599 (I505909,I505844);
nor I_29600 (I505926,I505525,I505909);
and I_29601 (I505943,I505844,I505926);
or I_29602 (I505960,I505748,I505943);
DFFARX1 I_29603  ( .D(I505960), .CLK(I2702), .RSTB(I505457), .Q(I505434) );
nand I_29604 (I505431,I505844,I505590);
DFFARX1 I_29605  ( .D(I505844), .CLK(I2702), .RSTB(I505457), .Q(I505422) );
not I_29606 (I506052,I2709);
nand I_29607 (I506069,I236182,I236185);
and I_29608 (I506086,I506069,I236176);
DFFARX1 I_29609  ( .D(I506086), .CLK(I2702), .RSTB(I506052), .Q(I506103) );
nor I_29610 (I506120,I236200,I236185);
nor I_29611 (I506137,I506120,I506103);
not I_29612 (I506035,I506120);
DFFARX1 I_29613  ( .D(I236179), .CLK(I2702), .RSTB(I506052), .Q(I506168) );
not I_29614 (I506185,I506168);
nor I_29615 (I506202,I506120,I506185);
nand I_29616 (I506038,I506168,I506137);
DFFARX1 I_29617  ( .D(I506168), .CLK(I2702), .RSTB(I506052), .Q(I506020) );
nand I_29618 (I506247,I236197,I236188);
and I_29619 (I506264,I506247,I236173);
DFFARX1 I_29620  ( .D(I506264), .CLK(I2702), .RSTB(I506052), .Q(I506281) );
nor I_29621 (I506041,I506281,I506103);
nand I_29622 (I506032,I506281,I506202);
DFFARX1 I_29623  ( .D(I236203), .CLK(I2702), .RSTB(I506052), .Q(I506326) );
and I_29624 (I506343,I506326,I236194);
DFFARX1 I_29625  ( .D(I506343), .CLK(I2702), .RSTB(I506052), .Q(I506360) );
not I_29626 (I506023,I506360);
nand I_29627 (I506391,I506343,I506281);
and I_29628 (I506408,I506103,I506391);
DFFARX1 I_29629  ( .D(I506408), .CLK(I2702), .RSTB(I506052), .Q(I506014) );
DFFARX1 I_29630  ( .D(I236191), .CLK(I2702), .RSTB(I506052), .Q(I506439) );
nand I_29631 (I506456,I506439,I506103);
and I_29632 (I506473,I506281,I506456);
DFFARX1 I_29633  ( .D(I506473), .CLK(I2702), .RSTB(I506052), .Q(I506044) );
not I_29634 (I506504,I506439);
nor I_29635 (I506521,I506120,I506504);
and I_29636 (I506538,I506439,I506521);
or I_29637 (I506555,I506343,I506538);
DFFARX1 I_29638  ( .D(I506555), .CLK(I2702), .RSTB(I506052), .Q(I506029) );
nand I_29639 (I506026,I506439,I506185);
DFFARX1 I_29640  ( .D(I506439), .CLK(I2702), .RSTB(I506052), .Q(I506017) );
not I_29641 (I506647,I2709);
nand I_29642 (I506664,I395175,I395187);
and I_29643 (I506681,I506664,I395169);
DFFARX1 I_29644  ( .D(I506681), .CLK(I2702), .RSTB(I506647), .Q(I506698) );
nor I_29645 (I506715,I395181,I395187);
nor I_29646 (I506732,I506715,I506698);
not I_29647 (I506630,I506715);
DFFARX1 I_29648  ( .D(I395166), .CLK(I2702), .RSTB(I506647), .Q(I506763) );
not I_29649 (I506780,I506763);
nor I_29650 (I506797,I506715,I506780);
nand I_29651 (I506633,I506763,I506732);
DFFARX1 I_29652  ( .D(I506763), .CLK(I2702), .RSTB(I506647), .Q(I506615) );
nand I_29653 (I506842,I395157,I395172);
and I_29654 (I506859,I506842,I395163);
DFFARX1 I_29655  ( .D(I506859), .CLK(I2702), .RSTB(I506647), .Q(I506876) );
nor I_29656 (I506636,I506876,I506698);
nand I_29657 (I506627,I506876,I506797);
DFFARX1 I_29658  ( .D(I395184), .CLK(I2702), .RSTB(I506647), .Q(I506921) );
and I_29659 (I506938,I506921,I395178);
DFFARX1 I_29660  ( .D(I506938), .CLK(I2702), .RSTB(I506647), .Q(I506955) );
not I_29661 (I506618,I506955);
nand I_29662 (I506986,I506938,I506876);
and I_29663 (I507003,I506698,I506986);
DFFARX1 I_29664  ( .D(I507003), .CLK(I2702), .RSTB(I506647), .Q(I506609) );
DFFARX1 I_29665  ( .D(I395160), .CLK(I2702), .RSTB(I506647), .Q(I507034) );
nand I_29666 (I507051,I507034,I506698);
and I_29667 (I507068,I506876,I507051);
DFFARX1 I_29668  ( .D(I507068), .CLK(I2702), .RSTB(I506647), .Q(I506639) );
not I_29669 (I507099,I507034);
nor I_29670 (I507116,I506715,I507099);
and I_29671 (I507133,I507034,I507116);
or I_29672 (I507150,I506938,I507133);
DFFARX1 I_29673  ( .D(I507150), .CLK(I2702), .RSTB(I506647), .Q(I506624) );
nand I_29674 (I506621,I507034,I506780);
DFFARX1 I_29675  ( .D(I507034), .CLK(I2702), .RSTB(I506647), .Q(I506612) );
not I_29676 (I507242,I2709);
nand I_29677 (I507259,I397113,I397125);
and I_29678 (I507276,I507259,I397107);
DFFARX1 I_29679  ( .D(I507276), .CLK(I2702), .RSTB(I507242), .Q(I507293) );
nor I_29680 (I507310,I397119,I397125);
nor I_29681 (I507327,I507310,I507293);
not I_29682 (I507225,I507310);
DFFARX1 I_29683  ( .D(I397104), .CLK(I2702), .RSTB(I507242), .Q(I507358) );
not I_29684 (I507375,I507358);
nor I_29685 (I507392,I507310,I507375);
nand I_29686 (I507228,I507358,I507327);
DFFARX1 I_29687  ( .D(I507358), .CLK(I2702), .RSTB(I507242), .Q(I507210) );
nand I_29688 (I507437,I397095,I397110);
and I_29689 (I507454,I507437,I397101);
DFFARX1 I_29690  ( .D(I507454), .CLK(I2702), .RSTB(I507242), .Q(I507471) );
nor I_29691 (I507231,I507471,I507293);
nand I_29692 (I507222,I507471,I507392);
DFFARX1 I_29693  ( .D(I397122), .CLK(I2702), .RSTB(I507242), .Q(I507516) );
and I_29694 (I507533,I507516,I397116);
DFFARX1 I_29695  ( .D(I507533), .CLK(I2702), .RSTB(I507242), .Q(I507550) );
not I_29696 (I507213,I507550);
nand I_29697 (I507581,I507533,I507471);
and I_29698 (I507598,I507293,I507581);
DFFARX1 I_29699  ( .D(I507598), .CLK(I2702), .RSTB(I507242), .Q(I507204) );
DFFARX1 I_29700  ( .D(I397098), .CLK(I2702), .RSTB(I507242), .Q(I507629) );
nand I_29701 (I507646,I507629,I507293);
and I_29702 (I507663,I507471,I507646);
DFFARX1 I_29703  ( .D(I507663), .CLK(I2702), .RSTB(I507242), .Q(I507234) );
not I_29704 (I507694,I507629);
nor I_29705 (I507711,I507310,I507694);
and I_29706 (I507728,I507629,I507711);
or I_29707 (I507745,I507533,I507728);
DFFARX1 I_29708  ( .D(I507745), .CLK(I2702), .RSTB(I507242), .Q(I507219) );
nand I_29709 (I507216,I507629,I507375);
DFFARX1 I_29710  ( .D(I507629), .CLK(I2702), .RSTB(I507242), .Q(I507207) );
not I_29711 (I507837,I2709);
nand I_29712 (I507854,I335743,I335755);
and I_29713 (I507871,I507854,I335737);
DFFARX1 I_29714  ( .D(I507871), .CLK(I2702), .RSTB(I507837), .Q(I507888) );
nor I_29715 (I507905,I335749,I335755);
nor I_29716 (I507922,I507905,I507888);
not I_29717 (I507820,I507905);
DFFARX1 I_29718  ( .D(I335734), .CLK(I2702), .RSTB(I507837), .Q(I507953) );
not I_29719 (I507970,I507953);
nor I_29720 (I507987,I507905,I507970);
nand I_29721 (I507823,I507953,I507922);
DFFARX1 I_29722  ( .D(I507953), .CLK(I2702), .RSTB(I507837), .Q(I507805) );
nand I_29723 (I508032,I335725,I335740);
and I_29724 (I508049,I508032,I335731);
DFFARX1 I_29725  ( .D(I508049), .CLK(I2702), .RSTB(I507837), .Q(I508066) );
nor I_29726 (I507826,I508066,I507888);
nand I_29727 (I507817,I508066,I507987);
DFFARX1 I_29728  ( .D(I335752), .CLK(I2702), .RSTB(I507837), .Q(I508111) );
and I_29729 (I508128,I508111,I335746);
DFFARX1 I_29730  ( .D(I508128), .CLK(I2702), .RSTB(I507837), .Q(I508145) );
not I_29731 (I507808,I508145);
nand I_29732 (I508176,I508128,I508066);
and I_29733 (I508193,I507888,I508176);
DFFARX1 I_29734  ( .D(I508193), .CLK(I2702), .RSTB(I507837), .Q(I507799) );
DFFARX1 I_29735  ( .D(I335728), .CLK(I2702), .RSTB(I507837), .Q(I508224) );
nand I_29736 (I508241,I508224,I507888);
and I_29737 (I508258,I508066,I508241);
DFFARX1 I_29738  ( .D(I508258), .CLK(I2702), .RSTB(I507837), .Q(I507829) );
not I_29739 (I508289,I508224);
nor I_29740 (I508306,I507905,I508289);
and I_29741 (I508323,I508224,I508306);
or I_29742 (I508340,I508128,I508323);
DFFARX1 I_29743  ( .D(I508340), .CLK(I2702), .RSTB(I507837), .Q(I507814) );
nand I_29744 (I507811,I508224,I507970);
DFFARX1 I_29745  ( .D(I508224), .CLK(I2702), .RSTB(I507837), .Q(I507802) );
not I_29746 (I508432,I2709);
nand I_29747 (I508449,I406157,I406169);
and I_29748 (I508466,I508449,I406151);
DFFARX1 I_29749  ( .D(I508466), .CLK(I2702), .RSTB(I508432), .Q(I508483) );
nor I_29750 (I508500,I406163,I406169);
nor I_29751 (I508517,I508500,I508483);
not I_29752 (I508415,I508500);
DFFARX1 I_29753  ( .D(I406148), .CLK(I2702), .RSTB(I508432), .Q(I508548) );
not I_29754 (I508565,I508548);
nor I_29755 (I508582,I508500,I508565);
nand I_29756 (I508418,I508548,I508517);
DFFARX1 I_29757  ( .D(I508548), .CLK(I2702), .RSTB(I508432), .Q(I508400) );
nand I_29758 (I508627,I406139,I406154);
and I_29759 (I508644,I508627,I406145);
DFFARX1 I_29760  ( .D(I508644), .CLK(I2702), .RSTB(I508432), .Q(I508661) );
nor I_29761 (I508421,I508661,I508483);
nand I_29762 (I508412,I508661,I508582);
DFFARX1 I_29763  ( .D(I406166), .CLK(I2702), .RSTB(I508432), .Q(I508706) );
and I_29764 (I508723,I508706,I406160);
DFFARX1 I_29765  ( .D(I508723), .CLK(I2702), .RSTB(I508432), .Q(I508740) );
not I_29766 (I508403,I508740);
nand I_29767 (I508771,I508723,I508661);
and I_29768 (I508788,I508483,I508771);
DFFARX1 I_29769  ( .D(I508788), .CLK(I2702), .RSTB(I508432), .Q(I508394) );
DFFARX1 I_29770  ( .D(I406142), .CLK(I2702), .RSTB(I508432), .Q(I508819) );
nand I_29771 (I508836,I508819,I508483);
and I_29772 (I508853,I508661,I508836);
DFFARX1 I_29773  ( .D(I508853), .CLK(I2702), .RSTB(I508432), .Q(I508424) );
not I_29774 (I508884,I508819);
nor I_29775 (I508901,I508500,I508884);
and I_29776 (I508918,I508819,I508901);
or I_29777 (I508935,I508723,I508918);
DFFARX1 I_29778  ( .D(I508935), .CLK(I2702), .RSTB(I508432), .Q(I508409) );
nand I_29779 (I508406,I508819,I508565);
DFFARX1 I_29780  ( .D(I508819), .CLK(I2702), .RSTB(I508432), .Q(I508397) );
not I_29781 (I509027,I2709);
nand I_29782 (I509044,I614951,I614942);
and I_29783 (I509061,I509044,I614960);
DFFARX1 I_29784  ( .D(I509061), .CLK(I2702), .RSTB(I509027), .Q(I509078) );
nor I_29785 (I509095,I614957,I614942);
nor I_29786 (I509112,I509095,I509078);
not I_29787 (I509010,I509095);
DFFARX1 I_29788  ( .D(I614939), .CLK(I2702), .RSTB(I509027), .Q(I509143) );
not I_29789 (I509160,I509143);
nor I_29790 (I509177,I509095,I509160);
nand I_29791 (I509013,I509143,I509112);
DFFARX1 I_29792  ( .D(I509143), .CLK(I2702), .RSTB(I509027), .Q(I508995) );
nand I_29793 (I509222,I614948,I614963);
and I_29794 (I509239,I509222,I614954);
DFFARX1 I_29795  ( .D(I509239), .CLK(I2702), .RSTB(I509027), .Q(I509256) );
nor I_29796 (I509016,I509256,I509078);
nand I_29797 (I509007,I509256,I509177);
DFFARX1 I_29798  ( .D(I614936), .CLK(I2702), .RSTB(I509027), .Q(I509301) );
and I_29799 (I509318,I509301,I614945);
DFFARX1 I_29800  ( .D(I509318), .CLK(I2702), .RSTB(I509027), .Q(I509335) );
not I_29801 (I508998,I509335);
nand I_29802 (I509366,I509318,I509256);
and I_29803 (I509383,I509078,I509366);
DFFARX1 I_29804  ( .D(I509383), .CLK(I2702), .RSTB(I509027), .Q(I508989) );
DFFARX1 I_29805  ( .D(I614933), .CLK(I2702), .RSTB(I509027), .Q(I509414) );
nand I_29806 (I509431,I509414,I509078);
and I_29807 (I509448,I509256,I509431);
DFFARX1 I_29808  ( .D(I509448), .CLK(I2702), .RSTB(I509027), .Q(I509019) );
not I_29809 (I509479,I509414);
nor I_29810 (I509496,I509095,I509479);
and I_29811 (I509513,I509414,I509496);
or I_29812 (I509530,I509318,I509513);
DFFARX1 I_29813  ( .D(I509530), .CLK(I2702), .RSTB(I509027), .Q(I509004) );
nand I_29814 (I509001,I509414,I509160);
DFFARX1 I_29815  ( .D(I509414), .CLK(I2702), .RSTB(I509027), .Q(I508992) );
not I_29816 (I509622,I2709);
nand I_29817 (I509639,I38058,I38064);
and I_29818 (I509656,I509639,I38061);
DFFARX1 I_29819  ( .D(I509656), .CLK(I2702), .RSTB(I509622), .Q(I509673) );
nor I_29820 (I509690,I38085,I38064);
nor I_29821 (I509707,I509690,I509673);
not I_29822 (I509605,I509690);
DFFARX1 I_29823  ( .D(I38076), .CLK(I2702), .RSTB(I509622), .Q(I509738) );
not I_29824 (I509755,I509738);
nor I_29825 (I509772,I509690,I509755);
nand I_29826 (I509608,I509738,I509707);
DFFARX1 I_29827  ( .D(I509738), .CLK(I2702), .RSTB(I509622), .Q(I509590) );
nand I_29828 (I509817,I38079,I38082);
and I_29829 (I509834,I509817,I38055);
DFFARX1 I_29830  ( .D(I509834), .CLK(I2702), .RSTB(I509622), .Q(I509851) );
nor I_29831 (I509611,I509851,I509673);
nand I_29832 (I509602,I509851,I509772);
DFFARX1 I_29833  ( .D(I38073), .CLK(I2702), .RSTB(I509622), .Q(I509896) );
and I_29834 (I509913,I509896,I38067);
DFFARX1 I_29835  ( .D(I509913), .CLK(I2702), .RSTB(I509622), .Q(I509930) );
not I_29836 (I509593,I509930);
nand I_29837 (I509961,I509913,I509851);
and I_29838 (I509978,I509673,I509961);
DFFARX1 I_29839  ( .D(I509978), .CLK(I2702), .RSTB(I509622), .Q(I509584) );
DFFARX1 I_29840  ( .D(I38070), .CLK(I2702), .RSTB(I509622), .Q(I510009) );
nand I_29841 (I510026,I510009,I509673);
and I_29842 (I510043,I509851,I510026);
DFFARX1 I_29843  ( .D(I510043), .CLK(I2702), .RSTB(I509622), .Q(I509614) );
not I_29844 (I510074,I510009);
nor I_29845 (I510091,I509690,I510074);
and I_29846 (I510108,I510009,I510091);
or I_29847 (I510125,I509913,I510108);
DFFARX1 I_29848  ( .D(I510125), .CLK(I2702), .RSTB(I509622), .Q(I509599) );
nand I_29849 (I509596,I510009,I509755);
DFFARX1 I_29850  ( .D(I510009), .CLK(I2702), .RSTB(I509622), .Q(I509587) );
not I_29851 (I510217,I2709);
nand I_29852 (I510234,I333159,I333171);
and I_29853 (I510251,I510234,I333153);
DFFARX1 I_29854  ( .D(I510251), .CLK(I2702), .RSTB(I510217), .Q(I510268) );
nor I_29855 (I510285,I333165,I333171);
nor I_29856 (I510302,I510285,I510268);
not I_29857 (I510200,I510285);
DFFARX1 I_29858  ( .D(I333150), .CLK(I2702), .RSTB(I510217), .Q(I510333) );
not I_29859 (I510350,I510333);
nor I_29860 (I510367,I510285,I510350);
nand I_29861 (I510203,I510333,I510302);
DFFARX1 I_29862  ( .D(I510333), .CLK(I2702), .RSTB(I510217), .Q(I510185) );
nand I_29863 (I510412,I333141,I333156);
and I_29864 (I510429,I510412,I333147);
DFFARX1 I_29865  ( .D(I510429), .CLK(I2702), .RSTB(I510217), .Q(I510446) );
nor I_29866 (I510206,I510446,I510268);
nand I_29867 (I510197,I510446,I510367);
DFFARX1 I_29868  ( .D(I333168), .CLK(I2702), .RSTB(I510217), .Q(I510491) );
and I_29869 (I510508,I510491,I333162);
DFFARX1 I_29870  ( .D(I510508), .CLK(I2702), .RSTB(I510217), .Q(I510525) );
not I_29871 (I510188,I510525);
nand I_29872 (I510556,I510508,I510446);
and I_29873 (I510573,I510268,I510556);
DFFARX1 I_29874  ( .D(I510573), .CLK(I2702), .RSTB(I510217), .Q(I510179) );
DFFARX1 I_29875  ( .D(I333144), .CLK(I2702), .RSTB(I510217), .Q(I510604) );
nand I_29876 (I510621,I510604,I510268);
and I_29877 (I510638,I510446,I510621);
DFFARX1 I_29878  ( .D(I510638), .CLK(I2702), .RSTB(I510217), .Q(I510209) );
not I_29879 (I510669,I510604);
nor I_29880 (I510686,I510285,I510669);
and I_29881 (I510703,I510604,I510686);
or I_29882 (I510720,I510508,I510703);
DFFARX1 I_29883  ( .D(I510720), .CLK(I2702), .RSTB(I510217), .Q(I510194) );
nand I_29884 (I510191,I510604,I510350);
DFFARX1 I_29885  ( .D(I510604), .CLK(I2702), .RSTB(I510217), .Q(I510182) );
not I_29886 (I510812,I2709);
nand I_29887 (I510829,I48156,I48162);
and I_29888 (I510846,I510829,I48159);
DFFARX1 I_29889  ( .D(I510846), .CLK(I2702), .RSTB(I510812), .Q(I510863) );
nor I_29890 (I510880,I48183,I48162);
nor I_29891 (I510897,I510880,I510863);
not I_29892 (I510795,I510880);
DFFARX1 I_29893  ( .D(I48174), .CLK(I2702), .RSTB(I510812), .Q(I510928) );
not I_29894 (I510945,I510928);
nor I_29895 (I510962,I510880,I510945);
nand I_29896 (I510798,I510928,I510897);
DFFARX1 I_29897  ( .D(I510928), .CLK(I2702), .RSTB(I510812), .Q(I510780) );
nand I_29898 (I511007,I48177,I48180);
and I_29899 (I511024,I511007,I48153);
DFFARX1 I_29900  ( .D(I511024), .CLK(I2702), .RSTB(I510812), .Q(I511041) );
nor I_29901 (I510801,I511041,I510863);
nand I_29902 (I510792,I511041,I510962);
DFFARX1 I_29903  ( .D(I48171), .CLK(I2702), .RSTB(I510812), .Q(I511086) );
and I_29904 (I511103,I511086,I48165);
DFFARX1 I_29905  ( .D(I511103), .CLK(I2702), .RSTB(I510812), .Q(I511120) );
not I_29906 (I510783,I511120);
nand I_29907 (I511151,I511103,I511041);
and I_29908 (I511168,I510863,I511151);
DFFARX1 I_29909  ( .D(I511168), .CLK(I2702), .RSTB(I510812), .Q(I510774) );
DFFARX1 I_29910  ( .D(I48168), .CLK(I2702), .RSTB(I510812), .Q(I511199) );
nand I_29911 (I511216,I511199,I510863);
and I_29912 (I511233,I511041,I511216);
DFFARX1 I_29913  ( .D(I511233), .CLK(I2702), .RSTB(I510812), .Q(I510804) );
not I_29914 (I511264,I511199);
nor I_29915 (I511281,I510880,I511264);
and I_29916 (I511298,I511199,I511281);
or I_29917 (I511315,I511103,I511298);
DFFARX1 I_29918  ( .D(I511315), .CLK(I2702), .RSTB(I510812), .Q(I510789) );
nand I_29919 (I510786,I511199,I510945);
DFFARX1 I_29920  ( .D(I511199), .CLK(I2702), .RSTB(I510812), .Q(I510777) );
not I_29921 (I511407,I2709);
nand I_29922 (I511424,I25155,I25161);
and I_29923 (I511441,I511424,I25158);
DFFARX1 I_29924  ( .D(I511441), .CLK(I2702), .RSTB(I511407), .Q(I511458) );
nor I_29925 (I511475,I25182,I25161);
nor I_29926 (I511492,I511475,I511458);
not I_29927 (I511390,I511475);
DFFARX1 I_29928  ( .D(I25173), .CLK(I2702), .RSTB(I511407), .Q(I511523) );
not I_29929 (I511540,I511523);
nor I_29930 (I511557,I511475,I511540);
nand I_29931 (I511393,I511523,I511492);
DFFARX1 I_29932  ( .D(I511523), .CLK(I2702), .RSTB(I511407), .Q(I511375) );
nand I_29933 (I511602,I25176,I25179);
and I_29934 (I511619,I511602,I25152);
DFFARX1 I_29935  ( .D(I511619), .CLK(I2702), .RSTB(I511407), .Q(I511636) );
nor I_29936 (I511396,I511636,I511458);
nand I_29937 (I511387,I511636,I511557);
DFFARX1 I_29938  ( .D(I25170), .CLK(I2702), .RSTB(I511407), .Q(I511681) );
and I_29939 (I511698,I511681,I25164);
DFFARX1 I_29940  ( .D(I511698), .CLK(I2702), .RSTB(I511407), .Q(I511715) );
not I_29941 (I511378,I511715);
nand I_29942 (I511746,I511698,I511636);
and I_29943 (I511763,I511458,I511746);
DFFARX1 I_29944  ( .D(I511763), .CLK(I2702), .RSTB(I511407), .Q(I511369) );
DFFARX1 I_29945  ( .D(I25167), .CLK(I2702), .RSTB(I511407), .Q(I511794) );
nand I_29946 (I511811,I511794,I511458);
and I_29947 (I511828,I511636,I511811);
DFFARX1 I_29948  ( .D(I511828), .CLK(I2702), .RSTB(I511407), .Q(I511399) );
not I_29949 (I511859,I511794);
nor I_29950 (I511876,I511475,I511859);
and I_29951 (I511893,I511794,I511876);
or I_29952 (I511910,I511698,I511893);
DFFARX1 I_29953  ( .D(I511910), .CLK(I2702), .RSTB(I511407), .Q(I511384) );
nand I_29954 (I511381,I511794,I511540);
DFFARX1 I_29955  ( .D(I511794), .CLK(I2702), .RSTB(I511407), .Q(I511372) );
not I_29956 (I512002,I2709);
nand I_29957 (I512019,I30765,I30771);
and I_29958 (I512036,I512019,I30768);
DFFARX1 I_29959  ( .D(I512036), .CLK(I2702), .RSTB(I512002), .Q(I512053) );
nor I_29960 (I512070,I30792,I30771);
nor I_29961 (I512087,I512070,I512053);
not I_29962 (I511985,I512070);
DFFARX1 I_29963  ( .D(I30783), .CLK(I2702), .RSTB(I512002), .Q(I512118) );
not I_29964 (I512135,I512118);
nor I_29965 (I512152,I512070,I512135);
nand I_29966 (I511988,I512118,I512087);
DFFARX1 I_29967  ( .D(I512118), .CLK(I2702), .RSTB(I512002), .Q(I511970) );
nand I_29968 (I512197,I30786,I30789);
and I_29969 (I512214,I512197,I30762);
DFFARX1 I_29970  ( .D(I512214), .CLK(I2702), .RSTB(I512002), .Q(I512231) );
nor I_29971 (I511991,I512231,I512053);
nand I_29972 (I511982,I512231,I512152);
DFFARX1 I_29973  ( .D(I30780), .CLK(I2702), .RSTB(I512002), .Q(I512276) );
and I_29974 (I512293,I512276,I30774);
DFFARX1 I_29975  ( .D(I512293), .CLK(I2702), .RSTB(I512002), .Q(I512310) );
not I_29976 (I511973,I512310);
nand I_29977 (I512341,I512293,I512231);
and I_29978 (I512358,I512053,I512341);
DFFARX1 I_29979  ( .D(I512358), .CLK(I2702), .RSTB(I512002), .Q(I511964) );
DFFARX1 I_29980  ( .D(I30777), .CLK(I2702), .RSTB(I512002), .Q(I512389) );
nand I_29981 (I512406,I512389,I512053);
and I_29982 (I512423,I512231,I512406);
DFFARX1 I_29983  ( .D(I512423), .CLK(I2702), .RSTB(I512002), .Q(I511994) );
not I_29984 (I512454,I512389);
nor I_29985 (I512471,I512070,I512454);
and I_29986 (I512488,I512389,I512471);
or I_29987 (I512505,I512293,I512488);
DFFARX1 I_29988  ( .D(I512505), .CLK(I2702), .RSTB(I512002), .Q(I511979) );
nand I_29989 (I511976,I512389,I512135);
DFFARX1 I_29990  ( .D(I512389), .CLK(I2702), .RSTB(I512002), .Q(I511967) );
not I_29991 (I512597,I2709);
nand I_29992 (I512614,I712338,I712344);
and I_29993 (I512631,I512614,I712335);
DFFARX1 I_29994  ( .D(I512631), .CLK(I2702), .RSTB(I512597), .Q(I512648) );
nor I_29995 (I512665,I712347,I712344);
nor I_29996 (I512682,I512665,I512648);
not I_29997 (I512580,I512665);
DFFARX1 I_29998  ( .D(I712326), .CLK(I2702), .RSTB(I512597), .Q(I512713) );
not I_29999 (I512730,I512713);
nor I_30000 (I512747,I512665,I512730);
nand I_30001 (I512583,I512713,I512682);
DFFARX1 I_30002  ( .D(I512713), .CLK(I2702), .RSTB(I512597), .Q(I512565) );
nand I_30003 (I512792,I712350,I712332);
and I_30004 (I512809,I512792,I712341);
DFFARX1 I_30005  ( .D(I512809), .CLK(I2702), .RSTB(I512597), .Q(I512826) );
nor I_30006 (I512586,I512826,I512648);
nand I_30007 (I512577,I512826,I512747);
DFFARX1 I_30008  ( .D(I712356), .CLK(I2702), .RSTB(I512597), .Q(I512871) );
and I_30009 (I512888,I512871,I712329);
DFFARX1 I_30010  ( .D(I512888), .CLK(I2702), .RSTB(I512597), .Q(I512905) );
not I_30011 (I512568,I512905);
nand I_30012 (I512936,I512888,I512826);
and I_30013 (I512953,I512648,I512936);
DFFARX1 I_30014  ( .D(I512953), .CLK(I2702), .RSTB(I512597), .Q(I512559) );
DFFARX1 I_30015  ( .D(I712353), .CLK(I2702), .RSTB(I512597), .Q(I512984) );
nand I_30016 (I513001,I512984,I512648);
and I_30017 (I513018,I512826,I513001);
DFFARX1 I_30018  ( .D(I513018), .CLK(I2702), .RSTB(I512597), .Q(I512589) );
not I_30019 (I513049,I512984);
nor I_30020 (I513066,I512665,I513049);
and I_30021 (I513083,I512984,I513066);
or I_30022 (I513100,I512888,I513083);
DFFARX1 I_30023  ( .D(I513100), .CLK(I2702), .RSTB(I512597), .Q(I512574) );
nand I_30024 (I512571,I512984,I512730);
DFFARX1 I_30025  ( .D(I512984), .CLK(I2702), .RSTB(I512597), .Q(I512562) );
not I_30026 (I513192,I2709);
nand I_30027 (I513209,I243322,I243325);
and I_30028 (I513226,I513209,I243316);
DFFARX1 I_30029  ( .D(I513226), .CLK(I2702), .RSTB(I513192), .Q(I513243) );
nor I_30030 (I513260,I243340,I243325);
nor I_30031 (I513277,I513260,I513243);
not I_30032 (I513175,I513260);
DFFARX1 I_30033  ( .D(I243319), .CLK(I2702), .RSTB(I513192), .Q(I513308) );
not I_30034 (I513325,I513308);
nor I_30035 (I513342,I513260,I513325);
nand I_30036 (I513178,I513308,I513277);
DFFARX1 I_30037  ( .D(I513308), .CLK(I2702), .RSTB(I513192), .Q(I513160) );
nand I_30038 (I513387,I243337,I243328);
and I_30039 (I513404,I513387,I243313);
DFFARX1 I_30040  ( .D(I513404), .CLK(I2702), .RSTB(I513192), .Q(I513421) );
nor I_30041 (I513181,I513421,I513243);
nand I_30042 (I513172,I513421,I513342);
DFFARX1 I_30043  ( .D(I243343), .CLK(I2702), .RSTB(I513192), .Q(I513466) );
and I_30044 (I513483,I513466,I243334);
DFFARX1 I_30045  ( .D(I513483), .CLK(I2702), .RSTB(I513192), .Q(I513500) );
not I_30046 (I513163,I513500);
nand I_30047 (I513531,I513483,I513421);
and I_30048 (I513548,I513243,I513531);
DFFARX1 I_30049  ( .D(I513548), .CLK(I2702), .RSTB(I513192), .Q(I513154) );
DFFARX1 I_30050  ( .D(I243331), .CLK(I2702), .RSTB(I513192), .Q(I513579) );
nand I_30051 (I513596,I513579,I513243);
and I_30052 (I513613,I513421,I513596);
DFFARX1 I_30053  ( .D(I513613), .CLK(I2702), .RSTB(I513192), .Q(I513184) );
not I_30054 (I513644,I513579);
nor I_30055 (I513661,I513260,I513644);
and I_30056 (I513678,I513579,I513661);
or I_30057 (I513695,I513483,I513678);
DFFARX1 I_30058  ( .D(I513695), .CLK(I2702), .RSTB(I513192), .Q(I513169) );
nand I_30059 (I513166,I513579,I513325);
DFFARX1 I_30060  ( .D(I513579), .CLK(I2702), .RSTB(I513192), .Q(I513157) );
not I_30061 (I513787,I2709);
nand I_30062 (I513804,I449482,I449485);
and I_30063 (I513821,I513804,I449479);
DFFARX1 I_30064  ( .D(I513821), .CLK(I2702), .RSTB(I513787), .Q(I513838) );
nor I_30065 (I513855,I449476,I449485);
nor I_30066 (I513872,I513855,I513838);
not I_30067 (I513770,I513855);
DFFARX1 I_30068  ( .D(I449458), .CLK(I2702), .RSTB(I513787), .Q(I513903) );
not I_30069 (I513920,I513903);
nor I_30070 (I513937,I513855,I513920);
nand I_30071 (I513773,I513903,I513872);
DFFARX1 I_30072  ( .D(I513903), .CLK(I2702), .RSTB(I513787), .Q(I513755) );
nand I_30073 (I513982,I449467,I449464);
and I_30074 (I513999,I513982,I449473);
DFFARX1 I_30075  ( .D(I513999), .CLK(I2702), .RSTB(I513787), .Q(I514016) );
nor I_30076 (I513776,I514016,I513838);
nand I_30077 (I513767,I514016,I513937);
DFFARX1 I_30078  ( .D(I449455), .CLK(I2702), .RSTB(I513787), .Q(I514061) );
and I_30079 (I514078,I514061,I449470);
DFFARX1 I_30080  ( .D(I514078), .CLK(I2702), .RSTB(I513787), .Q(I514095) );
not I_30081 (I513758,I514095);
nand I_30082 (I514126,I514078,I514016);
and I_30083 (I514143,I513838,I514126);
DFFARX1 I_30084  ( .D(I514143), .CLK(I2702), .RSTB(I513787), .Q(I513749) );
DFFARX1 I_30085  ( .D(I449461), .CLK(I2702), .RSTB(I513787), .Q(I514174) );
nand I_30086 (I514191,I514174,I513838);
and I_30087 (I514208,I514016,I514191);
DFFARX1 I_30088  ( .D(I514208), .CLK(I2702), .RSTB(I513787), .Q(I513779) );
not I_30089 (I514239,I514174);
nor I_30090 (I514256,I513855,I514239);
and I_30091 (I514273,I514174,I514256);
or I_30092 (I514290,I514078,I514273);
DFFARX1 I_30093  ( .D(I514290), .CLK(I2702), .RSTB(I513787), .Q(I513764) );
nand I_30094 (I513761,I514174,I513920);
DFFARX1 I_30095  ( .D(I514174), .CLK(I2702), .RSTB(I513787), .Q(I513752) );
not I_30096 (I514382,I2709);
nand I_30097 (I514399,I212983,I212980);
and I_30098 (I514416,I514399,I212977);
DFFARX1 I_30099  ( .D(I514416), .CLK(I2702), .RSTB(I514382), .Q(I514433) );
nor I_30100 (I514450,I212968,I212980);
nor I_30101 (I514467,I514450,I514433);
not I_30102 (I514365,I514450);
DFFARX1 I_30103  ( .D(I212986), .CLK(I2702), .RSTB(I514382), .Q(I514498) );
not I_30104 (I514515,I514498);
nor I_30105 (I514532,I514450,I514515);
nand I_30106 (I514368,I514498,I514467);
DFFARX1 I_30107  ( .D(I514498), .CLK(I2702), .RSTB(I514382), .Q(I514350) );
nand I_30108 (I514577,I212971,I212995);
and I_30109 (I514594,I514577,I212974);
DFFARX1 I_30110  ( .D(I514594), .CLK(I2702), .RSTB(I514382), .Q(I514611) );
nor I_30111 (I514371,I514611,I514433);
nand I_30112 (I514362,I514611,I514532);
DFFARX1 I_30113  ( .D(I212992), .CLK(I2702), .RSTB(I514382), .Q(I514656) );
and I_30114 (I514673,I514656,I212989);
DFFARX1 I_30115  ( .D(I514673), .CLK(I2702), .RSTB(I514382), .Q(I514690) );
not I_30116 (I514353,I514690);
nand I_30117 (I514721,I514673,I514611);
and I_30118 (I514738,I514433,I514721);
DFFARX1 I_30119  ( .D(I514738), .CLK(I2702), .RSTB(I514382), .Q(I514344) );
DFFARX1 I_30120  ( .D(I212998), .CLK(I2702), .RSTB(I514382), .Q(I514769) );
nand I_30121 (I514786,I514769,I514433);
and I_30122 (I514803,I514611,I514786);
DFFARX1 I_30123  ( .D(I514803), .CLK(I2702), .RSTB(I514382), .Q(I514374) );
not I_30124 (I514834,I514769);
nor I_30125 (I514851,I514450,I514834);
and I_30126 (I514868,I514769,I514851);
or I_30127 (I514885,I514673,I514868);
DFFARX1 I_30128  ( .D(I514885), .CLK(I2702), .RSTB(I514382), .Q(I514359) );
nand I_30129 (I514356,I514769,I514515);
DFFARX1 I_30130  ( .D(I514769), .CLK(I2702), .RSTB(I514382), .Q(I514347) );
not I_30131 (I514977,I2709);
nand I_30132 (I514994,I81414,I81426);
and I_30133 (I515011,I514994,I81435);
DFFARX1 I_30134  ( .D(I515011), .CLK(I2702), .RSTB(I514977), .Q(I515028) );
nor I_30135 (I515045,I81429,I81426);
nor I_30136 (I515062,I515045,I515028);
not I_30137 (I514960,I515045);
DFFARX1 I_30138  ( .D(I81423), .CLK(I2702), .RSTB(I514977), .Q(I515093) );
not I_30139 (I515110,I515093);
nor I_30140 (I515127,I515045,I515110);
nand I_30141 (I514963,I515093,I515062);
DFFARX1 I_30142  ( .D(I515093), .CLK(I2702), .RSTB(I514977), .Q(I514945) );
nand I_30143 (I515172,I81420,I81417);
and I_30144 (I515189,I515172,I81408);
DFFARX1 I_30145  ( .D(I515189), .CLK(I2702), .RSTB(I514977), .Q(I515206) );
nor I_30146 (I514966,I515206,I515028);
nand I_30147 (I514957,I515206,I515127);
DFFARX1 I_30148  ( .D(I81432), .CLK(I2702), .RSTB(I514977), .Q(I515251) );
and I_30149 (I515268,I515251,I81411);
DFFARX1 I_30150  ( .D(I515268), .CLK(I2702), .RSTB(I514977), .Q(I515285) );
not I_30151 (I514948,I515285);
nand I_30152 (I515316,I515268,I515206);
and I_30153 (I515333,I515028,I515316);
DFFARX1 I_30154  ( .D(I515333), .CLK(I2702), .RSTB(I514977), .Q(I514939) );
DFFARX1 I_30155  ( .D(I81405), .CLK(I2702), .RSTB(I514977), .Q(I515364) );
nand I_30156 (I515381,I515364,I515028);
and I_30157 (I515398,I515206,I515381);
DFFARX1 I_30158  ( .D(I515398), .CLK(I2702), .RSTB(I514977), .Q(I514969) );
not I_30159 (I515429,I515364);
nor I_30160 (I515446,I515045,I515429);
and I_30161 (I515463,I515364,I515446);
or I_30162 (I515480,I515268,I515463);
DFFARX1 I_30163  ( .D(I515480), .CLK(I2702), .RSTB(I514977), .Q(I514954) );
nand I_30164 (I514951,I515364,I515110);
DFFARX1 I_30165  ( .D(I515364), .CLK(I2702), .RSTB(I514977), .Q(I514942) );
not I_30166 (I515572,I2709);
nand I_30167 (I515589,I189951,I189963);
and I_30168 (I515606,I515589,I189942);
DFFARX1 I_30169  ( .D(I515606), .CLK(I2702), .RSTB(I515572), .Q(I515623) );
nor I_30170 (I515640,I189933,I189963);
nor I_30171 (I515657,I515640,I515623);
not I_30172 (I515555,I515640);
DFFARX1 I_30173  ( .D(I189945), .CLK(I2702), .RSTB(I515572), .Q(I515688) );
not I_30174 (I515705,I515688);
nor I_30175 (I515722,I515640,I515705);
nand I_30176 (I515558,I515688,I515657);
DFFARX1 I_30177  ( .D(I515688), .CLK(I2702), .RSTB(I515572), .Q(I515540) );
nand I_30178 (I515767,I189960,I189948);
and I_30179 (I515784,I515767,I189936);
DFFARX1 I_30180  ( .D(I515784), .CLK(I2702), .RSTB(I515572), .Q(I515801) );
nor I_30181 (I515561,I515801,I515623);
nand I_30182 (I515552,I515801,I515722);
DFFARX1 I_30183  ( .D(I189954), .CLK(I2702), .RSTB(I515572), .Q(I515846) );
and I_30184 (I515863,I515846,I189939);
DFFARX1 I_30185  ( .D(I515863), .CLK(I2702), .RSTB(I515572), .Q(I515880) );
not I_30186 (I515543,I515880);
nand I_30187 (I515911,I515863,I515801);
and I_30188 (I515928,I515623,I515911);
DFFARX1 I_30189  ( .D(I515928), .CLK(I2702), .RSTB(I515572), .Q(I515534) );
DFFARX1 I_30190  ( .D(I189957), .CLK(I2702), .RSTB(I515572), .Q(I515959) );
nand I_30191 (I515976,I515959,I515623);
and I_30192 (I515993,I515801,I515976);
DFFARX1 I_30193  ( .D(I515993), .CLK(I2702), .RSTB(I515572), .Q(I515564) );
not I_30194 (I516024,I515959);
nor I_30195 (I516041,I515640,I516024);
and I_30196 (I516058,I515959,I516041);
or I_30197 (I516075,I515863,I516058);
DFFARX1 I_30198  ( .D(I516075), .CLK(I2702), .RSTB(I515572), .Q(I515549) );
nand I_30199 (I515546,I515959,I515705);
DFFARX1 I_30200  ( .D(I515959), .CLK(I2702), .RSTB(I515572), .Q(I515537) );
not I_30201 (I516167,I2709);
nand I_30202 (I516184,I280119,I280125);
and I_30203 (I516201,I516184,I280107);
DFFARX1 I_30204  ( .D(I516201), .CLK(I2702), .RSTB(I516167), .Q(I516218) );
nor I_30205 (I516235,I280101,I280125);
nor I_30206 (I516252,I516235,I516218);
not I_30207 (I516150,I516235);
DFFARX1 I_30208  ( .D(I280131), .CLK(I2702), .RSTB(I516167), .Q(I516283) );
not I_30209 (I516300,I516283);
nor I_30210 (I516317,I516235,I516300);
nand I_30211 (I516153,I516283,I516252);
DFFARX1 I_30212  ( .D(I516283), .CLK(I2702), .RSTB(I516167), .Q(I516135) );
nand I_30213 (I516362,I280122,I280113);
and I_30214 (I516379,I516362,I280116);
DFFARX1 I_30215  ( .D(I516379), .CLK(I2702), .RSTB(I516167), .Q(I516396) );
nor I_30216 (I516156,I516396,I516218);
nand I_30217 (I516147,I516396,I516317);
DFFARX1 I_30218  ( .D(I280128), .CLK(I2702), .RSTB(I516167), .Q(I516441) );
and I_30219 (I516458,I516441,I280104);
DFFARX1 I_30220  ( .D(I516458), .CLK(I2702), .RSTB(I516167), .Q(I516475) );
not I_30221 (I516138,I516475);
nand I_30222 (I516506,I516458,I516396);
and I_30223 (I516523,I516218,I516506);
DFFARX1 I_30224  ( .D(I516523), .CLK(I2702), .RSTB(I516167), .Q(I516129) );
DFFARX1 I_30225  ( .D(I280110), .CLK(I2702), .RSTB(I516167), .Q(I516554) );
nand I_30226 (I516571,I516554,I516218);
and I_30227 (I516588,I516396,I516571);
DFFARX1 I_30228  ( .D(I516588), .CLK(I2702), .RSTB(I516167), .Q(I516159) );
not I_30229 (I516619,I516554);
nor I_30230 (I516636,I516235,I516619);
and I_30231 (I516653,I516554,I516636);
or I_30232 (I516670,I516458,I516653);
DFFARX1 I_30233  ( .D(I516670), .CLK(I2702), .RSTB(I516167), .Q(I516144) );
nand I_30234 (I516141,I516554,I516300);
DFFARX1 I_30235  ( .D(I516554), .CLK(I2702), .RSTB(I516167), .Q(I516132) );
not I_30236 (I516762,I2709);
nand I_30237 (I516779,I486474,I486477);
and I_30238 (I516796,I516779,I486471);
DFFARX1 I_30239  ( .D(I516796), .CLK(I2702), .RSTB(I516762), .Q(I516813) );
nor I_30240 (I516830,I486468,I486477);
nor I_30241 (I516847,I516830,I516813);
not I_30242 (I516745,I516830);
DFFARX1 I_30243  ( .D(I486450), .CLK(I2702), .RSTB(I516762), .Q(I516878) );
not I_30244 (I516895,I516878);
nor I_30245 (I516912,I516830,I516895);
nand I_30246 (I516748,I516878,I516847);
DFFARX1 I_30247  ( .D(I516878), .CLK(I2702), .RSTB(I516762), .Q(I516730) );
nand I_30248 (I516957,I486459,I486456);
and I_30249 (I516974,I516957,I486465);
DFFARX1 I_30250  ( .D(I516974), .CLK(I2702), .RSTB(I516762), .Q(I516991) );
nor I_30251 (I516751,I516991,I516813);
nand I_30252 (I516742,I516991,I516912);
DFFARX1 I_30253  ( .D(I486447), .CLK(I2702), .RSTB(I516762), .Q(I517036) );
and I_30254 (I517053,I517036,I486462);
DFFARX1 I_30255  ( .D(I517053), .CLK(I2702), .RSTB(I516762), .Q(I517070) );
not I_30256 (I516733,I517070);
nand I_30257 (I517101,I517053,I516991);
and I_30258 (I517118,I516813,I517101);
DFFARX1 I_30259  ( .D(I517118), .CLK(I2702), .RSTB(I516762), .Q(I516724) );
DFFARX1 I_30260  ( .D(I486453), .CLK(I2702), .RSTB(I516762), .Q(I517149) );
nand I_30261 (I517166,I517149,I516813);
and I_30262 (I517183,I516991,I517166);
DFFARX1 I_30263  ( .D(I517183), .CLK(I2702), .RSTB(I516762), .Q(I516754) );
not I_30264 (I517214,I517149);
nor I_30265 (I517231,I516830,I517214);
and I_30266 (I517248,I517149,I517231);
or I_30267 (I517265,I517053,I517248);
DFFARX1 I_30268  ( .D(I517265), .CLK(I2702), .RSTB(I516762), .Q(I516739) );
nand I_30269 (I516736,I517149,I516895);
DFFARX1 I_30270  ( .D(I517149), .CLK(I2702), .RSTB(I516762), .Q(I516727) );
not I_30271 (I517357,I2709);
nand I_30272 (I517374,I136324,I136336);
and I_30273 (I517391,I517374,I136345);
DFFARX1 I_30274  ( .D(I517391), .CLK(I2702), .RSTB(I517357), .Q(I517408) );
nor I_30275 (I517425,I136339,I136336);
nor I_30276 (I517442,I517425,I517408);
not I_30277 (I517340,I517425);
DFFARX1 I_30278  ( .D(I136333), .CLK(I2702), .RSTB(I517357), .Q(I517473) );
not I_30279 (I517490,I517473);
nor I_30280 (I517507,I517425,I517490);
nand I_30281 (I517343,I517473,I517442);
DFFARX1 I_30282  ( .D(I517473), .CLK(I2702), .RSTB(I517357), .Q(I517325) );
nand I_30283 (I517552,I136330,I136327);
and I_30284 (I517569,I517552,I136318);
DFFARX1 I_30285  ( .D(I517569), .CLK(I2702), .RSTB(I517357), .Q(I517586) );
nor I_30286 (I517346,I517586,I517408);
nand I_30287 (I517337,I517586,I517507);
DFFARX1 I_30288  ( .D(I136342), .CLK(I2702), .RSTB(I517357), .Q(I517631) );
and I_30289 (I517648,I517631,I136321);
DFFARX1 I_30290  ( .D(I517648), .CLK(I2702), .RSTB(I517357), .Q(I517665) );
not I_30291 (I517328,I517665);
nand I_30292 (I517696,I517648,I517586);
and I_30293 (I517713,I517408,I517696);
DFFARX1 I_30294  ( .D(I517713), .CLK(I2702), .RSTB(I517357), .Q(I517319) );
DFFARX1 I_30295  ( .D(I136315), .CLK(I2702), .RSTB(I517357), .Q(I517744) );
nand I_30296 (I517761,I517744,I517408);
and I_30297 (I517778,I517586,I517761);
DFFARX1 I_30298  ( .D(I517778), .CLK(I2702), .RSTB(I517357), .Q(I517349) );
not I_30299 (I517809,I517744);
nor I_30300 (I517826,I517425,I517809);
and I_30301 (I517843,I517744,I517826);
or I_30302 (I517860,I517648,I517843);
DFFARX1 I_30303  ( .D(I517860), .CLK(I2702), .RSTB(I517357), .Q(I517334) );
nand I_30304 (I517331,I517744,I517490);
DFFARX1 I_30305  ( .D(I517744), .CLK(I2702), .RSTB(I517357), .Q(I517322) );
not I_30306 (I517952,I2709);
nand I_30307 (I517969,I270174,I270180);
and I_30308 (I517986,I517969,I270162);
DFFARX1 I_30309  ( .D(I517986), .CLK(I2702), .RSTB(I517952), .Q(I518003) );
nor I_30310 (I518020,I270156,I270180);
nor I_30311 (I518037,I518020,I518003);
not I_30312 (I517935,I518020);
DFFARX1 I_30313  ( .D(I270186), .CLK(I2702), .RSTB(I517952), .Q(I518068) );
not I_30314 (I518085,I518068);
nor I_30315 (I518102,I518020,I518085);
nand I_30316 (I517938,I518068,I518037);
DFFARX1 I_30317  ( .D(I518068), .CLK(I2702), .RSTB(I517952), .Q(I517920) );
nand I_30318 (I518147,I270177,I270168);
and I_30319 (I518164,I518147,I270171);
DFFARX1 I_30320  ( .D(I518164), .CLK(I2702), .RSTB(I517952), .Q(I518181) );
nor I_30321 (I517941,I518181,I518003);
nand I_30322 (I517932,I518181,I518102);
DFFARX1 I_30323  ( .D(I270183), .CLK(I2702), .RSTB(I517952), .Q(I518226) );
and I_30324 (I518243,I518226,I270159);
DFFARX1 I_30325  ( .D(I518243), .CLK(I2702), .RSTB(I517952), .Q(I518260) );
not I_30326 (I517923,I518260);
nand I_30327 (I518291,I518243,I518181);
and I_30328 (I518308,I518003,I518291);
DFFARX1 I_30329  ( .D(I518308), .CLK(I2702), .RSTB(I517952), .Q(I517914) );
DFFARX1 I_30330  ( .D(I270165), .CLK(I2702), .RSTB(I517952), .Q(I518339) );
nand I_30331 (I518356,I518339,I518003);
and I_30332 (I518373,I518181,I518356);
DFFARX1 I_30333  ( .D(I518373), .CLK(I2702), .RSTB(I517952), .Q(I517944) );
not I_30334 (I518404,I518339);
nor I_30335 (I518421,I518020,I518404);
and I_30336 (I518438,I518339,I518421);
or I_30337 (I518455,I518243,I518438);
DFFARX1 I_30338  ( .D(I518455), .CLK(I2702), .RSTB(I517952), .Q(I517929) );
nand I_30339 (I517926,I518339,I518085);
DFFARX1 I_30340  ( .D(I518339), .CLK(I2702), .RSTB(I517952), .Q(I517917) );
not I_30341 (I518547,I2709);
nand I_30342 (I518564,I153486,I153498);
and I_30343 (I518581,I518564,I153477);
DFFARX1 I_30344  ( .D(I518581), .CLK(I2702), .RSTB(I518547), .Q(I518598) );
nor I_30345 (I518615,I153468,I153498);
nor I_30346 (I518632,I518615,I518598);
not I_30347 (I518530,I518615);
DFFARX1 I_30348  ( .D(I153480), .CLK(I2702), .RSTB(I518547), .Q(I518663) );
not I_30349 (I518680,I518663);
nor I_30350 (I518697,I518615,I518680);
nand I_30351 (I518533,I518663,I518632);
DFFARX1 I_30352  ( .D(I518663), .CLK(I2702), .RSTB(I518547), .Q(I518515) );
nand I_30353 (I518742,I153495,I153483);
and I_30354 (I518759,I518742,I153471);
DFFARX1 I_30355  ( .D(I518759), .CLK(I2702), .RSTB(I518547), .Q(I518776) );
nor I_30356 (I518536,I518776,I518598);
nand I_30357 (I518527,I518776,I518697);
DFFARX1 I_30358  ( .D(I153489), .CLK(I2702), .RSTB(I518547), .Q(I518821) );
and I_30359 (I518838,I518821,I153474);
DFFARX1 I_30360  ( .D(I518838), .CLK(I2702), .RSTB(I518547), .Q(I518855) );
not I_30361 (I518518,I518855);
nand I_30362 (I518886,I518838,I518776);
and I_30363 (I518903,I518598,I518886);
DFFARX1 I_30364  ( .D(I518903), .CLK(I2702), .RSTB(I518547), .Q(I518509) );
DFFARX1 I_30365  ( .D(I153492), .CLK(I2702), .RSTB(I518547), .Q(I518934) );
nand I_30366 (I518951,I518934,I518598);
and I_30367 (I518968,I518776,I518951);
DFFARX1 I_30368  ( .D(I518968), .CLK(I2702), .RSTB(I518547), .Q(I518539) );
not I_30369 (I518999,I518934);
nor I_30370 (I519016,I518615,I518999);
and I_30371 (I519033,I518934,I519016);
or I_30372 (I519050,I518838,I519033);
DFFARX1 I_30373  ( .D(I519050), .CLK(I2702), .RSTB(I518547), .Q(I518524) );
nand I_30374 (I518521,I518934,I518680);
DFFARX1 I_30375  ( .D(I518934), .CLK(I2702), .RSTB(I518547), .Q(I518512) );
not I_30376 (I519142,I2709);
nand I_30377 (I519159,I305313,I305319);
and I_30378 (I519176,I519159,I305301);
DFFARX1 I_30379  ( .D(I519176), .CLK(I2702), .RSTB(I519142), .Q(I519193) );
nor I_30380 (I519210,I305295,I305319);
nor I_30381 (I519227,I519210,I519193);
not I_30382 (I519125,I519210);
DFFARX1 I_30383  ( .D(I305325), .CLK(I2702), .RSTB(I519142), .Q(I519258) );
not I_30384 (I519275,I519258);
nor I_30385 (I519292,I519210,I519275);
nand I_30386 (I519128,I519258,I519227);
DFFARX1 I_30387  ( .D(I519258), .CLK(I2702), .RSTB(I519142), .Q(I519110) );
nand I_30388 (I519337,I305316,I305307);
and I_30389 (I519354,I519337,I305310);
DFFARX1 I_30390  ( .D(I519354), .CLK(I2702), .RSTB(I519142), .Q(I519371) );
nor I_30391 (I519131,I519371,I519193);
nand I_30392 (I519122,I519371,I519292);
DFFARX1 I_30393  ( .D(I305322), .CLK(I2702), .RSTB(I519142), .Q(I519416) );
and I_30394 (I519433,I519416,I305298);
DFFARX1 I_30395  ( .D(I519433), .CLK(I2702), .RSTB(I519142), .Q(I519450) );
not I_30396 (I519113,I519450);
nand I_30397 (I519481,I519433,I519371);
and I_30398 (I519498,I519193,I519481);
DFFARX1 I_30399  ( .D(I519498), .CLK(I2702), .RSTB(I519142), .Q(I519104) );
DFFARX1 I_30400  ( .D(I305304), .CLK(I2702), .RSTB(I519142), .Q(I519529) );
nand I_30401 (I519546,I519529,I519193);
and I_30402 (I519563,I519371,I519546);
DFFARX1 I_30403  ( .D(I519563), .CLK(I2702), .RSTB(I519142), .Q(I519134) );
not I_30404 (I519594,I519529);
nor I_30405 (I519611,I519210,I519594);
and I_30406 (I519628,I519529,I519611);
or I_30407 (I519645,I519433,I519628);
DFFARX1 I_30408  ( .D(I519645), .CLK(I2702), .RSTB(I519142), .Q(I519119) );
nand I_30409 (I519116,I519529,I519275);
DFFARX1 I_30410  ( .D(I519529), .CLK(I2702), .RSTB(I519142), .Q(I519107) );
not I_30411 (I519737,I2709);
nand I_30412 (I519754,I693842,I693848);
and I_30413 (I519771,I519754,I693839);
DFFARX1 I_30414  ( .D(I519771), .CLK(I2702), .RSTB(I519737), .Q(I519788) );
nor I_30415 (I519805,I693851,I693848);
nor I_30416 (I519822,I519805,I519788);
not I_30417 (I519720,I519805);
DFFARX1 I_30418  ( .D(I693830), .CLK(I2702), .RSTB(I519737), .Q(I519853) );
not I_30419 (I519870,I519853);
nor I_30420 (I519887,I519805,I519870);
nand I_30421 (I519723,I519853,I519822);
DFFARX1 I_30422  ( .D(I519853), .CLK(I2702), .RSTB(I519737), .Q(I519705) );
nand I_30423 (I519932,I693854,I693836);
and I_30424 (I519949,I519932,I693845);
DFFARX1 I_30425  ( .D(I519949), .CLK(I2702), .RSTB(I519737), .Q(I519966) );
nor I_30426 (I519726,I519966,I519788);
nand I_30427 (I519717,I519966,I519887);
DFFARX1 I_30428  ( .D(I693860), .CLK(I2702), .RSTB(I519737), .Q(I520011) );
and I_30429 (I520028,I520011,I693833);
DFFARX1 I_30430  ( .D(I520028), .CLK(I2702), .RSTB(I519737), .Q(I520045) );
not I_30431 (I519708,I520045);
nand I_30432 (I520076,I520028,I519966);
and I_30433 (I520093,I519788,I520076);
DFFARX1 I_30434  ( .D(I520093), .CLK(I2702), .RSTB(I519737), .Q(I519699) );
DFFARX1 I_30435  ( .D(I693857), .CLK(I2702), .RSTB(I519737), .Q(I520124) );
nand I_30436 (I520141,I520124,I519788);
and I_30437 (I520158,I519966,I520141);
DFFARX1 I_30438  ( .D(I520158), .CLK(I2702), .RSTB(I519737), .Q(I519729) );
not I_30439 (I520189,I520124);
nor I_30440 (I520206,I519805,I520189);
and I_30441 (I520223,I520124,I520206);
or I_30442 (I520240,I520028,I520223);
DFFARX1 I_30443  ( .D(I520240), .CLK(I2702), .RSTB(I519737), .Q(I519714) );
nand I_30444 (I519711,I520124,I519870);
DFFARX1 I_30445  ( .D(I520124), .CLK(I2702), .RSTB(I519737), .Q(I519702) );
not I_30446 (I520332,I2709);
nand I_30447 (I520349,I57512,I57524);
and I_30448 (I520366,I520349,I57533);
DFFARX1 I_30449  ( .D(I520366), .CLK(I2702), .RSTB(I520332), .Q(I520383) );
nor I_30450 (I520400,I57527,I57524);
nor I_30451 (I520417,I520400,I520383);
not I_30452 (I520315,I520400);
DFFARX1 I_30453  ( .D(I57521), .CLK(I2702), .RSTB(I520332), .Q(I520448) );
not I_30454 (I520465,I520448);
nor I_30455 (I520482,I520400,I520465);
nand I_30456 (I520318,I520448,I520417);
DFFARX1 I_30457  ( .D(I520448), .CLK(I2702), .RSTB(I520332), .Q(I520300) );
nand I_30458 (I520527,I57518,I57515);
and I_30459 (I520544,I520527,I57506);
DFFARX1 I_30460  ( .D(I520544), .CLK(I2702), .RSTB(I520332), .Q(I520561) );
nor I_30461 (I520321,I520561,I520383);
nand I_30462 (I520312,I520561,I520482);
DFFARX1 I_30463  ( .D(I57530), .CLK(I2702), .RSTB(I520332), .Q(I520606) );
and I_30464 (I520623,I520606,I57509);
DFFARX1 I_30465  ( .D(I520623), .CLK(I2702), .RSTB(I520332), .Q(I520640) );
not I_30466 (I520303,I520640);
nand I_30467 (I520671,I520623,I520561);
and I_30468 (I520688,I520383,I520671);
DFFARX1 I_30469  ( .D(I520688), .CLK(I2702), .RSTB(I520332), .Q(I520294) );
DFFARX1 I_30470  ( .D(I57503), .CLK(I2702), .RSTB(I520332), .Q(I520719) );
nand I_30471 (I520736,I520719,I520383);
and I_30472 (I520753,I520561,I520736);
DFFARX1 I_30473  ( .D(I520753), .CLK(I2702), .RSTB(I520332), .Q(I520324) );
not I_30474 (I520784,I520719);
nor I_30475 (I520801,I520400,I520784);
and I_30476 (I520818,I520719,I520801);
or I_30477 (I520835,I520623,I520818);
DFFARX1 I_30478  ( .D(I520835), .CLK(I2702), .RSTB(I520332), .Q(I520309) );
nand I_30479 (I520306,I520719,I520465);
DFFARX1 I_30480  ( .D(I520719), .CLK(I2702), .RSTB(I520332), .Q(I520297) );
not I_30481 (I520927,I2709);
nand I_30482 (I520944,I440234,I440237);
and I_30483 (I520961,I520944,I440231);
DFFARX1 I_30484  ( .D(I520961), .CLK(I2702), .RSTB(I520927), .Q(I520978) );
nor I_30485 (I520995,I440228,I440237);
nor I_30486 (I521012,I520995,I520978);
not I_30487 (I520910,I520995);
DFFARX1 I_30488  ( .D(I440210), .CLK(I2702), .RSTB(I520927), .Q(I521043) );
not I_30489 (I521060,I521043);
nor I_30490 (I521077,I520995,I521060);
nand I_30491 (I520913,I521043,I521012);
DFFARX1 I_30492  ( .D(I521043), .CLK(I2702), .RSTB(I520927), .Q(I520895) );
nand I_30493 (I521122,I440219,I440216);
and I_30494 (I521139,I521122,I440225);
DFFARX1 I_30495  ( .D(I521139), .CLK(I2702), .RSTB(I520927), .Q(I521156) );
nor I_30496 (I520916,I521156,I520978);
nand I_30497 (I520907,I521156,I521077);
DFFARX1 I_30498  ( .D(I440207), .CLK(I2702), .RSTB(I520927), .Q(I521201) );
and I_30499 (I521218,I521201,I440222);
DFFARX1 I_30500  ( .D(I521218), .CLK(I2702), .RSTB(I520927), .Q(I521235) );
not I_30501 (I520898,I521235);
nand I_30502 (I521266,I521218,I521156);
and I_30503 (I521283,I520978,I521266);
DFFARX1 I_30504  ( .D(I521283), .CLK(I2702), .RSTB(I520927), .Q(I520889) );
DFFARX1 I_30505  ( .D(I440213), .CLK(I2702), .RSTB(I520927), .Q(I521314) );
nand I_30506 (I521331,I521314,I520978);
and I_30507 (I521348,I521156,I521331);
DFFARX1 I_30508  ( .D(I521348), .CLK(I2702), .RSTB(I520927), .Q(I520919) );
not I_30509 (I521379,I521314);
nor I_30510 (I521396,I520995,I521379);
and I_30511 (I521413,I521314,I521396);
or I_30512 (I521430,I521218,I521413);
DFFARX1 I_30513  ( .D(I521430), .CLK(I2702), .RSTB(I520927), .Q(I520904) );
nand I_30514 (I520901,I521314,I521060);
DFFARX1 I_30515  ( .D(I521314), .CLK(I2702), .RSTB(I520927), .Q(I520892) );
not I_30516 (I521522,I2709);
nand I_30517 (I521539,I672190,I672181);
and I_30518 (I521556,I521539,I672199);
DFFARX1 I_30519  ( .D(I521556), .CLK(I2702), .RSTB(I521522), .Q(I521573) );
nor I_30520 (I521590,I672196,I672181);
nor I_30521 (I521607,I521590,I521573);
not I_30522 (I521505,I521590);
DFFARX1 I_30523  ( .D(I672178), .CLK(I2702), .RSTB(I521522), .Q(I521638) );
not I_30524 (I521655,I521638);
nor I_30525 (I521672,I521590,I521655);
nand I_30526 (I521508,I521638,I521607);
DFFARX1 I_30527  ( .D(I521638), .CLK(I2702), .RSTB(I521522), .Q(I521490) );
nand I_30528 (I521717,I672187,I672202);
and I_30529 (I521734,I521717,I672193);
DFFARX1 I_30530  ( .D(I521734), .CLK(I2702), .RSTB(I521522), .Q(I521751) );
nor I_30531 (I521511,I521751,I521573);
nand I_30532 (I521502,I521751,I521672);
DFFARX1 I_30533  ( .D(I672175), .CLK(I2702), .RSTB(I521522), .Q(I521796) );
and I_30534 (I521813,I521796,I672184);
DFFARX1 I_30535  ( .D(I521813), .CLK(I2702), .RSTB(I521522), .Q(I521830) );
not I_30536 (I521493,I521830);
nand I_30537 (I521861,I521813,I521751);
and I_30538 (I521878,I521573,I521861);
DFFARX1 I_30539  ( .D(I521878), .CLK(I2702), .RSTB(I521522), .Q(I521484) );
DFFARX1 I_30540  ( .D(I672172), .CLK(I2702), .RSTB(I521522), .Q(I521909) );
nand I_30541 (I521926,I521909,I521573);
and I_30542 (I521943,I521751,I521926);
DFFARX1 I_30543  ( .D(I521943), .CLK(I2702), .RSTB(I521522), .Q(I521514) );
not I_30544 (I521974,I521909);
nor I_30545 (I521991,I521590,I521974);
and I_30546 (I522008,I521909,I521991);
or I_30547 (I522025,I521813,I522008);
DFFARX1 I_30548  ( .D(I522025), .CLK(I2702), .RSTB(I521522), .Q(I521499) );
nand I_30549 (I521496,I521909,I521655);
DFFARX1 I_30550  ( .D(I521909), .CLK(I2702), .RSTB(I521522), .Q(I521487) );
not I_30551 (I522117,I2709);
nand I_30552 (I522134,I723320,I723326);
and I_30553 (I522151,I522134,I723317);
DFFARX1 I_30554  ( .D(I522151), .CLK(I2702), .RSTB(I522117), .Q(I522168) );
nor I_30555 (I522185,I723329,I723326);
nor I_30556 (I522202,I522185,I522168);
not I_30557 (I522100,I522185);
DFFARX1 I_30558  ( .D(I723308), .CLK(I2702), .RSTB(I522117), .Q(I522233) );
not I_30559 (I522250,I522233);
nor I_30560 (I522267,I522185,I522250);
nand I_30561 (I522103,I522233,I522202);
DFFARX1 I_30562  ( .D(I522233), .CLK(I2702), .RSTB(I522117), .Q(I522085) );
nand I_30563 (I522312,I723332,I723314);
and I_30564 (I522329,I522312,I723323);
DFFARX1 I_30565  ( .D(I522329), .CLK(I2702), .RSTB(I522117), .Q(I522346) );
nor I_30566 (I522106,I522346,I522168);
nand I_30567 (I522097,I522346,I522267);
DFFARX1 I_30568  ( .D(I723338), .CLK(I2702), .RSTB(I522117), .Q(I522391) );
and I_30569 (I522408,I522391,I723311);
DFFARX1 I_30570  ( .D(I522408), .CLK(I2702), .RSTB(I522117), .Q(I522425) );
not I_30571 (I522088,I522425);
nand I_30572 (I522456,I522408,I522346);
and I_30573 (I522473,I522168,I522456);
DFFARX1 I_30574  ( .D(I522473), .CLK(I2702), .RSTB(I522117), .Q(I522079) );
DFFARX1 I_30575  ( .D(I723335), .CLK(I2702), .RSTB(I522117), .Q(I522504) );
nand I_30576 (I522521,I522504,I522168);
and I_30577 (I522538,I522346,I522521);
DFFARX1 I_30578  ( .D(I522538), .CLK(I2702), .RSTB(I522117), .Q(I522109) );
not I_30579 (I522569,I522504);
nor I_30580 (I522586,I522185,I522569);
and I_30581 (I522603,I522504,I522586);
or I_30582 (I522620,I522408,I522603);
DFFARX1 I_30583  ( .D(I522620), .CLK(I2702), .RSTB(I522117), .Q(I522094) );
nand I_30584 (I522091,I522504,I522250);
DFFARX1 I_30585  ( .D(I522504), .CLK(I2702), .RSTB(I522117), .Q(I522082) );
not I_30586 (I522712,I2709);
nand I_30587 (I522729,I59450,I59462);
and I_30588 (I522746,I522729,I59471);
DFFARX1 I_30589  ( .D(I522746), .CLK(I2702), .RSTB(I522712), .Q(I522763) );
nor I_30590 (I522780,I59465,I59462);
nor I_30591 (I522797,I522780,I522763);
not I_30592 (I522695,I522780);
DFFARX1 I_30593  ( .D(I59459), .CLK(I2702), .RSTB(I522712), .Q(I522828) );
not I_30594 (I522845,I522828);
nor I_30595 (I522862,I522780,I522845);
nand I_30596 (I522698,I522828,I522797);
DFFARX1 I_30597  ( .D(I522828), .CLK(I2702), .RSTB(I522712), .Q(I522680) );
nand I_30598 (I522907,I59456,I59453);
and I_30599 (I522924,I522907,I59444);
DFFARX1 I_30600  ( .D(I522924), .CLK(I2702), .RSTB(I522712), .Q(I522941) );
nor I_30601 (I522701,I522941,I522763);
nand I_30602 (I522692,I522941,I522862);
DFFARX1 I_30603  ( .D(I59468), .CLK(I2702), .RSTB(I522712), .Q(I522986) );
and I_30604 (I523003,I522986,I59447);
DFFARX1 I_30605  ( .D(I523003), .CLK(I2702), .RSTB(I522712), .Q(I523020) );
not I_30606 (I522683,I523020);
nand I_30607 (I523051,I523003,I522941);
and I_30608 (I523068,I522763,I523051);
DFFARX1 I_30609  ( .D(I523068), .CLK(I2702), .RSTB(I522712), .Q(I522674) );
DFFARX1 I_30610  ( .D(I59441), .CLK(I2702), .RSTB(I522712), .Q(I523099) );
nand I_30611 (I523116,I523099,I522763);
and I_30612 (I523133,I522941,I523116);
DFFARX1 I_30613  ( .D(I523133), .CLK(I2702), .RSTB(I522712), .Q(I522704) );
not I_30614 (I523164,I523099);
nor I_30615 (I523181,I522780,I523164);
and I_30616 (I523198,I523099,I523181);
or I_30617 (I523215,I523003,I523198);
DFFARX1 I_30618  ( .D(I523215), .CLK(I2702), .RSTB(I522712), .Q(I522689) );
nand I_30619 (I522686,I523099,I522845);
DFFARX1 I_30620  ( .D(I523099), .CLK(I2702), .RSTB(I522712), .Q(I522677) );
not I_30621 (I523307,I2709);
nand I_30622 (I523324,I720430,I720436);
and I_30623 (I523341,I523324,I720427);
DFFARX1 I_30624  ( .D(I523341), .CLK(I2702), .RSTB(I523307), .Q(I523358) );
nor I_30625 (I523375,I720439,I720436);
nor I_30626 (I523392,I523375,I523358);
not I_30627 (I523290,I523375);
DFFARX1 I_30628  ( .D(I720418), .CLK(I2702), .RSTB(I523307), .Q(I523423) );
not I_30629 (I523440,I523423);
nor I_30630 (I523457,I523375,I523440);
nand I_30631 (I523293,I523423,I523392);
DFFARX1 I_30632  ( .D(I523423), .CLK(I2702), .RSTB(I523307), .Q(I523275) );
nand I_30633 (I523502,I720442,I720424);
and I_30634 (I523519,I523502,I720433);
DFFARX1 I_30635  ( .D(I523519), .CLK(I2702), .RSTB(I523307), .Q(I523536) );
nor I_30636 (I523296,I523536,I523358);
nand I_30637 (I523287,I523536,I523457);
DFFARX1 I_30638  ( .D(I720448), .CLK(I2702), .RSTB(I523307), .Q(I523581) );
and I_30639 (I523598,I523581,I720421);
DFFARX1 I_30640  ( .D(I523598), .CLK(I2702), .RSTB(I523307), .Q(I523615) );
not I_30641 (I523278,I523615);
nand I_30642 (I523646,I523598,I523536);
and I_30643 (I523663,I523358,I523646);
DFFARX1 I_30644  ( .D(I523663), .CLK(I2702), .RSTB(I523307), .Q(I523269) );
DFFARX1 I_30645  ( .D(I720445), .CLK(I2702), .RSTB(I523307), .Q(I523694) );
nand I_30646 (I523711,I523694,I523358);
and I_30647 (I523728,I523536,I523711);
DFFARX1 I_30648  ( .D(I523728), .CLK(I2702), .RSTB(I523307), .Q(I523299) );
not I_30649 (I523759,I523694);
nor I_30650 (I523776,I523375,I523759);
and I_30651 (I523793,I523694,I523776);
or I_30652 (I523810,I523598,I523793);
DFFARX1 I_30653  ( .D(I523810), .CLK(I2702), .RSTB(I523307), .Q(I523284) );
nand I_30654 (I523281,I523694,I523440);
DFFARX1 I_30655  ( .D(I523694), .CLK(I2702), .RSTB(I523307), .Q(I523272) );
not I_30656 (I523902,I2709);
nand I_30657 (I523919,I179343,I179355);
and I_30658 (I523936,I523919,I179334);
DFFARX1 I_30659  ( .D(I523936), .CLK(I2702), .RSTB(I523902), .Q(I523953) );
nor I_30660 (I523970,I179325,I179355);
nor I_30661 (I523987,I523970,I523953);
not I_30662 (I523885,I523970);
DFFARX1 I_30663  ( .D(I179337), .CLK(I2702), .RSTB(I523902), .Q(I524018) );
not I_30664 (I524035,I524018);
nor I_30665 (I524052,I523970,I524035);
nand I_30666 (I523888,I524018,I523987);
DFFARX1 I_30667  ( .D(I524018), .CLK(I2702), .RSTB(I523902), .Q(I523870) );
nand I_30668 (I524097,I179352,I179340);
and I_30669 (I524114,I524097,I179328);
DFFARX1 I_30670  ( .D(I524114), .CLK(I2702), .RSTB(I523902), .Q(I524131) );
nor I_30671 (I523891,I524131,I523953);
nand I_30672 (I523882,I524131,I524052);
DFFARX1 I_30673  ( .D(I179346), .CLK(I2702), .RSTB(I523902), .Q(I524176) );
and I_30674 (I524193,I524176,I179331);
DFFARX1 I_30675  ( .D(I524193), .CLK(I2702), .RSTB(I523902), .Q(I524210) );
not I_30676 (I523873,I524210);
nand I_30677 (I524241,I524193,I524131);
and I_30678 (I524258,I523953,I524241);
DFFARX1 I_30679  ( .D(I524258), .CLK(I2702), .RSTB(I523902), .Q(I523864) );
DFFARX1 I_30680  ( .D(I179349), .CLK(I2702), .RSTB(I523902), .Q(I524289) );
nand I_30681 (I524306,I524289,I523953);
and I_30682 (I524323,I524131,I524306);
DFFARX1 I_30683  ( .D(I524323), .CLK(I2702), .RSTB(I523902), .Q(I523894) );
not I_30684 (I524354,I524289);
nor I_30685 (I524371,I523970,I524354);
and I_30686 (I524388,I524289,I524371);
or I_30687 (I524405,I524193,I524388);
DFFARX1 I_30688  ( .D(I524405), .CLK(I2702), .RSTB(I523902), .Q(I523879) );
nand I_30689 (I523876,I524289,I524035);
DFFARX1 I_30690  ( .D(I524289), .CLK(I2702), .RSTB(I523902), .Q(I523867) );
not I_30691 (I524497,I2709);
nand I_30692 (I524514,I278793,I278799);
and I_30693 (I524531,I524514,I278781);
DFFARX1 I_30694  ( .D(I524531), .CLK(I2702), .RSTB(I524497), .Q(I524548) );
nor I_30695 (I524565,I278775,I278799);
nor I_30696 (I524582,I524565,I524548);
not I_30697 (I524480,I524565);
DFFARX1 I_30698  ( .D(I278805), .CLK(I2702), .RSTB(I524497), .Q(I524613) );
not I_30699 (I524630,I524613);
nor I_30700 (I524647,I524565,I524630);
nand I_30701 (I524483,I524613,I524582);
DFFARX1 I_30702  ( .D(I524613), .CLK(I2702), .RSTB(I524497), .Q(I524465) );
nand I_30703 (I524692,I278796,I278787);
and I_30704 (I524709,I524692,I278790);
DFFARX1 I_30705  ( .D(I524709), .CLK(I2702), .RSTB(I524497), .Q(I524726) );
nor I_30706 (I524486,I524726,I524548);
nand I_30707 (I524477,I524726,I524647);
DFFARX1 I_30708  ( .D(I278802), .CLK(I2702), .RSTB(I524497), .Q(I524771) );
and I_30709 (I524788,I524771,I278778);
DFFARX1 I_30710  ( .D(I524788), .CLK(I2702), .RSTB(I524497), .Q(I524805) );
not I_30711 (I524468,I524805);
nand I_30712 (I524836,I524788,I524726);
and I_30713 (I524853,I524548,I524836);
DFFARX1 I_30714  ( .D(I524853), .CLK(I2702), .RSTB(I524497), .Q(I524459) );
DFFARX1 I_30715  ( .D(I278784), .CLK(I2702), .RSTB(I524497), .Q(I524884) );
nand I_30716 (I524901,I524884,I524548);
and I_30717 (I524918,I524726,I524901);
DFFARX1 I_30718  ( .D(I524918), .CLK(I2702), .RSTB(I524497), .Q(I524489) );
not I_30719 (I524949,I524884);
nor I_30720 (I524966,I524565,I524949);
and I_30721 (I524983,I524884,I524966);
or I_30722 (I525000,I524788,I524983);
DFFARX1 I_30723  ( .D(I525000), .CLK(I2702), .RSTB(I524497), .Q(I524474) );
nand I_30724 (I524471,I524884,I524630);
DFFARX1 I_30725  ( .D(I524884), .CLK(I2702), .RSTB(I524497), .Q(I524462) );
not I_30726 (I525092,I2709);
nand I_30727 (I525109,I618096,I618087);
and I_30728 (I525126,I525109,I618105);
DFFARX1 I_30729  ( .D(I525126), .CLK(I2702), .RSTB(I525092), .Q(I525143) );
nor I_30730 (I525160,I618102,I618087);
nor I_30731 (I525177,I525160,I525143);
not I_30732 (I525075,I525160);
DFFARX1 I_30733  ( .D(I618084), .CLK(I2702), .RSTB(I525092), .Q(I525208) );
not I_30734 (I525225,I525208);
nor I_30735 (I525242,I525160,I525225);
nand I_30736 (I525078,I525208,I525177);
DFFARX1 I_30737  ( .D(I525208), .CLK(I2702), .RSTB(I525092), .Q(I525060) );
nand I_30738 (I525287,I618093,I618108);
and I_30739 (I525304,I525287,I618099);
DFFARX1 I_30740  ( .D(I525304), .CLK(I2702), .RSTB(I525092), .Q(I525321) );
nor I_30741 (I525081,I525321,I525143);
nand I_30742 (I525072,I525321,I525242);
DFFARX1 I_30743  ( .D(I618081), .CLK(I2702), .RSTB(I525092), .Q(I525366) );
and I_30744 (I525383,I525366,I618090);
DFFARX1 I_30745  ( .D(I525383), .CLK(I2702), .RSTB(I525092), .Q(I525400) );
not I_30746 (I525063,I525400);
nand I_30747 (I525431,I525383,I525321);
and I_30748 (I525448,I525143,I525431);
DFFARX1 I_30749  ( .D(I525448), .CLK(I2702), .RSTB(I525092), .Q(I525054) );
DFFARX1 I_30750  ( .D(I618078), .CLK(I2702), .RSTB(I525092), .Q(I525479) );
nand I_30751 (I525496,I525479,I525143);
and I_30752 (I525513,I525321,I525496);
DFFARX1 I_30753  ( .D(I525513), .CLK(I2702), .RSTB(I525092), .Q(I525084) );
not I_30754 (I525544,I525479);
nor I_30755 (I525561,I525160,I525544);
and I_30756 (I525578,I525479,I525561);
or I_30757 (I525595,I525383,I525578);
DFFARX1 I_30758  ( .D(I525595), .CLK(I2702), .RSTB(I525092), .Q(I525069) );
nand I_30759 (I525066,I525479,I525225);
DFFARX1 I_30760  ( .D(I525479), .CLK(I2702), .RSTB(I525092), .Q(I525057) );
not I_30761 (I525687,I2709);
nand I_30762 (I525704,I453528,I453531);
and I_30763 (I525721,I525704,I453525);
DFFARX1 I_30764  ( .D(I525721), .CLK(I2702), .RSTB(I525687), .Q(I525738) );
nor I_30765 (I525755,I453522,I453531);
nor I_30766 (I525772,I525755,I525738);
not I_30767 (I525670,I525755);
DFFARX1 I_30768  ( .D(I453504), .CLK(I2702), .RSTB(I525687), .Q(I525803) );
not I_30769 (I525820,I525803);
nor I_30770 (I525837,I525755,I525820);
nand I_30771 (I525673,I525803,I525772);
DFFARX1 I_30772  ( .D(I525803), .CLK(I2702), .RSTB(I525687), .Q(I525655) );
nand I_30773 (I525882,I453513,I453510);
and I_30774 (I525899,I525882,I453519);
DFFARX1 I_30775  ( .D(I525899), .CLK(I2702), .RSTB(I525687), .Q(I525916) );
nor I_30776 (I525676,I525916,I525738);
nand I_30777 (I525667,I525916,I525837);
DFFARX1 I_30778  ( .D(I453501), .CLK(I2702), .RSTB(I525687), .Q(I525961) );
and I_30779 (I525978,I525961,I453516);
DFFARX1 I_30780  ( .D(I525978), .CLK(I2702), .RSTB(I525687), .Q(I525995) );
not I_30781 (I525658,I525995);
nand I_30782 (I526026,I525978,I525916);
and I_30783 (I526043,I525738,I526026);
DFFARX1 I_30784  ( .D(I526043), .CLK(I2702), .RSTB(I525687), .Q(I525649) );
DFFARX1 I_30785  ( .D(I453507), .CLK(I2702), .RSTB(I525687), .Q(I526074) );
nand I_30786 (I526091,I526074,I525738);
and I_30787 (I526108,I525916,I526091);
DFFARX1 I_30788  ( .D(I526108), .CLK(I2702), .RSTB(I525687), .Q(I525679) );
not I_30789 (I526139,I526074);
nor I_30790 (I526156,I525755,I526139);
and I_30791 (I526173,I526074,I526156);
or I_30792 (I526190,I525978,I526173);
DFFARX1 I_30793  ( .D(I526190), .CLK(I2702), .RSTB(I525687), .Q(I525664) );
nand I_30794 (I525661,I526074,I525820);
DFFARX1 I_30795  ( .D(I526074), .CLK(I2702), .RSTB(I525687), .Q(I525652) );
not I_30796 (I526282,I2709);
nand I_30797 (I526299,I10008,I10014);
and I_30798 (I526316,I526299,I10011);
DFFARX1 I_30799  ( .D(I526316), .CLK(I2702), .RSTB(I526282), .Q(I526333) );
nor I_30800 (I526350,I10035,I10014);
nor I_30801 (I526367,I526350,I526333);
not I_30802 (I526265,I526350);
DFFARX1 I_30803  ( .D(I10026), .CLK(I2702), .RSTB(I526282), .Q(I526398) );
not I_30804 (I526415,I526398);
nor I_30805 (I526432,I526350,I526415);
nand I_30806 (I526268,I526398,I526367);
DFFARX1 I_30807  ( .D(I526398), .CLK(I2702), .RSTB(I526282), .Q(I526250) );
nand I_30808 (I526477,I10029,I10032);
and I_30809 (I526494,I526477,I10005);
DFFARX1 I_30810  ( .D(I526494), .CLK(I2702), .RSTB(I526282), .Q(I526511) );
nor I_30811 (I526271,I526511,I526333);
nand I_30812 (I526262,I526511,I526432);
DFFARX1 I_30813  ( .D(I10023), .CLK(I2702), .RSTB(I526282), .Q(I526556) );
and I_30814 (I526573,I526556,I10017);
DFFARX1 I_30815  ( .D(I526573), .CLK(I2702), .RSTB(I526282), .Q(I526590) );
not I_30816 (I526253,I526590);
nand I_30817 (I526621,I526573,I526511);
and I_30818 (I526638,I526333,I526621);
DFFARX1 I_30819  ( .D(I526638), .CLK(I2702), .RSTB(I526282), .Q(I526244) );
DFFARX1 I_30820  ( .D(I10020), .CLK(I2702), .RSTB(I526282), .Q(I526669) );
nand I_30821 (I526686,I526669,I526333);
and I_30822 (I526703,I526511,I526686);
DFFARX1 I_30823  ( .D(I526703), .CLK(I2702), .RSTB(I526282), .Q(I526274) );
not I_30824 (I526734,I526669);
nor I_30825 (I526751,I526350,I526734);
and I_30826 (I526768,I526669,I526751);
or I_30827 (I526785,I526573,I526768);
DFFARX1 I_30828  ( .D(I526785), .CLK(I2702), .RSTB(I526282), .Q(I526259) );
nand I_30829 (I526256,I526669,I526415);
DFFARX1 I_30830  ( .D(I526669), .CLK(I2702), .RSTB(I526282), .Q(I526247) );
not I_30831 (I526877,I2709);
nand I_30832 (I526894,I410679,I410691);
and I_30833 (I526911,I526894,I410673);
DFFARX1 I_30834  ( .D(I526911), .CLK(I2702), .RSTB(I526877), .Q(I526928) );
nor I_30835 (I526945,I410685,I410691);
nor I_30836 (I526962,I526945,I526928);
not I_30837 (I526860,I526945);
DFFARX1 I_30838  ( .D(I410670), .CLK(I2702), .RSTB(I526877), .Q(I526993) );
not I_30839 (I527010,I526993);
nor I_30840 (I527027,I526945,I527010);
nand I_30841 (I526863,I526993,I526962);
DFFARX1 I_30842  ( .D(I526993), .CLK(I2702), .RSTB(I526877), .Q(I526845) );
nand I_30843 (I527072,I410661,I410676);
and I_30844 (I527089,I527072,I410667);
DFFARX1 I_30845  ( .D(I527089), .CLK(I2702), .RSTB(I526877), .Q(I527106) );
nor I_30846 (I526866,I527106,I526928);
nand I_30847 (I526857,I527106,I527027);
DFFARX1 I_30848  ( .D(I410688), .CLK(I2702), .RSTB(I526877), .Q(I527151) );
and I_30849 (I527168,I527151,I410682);
DFFARX1 I_30850  ( .D(I527168), .CLK(I2702), .RSTB(I526877), .Q(I527185) );
not I_30851 (I526848,I527185);
nand I_30852 (I527216,I527168,I527106);
and I_30853 (I527233,I526928,I527216);
DFFARX1 I_30854  ( .D(I527233), .CLK(I2702), .RSTB(I526877), .Q(I526839) );
DFFARX1 I_30855  ( .D(I410664), .CLK(I2702), .RSTB(I526877), .Q(I527264) );
nand I_30856 (I527281,I527264,I526928);
and I_30857 (I527298,I527106,I527281);
DFFARX1 I_30858  ( .D(I527298), .CLK(I2702), .RSTB(I526877), .Q(I526869) );
not I_30859 (I527329,I527264);
nor I_30860 (I527346,I526945,I527329);
and I_30861 (I527363,I527264,I527346);
or I_30862 (I527380,I527168,I527363);
DFFARX1 I_30863  ( .D(I527380), .CLK(I2702), .RSTB(I526877), .Q(I526854) );
nand I_30864 (I526851,I527264,I527010);
DFFARX1 I_30865  ( .D(I527264), .CLK(I2702), .RSTB(I526877), .Q(I526842) );
not I_30866 (I527472,I2709);
nand I_30867 (I527489,I593494,I593485);
and I_30868 (I527506,I527489,I593503);
DFFARX1 I_30869  ( .D(I527506), .CLK(I2702), .RSTB(I527472), .Q(I527523) );
nor I_30870 (I527540,I593482,I593485);
nor I_30871 (I527557,I527540,I527523);
not I_30872 (I527455,I527540);
DFFARX1 I_30873  ( .D(I593491), .CLK(I2702), .RSTB(I527472), .Q(I527588) );
not I_30874 (I527605,I527588);
nor I_30875 (I527622,I527540,I527605);
nand I_30876 (I527458,I527588,I527557);
DFFARX1 I_30877  ( .D(I527588), .CLK(I2702), .RSTB(I527472), .Q(I527440) );
nand I_30878 (I527667,I593506,I593488);
and I_30879 (I527684,I527667,I593509);
DFFARX1 I_30880  ( .D(I527684), .CLK(I2702), .RSTB(I527472), .Q(I527701) );
nor I_30881 (I527461,I527701,I527523);
nand I_30882 (I527452,I527701,I527622);
DFFARX1 I_30883  ( .D(I593497), .CLK(I2702), .RSTB(I527472), .Q(I527746) );
and I_30884 (I527763,I527746,I593479);
DFFARX1 I_30885  ( .D(I527763), .CLK(I2702), .RSTB(I527472), .Q(I527780) );
not I_30886 (I527443,I527780);
nand I_30887 (I527811,I527763,I527701);
and I_30888 (I527828,I527523,I527811);
DFFARX1 I_30889  ( .D(I527828), .CLK(I2702), .RSTB(I527472), .Q(I527434) );
DFFARX1 I_30890  ( .D(I593500), .CLK(I2702), .RSTB(I527472), .Q(I527859) );
nand I_30891 (I527876,I527859,I527523);
and I_30892 (I527893,I527701,I527876);
DFFARX1 I_30893  ( .D(I527893), .CLK(I2702), .RSTB(I527472), .Q(I527464) );
not I_30894 (I527924,I527859);
nor I_30895 (I527941,I527540,I527924);
and I_30896 (I527958,I527859,I527941);
or I_30897 (I527975,I527763,I527958);
DFFARX1 I_30898  ( .D(I527975), .CLK(I2702), .RSTB(I527472), .Q(I527449) );
nand I_30899 (I527446,I527859,I527605);
DFFARX1 I_30900  ( .D(I527859), .CLK(I2702), .RSTB(I527472), .Q(I527437) );
not I_30901 (I528067,I2709);
nand I_30902 (I528084,I360937,I360949);
and I_30903 (I528101,I528084,I360931);
DFFARX1 I_30904  ( .D(I528101), .CLK(I2702), .RSTB(I528067), .Q(I528118) );
nor I_30905 (I528135,I360943,I360949);
nor I_30906 (I528152,I528135,I528118);
not I_30907 (I528050,I528135);
DFFARX1 I_30908  ( .D(I360928), .CLK(I2702), .RSTB(I528067), .Q(I528183) );
not I_30909 (I528200,I528183);
nor I_30910 (I528217,I528135,I528200);
nand I_30911 (I528053,I528183,I528152);
DFFARX1 I_30912  ( .D(I528183), .CLK(I2702), .RSTB(I528067), .Q(I528035) );
nand I_30913 (I528262,I360919,I360934);
and I_30914 (I528279,I528262,I360925);
DFFARX1 I_30915  ( .D(I528279), .CLK(I2702), .RSTB(I528067), .Q(I528296) );
nor I_30916 (I528056,I528296,I528118);
nand I_30917 (I528047,I528296,I528217);
DFFARX1 I_30918  ( .D(I360946), .CLK(I2702), .RSTB(I528067), .Q(I528341) );
and I_30919 (I528358,I528341,I360940);
DFFARX1 I_30920  ( .D(I528358), .CLK(I2702), .RSTB(I528067), .Q(I528375) );
not I_30921 (I528038,I528375);
nand I_30922 (I528406,I528358,I528296);
and I_30923 (I528423,I528118,I528406);
DFFARX1 I_30924  ( .D(I528423), .CLK(I2702), .RSTB(I528067), .Q(I528029) );
DFFARX1 I_30925  ( .D(I360922), .CLK(I2702), .RSTB(I528067), .Q(I528454) );
nand I_30926 (I528471,I528454,I528118);
and I_30927 (I528488,I528296,I528471);
DFFARX1 I_30928  ( .D(I528488), .CLK(I2702), .RSTB(I528067), .Q(I528059) );
not I_30929 (I528519,I528454);
nor I_30930 (I528536,I528135,I528519);
and I_30931 (I528553,I528454,I528536);
or I_30932 (I528570,I528358,I528553);
DFFARX1 I_30933  ( .D(I528570), .CLK(I2702), .RSTB(I528067), .Q(I528044) );
nand I_30934 (I528041,I528454,I528200);
DFFARX1 I_30935  ( .D(I528454), .CLK(I2702), .RSTB(I528067), .Q(I528032) );
not I_30936 (I528662,I2709);
nand I_30937 (I528679,I603609,I603600);
and I_30938 (I528696,I528679,I603618);
DFFARX1 I_30939  ( .D(I528696), .CLK(I2702), .RSTB(I528662), .Q(I528713) );
nor I_30940 (I528730,I603597,I603600);
nor I_30941 (I528747,I528730,I528713);
not I_30942 (I528645,I528730);
DFFARX1 I_30943  ( .D(I603606), .CLK(I2702), .RSTB(I528662), .Q(I528778) );
not I_30944 (I528795,I528778);
nor I_30945 (I528812,I528730,I528795);
nand I_30946 (I528648,I528778,I528747);
DFFARX1 I_30947  ( .D(I528778), .CLK(I2702), .RSTB(I528662), .Q(I528630) );
nand I_30948 (I528857,I603621,I603603);
and I_30949 (I528874,I528857,I603624);
DFFARX1 I_30950  ( .D(I528874), .CLK(I2702), .RSTB(I528662), .Q(I528891) );
nor I_30951 (I528651,I528891,I528713);
nand I_30952 (I528642,I528891,I528812);
DFFARX1 I_30953  ( .D(I603612), .CLK(I2702), .RSTB(I528662), .Q(I528936) );
and I_30954 (I528953,I528936,I603594);
DFFARX1 I_30955  ( .D(I528953), .CLK(I2702), .RSTB(I528662), .Q(I528970) );
not I_30956 (I528633,I528970);
nand I_30957 (I529001,I528953,I528891);
and I_30958 (I529018,I528713,I529001);
DFFARX1 I_30959  ( .D(I529018), .CLK(I2702), .RSTB(I528662), .Q(I528624) );
DFFARX1 I_30960  ( .D(I603615), .CLK(I2702), .RSTB(I528662), .Q(I529049) );
nand I_30961 (I529066,I529049,I528713);
and I_30962 (I529083,I528891,I529066);
DFFARX1 I_30963  ( .D(I529083), .CLK(I2702), .RSTB(I528662), .Q(I528654) );
not I_30964 (I529114,I529049);
nor I_30965 (I529131,I528730,I529114);
and I_30966 (I529148,I529049,I529131);
or I_30967 (I529165,I528953,I529148);
DFFARX1 I_30968  ( .D(I529165), .CLK(I2702), .RSTB(I528662), .Q(I528639) );
nand I_30969 (I528636,I529049,I528795);
DFFARX1 I_30970  ( .D(I529049), .CLK(I2702), .RSTB(I528662), .Q(I528627) );
not I_30971 (I529257,I2709);
nand I_30972 (I529274,I494396,I494369);
and I_30973 (I529291,I529274,I494372);
DFFARX1 I_30974  ( .D(I529291), .CLK(I2702), .RSTB(I529257), .Q(I529308) );
nor I_30975 (I529325,I494381,I494369);
nor I_30976 (I529342,I529325,I529308);
not I_30977 (I529240,I529325);
DFFARX1 I_30978  ( .D(I494378), .CLK(I2702), .RSTB(I529257), .Q(I529373) );
not I_30979 (I529390,I529373);
nor I_30980 (I529407,I529325,I529390);
nand I_30981 (I529243,I529373,I529342);
DFFARX1 I_30982  ( .D(I529373), .CLK(I2702), .RSTB(I529257), .Q(I529225) );
nand I_30983 (I529452,I494375,I494384);
and I_30984 (I529469,I529452,I494393);
DFFARX1 I_30985  ( .D(I529469), .CLK(I2702), .RSTB(I529257), .Q(I529486) );
nor I_30986 (I529246,I529486,I529308);
nand I_30987 (I529237,I529486,I529407);
DFFARX1 I_30988  ( .D(I494399), .CLK(I2702), .RSTB(I529257), .Q(I529531) );
and I_30989 (I529548,I529531,I494390);
DFFARX1 I_30990  ( .D(I529548), .CLK(I2702), .RSTB(I529257), .Q(I529565) );
not I_30991 (I529228,I529565);
nand I_30992 (I529596,I529548,I529486);
and I_30993 (I529613,I529308,I529596);
DFFARX1 I_30994  ( .D(I529613), .CLK(I2702), .RSTB(I529257), .Q(I529219) );
DFFARX1 I_30995  ( .D(I494387), .CLK(I2702), .RSTB(I529257), .Q(I529644) );
nand I_30996 (I529661,I529644,I529308);
and I_30997 (I529678,I529486,I529661);
DFFARX1 I_30998  ( .D(I529678), .CLK(I2702), .RSTB(I529257), .Q(I529249) );
not I_30999 (I529709,I529644);
nor I_31000 (I529726,I529325,I529709);
and I_31001 (I529743,I529644,I529726);
or I_31002 (I529760,I529548,I529743);
DFFARX1 I_31003  ( .D(I529760), .CLK(I2702), .RSTB(I529257), .Q(I529234) );
nand I_31004 (I529231,I529644,I529390);
DFFARX1 I_31005  ( .D(I529644), .CLK(I2702), .RSTB(I529257), .Q(I529222) );
not I_31006 (I529852,I2709);
nand I_31007 (I529869,I135678,I135690);
and I_31008 (I529886,I529869,I135699);
DFFARX1 I_31009  ( .D(I529886), .CLK(I2702), .RSTB(I529852), .Q(I529903) );
nor I_31010 (I529920,I135693,I135690);
nor I_31011 (I529937,I529920,I529903);
not I_31012 (I529835,I529920);
DFFARX1 I_31013  ( .D(I135687), .CLK(I2702), .RSTB(I529852), .Q(I529968) );
not I_31014 (I529985,I529968);
nor I_31015 (I530002,I529920,I529985);
nand I_31016 (I529838,I529968,I529937);
DFFARX1 I_31017  ( .D(I529968), .CLK(I2702), .RSTB(I529852), .Q(I529820) );
nand I_31018 (I530047,I135684,I135681);
and I_31019 (I530064,I530047,I135672);
DFFARX1 I_31020  ( .D(I530064), .CLK(I2702), .RSTB(I529852), .Q(I530081) );
nor I_31021 (I529841,I530081,I529903);
nand I_31022 (I529832,I530081,I530002);
DFFARX1 I_31023  ( .D(I135696), .CLK(I2702), .RSTB(I529852), .Q(I530126) );
and I_31024 (I530143,I530126,I135675);
DFFARX1 I_31025  ( .D(I530143), .CLK(I2702), .RSTB(I529852), .Q(I530160) );
not I_31026 (I529823,I530160);
nand I_31027 (I530191,I530143,I530081);
and I_31028 (I530208,I529903,I530191);
DFFARX1 I_31029  ( .D(I530208), .CLK(I2702), .RSTB(I529852), .Q(I529814) );
DFFARX1 I_31030  ( .D(I135669), .CLK(I2702), .RSTB(I529852), .Q(I530239) );
nand I_31031 (I530256,I530239,I529903);
and I_31032 (I530273,I530081,I530256);
DFFARX1 I_31033  ( .D(I530273), .CLK(I2702), .RSTB(I529852), .Q(I529844) );
not I_31034 (I530304,I530239);
nor I_31035 (I530321,I529920,I530304);
and I_31036 (I530338,I530239,I530321);
or I_31037 (I530355,I530143,I530338);
DFFARX1 I_31038  ( .D(I530355), .CLK(I2702), .RSTB(I529852), .Q(I529829) );
nand I_31039 (I529826,I530239,I529985);
DFFARX1 I_31040  ( .D(I530239), .CLK(I2702), .RSTB(I529852), .Q(I529817) );
not I_31041 (I530447,I2709);
nand I_31042 (I530464,I27960,I27966);
and I_31043 (I530481,I530464,I27963);
DFFARX1 I_31044  ( .D(I530481), .CLK(I2702), .RSTB(I530447), .Q(I530498) );
nor I_31045 (I530515,I27987,I27966);
nor I_31046 (I530532,I530515,I530498);
not I_31047 (I530430,I530515);
DFFARX1 I_31048  ( .D(I27978), .CLK(I2702), .RSTB(I530447), .Q(I530563) );
not I_31049 (I530580,I530563);
nor I_31050 (I530597,I530515,I530580);
nand I_31051 (I530433,I530563,I530532);
DFFARX1 I_31052  ( .D(I530563), .CLK(I2702), .RSTB(I530447), .Q(I530415) );
nand I_31053 (I530642,I27981,I27984);
and I_31054 (I530659,I530642,I27957);
DFFARX1 I_31055  ( .D(I530659), .CLK(I2702), .RSTB(I530447), .Q(I530676) );
nor I_31056 (I530436,I530676,I530498);
nand I_31057 (I530427,I530676,I530597);
DFFARX1 I_31058  ( .D(I27975), .CLK(I2702), .RSTB(I530447), .Q(I530721) );
and I_31059 (I530738,I530721,I27969);
DFFARX1 I_31060  ( .D(I530738), .CLK(I2702), .RSTB(I530447), .Q(I530755) );
not I_31061 (I530418,I530755);
nand I_31062 (I530786,I530738,I530676);
and I_31063 (I530803,I530498,I530786);
DFFARX1 I_31064  ( .D(I530803), .CLK(I2702), .RSTB(I530447), .Q(I530409) );
DFFARX1 I_31065  ( .D(I27972), .CLK(I2702), .RSTB(I530447), .Q(I530834) );
nand I_31066 (I530851,I530834,I530498);
and I_31067 (I530868,I530676,I530851);
DFFARX1 I_31068  ( .D(I530868), .CLK(I2702), .RSTB(I530447), .Q(I530439) );
not I_31069 (I530899,I530834);
nor I_31070 (I530916,I530515,I530899);
and I_31071 (I530933,I530834,I530916);
or I_31072 (I530950,I530738,I530933);
DFFARX1 I_31073  ( .D(I530950), .CLK(I2702), .RSTB(I530447), .Q(I530424) );
nand I_31074 (I530421,I530834,I530580);
DFFARX1 I_31075  ( .D(I530834), .CLK(I2702), .RSTB(I530447), .Q(I530412) );
not I_31076 (I531042,I2709);
nand I_31077 (I531059,I58158,I58170);
and I_31078 (I531076,I531059,I58179);
DFFARX1 I_31079  ( .D(I531076), .CLK(I2702), .RSTB(I531042), .Q(I531093) );
nor I_31080 (I531110,I58173,I58170);
nor I_31081 (I531127,I531110,I531093);
not I_31082 (I531025,I531110);
DFFARX1 I_31083  ( .D(I58167), .CLK(I2702), .RSTB(I531042), .Q(I531158) );
not I_31084 (I531175,I531158);
nor I_31085 (I531192,I531110,I531175);
nand I_31086 (I531028,I531158,I531127);
DFFARX1 I_31087  ( .D(I531158), .CLK(I2702), .RSTB(I531042), .Q(I531010) );
nand I_31088 (I531237,I58164,I58161);
and I_31089 (I531254,I531237,I58152);
DFFARX1 I_31090  ( .D(I531254), .CLK(I2702), .RSTB(I531042), .Q(I531271) );
nor I_31091 (I531031,I531271,I531093);
nand I_31092 (I531022,I531271,I531192);
DFFARX1 I_31093  ( .D(I58176), .CLK(I2702), .RSTB(I531042), .Q(I531316) );
and I_31094 (I531333,I531316,I58155);
DFFARX1 I_31095  ( .D(I531333), .CLK(I2702), .RSTB(I531042), .Q(I531350) );
not I_31096 (I531013,I531350);
nand I_31097 (I531381,I531333,I531271);
and I_31098 (I531398,I531093,I531381);
DFFARX1 I_31099  ( .D(I531398), .CLK(I2702), .RSTB(I531042), .Q(I531004) );
DFFARX1 I_31100  ( .D(I58149), .CLK(I2702), .RSTB(I531042), .Q(I531429) );
nand I_31101 (I531446,I531429,I531093);
and I_31102 (I531463,I531271,I531446);
DFFARX1 I_31103  ( .D(I531463), .CLK(I2702), .RSTB(I531042), .Q(I531034) );
not I_31104 (I531494,I531429);
nor I_31105 (I531511,I531110,I531494);
and I_31106 (I531528,I531429,I531511);
or I_31107 (I531545,I531333,I531528);
DFFARX1 I_31108  ( .D(I531545), .CLK(I2702), .RSTB(I531042), .Q(I531019) );
nand I_31109 (I531016,I531429,I531175);
DFFARX1 I_31110  ( .D(I531429), .CLK(I2702), .RSTB(I531042), .Q(I531007) );
not I_31111 (I531637,I2709);
nand I_31112 (I531654,I451216,I451219);
and I_31113 (I531671,I531654,I451213);
DFFARX1 I_31114  ( .D(I531671), .CLK(I2702), .RSTB(I531637), .Q(I531688) );
nor I_31115 (I531705,I451210,I451219);
nor I_31116 (I531722,I531705,I531688);
not I_31117 (I531620,I531705);
DFFARX1 I_31118  ( .D(I451192), .CLK(I2702), .RSTB(I531637), .Q(I531753) );
not I_31119 (I531770,I531753);
nor I_31120 (I531787,I531705,I531770);
nand I_31121 (I531623,I531753,I531722);
DFFARX1 I_31122  ( .D(I531753), .CLK(I2702), .RSTB(I531637), .Q(I531605) );
nand I_31123 (I531832,I451201,I451198);
and I_31124 (I531849,I531832,I451207);
DFFARX1 I_31125  ( .D(I531849), .CLK(I2702), .RSTB(I531637), .Q(I531866) );
nor I_31126 (I531626,I531866,I531688);
nand I_31127 (I531617,I531866,I531787);
DFFARX1 I_31128  ( .D(I451189), .CLK(I2702), .RSTB(I531637), .Q(I531911) );
and I_31129 (I531928,I531911,I451204);
DFFARX1 I_31130  ( .D(I531928), .CLK(I2702), .RSTB(I531637), .Q(I531945) );
not I_31131 (I531608,I531945);
nand I_31132 (I531976,I531928,I531866);
and I_31133 (I531993,I531688,I531976);
DFFARX1 I_31134  ( .D(I531993), .CLK(I2702), .RSTB(I531637), .Q(I531599) );
DFFARX1 I_31135  ( .D(I451195), .CLK(I2702), .RSTB(I531637), .Q(I532024) );
nand I_31136 (I532041,I532024,I531688);
and I_31137 (I532058,I531866,I532041);
DFFARX1 I_31138  ( .D(I532058), .CLK(I2702), .RSTB(I531637), .Q(I531629) );
not I_31139 (I532089,I532024);
nor I_31140 (I532106,I531705,I532089);
and I_31141 (I532123,I532024,I532106);
or I_31142 (I532140,I531928,I532123);
DFFARX1 I_31143  ( .D(I532140), .CLK(I2702), .RSTB(I531637), .Q(I531614) );
nand I_31144 (I531611,I532024,I531770);
DFFARX1 I_31145  ( .D(I532024), .CLK(I2702), .RSTB(I531637), .Q(I531602) );
not I_31146 (I532232,I2709);
nand I_31147 (I532249,I83352,I83364);
and I_31148 (I532266,I532249,I83373);
DFFARX1 I_31149  ( .D(I532266), .CLK(I2702), .RSTB(I532232), .Q(I532283) );
nor I_31150 (I532300,I83367,I83364);
nor I_31151 (I532317,I532300,I532283);
not I_31152 (I532215,I532300);
DFFARX1 I_31153  ( .D(I83361), .CLK(I2702), .RSTB(I532232), .Q(I532348) );
not I_31154 (I532365,I532348);
nor I_31155 (I532382,I532300,I532365);
nand I_31156 (I532218,I532348,I532317);
DFFARX1 I_31157  ( .D(I532348), .CLK(I2702), .RSTB(I532232), .Q(I532200) );
nand I_31158 (I532427,I83358,I83355);
and I_31159 (I532444,I532427,I83346);
DFFARX1 I_31160  ( .D(I532444), .CLK(I2702), .RSTB(I532232), .Q(I532461) );
nor I_31161 (I532221,I532461,I532283);
nand I_31162 (I532212,I532461,I532382);
DFFARX1 I_31163  ( .D(I83370), .CLK(I2702), .RSTB(I532232), .Q(I532506) );
and I_31164 (I532523,I532506,I83349);
DFFARX1 I_31165  ( .D(I532523), .CLK(I2702), .RSTB(I532232), .Q(I532540) );
not I_31166 (I532203,I532540);
nand I_31167 (I532571,I532523,I532461);
and I_31168 (I532588,I532283,I532571);
DFFARX1 I_31169  ( .D(I532588), .CLK(I2702), .RSTB(I532232), .Q(I532194) );
DFFARX1 I_31170  ( .D(I83343), .CLK(I2702), .RSTB(I532232), .Q(I532619) );
nand I_31171 (I532636,I532619,I532283);
and I_31172 (I532653,I532461,I532636);
DFFARX1 I_31173  ( .D(I532653), .CLK(I2702), .RSTB(I532232), .Q(I532224) );
not I_31174 (I532684,I532619);
nor I_31175 (I532701,I532300,I532684);
and I_31176 (I532718,I532619,I532701);
or I_31177 (I532735,I532523,I532718);
DFFARX1 I_31178  ( .D(I532735), .CLK(I2702), .RSTB(I532232), .Q(I532209) );
nand I_31179 (I532206,I532619,I532365);
DFFARX1 I_31180  ( .D(I532619), .CLK(I2702), .RSTB(I532232), .Q(I532197) );
not I_31181 (I532827,I2709);
nand I_31182 (I532844,I405511,I405523);
and I_31183 (I532861,I532844,I405505);
DFFARX1 I_31184  ( .D(I532861), .CLK(I2702), .RSTB(I532827), .Q(I532878) );
nor I_31185 (I532895,I405517,I405523);
nor I_31186 (I532912,I532895,I532878);
not I_31187 (I532810,I532895);
DFFARX1 I_31188  ( .D(I405502), .CLK(I2702), .RSTB(I532827), .Q(I532943) );
not I_31189 (I532960,I532943);
nor I_31190 (I532977,I532895,I532960);
nand I_31191 (I532813,I532943,I532912);
DFFARX1 I_31192  ( .D(I532943), .CLK(I2702), .RSTB(I532827), .Q(I532795) );
nand I_31193 (I533022,I405493,I405508);
and I_31194 (I533039,I533022,I405499);
DFFARX1 I_31195  ( .D(I533039), .CLK(I2702), .RSTB(I532827), .Q(I533056) );
nor I_31196 (I532816,I533056,I532878);
nand I_31197 (I532807,I533056,I532977);
DFFARX1 I_31198  ( .D(I405520), .CLK(I2702), .RSTB(I532827), .Q(I533101) );
and I_31199 (I533118,I533101,I405514);
DFFARX1 I_31200  ( .D(I533118), .CLK(I2702), .RSTB(I532827), .Q(I533135) );
not I_31201 (I532798,I533135);
nand I_31202 (I533166,I533118,I533056);
and I_31203 (I533183,I532878,I533166);
DFFARX1 I_31204  ( .D(I533183), .CLK(I2702), .RSTB(I532827), .Q(I532789) );
DFFARX1 I_31205  ( .D(I405496), .CLK(I2702), .RSTB(I532827), .Q(I533214) );
nand I_31206 (I533231,I533214,I532878);
and I_31207 (I533248,I533056,I533231);
DFFARX1 I_31208  ( .D(I533248), .CLK(I2702), .RSTB(I532827), .Q(I532819) );
not I_31209 (I533279,I533214);
nor I_31210 (I533296,I532895,I533279);
and I_31211 (I533313,I533214,I533296);
or I_31212 (I533330,I533118,I533313);
DFFARX1 I_31213  ( .D(I533330), .CLK(I2702), .RSTB(I532827), .Q(I532804) );
nand I_31214 (I532801,I533214,I532960);
DFFARX1 I_31215  ( .D(I533214), .CLK(I2702), .RSTB(I532827), .Q(I532792) );
not I_31216 (I533422,I2709);
nand I_31217 (I533439,I2263,I2695);
and I_31218 (I533456,I533439,I1239);
DFFARX1 I_31219  ( .D(I533456), .CLK(I2702), .RSTB(I533422), .Q(I533473) );
nor I_31220 (I533490,I2359,I2695);
nor I_31221 (I533507,I533490,I533473);
not I_31222 (I533405,I533490);
DFFARX1 I_31223  ( .D(I1767), .CLK(I2702), .RSTB(I533422), .Q(I533538) );
not I_31224 (I533555,I533538);
nor I_31225 (I533572,I533490,I533555);
nand I_31226 (I533408,I533538,I533507);
DFFARX1 I_31227  ( .D(I533538), .CLK(I2702), .RSTB(I533422), .Q(I533390) );
nand I_31228 (I533617,I1815,I1511);
and I_31229 (I533634,I533617,I1711);
DFFARX1 I_31230  ( .D(I533634), .CLK(I2702), .RSTB(I533422), .Q(I533651) );
nor I_31231 (I533411,I533651,I533473);
nand I_31232 (I533402,I533651,I533572);
DFFARX1 I_31233  ( .D(I1639), .CLK(I2702), .RSTB(I533422), .Q(I533696) );
and I_31234 (I533713,I533696,I2567);
DFFARX1 I_31235  ( .D(I533713), .CLK(I2702), .RSTB(I533422), .Q(I533730) );
not I_31236 (I533393,I533730);
nand I_31237 (I533761,I533713,I533651);
and I_31238 (I533778,I533473,I533761);
DFFARX1 I_31239  ( .D(I533778), .CLK(I2702), .RSTB(I533422), .Q(I533384) );
DFFARX1 I_31240  ( .D(I1407), .CLK(I2702), .RSTB(I533422), .Q(I533809) );
nand I_31241 (I533826,I533809,I533473);
and I_31242 (I533843,I533651,I533826);
DFFARX1 I_31243  ( .D(I533843), .CLK(I2702), .RSTB(I533422), .Q(I533414) );
not I_31244 (I533874,I533809);
nor I_31245 (I533891,I533490,I533874);
and I_31246 (I533908,I533809,I533891);
or I_31247 (I533925,I533713,I533908);
DFFARX1 I_31248  ( .D(I533925), .CLK(I2702), .RSTB(I533422), .Q(I533399) );
nand I_31249 (I533396,I533809,I533555);
DFFARX1 I_31250  ( .D(I533809), .CLK(I2702), .RSTB(I533422), .Q(I533387) );
not I_31251 (I534017,I2709);
nand I_31252 (I534034,I436766,I436769);
and I_31253 (I534051,I534034,I436763);
DFFARX1 I_31254  ( .D(I534051), .CLK(I2702), .RSTB(I534017), .Q(I534068) );
nor I_31255 (I534085,I436760,I436769);
nor I_31256 (I534102,I534085,I534068);
not I_31257 (I534000,I534085);
DFFARX1 I_31258  ( .D(I436742), .CLK(I2702), .RSTB(I534017), .Q(I534133) );
not I_31259 (I534150,I534133);
nor I_31260 (I534167,I534085,I534150);
nand I_31261 (I534003,I534133,I534102);
DFFARX1 I_31262  ( .D(I534133), .CLK(I2702), .RSTB(I534017), .Q(I533985) );
nand I_31263 (I534212,I436751,I436748);
and I_31264 (I534229,I534212,I436757);
DFFARX1 I_31265  ( .D(I534229), .CLK(I2702), .RSTB(I534017), .Q(I534246) );
nor I_31266 (I534006,I534246,I534068);
nand I_31267 (I533997,I534246,I534167);
DFFARX1 I_31268  ( .D(I436739), .CLK(I2702), .RSTB(I534017), .Q(I534291) );
and I_31269 (I534308,I534291,I436754);
DFFARX1 I_31270  ( .D(I534308), .CLK(I2702), .RSTB(I534017), .Q(I534325) );
not I_31271 (I533988,I534325);
nand I_31272 (I534356,I534308,I534246);
and I_31273 (I534373,I534068,I534356);
DFFARX1 I_31274  ( .D(I534373), .CLK(I2702), .RSTB(I534017), .Q(I533979) );
DFFARX1 I_31275  ( .D(I436745), .CLK(I2702), .RSTB(I534017), .Q(I534404) );
nand I_31276 (I534421,I534404,I534068);
and I_31277 (I534438,I534246,I534421);
DFFARX1 I_31278  ( .D(I534438), .CLK(I2702), .RSTB(I534017), .Q(I534009) );
not I_31279 (I534469,I534404);
nor I_31280 (I534486,I534085,I534469);
and I_31281 (I534503,I534404,I534486);
or I_31282 (I534520,I534308,I534503);
DFFARX1 I_31283  ( .D(I534520), .CLK(I2702), .RSTB(I534017), .Q(I533994) );
nand I_31284 (I533991,I534404,I534150);
DFFARX1 I_31285  ( .D(I534404), .CLK(I2702), .RSTB(I534017), .Q(I533982) );
not I_31286 (I534612,I2709);
nand I_31287 (I534629,I246306,I246312);
and I_31288 (I534646,I534629,I246294);
DFFARX1 I_31289  ( .D(I534646), .CLK(I2702), .RSTB(I534612), .Q(I534663) );
nor I_31290 (I534680,I246288,I246312);
nor I_31291 (I534697,I534680,I534663);
not I_31292 (I534595,I534680);
DFFARX1 I_31293  ( .D(I246318), .CLK(I2702), .RSTB(I534612), .Q(I534728) );
not I_31294 (I534745,I534728);
nor I_31295 (I534762,I534680,I534745);
nand I_31296 (I534598,I534728,I534697);
DFFARX1 I_31297  ( .D(I534728), .CLK(I2702), .RSTB(I534612), .Q(I534580) );
nand I_31298 (I534807,I246309,I246300);
and I_31299 (I534824,I534807,I246303);
DFFARX1 I_31300  ( .D(I534824), .CLK(I2702), .RSTB(I534612), .Q(I534841) );
nor I_31301 (I534601,I534841,I534663);
nand I_31302 (I534592,I534841,I534762);
DFFARX1 I_31303  ( .D(I246315), .CLK(I2702), .RSTB(I534612), .Q(I534886) );
and I_31304 (I534903,I534886,I246291);
DFFARX1 I_31305  ( .D(I534903), .CLK(I2702), .RSTB(I534612), .Q(I534920) );
not I_31306 (I534583,I534920);
nand I_31307 (I534951,I534903,I534841);
and I_31308 (I534968,I534663,I534951);
DFFARX1 I_31309  ( .D(I534968), .CLK(I2702), .RSTB(I534612), .Q(I534574) );
DFFARX1 I_31310  ( .D(I246297), .CLK(I2702), .RSTB(I534612), .Q(I534999) );
nand I_31311 (I535016,I534999,I534663);
and I_31312 (I535033,I534841,I535016);
DFFARX1 I_31313  ( .D(I535033), .CLK(I2702), .RSTB(I534612), .Q(I534604) );
not I_31314 (I535064,I534999);
nor I_31315 (I535081,I534680,I535064);
and I_31316 (I535098,I534999,I535081);
or I_31317 (I535115,I534903,I535098);
DFFARX1 I_31318  ( .D(I535115), .CLK(I2702), .RSTB(I534612), .Q(I534589) );
nand I_31319 (I534586,I534999,I534745);
DFFARX1 I_31320  ( .D(I534999), .CLK(I2702), .RSTB(I534612), .Q(I534577) );
not I_31321 (I535207,I2709);
nand I_31322 (I535224,I140889,I140901);
and I_31323 (I535241,I535224,I140880);
DFFARX1 I_31324  ( .D(I535241), .CLK(I2702), .RSTB(I535207), .Q(I535258) );
nor I_31325 (I535275,I140871,I140901);
nor I_31326 (I535292,I535275,I535258);
not I_31327 (I535190,I535275);
DFFARX1 I_31328  ( .D(I140883), .CLK(I2702), .RSTB(I535207), .Q(I535323) );
not I_31329 (I535340,I535323);
nor I_31330 (I535357,I535275,I535340);
nand I_31331 (I535193,I535323,I535292);
DFFARX1 I_31332  ( .D(I535323), .CLK(I2702), .RSTB(I535207), .Q(I535175) );
nand I_31333 (I535402,I140898,I140886);
and I_31334 (I535419,I535402,I140874);
DFFARX1 I_31335  ( .D(I535419), .CLK(I2702), .RSTB(I535207), .Q(I535436) );
nor I_31336 (I535196,I535436,I535258);
nand I_31337 (I535187,I535436,I535357);
DFFARX1 I_31338  ( .D(I140892), .CLK(I2702), .RSTB(I535207), .Q(I535481) );
and I_31339 (I535498,I535481,I140877);
DFFARX1 I_31340  ( .D(I535498), .CLK(I2702), .RSTB(I535207), .Q(I535515) );
not I_31341 (I535178,I535515);
nand I_31342 (I535546,I535498,I535436);
and I_31343 (I535563,I535258,I535546);
DFFARX1 I_31344  ( .D(I535563), .CLK(I2702), .RSTB(I535207), .Q(I535169) );
DFFARX1 I_31345  ( .D(I140895), .CLK(I2702), .RSTB(I535207), .Q(I535594) );
nand I_31346 (I535611,I535594,I535258);
and I_31347 (I535628,I535436,I535611);
DFFARX1 I_31348  ( .D(I535628), .CLK(I2702), .RSTB(I535207), .Q(I535199) );
not I_31349 (I535659,I535594);
nor I_31350 (I535676,I535275,I535659);
and I_31351 (I535693,I535594,I535676);
or I_31352 (I535710,I535498,I535693);
DFFARX1 I_31353  ( .D(I535710), .CLK(I2702), .RSTB(I535207), .Q(I535184) );
nand I_31354 (I535181,I535594,I535340);
DFFARX1 I_31355  ( .D(I535594), .CLK(I2702), .RSTB(I535207), .Q(I535172) );
not I_31356 (I535802,I2709);
nand I_31357 (I535819,I32448,I32454);
and I_31358 (I535836,I535819,I32451);
DFFARX1 I_31359  ( .D(I535836), .CLK(I2702), .RSTB(I535802), .Q(I535853) );
nor I_31360 (I535870,I32475,I32454);
nor I_31361 (I535887,I535870,I535853);
not I_31362 (I535785,I535870);
DFFARX1 I_31363  ( .D(I32466), .CLK(I2702), .RSTB(I535802), .Q(I535918) );
not I_31364 (I535935,I535918);
nor I_31365 (I535952,I535870,I535935);
nand I_31366 (I535788,I535918,I535887);
DFFARX1 I_31367  ( .D(I535918), .CLK(I2702), .RSTB(I535802), .Q(I535770) );
nand I_31368 (I535997,I32469,I32472);
and I_31369 (I536014,I535997,I32445);
DFFARX1 I_31370  ( .D(I536014), .CLK(I2702), .RSTB(I535802), .Q(I536031) );
nor I_31371 (I535791,I536031,I535853);
nand I_31372 (I535782,I536031,I535952);
DFFARX1 I_31373  ( .D(I32463), .CLK(I2702), .RSTB(I535802), .Q(I536076) );
and I_31374 (I536093,I536076,I32457);
DFFARX1 I_31375  ( .D(I536093), .CLK(I2702), .RSTB(I535802), .Q(I536110) );
not I_31376 (I535773,I536110);
nand I_31377 (I536141,I536093,I536031);
and I_31378 (I536158,I535853,I536141);
DFFARX1 I_31379  ( .D(I536158), .CLK(I2702), .RSTB(I535802), .Q(I535764) );
DFFARX1 I_31380  ( .D(I32460), .CLK(I2702), .RSTB(I535802), .Q(I536189) );
nand I_31381 (I536206,I536189,I535853);
and I_31382 (I536223,I536031,I536206);
DFFARX1 I_31383  ( .D(I536223), .CLK(I2702), .RSTB(I535802), .Q(I535794) );
not I_31384 (I536254,I536189);
nor I_31385 (I536271,I535870,I536254);
and I_31386 (I536288,I536189,I536271);
or I_31387 (I536305,I536093,I536288);
DFFARX1 I_31388  ( .D(I536305), .CLK(I2702), .RSTB(I535802), .Q(I535779) );
nand I_31389 (I535776,I536189,I535935);
DFFARX1 I_31390  ( .D(I536189), .CLK(I2702), .RSTB(I535802), .Q(I535767) );
not I_31391 (I536397,I2709);
nand I_31392 (I536414,I71724,I71736);
and I_31393 (I536431,I536414,I71745);
DFFARX1 I_31394  ( .D(I536431), .CLK(I2702), .RSTB(I536397), .Q(I536448) );
nor I_31395 (I536465,I71739,I71736);
nor I_31396 (I536482,I536465,I536448);
not I_31397 (I536380,I536465);
DFFARX1 I_31398  ( .D(I71733), .CLK(I2702), .RSTB(I536397), .Q(I536513) );
not I_31399 (I536530,I536513);
nor I_31400 (I536547,I536465,I536530);
nand I_31401 (I536383,I536513,I536482);
DFFARX1 I_31402  ( .D(I536513), .CLK(I2702), .RSTB(I536397), .Q(I536365) );
nand I_31403 (I536592,I71730,I71727);
and I_31404 (I536609,I536592,I71718);
DFFARX1 I_31405  ( .D(I536609), .CLK(I2702), .RSTB(I536397), .Q(I536626) );
nor I_31406 (I536386,I536626,I536448);
nand I_31407 (I536377,I536626,I536547);
DFFARX1 I_31408  ( .D(I71742), .CLK(I2702), .RSTB(I536397), .Q(I536671) );
and I_31409 (I536688,I536671,I71721);
DFFARX1 I_31410  ( .D(I536688), .CLK(I2702), .RSTB(I536397), .Q(I536705) );
not I_31411 (I536368,I536705);
nand I_31412 (I536736,I536688,I536626);
and I_31413 (I536753,I536448,I536736);
DFFARX1 I_31414  ( .D(I536753), .CLK(I2702), .RSTB(I536397), .Q(I536359) );
DFFARX1 I_31415  ( .D(I71715), .CLK(I2702), .RSTB(I536397), .Q(I536784) );
nand I_31416 (I536801,I536784,I536448);
and I_31417 (I536818,I536626,I536801);
DFFARX1 I_31418  ( .D(I536818), .CLK(I2702), .RSTB(I536397), .Q(I536389) );
not I_31419 (I536849,I536784);
nor I_31420 (I536866,I536465,I536849);
and I_31421 (I536883,I536784,I536866);
or I_31422 (I536900,I536688,I536883);
DFFARX1 I_31423  ( .D(I536900), .CLK(I2702), .RSTB(I536397), .Q(I536374) );
nand I_31424 (I536371,I536784,I536530);
DFFARX1 I_31425  ( .D(I536784), .CLK(I2702), .RSTB(I536397), .Q(I536362) );
not I_31426 (I536992,I2709);
nand I_31427 (I537009,I232612,I232615);
and I_31428 (I537026,I537009,I232606);
DFFARX1 I_31429  ( .D(I537026), .CLK(I2702), .RSTB(I536992), .Q(I537043) );
nor I_31430 (I537060,I232630,I232615);
nor I_31431 (I537077,I537060,I537043);
not I_31432 (I536975,I537060);
DFFARX1 I_31433  ( .D(I232609), .CLK(I2702), .RSTB(I536992), .Q(I537108) );
not I_31434 (I537125,I537108);
nor I_31435 (I537142,I537060,I537125);
nand I_31436 (I536978,I537108,I537077);
DFFARX1 I_31437  ( .D(I537108), .CLK(I2702), .RSTB(I536992), .Q(I536960) );
nand I_31438 (I537187,I232627,I232618);
and I_31439 (I537204,I537187,I232603);
DFFARX1 I_31440  ( .D(I537204), .CLK(I2702), .RSTB(I536992), .Q(I537221) );
nor I_31441 (I536981,I537221,I537043);
nand I_31442 (I536972,I537221,I537142);
DFFARX1 I_31443  ( .D(I232633), .CLK(I2702), .RSTB(I536992), .Q(I537266) );
and I_31444 (I537283,I537266,I232624);
DFFARX1 I_31445  ( .D(I537283), .CLK(I2702), .RSTB(I536992), .Q(I537300) );
not I_31446 (I536963,I537300);
nand I_31447 (I537331,I537283,I537221);
and I_31448 (I537348,I537043,I537331);
DFFARX1 I_31449  ( .D(I537348), .CLK(I2702), .RSTB(I536992), .Q(I536954) );
DFFARX1 I_31450  ( .D(I232621), .CLK(I2702), .RSTB(I536992), .Q(I537379) );
nand I_31451 (I537396,I537379,I537043);
and I_31452 (I537413,I537221,I537396);
DFFARX1 I_31453  ( .D(I537413), .CLK(I2702), .RSTB(I536992), .Q(I536984) );
not I_31454 (I537444,I537379);
nor I_31455 (I537461,I537060,I537444);
and I_31456 (I537478,I537379,I537461);
or I_31457 (I537495,I537283,I537478);
DFFARX1 I_31458  ( .D(I537495), .CLK(I2702), .RSTB(I536992), .Q(I536969) );
nand I_31459 (I536966,I537379,I537125);
DFFARX1 I_31460  ( .D(I537379), .CLK(I2702), .RSTB(I536992), .Q(I536957) );
not I_31461 (I537587,I2709);
nand I_31462 (I537604,I445436,I445439);
and I_31463 (I537621,I537604,I445433);
DFFARX1 I_31464  ( .D(I537621), .CLK(I2702), .RSTB(I537587), .Q(I537638) );
nor I_31465 (I537655,I445430,I445439);
nor I_31466 (I537672,I537655,I537638);
not I_31467 (I537570,I537655);
DFFARX1 I_31468  ( .D(I445412), .CLK(I2702), .RSTB(I537587), .Q(I537703) );
not I_31469 (I537720,I537703);
nor I_31470 (I537737,I537655,I537720);
nand I_31471 (I537573,I537703,I537672);
DFFARX1 I_31472  ( .D(I537703), .CLK(I2702), .RSTB(I537587), .Q(I537555) );
nand I_31473 (I537782,I445421,I445418);
and I_31474 (I537799,I537782,I445427);
DFFARX1 I_31475  ( .D(I537799), .CLK(I2702), .RSTB(I537587), .Q(I537816) );
nor I_31476 (I537576,I537816,I537638);
nand I_31477 (I537567,I537816,I537737);
DFFARX1 I_31478  ( .D(I445409), .CLK(I2702), .RSTB(I537587), .Q(I537861) );
and I_31479 (I537878,I537861,I445424);
DFFARX1 I_31480  ( .D(I537878), .CLK(I2702), .RSTB(I537587), .Q(I537895) );
not I_31481 (I537558,I537895);
nand I_31482 (I537926,I537878,I537816);
and I_31483 (I537943,I537638,I537926);
DFFARX1 I_31484  ( .D(I537943), .CLK(I2702), .RSTB(I537587), .Q(I537549) );
DFFARX1 I_31485  ( .D(I445415), .CLK(I2702), .RSTB(I537587), .Q(I537974) );
nand I_31486 (I537991,I537974,I537638);
and I_31487 (I538008,I537816,I537991);
DFFARX1 I_31488  ( .D(I538008), .CLK(I2702), .RSTB(I537587), .Q(I537579) );
not I_31489 (I538039,I537974);
nor I_31490 (I538056,I537655,I538039);
and I_31491 (I538073,I537974,I538056);
or I_31492 (I538090,I537878,I538073);
DFFARX1 I_31493  ( .D(I538090), .CLK(I2702), .RSTB(I537587), .Q(I537564) );
nand I_31494 (I537561,I537974,I537720);
DFFARX1 I_31495  ( .D(I537974), .CLK(I2702), .RSTB(I537587), .Q(I537552) );
not I_31496 (I538182,I2709);
nand I_31497 (I538199,I197907,I197919);
and I_31498 (I538216,I538199,I197898);
DFFARX1 I_31499  ( .D(I538216), .CLK(I2702), .RSTB(I538182), .Q(I538233) );
nor I_31500 (I538250,I197889,I197919);
nor I_31501 (I538267,I538250,I538233);
not I_31502 (I538165,I538250);
DFFARX1 I_31503  ( .D(I197901), .CLK(I2702), .RSTB(I538182), .Q(I538298) );
not I_31504 (I538315,I538298);
nor I_31505 (I538332,I538250,I538315);
nand I_31506 (I538168,I538298,I538267);
DFFARX1 I_31507  ( .D(I538298), .CLK(I2702), .RSTB(I538182), .Q(I538150) );
nand I_31508 (I538377,I197916,I197904);
and I_31509 (I538394,I538377,I197892);
DFFARX1 I_31510  ( .D(I538394), .CLK(I2702), .RSTB(I538182), .Q(I538411) );
nor I_31511 (I538171,I538411,I538233);
nand I_31512 (I538162,I538411,I538332);
DFFARX1 I_31513  ( .D(I197910), .CLK(I2702), .RSTB(I538182), .Q(I538456) );
and I_31514 (I538473,I538456,I197895);
DFFARX1 I_31515  ( .D(I538473), .CLK(I2702), .RSTB(I538182), .Q(I538490) );
not I_31516 (I538153,I538490);
nand I_31517 (I538521,I538473,I538411);
and I_31518 (I538538,I538233,I538521);
DFFARX1 I_31519  ( .D(I538538), .CLK(I2702), .RSTB(I538182), .Q(I538144) );
DFFARX1 I_31520  ( .D(I197913), .CLK(I2702), .RSTB(I538182), .Q(I538569) );
nand I_31521 (I538586,I538569,I538233);
and I_31522 (I538603,I538411,I538586);
DFFARX1 I_31523  ( .D(I538603), .CLK(I2702), .RSTB(I538182), .Q(I538174) );
not I_31524 (I538634,I538569);
nor I_31525 (I538651,I538250,I538634);
and I_31526 (I538668,I538569,I538651);
or I_31527 (I538685,I538473,I538668);
DFFARX1 I_31528  ( .D(I538685), .CLK(I2702), .RSTB(I538182), .Q(I538159) );
nand I_31529 (I538156,I538569,I538315);
DFFARX1 I_31530  ( .D(I538569), .CLK(I2702), .RSTB(I538182), .Q(I538147) );
not I_31531 (I538777,I2709);
nand I_31532 (I538794,I187299,I187311);
and I_31533 (I538811,I538794,I187290);
DFFARX1 I_31534  ( .D(I538811), .CLK(I2702), .RSTB(I538777), .Q(I538828) );
nor I_31535 (I538845,I187281,I187311);
nor I_31536 (I538862,I538845,I538828);
not I_31537 (I538760,I538845);
DFFARX1 I_31538  ( .D(I187293), .CLK(I2702), .RSTB(I538777), .Q(I538893) );
not I_31539 (I538910,I538893);
nor I_31540 (I538927,I538845,I538910);
nand I_31541 (I538763,I538893,I538862);
DFFARX1 I_31542  ( .D(I538893), .CLK(I2702), .RSTB(I538777), .Q(I538745) );
nand I_31543 (I538972,I187308,I187296);
and I_31544 (I538989,I538972,I187284);
DFFARX1 I_31545  ( .D(I538989), .CLK(I2702), .RSTB(I538777), .Q(I539006) );
nor I_31546 (I538766,I539006,I538828);
nand I_31547 (I538757,I539006,I538927);
DFFARX1 I_31548  ( .D(I187302), .CLK(I2702), .RSTB(I538777), .Q(I539051) );
and I_31549 (I539068,I539051,I187287);
DFFARX1 I_31550  ( .D(I539068), .CLK(I2702), .RSTB(I538777), .Q(I539085) );
not I_31551 (I538748,I539085);
nand I_31552 (I539116,I539068,I539006);
and I_31553 (I539133,I538828,I539116);
DFFARX1 I_31554  ( .D(I539133), .CLK(I2702), .RSTB(I538777), .Q(I538739) );
DFFARX1 I_31555  ( .D(I187305), .CLK(I2702), .RSTB(I538777), .Q(I539164) );
nand I_31556 (I539181,I539164,I538828);
and I_31557 (I539198,I539006,I539181);
DFFARX1 I_31558  ( .D(I539198), .CLK(I2702), .RSTB(I538777), .Q(I538769) );
not I_31559 (I539229,I539164);
nor I_31560 (I539246,I538845,I539229);
and I_31561 (I539263,I539164,I539246);
or I_31562 (I539280,I539068,I539263);
DFFARX1 I_31563  ( .D(I539280), .CLK(I2702), .RSTB(I538777), .Q(I538754) );
nand I_31564 (I538751,I539164,I538910);
DFFARX1 I_31565  ( .D(I539164), .CLK(I2702), .RSTB(I538777), .Q(I538742) );
not I_31566 (I539372,I2709);
nand I_31567 (I539389,I686028,I686019);
and I_31568 (I539406,I539389,I686037);
DFFARX1 I_31569  ( .D(I539406), .CLK(I2702), .RSTB(I539372), .Q(I539423) );
nor I_31570 (I539440,I686034,I686019);
nor I_31571 (I539457,I539440,I539423);
not I_31572 (I539355,I539440);
DFFARX1 I_31573  ( .D(I686016), .CLK(I2702), .RSTB(I539372), .Q(I539488) );
not I_31574 (I539505,I539488);
nor I_31575 (I539522,I539440,I539505);
nand I_31576 (I539358,I539488,I539457);
DFFARX1 I_31577  ( .D(I539488), .CLK(I2702), .RSTB(I539372), .Q(I539340) );
nand I_31578 (I539567,I686025,I686040);
and I_31579 (I539584,I539567,I686031);
DFFARX1 I_31580  ( .D(I539584), .CLK(I2702), .RSTB(I539372), .Q(I539601) );
nor I_31581 (I539361,I539601,I539423);
nand I_31582 (I539352,I539601,I539522);
DFFARX1 I_31583  ( .D(I686013), .CLK(I2702), .RSTB(I539372), .Q(I539646) );
and I_31584 (I539663,I539646,I686022);
DFFARX1 I_31585  ( .D(I539663), .CLK(I2702), .RSTB(I539372), .Q(I539680) );
not I_31586 (I539343,I539680);
nand I_31587 (I539711,I539663,I539601);
and I_31588 (I539728,I539423,I539711);
DFFARX1 I_31589  ( .D(I539728), .CLK(I2702), .RSTB(I539372), .Q(I539334) );
DFFARX1 I_31590  ( .D(I686010), .CLK(I2702), .RSTB(I539372), .Q(I539759) );
nand I_31591 (I539776,I539759,I539423);
and I_31592 (I539793,I539601,I539776);
DFFARX1 I_31593  ( .D(I539793), .CLK(I2702), .RSTB(I539372), .Q(I539364) );
not I_31594 (I539824,I539759);
nor I_31595 (I539841,I539440,I539824);
and I_31596 (I539858,I539759,I539841);
or I_31597 (I539875,I539663,I539858);
DFFARX1 I_31598  ( .D(I539875), .CLK(I2702), .RSTB(I539372), .Q(I539349) );
nand I_31599 (I539346,I539759,I539505);
DFFARX1 I_31600  ( .D(I539759), .CLK(I2702), .RSTB(I539372), .Q(I539337) );
not I_31601 (I539967,I2709);
nand I_31602 (I539984,I275478,I275484);
and I_31603 (I540001,I539984,I275466);
DFFARX1 I_31604  ( .D(I540001), .CLK(I2702), .RSTB(I539967), .Q(I540018) );
nor I_31605 (I540035,I275460,I275484);
nor I_31606 (I540052,I540035,I540018);
not I_31607 (I539950,I540035);
DFFARX1 I_31608  ( .D(I275490), .CLK(I2702), .RSTB(I539967), .Q(I540083) );
not I_31609 (I540100,I540083);
nor I_31610 (I540117,I540035,I540100);
nand I_31611 (I539953,I540083,I540052);
DFFARX1 I_31612  ( .D(I540083), .CLK(I2702), .RSTB(I539967), .Q(I539935) );
nand I_31613 (I540162,I275481,I275472);
and I_31614 (I540179,I540162,I275475);
DFFARX1 I_31615  ( .D(I540179), .CLK(I2702), .RSTB(I539967), .Q(I540196) );
nor I_31616 (I539956,I540196,I540018);
nand I_31617 (I539947,I540196,I540117);
DFFARX1 I_31618  ( .D(I275487), .CLK(I2702), .RSTB(I539967), .Q(I540241) );
and I_31619 (I540258,I540241,I275463);
DFFARX1 I_31620  ( .D(I540258), .CLK(I2702), .RSTB(I539967), .Q(I540275) );
not I_31621 (I539938,I540275);
nand I_31622 (I540306,I540258,I540196);
and I_31623 (I540323,I540018,I540306);
DFFARX1 I_31624  ( .D(I540323), .CLK(I2702), .RSTB(I539967), .Q(I539929) );
DFFARX1 I_31625  ( .D(I275469), .CLK(I2702), .RSTB(I539967), .Q(I540354) );
nand I_31626 (I540371,I540354,I540018);
and I_31627 (I540388,I540196,I540371);
DFFARX1 I_31628  ( .D(I540388), .CLK(I2702), .RSTB(I539967), .Q(I539959) );
not I_31629 (I540419,I540354);
nor I_31630 (I540436,I540035,I540419);
and I_31631 (I540453,I540354,I540436);
or I_31632 (I540470,I540258,I540453);
DFFARX1 I_31633  ( .D(I540470), .CLK(I2702), .RSTB(I539967), .Q(I539944) );
nand I_31634 (I539941,I540354,I540100);
DFFARX1 I_31635  ( .D(I540354), .CLK(I2702), .RSTB(I539967), .Q(I539932) );
not I_31636 (I540562,I2709);
nand I_31637 (I540579,I430955,I430943);
and I_31638 (I540596,I540579,I430949);
DFFARX1 I_31639  ( .D(I540596), .CLK(I2702), .RSTB(I540562), .Q(I540613) );
nor I_31640 (I540630,I430940,I430943);
nor I_31641 (I540647,I540630,I540613);
not I_31642 (I540545,I540630);
DFFARX1 I_31643  ( .D(I430925), .CLK(I2702), .RSTB(I540562), .Q(I540678) );
not I_31644 (I540695,I540678);
nor I_31645 (I540712,I540630,I540695);
nand I_31646 (I540548,I540678,I540647);
DFFARX1 I_31647  ( .D(I540678), .CLK(I2702), .RSTB(I540562), .Q(I540530) );
nand I_31648 (I540757,I430934,I430952);
and I_31649 (I540774,I540757,I430946);
DFFARX1 I_31650  ( .D(I540774), .CLK(I2702), .RSTB(I540562), .Q(I540791) );
nor I_31651 (I540551,I540791,I540613);
nand I_31652 (I540542,I540791,I540712);
DFFARX1 I_31653  ( .D(I430937), .CLK(I2702), .RSTB(I540562), .Q(I540836) );
and I_31654 (I540853,I540836,I430931);
DFFARX1 I_31655  ( .D(I540853), .CLK(I2702), .RSTB(I540562), .Q(I540870) );
not I_31656 (I540533,I540870);
nand I_31657 (I540901,I540853,I540791);
and I_31658 (I540918,I540613,I540901);
DFFARX1 I_31659  ( .D(I540918), .CLK(I2702), .RSTB(I540562), .Q(I540524) );
DFFARX1 I_31660  ( .D(I430928), .CLK(I2702), .RSTB(I540562), .Q(I540949) );
nand I_31661 (I540966,I540949,I540613);
and I_31662 (I540983,I540791,I540966);
DFFARX1 I_31663  ( .D(I540983), .CLK(I2702), .RSTB(I540562), .Q(I540554) );
not I_31664 (I541014,I540949);
nor I_31665 (I541031,I540630,I541014);
and I_31666 (I541048,I540949,I541031);
or I_31667 (I541065,I540853,I541048);
DFFARX1 I_31668  ( .D(I541065), .CLK(I2702), .RSTB(I540562), .Q(I540539) );
nand I_31669 (I540536,I540949,I540695);
DFFARX1 I_31670  ( .D(I540949), .CLK(I2702), .RSTB(I540562), .Q(I540527) );
not I_31671 (I541157,I2709);
nand I_31672 (I541174,I672819,I672810);
and I_31673 (I541191,I541174,I672828);
DFFARX1 I_31674  ( .D(I541191), .CLK(I2702), .RSTB(I541157), .Q(I541208) );
nor I_31675 (I541225,I672825,I672810);
nor I_31676 (I541242,I541225,I541208);
not I_31677 (I541140,I541225);
DFFARX1 I_31678  ( .D(I672807), .CLK(I2702), .RSTB(I541157), .Q(I541273) );
not I_31679 (I541290,I541273);
nor I_31680 (I541307,I541225,I541290);
nand I_31681 (I541143,I541273,I541242);
DFFARX1 I_31682  ( .D(I541273), .CLK(I2702), .RSTB(I541157), .Q(I541125) );
nand I_31683 (I541352,I672816,I672831);
and I_31684 (I541369,I541352,I672822);
DFFARX1 I_31685  ( .D(I541369), .CLK(I2702), .RSTB(I541157), .Q(I541386) );
nor I_31686 (I541146,I541386,I541208);
nand I_31687 (I541137,I541386,I541307);
DFFARX1 I_31688  ( .D(I672804), .CLK(I2702), .RSTB(I541157), .Q(I541431) );
and I_31689 (I541448,I541431,I672813);
DFFARX1 I_31690  ( .D(I541448), .CLK(I2702), .RSTB(I541157), .Q(I541465) );
not I_31691 (I541128,I541465);
nand I_31692 (I541496,I541448,I541386);
and I_31693 (I541513,I541208,I541496);
DFFARX1 I_31694  ( .D(I541513), .CLK(I2702), .RSTB(I541157), .Q(I541119) );
DFFARX1 I_31695  ( .D(I672801), .CLK(I2702), .RSTB(I541157), .Q(I541544) );
nand I_31696 (I541561,I541544,I541208);
and I_31697 (I541578,I541386,I541561);
DFFARX1 I_31698  ( .D(I541578), .CLK(I2702), .RSTB(I541157), .Q(I541149) );
not I_31699 (I541609,I541544);
nor I_31700 (I541626,I541225,I541609);
and I_31701 (I541643,I541544,I541626);
or I_31702 (I541660,I541448,I541643);
DFFARX1 I_31703  ( .D(I541660), .CLK(I2702), .RSTB(I541157), .Q(I541134) );
nand I_31704 (I541131,I541544,I541290);
DFFARX1 I_31705  ( .D(I541544), .CLK(I2702), .RSTB(I541157), .Q(I541122) );
not I_31706 (I541752,I2709);
nand I_31707 (I541769,I97564,I97576);
and I_31708 (I541786,I541769,I97585);
DFFARX1 I_31709  ( .D(I541786), .CLK(I2702), .RSTB(I541752), .Q(I541803) );
nor I_31710 (I541820,I97579,I97576);
nor I_31711 (I541837,I541820,I541803);
not I_31712 (I541735,I541820);
DFFARX1 I_31713  ( .D(I97573), .CLK(I2702), .RSTB(I541752), .Q(I541868) );
not I_31714 (I541885,I541868);
nor I_31715 (I541902,I541820,I541885);
nand I_31716 (I541738,I541868,I541837);
DFFARX1 I_31717  ( .D(I541868), .CLK(I2702), .RSTB(I541752), .Q(I541720) );
nand I_31718 (I541947,I97570,I97567);
and I_31719 (I541964,I541947,I97558);
DFFARX1 I_31720  ( .D(I541964), .CLK(I2702), .RSTB(I541752), .Q(I541981) );
nor I_31721 (I541741,I541981,I541803);
nand I_31722 (I541732,I541981,I541902);
DFFARX1 I_31723  ( .D(I97582), .CLK(I2702), .RSTB(I541752), .Q(I542026) );
and I_31724 (I542043,I542026,I97561);
DFFARX1 I_31725  ( .D(I542043), .CLK(I2702), .RSTB(I541752), .Q(I542060) );
not I_31726 (I541723,I542060);
nand I_31727 (I542091,I542043,I541981);
and I_31728 (I542108,I541803,I542091);
DFFARX1 I_31729  ( .D(I542108), .CLK(I2702), .RSTB(I541752), .Q(I541714) );
DFFARX1 I_31730  ( .D(I97555), .CLK(I2702), .RSTB(I541752), .Q(I542139) );
nand I_31731 (I542156,I542139,I541803);
and I_31732 (I542173,I541981,I542156);
DFFARX1 I_31733  ( .D(I542173), .CLK(I2702), .RSTB(I541752), .Q(I541744) );
not I_31734 (I542204,I542139);
nor I_31735 (I542221,I541820,I542204);
and I_31736 (I542238,I542139,I542221);
or I_31737 (I542255,I542043,I542238);
DFFARX1 I_31738  ( .D(I542255), .CLK(I2702), .RSTB(I541752), .Q(I541729) );
nand I_31739 (I541726,I542139,I541885);
DFFARX1 I_31740  ( .D(I542139), .CLK(I2702), .RSTB(I541752), .Q(I541717) );
not I_31741 (I542347,I2709);
nand I_31742 (I542364,I240942,I240945);
and I_31743 (I542381,I542364,I240936);
DFFARX1 I_31744  ( .D(I542381), .CLK(I2702), .RSTB(I542347), .Q(I542398) );
nor I_31745 (I542415,I240960,I240945);
nor I_31746 (I542432,I542415,I542398);
not I_31747 (I542330,I542415);
DFFARX1 I_31748  ( .D(I240939), .CLK(I2702), .RSTB(I542347), .Q(I542463) );
not I_31749 (I542480,I542463);
nor I_31750 (I542497,I542415,I542480);
nand I_31751 (I542333,I542463,I542432);
DFFARX1 I_31752  ( .D(I542463), .CLK(I2702), .RSTB(I542347), .Q(I542315) );
nand I_31753 (I542542,I240957,I240948);
and I_31754 (I542559,I542542,I240933);
DFFARX1 I_31755  ( .D(I542559), .CLK(I2702), .RSTB(I542347), .Q(I542576) );
nor I_31756 (I542336,I542576,I542398);
nand I_31757 (I542327,I542576,I542497);
DFFARX1 I_31758  ( .D(I240963), .CLK(I2702), .RSTB(I542347), .Q(I542621) );
and I_31759 (I542638,I542621,I240954);
DFFARX1 I_31760  ( .D(I542638), .CLK(I2702), .RSTB(I542347), .Q(I542655) );
not I_31761 (I542318,I542655);
nand I_31762 (I542686,I542638,I542576);
and I_31763 (I542703,I542398,I542686);
DFFARX1 I_31764  ( .D(I542703), .CLK(I2702), .RSTB(I542347), .Q(I542309) );
DFFARX1 I_31765  ( .D(I240951), .CLK(I2702), .RSTB(I542347), .Q(I542734) );
nand I_31766 (I542751,I542734,I542398);
and I_31767 (I542768,I542576,I542751);
DFFARX1 I_31768  ( .D(I542768), .CLK(I2702), .RSTB(I542347), .Q(I542339) );
not I_31769 (I542799,I542734);
nor I_31770 (I542816,I542415,I542799);
and I_31771 (I542833,I542734,I542816);
or I_31772 (I542850,I542638,I542833);
DFFARX1 I_31773  ( .D(I542850), .CLK(I2702), .RSTB(I542347), .Q(I542324) );
nand I_31774 (I542321,I542734,I542480);
DFFARX1 I_31775  ( .D(I542734), .CLK(I2702), .RSTB(I542347), .Q(I542312) );
not I_31776 (I542942,I2709);
nand I_31777 (I542959,I80122,I80134);
and I_31778 (I542976,I542959,I80143);
DFFARX1 I_31779  ( .D(I542976), .CLK(I2702), .RSTB(I542942), .Q(I542993) );
nor I_31780 (I543010,I80137,I80134);
nor I_31781 (I543027,I543010,I542993);
not I_31782 (I542925,I543010);
DFFARX1 I_31783  ( .D(I80131), .CLK(I2702), .RSTB(I542942), .Q(I543058) );
not I_31784 (I543075,I543058);
nor I_31785 (I543092,I543010,I543075);
nand I_31786 (I542928,I543058,I543027);
DFFARX1 I_31787  ( .D(I543058), .CLK(I2702), .RSTB(I542942), .Q(I542910) );
nand I_31788 (I543137,I80128,I80125);
and I_31789 (I543154,I543137,I80116);
DFFARX1 I_31790  ( .D(I543154), .CLK(I2702), .RSTB(I542942), .Q(I543171) );
nor I_31791 (I542931,I543171,I542993);
nand I_31792 (I542922,I543171,I543092);
DFFARX1 I_31793  ( .D(I80140), .CLK(I2702), .RSTB(I542942), .Q(I543216) );
and I_31794 (I543233,I543216,I80119);
DFFARX1 I_31795  ( .D(I543233), .CLK(I2702), .RSTB(I542942), .Q(I543250) );
not I_31796 (I542913,I543250);
nand I_31797 (I543281,I543233,I543171);
and I_31798 (I543298,I542993,I543281);
DFFARX1 I_31799  ( .D(I543298), .CLK(I2702), .RSTB(I542942), .Q(I542904) );
DFFARX1 I_31800  ( .D(I80113), .CLK(I2702), .RSTB(I542942), .Q(I543329) );
nand I_31801 (I543346,I543329,I542993);
and I_31802 (I543363,I543171,I543346);
DFFARX1 I_31803  ( .D(I543363), .CLK(I2702), .RSTB(I542942), .Q(I542934) );
not I_31804 (I543394,I543329);
nor I_31805 (I543411,I543010,I543394);
and I_31806 (I543428,I543329,I543411);
or I_31807 (I543445,I543233,I543428);
DFFARX1 I_31808  ( .D(I543445), .CLK(I2702), .RSTB(I542942), .Q(I542919) );
nand I_31809 (I542916,I543329,I543075);
DFFARX1 I_31810  ( .D(I543329), .CLK(I2702), .RSTB(I542942), .Q(I542907) );
not I_31811 (I543537,I2709);
nand I_31812 (I543554,I446014,I446017);
and I_31813 (I543571,I543554,I446011);
DFFARX1 I_31814  ( .D(I543571), .CLK(I2702), .RSTB(I543537), .Q(I543588) );
nor I_31815 (I543605,I446008,I446017);
nor I_31816 (I543622,I543605,I543588);
not I_31817 (I543520,I543605);
DFFARX1 I_31818  ( .D(I445990), .CLK(I2702), .RSTB(I543537), .Q(I543653) );
not I_31819 (I543670,I543653);
nor I_31820 (I543687,I543605,I543670);
nand I_31821 (I543523,I543653,I543622);
DFFARX1 I_31822  ( .D(I543653), .CLK(I2702), .RSTB(I543537), .Q(I543505) );
nand I_31823 (I543732,I445999,I445996);
and I_31824 (I543749,I543732,I446005);
DFFARX1 I_31825  ( .D(I543749), .CLK(I2702), .RSTB(I543537), .Q(I543766) );
nor I_31826 (I543526,I543766,I543588);
nand I_31827 (I543517,I543766,I543687);
DFFARX1 I_31828  ( .D(I445987), .CLK(I2702), .RSTB(I543537), .Q(I543811) );
and I_31829 (I543828,I543811,I446002);
DFFARX1 I_31830  ( .D(I543828), .CLK(I2702), .RSTB(I543537), .Q(I543845) );
not I_31831 (I543508,I543845);
nand I_31832 (I543876,I543828,I543766);
and I_31833 (I543893,I543588,I543876);
DFFARX1 I_31834  ( .D(I543893), .CLK(I2702), .RSTB(I543537), .Q(I543499) );
DFFARX1 I_31835  ( .D(I445993), .CLK(I2702), .RSTB(I543537), .Q(I543924) );
nand I_31836 (I543941,I543924,I543588);
and I_31837 (I543958,I543766,I543941);
DFFARX1 I_31838  ( .D(I543958), .CLK(I2702), .RSTB(I543537), .Q(I543529) );
not I_31839 (I543989,I543924);
nor I_31840 (I544006,I543605,I543989);
and I_31841 (I544023,I543924,I544006);
or I_31842 (I544040,I543828,I544023);
DFFARX1 I_31843  ( .D(I544040), .CLK(I2702), .RSTB(I543537), .Q(I543514) );
nand I_31844 (I543511,I543924,I543670);
DFFARX1 I_31845  ( .D(I543924), .CLK(I2702), .RSTB(I543537), .Q(I543502) );
not I_31846 (I544132,I2709);
nand I_31847 (I544149,I129864,I129876);
and I_31848 (I544166,I544149,I129885);
DFFARX1 I_31849  ( .D(I544166), .CLK(I2702), .RSTB(I544132), .Q(I544183) );
nor I_31850 (I544200,I129879,I129876);
nor I_31851 (I544217,I544200,I544183);
not I_31852 (I544115,I544200);
DFFARX1 I_31853  ( .D(I129873), .CLK(I2702), .RSTB(I544132), .Q(I544248) );
not I_31854 (I544265,I544248);
nor I_31855 (I544282,I544200,I544265);
nand I_31856 (I544118,I544248,I544217);
DFFARX1 I_31857  ( .D(I544248), .CLK(I2702), .RSTB(I544132), .Q(I544100) );
nand I_31858 (I544327,I129870,I129867);
and I_31859 (I544344,I544327,I129858);
DFFARX1 I_31860  ( .D(I544344), .CLK(I2702), .RSTB(I544132), .Q(I544361) );
nor I_31861 (I544121,I544361,I544183);
nand I_31862 (I544112,I544361,I544282);
DFFARX1 I_31863  ( .D(I129882), .CLK(I2702), .RSTB(I544132), .Q(I544406) );
and I_31864 (I544423,I544406,I129861);
DFFARX1 I_31865  ( .D(I544423), .CLK(I2702), .RSTB(I544132), .Q(I544440) );
not I_31866 (I544103,I544440);
nand I_31867 (I544471,I544423,I544361);
and I_31868 (I544488,I544183,I544471);
DFFARX1 I_31869  ( .D(I544488), .CLK(I2702), .RSTB(I544132), .Q(I544094) );
DFFARX1 I_31870  ( .D(I129855), .CLK(I2702), .RSTB(I544132), .Q(I544519) );
nand I_31871 (I544536,I544519,I544183);
and I_31872 (I544553,I544361,I544536);
DFFARX1 I_31873  ( .D(I544553), .CLK(I2702), .RSTB(I544132), .Q(I544124) );
not I_31874 (I544584,I544519);
nor I_31875 (I544601,I544200,I544584);
and I_31876 (I544618,I544519,I544601);
or I_31877 (I544635,I544423,I544618);
DFFARX1 I_31878  ( .D(I544635), .CLK(I2702), .RSTB(I544132), .Q(I544109) );
nand I_31879 (I544106,I544519,I544265);
DFFARX1 I_31880  ( .D(I544519), .CLK(I2702), .RSTB(I544132), .Q(I544097) );
not I_31881 (I544727,I2709);
nand I_31882 (I544744,I389361,I389373);
and I_31883 (I544761,I544744,I389355);
DFFARX1 I_31884  ( .D(I544761), .CLK(I2702), .RSTB(I544727), .Q(I544778) );
nor I_31885 (I544795,I389367,I389373);
nor I_31886 (I544812,I544795,I544778);
not I_31887 (I544710,I544795);
DFFARX1 I_31888  ( .D(I389352), .CLK(I2702), .RSTB(I544727), .Q(I544843) );
not I_31889 (I544860,I544843);
nor I_31890 (I544877,I544795,I544860);
nand I_31891 (I544713,I544843,I544812);
DFFARX1 I_31892  ( .D(I544843), .CLK(I2702), .RSTB(I544727), .Q(I544695) );
nand I_31893 (I544922,I389343,I389358);
and I_31894 (I544939,I544922,I389349);
DFFARX1 I_31895  ( .D(I544939), .CLK(I2702), .RSTB(I544727), .Q(I544956) );
nor I_31896 (I544716,I544956,I544778);
nand I_31897 (I544707,I544956,I544877);
DFFARX1 I_31898  ( .D(I389370), .CLK(I2702), .RSTB(I544727), .Q(I545001) );
and I_31899 (I545018,I545001,I389364);
DFFARX1 I_31900  ( .D(I545018), .CLK(I2702), .RSTB(I544727), .Q(I545035) );
not I_31901 (I544698,I545035);
nand I_31902 (I545066,I545018,I544956);
and I_31903 (I545083,I544778,I545066);
DFFARX1 I_31904  ( .D(I545083), .CLK(I2702), .RSTB(I544727), .Q(I544689) );
DFFARX1 I_31905  ( .D(I389346), .CLK(I2702), .RSTB(I544727), .Q(I545114) );
nand I_31906 (I545131,I545114,I544778);
and I_31907 (I545148,I544956,I545131);
DFFARX1 I_31908  ( .D(I545148), .CLK(I2702), .RSTB(I544727), .Q(I544719) );
not I_31909 (I545179,I545114);
nor I_31910 (I545196,I544795,I545179);
and I_31911 (I545213,I545114,I545196);
or I_31912 (I545230,I545018,I545213);
DFFARX1 I_31913  ( .D(I545230), .CLK(I2702), .RSTB(I544727), .Q(I544704) );
nand I_31914 (I544701,I545114,I544860);
DFFARX1 I_31915  ( .D(I545114), .CLK(I2702), .RSTB(I544727), .Q(I544692) );
not I_31916 (I545322,I2709);
nand I_31917 (I545339,I180669,I180681);
and I_31918 (I545356,I545339,I180660);
DFFARX1 I_31919  ( .D(I545356), .CLK(I2702), .RSTB(I545322), .Q(I545373) );
nor I_31920 (I545390,I180651,I180681);
nor I_31921 (I545407,I545390,I545373);
not I_31922 (I545305,I545390);
DFFARX1 I_31923  ( .D(I180663), .CLK(I2702), .RSTB(I545322), .Q(I545438) );
not I_31924 (I545455,I545438);
nor I_31925 (I545472,I545390,I545455);
nand I_31926 (I545308,I545438,I545407);
DFFARX1 I_31927  ( .D(I545438), .CLK(I2702), .RSTB(I545322), .Q(I545290) );
nand I_31928 (I545517,I180678,I180666);
and I_31929 (I545534,I545517,I180654);
DFFARX1 I_31930  ( .D(I545534), .CLK(I2702), .RSTB(I545322), .Q(I545551) );
nor I_31931 (I545311,I545551,I545373);
nand I_31932 (I545302,I545551,I545472);
DFFARX1 I_31933  ( .D(I180672), .CLK(I2702), .RSTB(I545322), .Q(I545596) );
and I_31934 (I545613,I545596,I180657);
DFFARX1 I_31935  ( .D(I545613), .CLK(I2702), .RSTB(I545322), .Q(I545630) );
not I_31936 (I545293,I545630);
nand I_31937 (I545661,I545613,I545551);
and I_31938 (I545678,I545373,I545661);
DFFARX1 I_31939  ( .D(I545678), .CLK(I2702), .RSTB(I545322), .Q(I545284) );
DFFARX1 I_31940  ( .D(I180675), .CLK(I2702), .RSTB(I545322), .Q(I545709) );
nand I_31941 (I545726,I545709,I545373);
and I_31942 (I545743,I545551,I545726);
DFFARX1 I_31943  ( .D(I545743), .CLK(I2702), .RSTB(I545322), .Q(I545314) );
not I_31944 (I545774,I545709);
nor I_31945 (I545791,I545390,I545774);
and I_31946 (I545808,I545709,I545791);
or I_31947 (I545825,I545613,I545808);
DFFARX1 I_31948  ( .D(I545825), .CLK(I2702), .RSTB(I545322), .Q(I545299) );
nand I_31949 (I545296,I545709,I545455);
DFFARX1 I_31950  ( .D(I545709), .CLK(I2702), .RSTB(I545322), .Q(I545287) );
not I_31951 (I545917,I2709);
nand I_31952 (I545934,I369981,I369993);
and I_31953 (I545951,I545934,I369975);
DFFARX1 I_31954  ( .D(I545951), .CLK(I2702), .RSTB(I545917), .Q(I545968) );
nor I_31955 (I545985,I369987,I369993);
nor I_31956 (I546002,I545985,I545968);
not I_31957 (I545900,I545985);
DFFARX1 I_31958  ( .D(I369972), .CLK(I2702), .RSTB(I545917), .Q(I546033) );
not I_31959 (I546050,I546033);
nor I_31960 (I546067,I545985,I546050);
nand I_31961 (I545903,I546033,I546002);
DFFARX1 I_31962  ( .D(I546033), .CLK(I2702), .RSTB(I545917), .Q(I545885) );
nand I_31963 (I546112,I369963,I369978);
and I_31964 (I546129,I546112,I369969);
DFFARX1 I_31965  ( .D(I546129), .CLK(I2702), .RSTB(I545917), .Q(I546146) );
nor I_31966 (I545906,I546146,I545968);
nand I_31967 (I545897,I546146,I546067);
DFFARX1 I_31968  ( .D(I369990), .CLK(I2702), .RSTB(I545917), .Q(I546191) );
and I_31969 (I546208,I546191,I369984);
DFFARX1 I_31970  ( .D(I546208), .CLK(I2702), .RSTB(I545917), .Q(I546225) );
not I_31971 (I545888,I546225);
nand I_31972 (I546256,I546208,I546146);
and I_31973 (I546273,I545968,I546256);
DFFARX1 I_31974  ( .D(I546273), .CLK(I2702), .RSTB(I545917), .Q(I545879) );
DFFARX1 I_31975  ( .D(I369966), .CLK(I2702), .RSTB(I545917), .Q(I546304) );
nand I_31976 (I546321,I546304,I545968);
and I_31977 (I546338,I546146,I546321);
DFFARX1 I_31978  ( .D(I546338), .CLK(I2702), .RSTB(I545917), .Q(I545909) );
not I_31979 (I546369,I546304);
nor I_31980 (I546386,I545985,I546369);
and I_31981 (I546403,I546304,I546386);
or I_31982 (I546420,I546208,I546403);
DFFARX1 I_31983  ( .D(I546420), .CLK(I2702), .RSTB(I545917), .Q(I545894) );
nand I_31984 (I545891,I546304,I546050);
DFFARX1 I_31985  ( .D(I546304), .CLK(I2702), .RSTB(I545917), .Q(I545882) );
not I_31986 (I546512,I2709);
nand I_31987 (I546529,I296031,I296037);
and I_31988 (I546546,I546529,I296019);
DFFARX1 I_31989  ( .D(I546546), .CLK(I2702), .RSTB(I546512), .Q(I546563) );
nor I_31990 (I546580,I296013,I296037);
nor I_31991 (I546597,I546580,I546563);
not I_31992 (I546495,I546580);
DFFARX1 I_31993  ( .D(I296043), .CLK(I2702), .RSTB(I546512), .Q(I546628) );
not I_31994 (I546645,I546628);
nor I_31995 (I546662,I546580,I546645);
nand I_31996 (I546498,I546628,I546597);
DFFARX1 I_31997  ( .D(I546628), .CLK(I2702), .RSTB(I546512), .Q(I546480) );
nand I_31998 (I546707,I296034,I296025);
and I_31999 (I546724,I546707,I296028);
DFFARX1 I_32000  ( .D(I546724), .CLK(I2702), .RSTB(I546512), .Q(I546741) );
nor I_32001 (I546501,I546741,I546563);
nand I_32002 (I546492,I546741,I546662);
DFFARX1 I_32003  ( .D(I296040), .CLK(I2702), .RSTB(I546512), .Q(I546786) );
and I_32004 (I546803,I546786,I296016);
DFFARX1 I_32005  ( .D(I546803), .CLK(I2702), .RSTB(I546512), .Q(I546820) );
not I_32006 (I546483,I546820);
nand I_32007 (I546851,I546803,I546741);
and I_32008 (I546868,I546563,I546851);
DFFARX1 I_32009  ( .D(I546868), .CLK(I2702), .RSTB(I546512), .Q(I546474) );
DFFARX1 I_32010  ( .D(I296022), .CLK(I2702), .RSTB(I546512), .Q(I546899) );
nand I_32011 (I546916,I546899,I546563);
and I_32012 (I546933,I546741,I546916);
DFFARX1 I_32013  ( .D(I546933), .CLK(I2702), .RSTB(I546512), .Q(I546504) );
not I_32014 (I546964,I546899);
nor I_32015 (I546981,I546580,I546964);
and I_32016 (I546998,I546899,I546981);
or I_32017 (I547015,I546803,I546998);
DFFARX1 I_32018  ( .D(I547015), .CLK(I2702), .RSTB(I546512), .Q(I546489) );
nand I_32019 (I546486,I546899,I546645);
DFFARX1 I_32020  ( .D(I546899), .CLK(I2702), .RSTB(I546512), .Q(I546477) );
not I_32021 (I547107,I2709);
nand I_32022 (I547124,I223098,I223095);
and I_32023 (I547141,I547124,I223092);
DFFARX1 I_32024  ( .D(I547141), .CLK(I2702), .RSTB(I547107), .Q(I547158) );
nor I_32025 (I547175,I223083,I223095);
nor I_32026 (I547192,I547175,I547158);
not I_32027 (I547090,I547175);
DFFARX1 I_32028  ( .D(I223101), .CLK(I2702), .RSTB(I547107), .Q(I547223) );
not I_32029 (I547240,I547223);
nor I_32030 (I547257,I547175,I547240);
nand I_32031 (I547093,I547223,I547192);
DFFARX1 I_32032  ( .D(I547223), .CLK(I2702), .RSTB(I547107), .Q(I547075) );
nand I_32033 (I547302,I223086,I223110);
and I_32034 (I547319,I547302,I223089);
DFFARX1 I_32035  ( .D(I547319), .CLK(I2702), .RSTB(I547107), .Q(I547336) );
nor I_32036 (I547096,I547336,I547158);
nand I_32037 (I547087,I547336,I547257);
DFFARX1 I_32038  ( .D(I223107), .CLK(I2702), .RSTB(I547107), .Q(I547381) );
and I_32039 (I547398,I547381,I223104);
DFFARX1 I_32040  ( .D(I547398), .CLK(I2702), .RSTB(I547107), .Q(I547415) );
not I_32041 (I547078,I547415);
nand I_32042 (I547446,I547398,I547336);
and I_32043 (I547463,I547158,I547446);
DFFARX1 I_32044  ( .D(I547463), .CLK(I2702), .RSTB(I547107), .Q(I547069) );
DFFARX1 I_32045  ( .D(I223113), .CLK(I2702), .RSTB(I547107), .Q(I547494) );
nand I_32046 (I547511,I547494,I547158);
and I_32047 (I547528,I547336,I547511);
DFFARX1 I_32048  ( .D(I547528), .CLK(I2702), .RSTB(I547107), .Q(I547099) );
not I_32049 (I547559,I547494);
nor I_32050 (I547576,I547175,I547559);
and I_32051 (I547593,I547494,I547576);
or I_32052 (I547610,I547398,I547593);
DFFARX1 I_32053  ( .D(I547610), .CLK(I2702), .RSTB(I547107), .Q(I547084) );
nand I_32054 (I547081,I547494,I547240);
DFFARX1 I_32055  ( .D(I547494), .CLK(I2702), .RSTB(I547107), .Q(I547072) );
not I_32056 (I547702,I2709);
nand I_32057 (I547719,I615580,I615571);
and I_32058 (I547736,I547719,I615589);
DFFARX1 I_32059  ( .D(I547736), .CLK(I2702), .RSTB(I547702), .Q(I547753) );
nor I_32060 (I547770,I615586,I615571);
nor I_32061 (I547787,I547770,I547753);
not I_32062 (I547685,I547770);
DFFARX1 I_32063  ( .D(I615568), .CLK(I2702), .RSTB(I547702), .Q(I547818) );
not I_32064 (I547835,I547818);
nor I_32065 (I547852,I547770,I547835);
nand I_32066 (I547688,I547818,I547787);
DFFARX1 I_32067  ( .D(I547818), .CLK(I2702), .RSTB(I547702), .Q(I547670) );
nand I_32068 (I547897,I615577,I615592);
and I_32069 (I547914,I547897,I615583);
DFFARX1 I_32070  ( .D(I547914), .CLK(I2702), .RSTB(I547702), .Q(I547931) );
nor I_32071 (I547691,I547931,I547753);
nand I_32072 (I547682,I547931,I547852);
DFFARX1 I_32073  ( .D(I615565), .CLK(I2702), .RSTB(I547702), .Q(I547976) );
and I_32074 (I547993,I547976,I615574);
DFFARX1 I_32075  ( .D(I547993), .CLK(I2702), .RSTB(I547702), .Q(I548010) );
not I_32076 (I547673,I548010);
nand I_32077 (I548041,I547993,I547931);
and I_32078 (I548058,I547753,I548041);
DFFARX1 I_32079  ( .D(I548058), .CLK(I2702), .RSTB(I547702), .Q(I547664) );
DFFARX1 I_32080  ( .D(I615562), .CLK(I2702), .RSTB(I547702), .Q(I548089) );
nand I_32081 (I548106,I548089,I547753);
and I_32082 (I548123,I547931,I548106);
DFFARX1 I_32083  ( .D(I548123), .CLK(I2702), .RSTB(I547702), .Q(I547694) );
not I_32084 (I548154,I548089);
nor I_32085 (I548171,I547770,I548154);
and I_32086 (I548188,I548089,I548171);
or I_32087 (I548205,I547993,I548188);
DFFARX1 I_32088  ( .D(I548205), .CLK(I2702), .RSTB(I547702), .Q(I547679) );
nand I_32089 (I547676,I548089,I547835);
DFFARX1 I_32090  ( .D(I548089), .CLK(I2702), .RSTB(I547702), .Q(I547667) );
not I_32091 (I548297,I2709);
nand I_32092 (I548314,I474914,I474917);
and I_32093 (I548331,I548314,I474911);
DFFARX1 I_32094  ( .D(I548331), .CLK(I2702), .RSTB(I548297), .Q(I548348) );
nor I_32095 (I548365,I474908,I474917);
nor I_32096 (I548382,I548365,I548348);
not I_32097 (I548280,I548365);
DFFARX1 I_32098  ( .D(I474890), .CLK(I2702), .RSTB(I548297), .Q(I548413) );
not I_32099 (I548430,I548413);
nor I_32100 (I548447,I548365,I548430);
nand I_32101 (I548283,I548413,I548382);
DFFARX1 I_32102  ( .D(I548413), .CLK(I2702), .RSTB(I548297), .Q(I548265) );
nand I_32103 (I548492,I474899,I474896);
and I_32104 (I548509,I548492,I474905);
DFFARX1 I_32105  ( .D(I548509), .CLK(I2702), .RSTB(I548297), .Q(I548526) );
nor I_32106 (I548286,I548526,I548348);
nand I_32107 (I548277,I548526,I548447);
DFFARX1 I_32108  ( .D(I474887), .CLK(I2702), .RSTB(I548297), .Q(I548571) );
and I_32109 (I548588,I548571,I474902);
DFFARX1 I_32110  ( .D(I548588), .CLK(I2702), .RSTB(I548297), .Q(I548605) );
not I_32111 (I548268,I548605);
nand I_32112 (I548636,I548588,I548526);
and I_32113 (I548653,I548348,I548636);
DFFARX1 I_32114  ( .D(I548653), .CLK(I2702), .RSTB(I548297), .Q(I548259) );
DFFARX1 I_32115  ( .D(I474893), .CLK(I2702), .RSTB(I548297), .Q(I548684) );
nand I_32116 (I548701,I548684,I548348);
and I_32117 (I548718,I548526,I548701);
DFFARX1 I_32118  ( .D(I548718), .CLK(I2702), .RSTB(I548297), .Q(I548289) );
not I_32119 (I548749,I548684);
nor I_32120 (I548766,I548365,I548749);
and I_32121 (I548783,I548684,I548766);
or I_32122 (I548800,I548588,I548783);
DFFARX1 I_32123  ( .D(I548800), .CLK(I2702), .RSTB(I548297), .Q(I548274) );
nand I_32124 (I548271,I548684,I548430);
DFFARX1 I_32125  ( .D(I548684), .CLK(I2702), .RSTB(I548297), .Q(I548262) );
not I_32126 (I548892,I2709);
nand I_32127 (I548909,I462776,I462779);
and I_32128 (I548926,I548909,I462773);
DFFARX1 I_32129  ( .D(I548926), .CLK(I2702), .RSTB(I548892), .Q(I548943) );
nor I_32130 (I548960,I462770,I462779);
nor I_32131 (I548977,I548960,I548943);
not I_32132 (I548875,I548960);
DFFARX1 I_32133  ( .D(I462752), .CLK(I2702), .RSTB(I548892), .Q(I549008) );
not I_32134 (I549025,I549008);
nor I_32135 (I549042,I548960,I549025);
nand I_32136 (I548878,I549008,I548977);
DFFARX1 I_32137  ( .D(I549008), .CLK(I2702), .RSTB(I548892), .Q(I548860) );
nand I_32138 (I549087,I462761,I462758);
and I_32139 (I549104,I549087,I462767);
DFFARX1 I_32140  ( .D(I549104), .CLK(I2702), .RSTB(I548892), .Q(I549121) );
nor I_32141 (I548881,I549121,I548943);
nand I_32142 (I548872,I549121,I549042);
DFFARX1 I_32143  ( .D(I462749), .CLK(I2702), .RSTB(I548892), .Q(I549166) );
and I_32144 (I549183,I549166,I462764);
DFFARX1 I_32145  ( .D(I549183), .CLK(I2702), .RSTB(I548892), .Q(I549200) );
not I_32146 (I548863,I549200);
nand I_32147 (I549231,I549183,I549121);
and I_32148 (I549248,I548943,I549231);
DFFARX1 I_32149  ( .D(I549248), .CLK(I2702), .RSTB(I548892), .Q(I548854) );
DFFARX1 I_32150  ( .D(I462755), .CLK(I2702), .RSTB(I548892), .Q(I549279) );
nand I_32151 (I549296,I549279,I548943);
and I_32152 (I549313,I549121,I549296);
DFFARX1 I_32153  ( .D(I549313), .CLK(I2702), .RSTB(I548892), .Q(I548884) );
not I_32154 (I549344,I549279);
nor I_32155 (I549361,I548960,I549344);
and I_32156 (I549378,I549279,I549361);
or I_32157 (I549395,I549183,I549378);
DFFARX1 I_32158  ( .D(I549395), .CLK(I2702), .RSTB(I548892), .Q(I548869) );
nand I_32159 (I548866,I549279,I549025);
DFFARX1 I_32160  ( .D(I549279), .CLK(I2702), .RSTB(I548892), .Q(I548857) );
not I_32161 (I549487,I2709);
nand I_32162 (I549504,I699622,I699628);
and I_32163 (I549521,I549504,I699619);
DFFARX1 I_32164  ( .D(I549521), .CLK(I2702), .RSTB(I549487), .Q(I549538) );
nor I_32165 (I549555,I699631,I699628);
nor I_32166 (I549572,I549555,I549538);
not I_32167 (I549470,I549555);
DFFARX1 I_32168  ( .D(I699610), .CLK(I2702), .RSTB(I549487), .Q(I549603) );
not I_32169 (I549620,I549603);
nor I_32170 (I549637,I549555,I549620);
nand I_32171 (I549473,I549603,I549572);
DFFARX1 I_32172  ( .D(I549603), .CLK(I2702), .RSTB(I549487), .Q(I549455) );
nand I_32173 (I549682,I699634,I699616);
and I_32174 (I549699,I549682,I699625);
DFFARX1 I_32175  ( .D(I549699), .CLK(I2702), .RSTB(I549487), .Q(I549716) );
nor I_32176 (I549476,I549716,I549538);
nand I_32177 (I549467,I549716,I549637);
DFFARX1 I_32178  ( .D(I699640), .CLK(I2702), .RSTB(I549487), .Q(I549761) );
and I_32179 (I549778,I549761,I699613);
DFFARX1 I_32180  ( .D(I549778), .CLK(I2702), .RSTB(I549487), .Q(I549795) );
not I_32181 (I549458,I549795);
nand I_32182 (I549826,I549778,I549716);
and I_32183 (I549843,I549538,I549826);
DFFARX1 I_32184  ( .D(I549843), .CLK(I2702), .RSTB(I549487), .Q(I549449) );
DFFARX1 I_32185  ( .D(I699637), .CLK(I2702), .RSTB(I549487), .Q(I549874) );
nand I_32186 (I549891,I549874,I549538);
and I_32187 (I549908,I549716,I549891);
DFFARX1 I_32188  ( .D(I549908), .CLK(I2702), .RSTB(I549487), .Q(I549479) );
not I_32189 (I549939,I549874);
nor I_32190 (I549956,I549555,I549939);
and I_32191 (I549973,I549874,I549956);
or I_32192 (I549990,I549778,I549973);
DFFARX1 I_32193  ( .D(I549990), .CLK(I2702), .RSTB(I549487), .Q(I549464) );
nand I_32194 (I549461,I549874,I549620);
DFFARX1 I_32195  ( .D(I549874), .CLK(I2702), .RSTB(I549487), .Q(I549452) );
not I_32196 (I550082,I2709);
nand I_32197 (I550099,I583974,I583965);
and I_32198 (I550116,I550099,I583983);
DFFARX1 I_32199  ( .D(I550116), .CLK(I2702), .RSTB(I550082), .Q(I550133) );
nor I_32200 (I550150,I583962,I583965);
nor I_32201 (I550167,I550150,I550133);
not I_32202 (I550065,I550150);
DFFARX1 I_32203  ( .D(I583971), .CLK(I2702), .RSTB(I550082), .Q(I550198) );
not I_32204 (I550215,I550198);
nor I_32205 (I550232,I550150,I550215);
nand I_32206 (I550068,I550198,I550167);
DFFARX1 I_32207  ( .D(I550198), .CLK(I2702), .RSTB(I550082), .Q(I550050) );
nand I_32208 (I550277,I583986,I583968);
and I_32209 (I550294,I550277,I583989);
DFFARX1 I_32210  ( .D(I550294), .CLK(I2702), .RSTB(I550082), .Q(I550311) );
nor I_32211 (I550071,I550311,I550133);
nand I_32212 (I550062,I550311,I550232);
DFFARX1 I_32213  ( .D(I583977), .CLK(I2702), .RSTB(I550082), .Q(I550356) );
and I_32214 (I550373,I550356,I583959);
DFFARX1 I_32215  ( .D(I550373), .CLK(I2702), .RSTB(I550082), .Q(I550390) );
not I_32216 (I550053,I550390);
nand I_32217 (I550421,I550373,I550311);
and I_32218 (I550438,I550133,I550421);
DFFARX1 I_32219  ( .D(I550438), .CLK(I2702), .RSTB(I550082), .Q(I550044) );
DFFARX1 I_32220  ( .D(I583980), .CLK(I2702), .RSTB(I550082), .Q(I550469) );
nand I_32221 (I550486,I550469,I550133);
and I_32222 (I550503,I550311,I550486);
DFFARX1 I_32223  ( .D(I550503), .CLK(I2702), .RSTB(I550082), .Q(I550074) );
not I_32224 (I550534,I550469);
nor I_32225 (I550551,I550150,I550534);
and I_32226 (I550568,I550469,I550551);
or I_32227 (I550585,I550373,I550568);
DFFARX1 I_32228  ( .D(I550585), .CLK(I2702), .RSTB(I550082), .Q(I550059) );
nand I_32229 (I550056,I550469,I550215);
DFFARX1 I_32230  ( .D(I550469), .CLK(I2702), .RSTB(I550082), .Q(I550047) );
not I_32231 (I550677,I2709);
nand I_32232 (I550694,I428507,I428495);
and I_32233 (I550711,I550694,I428501);
DFFARX1 I_32234  ( .D(I550711), .CLK(I2702), .RSTB(I550677), .Q(I550728) );
nor I_32235 (I550745,I428492,I428495);
nor I_32236 (I550762,I550745,I550728);
not I_32237 (I550660,I550745);
DFFARX1 I_32238  ( .D(I428477), .CLK(I2702), .RSTB(I550677), .Q(I550793) );
not I_32239 (I550810,I550793);
nor I_32240 (I550827,I550745,I550810);
nand I_32241 (I550663,I550793,I550762);
DFFARX1 I_32242  ( .D(I550793), .CLK(I2702), .RSTB(I550677), .Q(I550645) );
nand I_32243 (I550872,I428486,I428504);
and I_32244 (I550889,I550872,I428498);
DFFARX1 I_32245  ( .D(I550889), .CLK(I2702), .RSTB(I550677), .Q(I550906) );
nor I_32246 (I550666,I550906,I550728);
nand I_32247 (I550657,I550906,I550827);
DFFARX1 I_32248  ( .D(I428489), .CLK(I2702), .RSTB(I550677), .Q(I550951) );
and I_32249 (I550968,I550951,I428483);
DFFARX1 I_32250  ( .D(I550968), .CLK(I2702), .RSTB(I550677), .Q(I550985) );
not I_32251 (I550648,I550985);
nand I_32252 (I551016,I550968,I550906);
and I_32253 (I551033,I550728,I551016);
DFFARX1 I_32254  ( .D(I551033), .CLK(I2702), .RSTB(I550677), .Q(I550639) );
DFFARX1 I_32255  ( .D(I428480), .CLK(I2702), .RSTB(I550677), .Q(I551064) );
nand I_32256 (I551081,I551064,I550728);
and I_32257 (I551098,I550906,I551081);
DFFARX1 I_32258  ( .D(I551098), .CLK(I2702), .RSTB(I550677), .Q(I550669) );
not I_32259 (I551129,I551064);
nor I_32260 (I551146,I550745,I551129);
and I_32261 (I551163,I551064,I551146);
or I_32262 (I551180,I550968,I551163);
DFFARX1 I_32263  ( .D(I551180), .CLK(I2702), .RSTB(I550677), .Q(I550654) );
nand I_32264 (I550651,I551064,I550810);
DFFARX1 I_32265  ( .D(I551064), .CLK(I2702), .RSTB(I550677), .Q(I550642) );
not I_32266 (I551272,I2709);
nand I_32267 (I551289,I650804,I650795);
and I_32268 (I551306,I551289,I650813);
DFFARX1 I_32269  ( .D(I551306), .CLK(I2702), .RSTB(I551272), .Q(I551323) );
nor I_32270 (I551340,I650810,I650795);
nor I_32271 (I551357,I551340,I551323);
not I_32272 (I551255,I551340);
DFFARX1 I_32273  ( .D(I650792), .CLK(I2702), .RSTB(I551272), .Q(I551388) );
not I_32274 (I551405,I551388);
nor I_32275 (I551422,I551340,I551405);
nand I_32276 (I551258,I551388,I551357);
DFFARX1 I_32277  ( .D(I551388), .CLK(I2702), .RSTB(I551272), .Q(I551240) );
nand I_32278 (I551467,I650801,I650816);
and I_32279 (I551484,I551467,I650807);
DFFARX1 I_32280  ( .D(I551484), .CLK(I2702), .RSTB(I551272), .Q(I551501) );
nor I_32281 (I551261,I551501,I551323);
nand I_32282 (I551252,I551501,I551422);
DFFARX1 I_32283  ( .D(I650789), .CLK(I2702), .RSTB(I551272), .Q(I551546) );
and I_32284 (I551563,I551546,I650798);
DFFARX1 I_32285  ( .D(I551563), .CLK(I2702), .RSTB(I551272), .Q(I551580) );
not I_32286 (I551243,I551580);
nand I_32287 (I551611,I551563,I551501);
and I_32288 (I551628,I551323,I551611);
DFFARX1 I_32289  ( .D(I551628), .CLK(I2702), .RSTB(I551272), .Q(I551234) );
DFFARX1 I_32290  ( .D(I650786), .CLK(I2702), .RSTB(I551272), .Q(I551659) );
nand I_32291 (I551676,I551659,I551323);
and I_32292 (I551693,I551501,I551676);
DFFARX1 I_32293  ( .D(I551693), .CLK(I2702), .RSTB(I551272), .Q(I551264) );
not I_32294 (I551724,I551659);
nor I_32295 (I551741,I551340,I551724);
and I_32296 (I551758,I551659,I551741);
or I_32297 (I551775,I551563,I551758);
DFFARX1 I_32298  ( .D(I551775), .CLK(I2702), .RSTB(I551272), .Q(I551249) );
nand I_32299 (I551246,I551659,I551405);
DFFARX1 I_32300  ( .D(I551659), .CLK(I2702), .RSTB(I551272), .Q(I551237) );
not I_32301 (I551867,I2709);
nand I_32302 (I551884,I382901,I382913);
and I_32303 (I551901,I551884,I382895);
DFFARX1 I_32304  ( .D(I551901), .CLK(I2702), .RSTB(I551867), .Q(I551918) );
nor I_32305 (I551935,I382907,I382913);
nor I_32306 (I551952,I551935,I551918);
not I_32307 (I551850,I551935);
DFFARX1 I_32308  ( .D(I382892), .CLK(I2702), .RSTB(I551867), .Q(I551983) );
not I_32309 (I552000,I551983);
nor I_32310 (I552017,I551935,I552000);
nand I_32311 (I551853,I551983,I551952);
DFFARX1 I_32312  ( .D(I551983), .CLK(I2702), .RSTB(I551867), .Q(I551835) );
nand I_32313 (I552062,I382883,I382898);
and I_32314 (I552079,I552062,I382889);
DFFARX1 I_32315  ( .D(I552079), .CLK(I2702), .RSTB(I551867), .Q(I552096) );
nor I_32316 (I551856,I552096,I551918);
nand I_32317 (I551847,I552096,I552017);
DFFARX1 I_32318  ( .D(I382910), .CLK(I2702), .RSTB(I551867), .Q(I552141) );
and I_32319 (I552158,I552141,I382904);
DFFARX1 I_32320  ( .D(I552158), .CLK(I2702), .RSTB(I551867), .Q(I552175) );
not I_32321 (I551838,I552175);
nand I_32322 (I552206,I552158,I552096);
and I_32323 (I552223,I551918,I552206);
DFFARX1 I_32324  ( .D(I552223), .CLK(I2702), .RSTB(I551867), .Q(I551829) );
DFFARX1 I_32325  ( .D(I382886), .CLK(I2702), .RSTB(I551867), .Q(I552254) );
nand I_32326 (I552271,I552254,I551918);
and I_32327 (I552288,I552096,I552271);
DFFARX1 I_32328  ( .D(I552288), .CLK(I2702), .RSTB(I551867), .Q(I551859) );
not I_32329 (I552319,I552254);
nor I_32330 (I552336,I551935,I552319);
and I_32331 (I552353,I552254,I552336);
or I_32332 (I552370,I552158,I552353);
DFFARX1 I_32333  ( .D(I552370), .CLK(I2702), .RSTB(I551867), .Q(I551844) );
nand I_32334 (I551841,I552254,I552000);
DFFARX1 I_32335  ( .D(I552254), .CLK(I2702), .RSTB(I551867), .Q(I551832) );
not I_32336 (I552462,I2709);
nand I_32337 (I552479,I102086,I102098);
and I_32338 (I552496,I552479,I102107);
DFFARX1 I_32339  ( .D(I552496), .CLK(I2702), .RSTB(I552462), .Q(I552513) );
nor I_32340 (I552530,I102101,I102098);
nor I_32341 (I552547,I552530,I552513);
not I_32342 (I552445,I552530);
DFFARX1 I_32343  ( .D(I102095), .CLK(I2702), .RSTB(I552462), .Q(I552578) );
not I_32344 (I552595,I552578);
nor I_32345 (I552612,I552530,I552595);
nand I_32346 (I552448,I552578,I552547);
DFFARX1 I_32347  ( .D(I552578), .CLK(I2702), .RSTB(I552462), .Q(I552430) );
nand I_32348 (I552657,I102092,I102089);
and I_32349 (I552674,I552657,I102080);
DFFARX1 I_32350  ( .D(I552674), .CLK(I2702), .RSTB(I552462), .Q(I552691) );
nor I_32351 (I552451,I552691,I552513);
nand I_32352 (I552442,I552691,I552612);
DFFARX1 I_32353  ( .D(I102104), .CLK(I2702), .RSTB(I552462), .Q(I552736) );
and I_32354 (I552753,I552736,I102083);
DFFARX1 I_32355  ( .D(I552753), .CLK(I2702), .RSTB(I552462), .Q(I552770) );
not I_32356 (I552433,I552770);
nand I_32357 (I552801,I552753,I552691);
and I_32358 (I552818,I552513,I552801);
DFFARX1 I_32359  ( .D(I552818), .CLK(I2702), .RSTB(I552462), .Q(I552424) );
DFFARX1 I_32360  ( .D(I102077), .CLK(I2702), .RSTB(I552462), .Q(I552849) );
nand I_32361 (I552866,I552849,I552513);
and I_32362 (I552883,I552691,I552866);
DFFARX1 I_32363  ( .D(I552883), .CLK(I2702), .RSTB(I552462), .Q(I552454) );
not I_32364 (I552914,I552849);
nor I_32365 (I552931,I552530,I552914);
and I_32366 (I552948,I552849,I552931);
or I_32367 (I552965,I552753,I552948);
DFFARX1 I_32368  ( .D(I552965), .CLK(I2702), .RSTB(I552462), .Q(I552439) );
nand I_32369 (I552436,I552849,I552595);
DFFARX1 I_32370  ( .D(I552849), .CLK(I2702), .RSTB(I552462), .Q(I552427) );
not I_32371 (I553057,I2709);
nand I_32372 (I553074,I6642,I6648);
and I_32373 (I553091,I553074,I6645);
DFFARX1 I_32374  ( .D(I553091), .CLK(I2702), .RSTB(I553057), .Q(I553108) );
nor I_32375 (I553125,I6669,I6648);
nor I_32376 (I553142,I553125,I553108);
not I_32377 (I553040,I553125);
DFFARX1 I_32378  ( .D(I6660), .CLK(I2702), .RSTB(I553057), .Q(I553173) );
not I_32379 (I553190,I553173);
nor I_32380 (I553207,I553125,I553190);
nand I_32381 (I553043,I553173,I553142);
DFFARX1 I_32382  ( .D(I553173), .CLK(I2702), .RSTB(I553057), .Q(I553025) );
nand I_32383 (I553252,I6663,I6666);
and I_32384 (I553269,I553252,I6639);
DFFARX1 I_32385  ( .D(I553269), .CLK(I2702), .RSTB(I553057), .Q(I553286) );
nor I_32386 (I553046,I553286,I553108);
nand I_32387 (I553037,I553286,I553207);
DFFARX1 I_32388  ( .D(I6657), .CLK(I2702), .RSTB(I553057), .Q(I553331) );
and I_32389 (I553348,I553331,I6651);
DFFARX1 I_32390  ( .D(I553348), .CLK(I2702), .RSTB(I553057), .Q(I553365) );
not I_32391 (I553028,I553365);
nand I_32392 (I553396,I553348,I553286);
and I_32393 (I553413,I553108,I553396);
DFFARX1 I_32394  ( .D(I553413), .CLK(I2702), .RSTB(I553057), .Q(I553019) );
DFFARX1 I_32395  ( .D(I6654), .CLK(I2702), .RSTB(I553057), .Q(I553444) );
nand I_32396 (I553461,I553444,I553108);
and I_32397 (I553478,I553286,I553461);
DFFARX1 I_32398  ( .D(I553478), .CLK(I2702), .RSTB(I553057), .Q(I553049) );
not I_32399 (I553509,I553444);
nor I_32400 (I553526,I553125,I553509);
and I_32401 (I553543,I553444,I553526);
or I_32402 (I553560,I553348,I553543);
DFFARX1 I_32403  ( .D(I553560), .CLK(I2702), .RSTB(I553057), .Q(I553034) );
nand I_32404 (I553031,I553444,I553190);
DFFARX1 I_32405  ( .D(I553444), .CLK(I2702), .RSTB(I553057), .Q(I553022) );
not I_32406 (I553652,I2709);
nand I_32407 (I553669,I274815,I274821);
and I_32408 (I553686,I553669,I274803);
DFFARX1 I_32409  ( .D(I553686), .CLK(I2702), .RSTB(I553652), .Q(I553703) );
nor I_32410 (I553720,I274797,I274821);
nor I_32411 (I553737,I553720,I553703);
not I_32412 (I553635,I553720);
DFFARX1 I_32413  ( .D(I274827), .CLK(I2702), .RSTB(I553652), .Q(I553768) );
not I_32414 (I553785,I553768);
nor I_32415 (I553802,I553720,I553785);
nand I_32416 (I553638,I553768,I553737);
DFFARX1 I_32417  ( .D(I553768), .CLK(I2702), .RSTB(I553652), .Q(I553620) );
nand I_32418 (I553847,I274818,I274809);
and I_32419 (I553864,I553847,I274812);
DFFARX1 I_32420  ( .D(I553864), .CLK(I2702), .RSTB(I553652), .Q(I553881) );
nor I_32421 (I553641,I553881,I553703);
nand I_32422 (I553632,I553881,I553802);
DFFARX1 I_32423  ( .D(I274824), .CLK(I2702), .RSTB(I553652), .Q(I553926) );
and I_32424 (I553943,I553926,I274800);
DFFARX1 I_32425  ( .D(I553943), .CLK(I2702), .RSTB(I553652), .Q(I553960) );
not I_32426 (I553623,I553960);
nand I_32427 (I553991,I553943,I553881);
and I_32428 (I554008,I553703,I553991);
DFFARX1 I_32429  ( .D(I554008), .CLK(I2702), .RSTB(I553652), .Q(I553614) );
DFFARX1 I_32430  ( .D(I274806), .CLK(I2702), .RSTB(I553652), .Q(I554039) );
nand I_32431 (I554056,I554039,I553703);
and I_32432 (I554073,I553881,I554056);
DFFARX1 I_32433  ( .D(I554073), .CLK(I2702), .RSTB(I553652), .Q(I553644) );
not I_32434 (I554104,I554039);
nor I_32435 (I554121,I553720,I554104);
and I_32436 (I554138,I554039,I554121);
or I_32437 (I554155,I553943,I554138);
DFFARX1 I_32438  ( .D(I554155), .CLK(I2702), .RSTB(I553652), .Q(I553629) );
nand I_32439 (I553626,I554039,I553785);
DFFARX1 I_32440  ( .D(I554039), .CLK(I2702), .RSTB(I553652), .Q(I553617) );
not I_32441 (I554247,I2709);
nand I_32442 (I554264,I431564,I431567);
and I_32443 (I554281,I554264,I431561);
DFFARX1 I_32444  ( .D(I554281), .CLK(I2702), .RSTB(I554247), .Q(I554298) );
nor I_32445 (I554315,I431558,I431567);
nor I_32446 (I554332,I554315,I554298);
not I_32447 (I554230,I554315);
DFFARX1 I_32448  ( .D(I431540), .CLK(I2702), .RSTB(I554247), .Q(I554363) );
not I_32449 (I554380,I554363);
nor I_32450 (I554397,I554315,I554380);
nand I_32451 (I554233,I554363,I554332);
DFFARX1 I_32452  ( .D(I554363), .CLK(I2702), .RSTB(I554247), .Q(I554215) );
nand I_32453 (I554442,I431549,I431546);
and I_32454 (I554459,I554442,I431555);
DFFARX1 I_32455  ( .D(I554459), .CLK(I2702), .RSTB(I554247), .Q(I554476) );
nor I_32456 (I554236,I554476,I554298);
nand I_32457 (I554227,I554476,I554397);
DFFARX1 I_32458  ( .D(I431537), .CLK(I2702), .RSTB(I554247), .Q(I554521) );
and I_32459 (I554538,I554521,I431552);
DFFARX1 I_32460  ( .D(I554538), .CLK(I2702), .RSTB(I554247), .Q(I554555) );
not I_32461 (I554218,I554555);
nand I_32462 (I554586,I554538,I554476);
and I_32463 (I554603,I554298,I554586);
DFFARX1 I_32464  ( .D(I554603), .CLK(I2702), .RSTB(I554247), .Q(I554209) );
DFFARX1 I_32465  ( .D(I431543), .CLK(I2702), .RSTB(I554247), .Q(I554634) );
nand I_32466 (I554651,I554634,I554298);
and I_32467 (I554668,I554476,I554651);
DFFARX1 I_32468  ( .D(I554668), .CLK(I2702), .RSTB(I554247), .Q(I554239) );
not I_32469 (I554699,I554634);
nor I_32470 (I554716,I554315,I554699);
and I_32471 (I554733,I554634,I554716);
or I_32472 (I554750,I554538,I554733);
DFFARX1 I_32473  ( .D(I554750), .CLK(I2702), .RSTB(I554247), .Q(I554224) );
nand I_32474 (I554221,I554634,I554380);
DFFARX1 I_32475  ( .D(I554634), .CLK(I2702), .RSTB(I554247), .Q(I554212) );
not I_32476 (I554842,I2709);
nand I_32477 (I554859,I363521,I363533);
and I_32478 (I554876,I554859,I363515);
DFFARX1 I_32479  ( .D(I554876), .CLK(I2702), .RSTB(I554842), .Q(I554893) );
nor I_32480 (I554910,I363527,I363533);
nor I_32481 (I554927,I554910,I554893);
not I_32482 (I554825,I554910);
DFFARX1 I_32483  ( .D(I363512), .CLK(I2702), .RSTB(I554842), .Q(I554958) );
not I_32484 (I554975,I554958);
nor I_32485 (I554992,I554910,I554975);
nand I_32486 (I554828,I554958,I554927);
DFFARX1 I_32487  ( .D(I554958), .CLK(I2702), .RSTB(I554842), .Q(I554810) );
nand I_32488 (I555037,I363503,I363518);
and I_32489 (I555054,I555037,I363509);
DFFARX1 I_32490  ( .D(I555054), .CLK(I2702), .RSTB(I554842), .Q(I555071) );
nor I_32491 (I554831,I555071,I554893);
nand I_32492 (I554822,I555071,I554992);
DFFARX1 I_32493  ( .D(I363530), .CLK(I2702), .RSTB(I554842), .Q(I555116) );
and I_32494 (I555133,I555116,I363524);
DFFARX1 I_32495  ( .D(I555133), .CLK(I2702), .RSTB(I554842), .Q(I555150) );
not I_32496 (I554813,I555150);
nand I_32497 (I555181,I555133,I555071);
and I_32498 (I555198,I554893,I555181);
DFFARX1 I_32499  ( .D(I555198), .CLK(I2702), .RSTB(I554842), .Q(I554804) );
DFFARX1 I_32500  ( .D(I363506), .CLK(I2702), .RSTB(I554842), .Q(I555229) );
nand I_32501 (I555246,I555229,I554893);
and I_32502 (I555263,I555071,I555246);
DFFARX1 I_32503  ( .D(I555263), .CLK(I2702), .RSTB(I554842), .Q(I554834) );
not I_32504 (I555294,I555229);
nor I_32505 (I555311,I554910,I555294);
and I_32506 (I555328,I555229,I555311);
or I_32507 (I555345,I555133,I555328);
DFFARX1 I_32508  ( .D(I555345), .CLK(I2702), .RSTB(I554842), .Q(I554819) );
nand I_32509 (I554816,I555229,I554975);
DFFARX1 I_32510  ( .D(I555229), .CLK(I2702), .RSTB(I554842), .Q(I554807) );
not I_32511 (I555437,I2709);
nand I_32512 (I555454,I667158,I667149);
and I_32513 (I555471,I555454,I667167);
DFFARX1 I_32514  ( .D(I555471), .CLK(I2702), .RSTB(I555437), .Q(I555488) );
nor I_32515 (I555505,I667164,I667149);
nor I_32516 (I555522,I555505,I555488);
not I_32517 (I555420,I555505);
DFFARX1 I_32518  ( .D(I667146), .CLK(I2702), .RSTB(I555437), .Q(I555553) );
not I_32519 (I555570,I555553);
nor I_32520 (I555587,I555505,I555570);
nand I_32521 (I555423,I555553,I555522);
DFFARX1 I_32522  ( .D(I555553), .CLK(I2702), .RSTB(I555437), .Q(I555405) );
nand I_32523 (I555632,I667155,I667170);
and I_32524 (I555649,I555632,I667161);
DFFARX1 I_32525  ( .D(I555649), .CLK(I2702), .RSTB(I555437), .Q(I555666) );
nor I_32526 (I555426,I555666,I555488);
nand I_32527 (I555417,I555666,I555587);
DFFARX1 I_32528  ( .D(I667143), .CLK(I2702), .RSTB(I555437), .Q(I555711) );
and I_32529 (I555728,I555711,I667152);
DFFARX1 I_32530  ( .D(I555728), .CLK(I2702), .RSTB(I555437), .Q(I555745) );
not I_32531 (I555408,I555745);
nand I_32532 (I555776,I555728,I555666);
and I_32533 (I555793,I555488,I555776);
DFFARX1 I_32534  ( .D(I555793), .CLK(I2702), .RSTB(I555437), .Q(I555399) );
DFFARX1 I_32535  ( .D(I667140), .CLK(I2702), .RSTB(I555437), .Q(I555824) );
nand I_32536 (I555841,I555824,I555488);
and I_32537 (I555858,I555666,I555841);
DFFARX1 I_32538  ( .D(I555858), .CLK(I2702), .RSTB(I555437), .Q(I555429) );
not I_32539 (I555889,I555824);
nor I_32540 (I555906,I555505,I555889);
and I_32541 (I555923,I555824,I555906);
or I_32542 (I555940,I555728,I555923);
DFFARX1 I_32543  ( .D(I555940), .CLK(I2702), .RSTB(I555437), .Q(I555414) );
nand I_32544 (I555411,I555824,I555570);
DFFARX1 I_32545  ( .D(I555824), .CLK(I2702), .RSTB(I555437), .Q(I555402) );
not I_32546 (I556032,I2709);
nand I_32547 (I556049,I437922,I437925);
and I_32548 (I556066,I556049,I437919);
DFFARX1 I_32549  ( .D(I556066), .CLK(I2702), .RSTB(I556032), .Q(I556083) );
nor I_32550 (I556100,I437916,I437925);
nor I_32551 (I556117,I556100,I556083);
not I_32552 (I556015,I556100);
DFFARX1 I_32553  ( .D(I437898), .CLK(I2702), .RSTB(I556032), .Q(I556148) );
not I_32554 (I556165,I556148);
nor I_32555 (I556182,I556100,I556165);
nand I_32556 (I556018,I556148,I556117);
DFFARX1 I_32557  ( .D(I556148), .CLK(I2702), .RSTB(I556032), .Q(I556000) );
nand I_32558 (I556227,I437907,I437904);
and I_32559 (I556244,I556227,I437913);
DFFARX1 I_32560  ( .D(I556244), .CLK(I2702), .RSTB(I556032), .Q(I556261) );
nor I_32561 (I556021,I556261,I556083);
nand I_32562 (I556012,I556261,I556182);
DFFARX1 I_32563  ( .D(I437895), .CLK(I2702), .RSTB(I556032), .Q(I556306) );
and I_32564 (I556323,I556306,I437910);
DFFARX1 I_32565  ( .D(I556323), .CLK(I2702), .RSTB(I556032), .Q(I556340) );
not I_32566 (I556003,I556340);
nand I_32567 (I556371,I556323,I556261);
and I_32568 (I556388,I556083,I556371);
DFFARX1 I_32569  ( .D(I556388), .CLK(I2702), .RSTB(I556032), .Q(I555994) );
DFFARX1 I_32570  ( .D(I437901), .CLK(I2702), .RSTB(I556032), .Q(I556419) );
nand I_32571 (I556436,I556419,I556083);
and I_32572 (I556453,I556261,I556436);
DFFARX1 I_32573  ( .D(I556453), .CLK(I2702), .RSTB(I556032), .Q(I556024) );
not I_32574 (I556484,I556419);
nor I_32575 (I556501,I556100,I556484);
and I_32576 (I556518,I556419,I556501);
or I_32577 (I556535,I556323,I556518);
DFFARX1 I_32578  ( .D(I556535), .CLK(I2702), .RSTB(I556032), .Q(I556009) );
nand I_32579 (I556006,I556419,I556165);
DFFARX1 I_32580  ( .D(I556419), .CLK(I2702), .RSTB(I556032), .Q(I555997) );
not I_32581 (I556627,I2709);
nand I_32582 (I556644,I495623,I495611);
and I_32583 (I556661,I556644,I495608);
DFFARX1 I_32584  ( .D(I556661), .CLK(I2702), .RSTB(I556627), .Q(I556678) );
nor I_32585 (I556695,I495602,I495611);
nor I_32586 (I556712,I556695,I556678);
not I_32587 (I556610,I556695);
DFFARX1 I_32588  ( .D(I495617), .CLK(I2702), .RSTB(I556627), .Q(I556743) );
not I_32589 (I556760,I556743);
nor I_32590 (I556777,I556695,I556760);
nand I_32591 (I556613,I556743,I556712);
DFFARX1 I_32592  ( .D(I556743), .CLK(I2702), .RSTB(I556627), .Q(I556595) );
nand I_32593 (I556822,I495614,I495620);
and I_32594 (I556839,I556822,I495605);
DFFARX1 I_32595  ( .D(I556839), .CLK(I2702), .RSTB(I556627), .Q(I556856) );
nor I_32596 (I556616,I556856,I556678);
nand I_32597 (I556607,I556856,I556777);
DFFARX1 I_32598  ( .D(I495593), .CLK(I2702), .RSTB(I556627), .Q(I556901) );
and I_32599 (I556918,I556901,I495596);
DFFARX1 I_32600  ( .D(I556918), .CLK(I2702), .RSTB(I556627), .Q(I556935) );
not I_32601 (I556598,I556935);
nand I_32602 (I556966,I556918,I556856);
and I_32603 (I556983,I556678,I556966);
DFFARX1 I_32604  ( .D(I556983), .CLK(I2702), .RSTB(I556627), .Q(I556589) );
DFFARX1 I_32605  ( .D(I495599), .CLK(I2702), .RSTB(I556627), .Q(I557014) );
nand I_32606 (I557031,I557014,I556678);
and I_32607 (I557048,I556856,I557031);
DFFARX1 I_32608  ( .D(I557048), .CLK(I2702), .RSTB(I556627), .Q(I556619) );
not I_32609 (I557079,I557014);
nor I_32610 (I557096,I556695,I557079);
and I_32611 (I557113,I557014,I557096);
or I_32612 (I557130,I556918,I557113);
DFFARX1 I_32613  ( .D(I557130), .CLK(I2702), .RSTB(I556627), .Q(I556604) );
nand I_32614 (I556601,I557014,I556760);
DFFARX1 I_32615  ( .D(I557014), .CLK(I2702), .RSTB(I556627), .Q(I556592) );
not I_32616 (I557222,I2709);
nand I_32617 (I557239,I254925,I254931);
and I_32618 (I557256,I557239,I254913);
DFFARX1 I_32619  ( .D(I557256), .CLK(I2702), .RSTB(I557222), .Q(I557273) );
nor I_32620 (I557290,I254907,I254931);
nor I_32621 (I557307,I557290,I557273);
not I_32622 (I557205,I557290);
DFFARX1 I_32623  ( .D(I254937), .CLK(I2702), .RSTB(I557222), .Q(I557338) );
not I_32624 (I557355,I557338);
nor I_32625 (I557372,I557290,I557355);
nand I_32626 (I557208,I557338,I557307);
DFFARX1 I_32627  ( .D(I557338), .CLK(I2702), .RSTB(I557222), .Q(I557190) );
nand I_32628 (I557417,I254928,I254919);
and I_32629 (I557434,I557417,I254922);
DFFARX1 I_32630  ( .D(I557434), .CLK(I2702), .RSTB(I557222), .Q(I557451) );
nor I_32631 (I557211,I557451,I557273);
nand I_32632 (I557202,I557451,I557372);
DFFARX1 I_32633  ( .D(I254934), .CLK(I2702), .RSTB(I557222), .Q(I557496) );
and I_32634 (I557513,I557496,I254910);
DFFARX1 I_32635  ( .D(I557513), .CLK(I2702), .RSTB(I557222), .Q(I557530) );
not I_32636 (I557193,I557530);
nand I_32637 (I557561,I557513,I557451);
and I_32638 (I557578,I557273,I557561);
DFFARX1 I_32639  ( .D(I557578), .CLK(I2702), .RSTB(I557222), .Q(I557184) );
DFFARX1 I_32640  ( .D(I254916), .CLK(I2702), .RSTB(I557222), .Q(I557609) );
nand I_32641 (I557626,I557609,I557273);
and I_32642 (I557643,I557451,I557626);
DFFARX1 I_32643  ( .D(I557643), .CLK(I2702), .RSTB(I557222), .Q(I557214) );
not I_32644 (I557674,I557609);
nor I_32645 (I557691,I557290,I557674);
and I_32646 (I557708,I557609,I557691);
or I_32647 (I557725,I557513,I557708);
DFFARX1 I_32648  ( .D(I557725), .CLK(I2702), .RSTB(I557222), .Q(I557199) );
nand I_32649 (I557196,I557609,I557355);
DFFARX1 I_32650  ( .D(I557609), .CLK(I2702), .RSTB(I557222), .Q(I557187) );
not I_32651 (I557817,I2709);
nand I_32652 (I557834,I177354,I177366);
and I_32653 (I557851,I557834,I177345);
DFFARX1 I_32654  ( .D(I557851), .CLK(I2702), .RSTB(I557817), .Q(I557868) );
nor I_32655 (I557885,I177336,I177366);
nor I_32656 (I557902,I557885,I557868);
not I_32657 (I557800,I557885);
DFFARX1 I_32658  ( .D(I177348), .CLK(I2702), .RSTB(I557817), .Q(I557933) );
not I_32659 (I557950,I557933);
nor I_32660 (I557967,I557885,I557950);
nand I_32661 (I557803,I557933,I557902);
DFFARX1 I_32662  ( .D(I557933), .CLK(I2702), .RSTB(I557817), .Q(I557785) );
nand I_32663 (I558012,I177363,I177351);
and I_32664 (I558029,I558012,I177339);
DFFARX1 I_32665  ( .D(I558029), .CLK(I2702), .RSTB(I557817), .Q(I558046) );
nor I_32666 (I557806,I558046,I557868);
nand I_32667 (I557797,I558046,I557967);
DFFARX1 I_32668  ( .D(I177357), .CLK(I2702), .RSTB(I557817), .Q(I558091) );
and I_32669 (I558108,I558091,I177342);
DFFARX1 I_32670  ( .D(I558108), .CLK(I2702), .RSTB(I557817), .Q(I558125) );
not I_32671 (I557788,I558125);
nand I_32672 (I558156,I558108,I558046);
and I_32673 (I558173,I557868,I558156);
DFFARX1 I_32674  ( .D(I558173), .CLK(I2702), .RSTB(I557817), .Q(I557779) );
DFFARX1 I_32675  ( .D(I177360), .CLK(I2702), .RSTB(I557817), .Q(I558204) );
nand I_32676 (I558221,I558204,I557868);
and I_32677 (I558238,I558046,I558221);
DFFARX1 I_32678  ( .D(I558238), .CLK(I2702), .RSTB(I557817), .Q(I557809) );
not I_32679 (I558269,I558204);
nor I_32680 (I558286,I557885,I558269);
and I_32681 (I558303,I558204,I558286);
or I_32682 (I558320,I558108,I558303);
DFFARX1 I_32683  ( .D(I558320), .CLK(I2702), .RSTB(I557817), .Q(I557794) );
nand I_32684 (I557791,I558204,I557950);
DFFARX1 I_32685  ( .D(I558204), .CLK(I2702), .RSTB(I557817), .Q(I557782) );
not I_32686 (I558412,I2709);
nand I_32687 (I558429,I145530,I145542);
and I_32688 (I558446,I558429,I145521);
DFFARX1 I_32689  ( .D(I558446), .CLK(I2702), .RSTB(I558412), .Q(I558463) );
nor I_32690 (I558480,I145512,I145542);
nor I_32691 (I558497,I558480,I558463);
not I_32692 (I558395,I558480);
DFFARX1 I_32693  ( .D(I145524), .CLK(I2702), .RSTB(I558412), .Q(I558528) );
not I_32694 (I558545,I558528);
nor I_32695 (I558562,I558480,I558545);
nand I_32696 (I558398,I558528,I558497);
DFFARX1 I_32697  ( .D(I558528), .CLK(I2702), .RSTB(I558412), .Q(I558380) );
nand I_32698 (I558607,I145539,I145527);
and I_32699 (I558624,I558607,I145515);
DFFARX1 I_32700  ( .D(I558624), .CLK(I2702), .RSTB(I558412), .Q(I558641) );
nor I_32701 (I558401,I558641,I558463);
nand I_32702 (I558392,I558641,I558562);
DFFARX1 I_32703  ( .D(I145533), .CLK(I2702), .RSTB(I558412), .Q(I558686) );
and I_32704 (I558703,I558686,I145518);
DFFARX1 I_32705  ( .D(I558703), .CLK(I2702), .RSTB(I558412), .Q(I558720) );
not I_32706 (I558383,I558720);
nand I_32707 (I558751,I558703,I558641);
and I_32708 (I558768,I558463,I558751);
DFFARX1 I_32709  ( .D(I558768), .CLK(I2702), .RSTB(I558412), .Q(I558374) );
DFFARX1 I_32710  ( .D(I145536), .CLK(I2702), .RSTB(I558412), .Q(I558799) );
nand I_32711 (I558816,I558799,I558463);
and I_32712 (I558833,I558641,I558816);
DFFARX1 I_32713  ( .D(I558833), .CLK(I2702), .RSTB(I558412), .Q(I558404) );
not I_32714 (I558864,I558799);
nor I_32715 (I558881,I558480,I558864);
and I_32716 (I558898,I558799,I558881);
or I_32717 (I558915,I558703,I558898);
DFFARX1 I_32718  ( .D(I558915), .CLK(I2702), .RSTB(I558412), .Q(I558389) );
nand I_32719 (I558386,I558799,I558545);
DFFARX1 I_32720  ( .D(I558799), .CLK(I2702), .RSTB(I558412), .Q(I558377) );
not I_32721 (I559007,I2709);
nand I_32722 (I559024,I674077,I674068);
and I_32723 (I559041,I559024,I674086);
DFFARX1 I_32724  ( .D(I559041), .CLK(I2702), .RSTB(I559007), .Q(I559058) );
nor I_32725 (I559075,I674083,I674068);
nor I_32726 (I559092,I559075,I559058);
not I_32727 (I558990,I559075);
DFFARX1 I_32728  ( .D(I674065), .CLK(I2702), .RSTB(I559007), .Q(I559123) );
not I_32729 (I559140,I559123);
nor I_32730 (I559157,I559075,I559140);
nand I_32731 (I558993,I559123,I559092);
DFFARX1 I_32732  ( .D(I559123), .CLK(I2702), .RSTB(I559007), .Q(I558975) );
nand I_32733 (I559202,I674074,I674089);
and I_32734 (I559219,I559202,I674080);
DFFARX1 I_32735  ( .D(I559219), .CLK(I2702), .RSTB(I559007), .Q(I559236) );
nor I_32736 (I558996,I559236,I559058);
nand I_32737 (I558987,I559236,I559157);
DFFARX1 I_32738  ( .D(I674062), .CLK(I2702), .RSTB(I559007), .Q(I559281) );
and I_32739 (I559298,I559281,I674071);
DFFARX1 I_32740  ( .D(I559298), .CLK(I2702), .RSTB(I559007), .Q(I559315) );
not I_32741 (I558978,I559315);
nand I_32742 (I559346,I559298,I559236);
and I_32743 (I559363,I559058,I559346);
DFFARX1 I_32744  ( .D(I559363), .CLK(I2702), .RSTB(I559007), .Q(I558969) );
DFFARX1 I_32745  ( .D(I674059), .CLK(I2702), .RSTB(I559007), .Q(I559394) );
nand I_32746 (I559411,I559394,I559058);
and I_32747 (I559428,I559236,I559411);
DFFARX1 I_32748  ( .D(I559428), .CLK(I2702), .RSTB(I559007), .Q(I558999) );
not I_32749 (I559459,I559394);
nor I_32750 (I559476,I559075,I559459);
and I_32751 (I559493,I559394,I559476);
or I_32752 (I559510,I559298,I559493);
DFFARX1 I_32753  ( .D(I559510), .CLK(I2702), .RSTB(I559007), .Q(I558984) );
nand I_32754 (I558981,I559394,I559140);
DFFARX1 I_32755  ( .D(I559394), .CLK(I2702), .RSTB(I559007), .Q(I558972) );
not I_32756 (I559602,I2709);
nand I_32757 (I559619,I172713,I172725);
and I_32758 (I559636,I559619,I172704);
DFFARX1 I_32759  ( .D(I559636), .CLK(I2702), .RSTB(I559602), .Q(I559653) );
nor I_32760 (I559670,I172695,I172725);
nor I_32761 (I559687,I559670,I559653);
not I_32762 (I559585,I559670);
DFFARX1 I_32763  ( .D(I172707), .CLK(I2702), .RSTB(I559602), .Q(I559718) );
not I_32764 (I559735,I559718);
nor I_32765 (I559752,I559670,I559735);
nand I_32766 (I559588,I559718,I559687);
DFFARX1 I_32767  ( .D(I559718), .CLK(I2702), .RSTB(I559602), .Q(I559570) );
nand I_32768 (I559797,I172722,I172710);
and I_32769 (I559814,I559797,I172698);
DFFARX1 I_32770  ( .D(I559814), .CLK(I2702), .RSTB(I559602), .Q(I559831) );
nor I_32771 (I559591,I559831,I559653);
nand I_32772 (I559582,I559831,I559752);
DFFARX1 I_32773  ( .D(I172716), .CLK(I2702), .RSTB(I559602), .Q(I559876) );
and I_32774 (I559893,I559876,I172701);
DFFARX1 I_32775  ( .D(I559893), .CLK(I2702), .RSTB(I559602), .Q(I559910) );
not I_32776 (I559573,I559910);
nand I_32777 (I559941,I559893,I559831);
and I_32778 (I559958,I559653,I559941);
DFFARX1 I_32779  ( .D(I559958), .CLK(I2702), .RSTB(I559602), .Q(I559564) );
DFFARX1 I_32780  ( .D(I172719), .CLK(I2702), .RSTB(I559602), .Q(I559989) );
nand I_32781 (I560006,I559989,I559653);
and I_32782 (I560023,I559831,I560006);
DFFARX1 I_32783  ( .D(I560023), .CLK(I2702), .RSTB(I559602), .Q(I559594) );
not I_32784 (I560054,I559989);
nor I_32785 (I560071,I559670,I560054);
and I_32786 (I560088,I559989,I560071);
or I_32787 (I560105,I559893,I560088);
DFFARX1 I_32788  ( .D(I560105), .CLK(I2702), .RSTB(I559602), .Q(I559579) );
nand I_32789 (I559576,I559989,I559735);
DFFARX1 I_32790  ( .D(I559989), .CLK(I2702), .RSTB(I559602), .Q(I559567) );
not I_32791 (I560197,I2709);
nand I_32792 (I560214,I66556,I66568);
and I_32793 (I560231,I560214,I66577);
DFFARX1 I_32794  ( .D(I560231), .CLK(I2702), .RSTB(I560197), .Q(I560248) );
nor I_32795 (I560265,I66571,I66568);
nor I_32796 (I560282,I560265,I560248);
not I_32797 (I560180,I560265);
DFFARX1 I_32798  ( .D(I66565), .CLK(I2702), .RSTB(I560197), .Q(I560313) );
not I_32799 (I560330,I560313);
nor I_32800 (I560347,I560265,I560330);
nand I_32801 (I560183,I560313,I560282);
DFFARX1 I_32802  ( .D(I560313), .CLK(I2702), .RSTB(I560197), .Q(I560165) );
nand I_32803 (I560392,I66562,I66559);
and I_32804 (I560409,I560392,I66550);
DFFARX1 I_32805  ( .D(I560409), .CLK(I2702), .RSTB(I560197), .Q(I560426) );
nor I_32806 (I560186,I560426,I560248);
nand I_32807 (I560177,I560426,I560347);
DFFARX1 I_32808  ( .D(I66574), .CLK(I2702), .RSTB(I560197), .Q(I560471) );
and I_32809 (I560488,I560471,I66553);
DFFARX1 I_32810  ( .D(I560488), .CLK(I2702), .RSTB(I560197), .Q(I560505) );
not I_32811 (I560168,I560505);
nand I_32812 (I560536,I560488,I560426);
and I_32813 (I560553,I560248,I560536);
DFFARX1 I_32814  ( .D(I560553), .CLK(I2702), .RSTB(I560197), .Q(I560159) );
DFFARX1 I_32815  ( .D(I66547), .CLK(I2702), .RSTB(I560197), .Q(I560584) );
nand I_32816 (I560601,I560584,I560248);
and I_32817 (I560618,I560426,I560601);
DFFARX1 I_32818  ( .D(I560618), .CLK(I2702), .RSTB(I560197), .Q(I560189) );
not I_32819 (I560649,I560584);
nor I_32820 (I560666,I560265,I560649);
and I_32821 (I560683,I560584,I560666);
or I_32822 (I560700,I560488,I560683);
DFFARX1 I_32823  ( .D(I560700), .CLK(I2702), .RSTB(I560197), .Q(I560174) );
nand I_32824 (I560171,I560584,I560330);
DFFARX1 I_32825  ( .D(I560584), .CLK(I2702), .RSTB(I560197), .Q(I560162) );
not I_32826 (I560792,I2709);
nand I_32827 (I560809,I653320,I653311);
and I_32828 (I560826,I560809,I653329);
DFFARX1 I_32829  ( .D(I560826), .CLK(I2702), .RSTB(I560792), .Q(I560843) );
nor I_32830 (I560860,I653326,I653311);
nor I_32831 (I560877,I560860,I560843);
not I_32832 (I560775,I560860);
DFFARX1 I_32833  ( .D(I653308), .CLK(I2702), .RSTB(I560792), .Q(I560908) );
not I_32834 (I560925,I560908);
nor I_32835 (I560942,I560860,I560925);
nand I_32836 (I560778,I560908,I560877);
DFFARX1 I_32837  ( .D(I560908), .CLK(I2702), .RSTB(I560792), .Q(I560760) );
nand I_32838 (I560987,I653317,I653332);
and I_32839 (I561004,I560987,I653323);
DFFARX1 I_32840  ( .D(I561004), .CLK(I2702), .RSTB(I560792), .Q(I561021) );
nor I_32841 (I560781,I561021,I560843);
nand I_32842 (I560772,I561021,I560942);
DFFARX1 I_32843  ( .D(I653305), .CLK(I2702), .RSTB(I560792), .Q(I561066) );
and I_32844 (I561083,I561066,I653314);
DFFARX1 I_32845  ( .D(I561083), .CLK(I2702), .RSTB(I560792), .Q(I561100) );
not I_32846 (I560763,I561100);
nand I_32847 (I561131,I561083,I561021);
and I_32848 (I561148,I560843,I561131);
DFFARX1 I_32849  ( .D(I561148), .CLK(I2702), .RSTB(I560792), .Q(I560754) );
DFFARX1 I_32850  ( .D(I653302), .CLK(I2702), .RSTB(I560792), .Q(I561179) );
nand I_32851 (I561196,I561179,I560843);
and I_32852 (I561213,I561021,I561196);
DFFARX1 I_32853  ( .D(I561213), .CLK(I2702), .RSTB(I560792), .Q(I560784) );
not I_32854 (I561244,I561179);
nor I_32855 (I561261,I560860,I561244);
and I_32856 (I561278,I561179,I561261);
or I_32857 (I561295,I561083,I561278);
DFFARX1 I_32858  ( .D(I561295), .CLK(I2702), .RSTB(I560792), .Q(I560769) );
nand I_32859 (I560766,I561179,I560925);
DFFARX1 I_32860  ( .D(I561179), .CLK(I2702), .RSTB(I560792), .Q(I560757) );
not I_32861 (I561387,I2709);
nand I_32862 (I561404,I430343,I430331);
and I_32863 (I561421,I561404,I430337);
DFFARX1 I_32864  ( .D(I561421), .CLK(I2702), .RSTB(I561387), .Q(I561438) );
nor I_32865 (I561455,I430328,I430331);
nor I_32866 (I561472,I561455,I561438);
not I_32867 (I561370,I561455);
DFFARX1 I_32868  ( .D(I430313), .CLK(I2702), .RSTB(I561387), .Q(I561503) );
not I_32869 (I561520,I561503);
nor I_32870 (I561537,I561455,I561520);
nand I_32871 (I561373,I561503,I561472);
DFFARX1 I_32872  ( .D(I561503), .CLK(I2702), .RSTB(I561387), .Q(I561355) );
nand I_32873 (I561582,I430322,I430340);
and I_32874 (I561599,I561582,I430334);
DFFARX1 I_32875  ( .D(I561599), .CLK(I2702), .RSTB(I561387), .Q(I561616) );
nor I_32876 (I561376,I561616,I561438);
nand I_32877 (I561367,I561616,I561537);
DFFARX1 I_32878  ( .D(I430325), .CLK(I2702), .RSTB(I561387), .Q(I561661) );
and I_32879 (I561678,I561661,I430319);
DFFARX1 I_32880  ( .D(I561678), .CLK(I2702), .RSTB(I561387), .Q(I561695) );
not I_32881 (I561358,I561695);
nand I_32882 (I561726,I561678,I561616);
and I_32883 (I561743,I561438,I561726);
DFFARX1 I_32884  ( .D(I561743), .CLK(I2702), .RSTB(I561387), .Q(I561349) );
DFFARX1 I_32885  ( .D(I430316), .CLK(I2702), .RSTB(I561387), .Q(I561774) );
nand I_32886 (I561791,I561774,I561438);
and I_32887 (I561808,I561616,I561791);
DFFARX1 I_32888  ( .D(I561808), .CLK(I2702), .RSTB(I561387), .Q(I561379) );
not I_32889 (I561839,I561774);
nor I_32890 (I561856,I561455,I561839);
and I_32891 (I561873,I561774,I561856);
or I_32892 (I561890,I561678,I561873);
DFFARX1 I_32893  ( .D(I561890), .CLK(I2702), .RSTB(I561387), .Q(I561364) );
nand I_32894 (I561361,I561774,I561520);
DFFARX1 I_32895  ( .D(I561774), .CLK(I2702), .RSTB(I561387), .Q(I561352) );
not I_32896 (I561982,I2709);
nand I_32897 (I561999,I310617,I310623);
and I_32898 (I562016,I561999,I310605);
DFFARX1 I_32899  ( .D(I562016), .CLK(I2702), .RSTB(I561982), .Q(I562033) );
nor I_32900 (I562050,I310599,I310623);
nor I_32901 (I562067,I562050,I562033);
not I_32902 (I561965,I562050);
DFFARX1 I_32903  ( .D(I310629), .CLK(I2702), .RSTB(I561982), .Q(I562098) );
not I_32904 (I562115,I562098);
nor I_32905 (I562132,I562050,I562115);
nand I_32906 (I561968,I562098,I562067);
DFFARX1 I_32907  ( .D(I562098), .CLK(I2702), .RSTB(I561982), .Q(I561950) );
nand I_32908 (I562177,I310620,I310611);
and I_32909 (I562194,I562177,I310614);
DFFARX1 I_32910  ( .D(I562194), .CLK(I2702), .RSTB(I561982), .Q(I562211) );
nor I_32911 (I561971,I562211,I562033);
nand I_32912 (I561962,I562211,I562132);
DFFARX1 I_32913  ( .D(I310626), .CLK(I2702), .RSTB(I561982), .Q(I562256) );
and I_32914 (I562273,I562256,I310602);
DFFARX1 I_32915  ( .D(I562273), .CLK(I2702), .RSTB(I561982), .Q(I562290) );
not I_32916 (I561953,I562290);
nand I_32917 (I562321,I562273,I562211);
and I_32918 (I562338,I562033,I562321);
DFFARX1 I_32919  ( .D(I562338), .CLK(I2702), .RSTB(I561982), .Q(I561944) );
DFFARX1 I_32920  ( .D(I310608), .CLK(I2702), .RSTB(I561982), .Q(I562369) );
nand I_32921 (I562386,I562369,I562033);
and I_32922 (I562403,I562211,I562386);
DFFARX1 I_32923  ( .D(I562403), .CLK(I2702), .RSTB(I561982), .Q(I561974) );
not I_32924 (I562434,I562369);
nor I_32925 (I562451,I562050,I562434);
and I_32926 (I562468,I562369,I562451);
or I_32927 (I562485,I562273,I562468);
DFFARX1 I_32928  ( .D(I562485), .CLK(I2702), .RSTB(I561982), .Q(I561959) );
nand I_32929 (I561956,I562369,I562115);
DFFARX1 I_32930  ( .D(I562369), .CLK(I2702), .RSTB(I561982), .Q(I561947) );
not I_32931 (I562577,I2709);
nand I_32932 (I562594,I132448,I132460);
and I_32933 (I562611,I562594,I132469);
DFFARX1 I_32934  ( .D(I562611), .CLK(I2702), .RSTB(I562577), .Q(I562628) );
nor I_32935 (I562645,I132463,I132460);
nor I_32936 (I562662,I562645,I562628);
not I_32937 (I562560,I562645);
DFFARX1 I_32938  ( .D(I132457), .CLK(I2702), .RSTB(I562577), .Q(I562693) );
not I_32939 (I562710,I562693);
nor I_32940 (I562727,I562645,I562710);
nand I_32941 (I562563,I562693,I562662);
DFFARX1 I_32942  ( .D(I562693), .CLK(I2702), .RSTB(I562577), .Q(I562545) );
nand I_32943 (I562772,I132454,I132451);
and I_32944 (I562789,I562772,I132442);
DFFARX1 I_32945  ( .D(I562789), .CLK(I2702), .RSTB(I562577), .Q(I562806) );
nor I_32946 (I562566,I562806,I562628);
nand I_32947 (I562557,I562806,I562727);
DFFARX1 I_32948  ( .D(I132466), .CLK(I2702), .RSTB(I562577), .Q(I562851) );
and I_32949 (I562868,I562851,I132445);
DFFARX1 I_32950  ( .D(I562868), .CLK(I2702), .RSTB(I562577), .Q(I562885) );
not I_32951 (I562548,I562885);
nand I_32952 (I562916,I562868,I562806);
and I_32953 (I562933,I562628,I562916);
DFFARX1 I_32954  ( .D(I562933), .CLK(I2702), .RSTB(I562577), .Q(I562539) );
DFFARX1 I_32955  ( .D(I132439), .CLK(I2702), .RSTB(I562577), .Q(I562964) );
nand I_32956 (I562981,I562964,I562628);
and I_32957 (I562998,I562806,I562981);
DFFARX1 I_32958  ( .D(I562998), .CLK(I2702), .RSTB(I562577), .Q(I562569) );
not I_32959 (I563029,I562964);
nor I_32960 (I563046,I562645,I563029);
and I_32961 (I563063,I562964,I563046);
or I_32962 (I563080,I562868,I563063);
DFFARX1 I_32963  ( .D(I563080), .CLK(I2702), .RSTB(I562577), .Q(I562554) );
nand I_32964 (I562551,I562964,I562710);
DFFARX1 I_32965  ( .D(I562964), .CLK(I2702), .RSTB(I562577), .Q(I562542) );
not I_32966 (I563172,I2709);
nand I_32967 (I563189,I368689,I368701);
and I_32968 (I563206,I563189,I368683);
DFFARX1 I_32969  ( .D(I563206), .CLK(I2702), .RSTB(I563172), .Q(I563223) );
nor I_32970 (I563240,I368695,I368701);
nor I_32971 (I563257,I563240,I563223);
not I_32972 (I563155,I563240);
DFFARX1 I_32973  ( .D(I368680), .CLK(I2702), .RSTB(I563172), .Q(I563288) );
not I_32974 (I563305,I563288);
nor I_32975 (I563322,I563240,I563305);
nand I_32976 (I563158,I563288,I563257);
DFFARX1 I_32977  ( .D(I563288), .CLK(I2702), .RSTB(I563172), .Q(I563140) );
nand I_32978 (I563367,I368671,I368686);
and I_32979 (I563384,I563367,I368677);
DFFARX1 I_32980  ( .D(I563384), .CLK(I2702), .RSTB(I563172), .Q(I563401) );
nor I_32981 (I563161,I563401,I563223);
nand I_32982 (I563152,I563401,I563322);
DFFARX1 I_32983  ( .D(I368698), .CLK(I2702), .RSTB(I563172), .Q(I563446) );
and I_32984 (I563463,I563446,I368692);
DFFARX1 I_32985  ( .D(I563463), .CLK(I2702), .RSTB(I563172), .Q(I563480) );
not I_32986 (I563143,I563480);
nand I_32987 (I563511,I563463,I563401);
and I_32988 (I563528,I563223,I563511);
DFFARX1 I_32989  ( .D(I563528), .CLK(I2702), .RSTB(I563172), .Q(I563134) );
DFFARX1 I_32990  ( .D(I368674), .CLK(I2702), .RSTB(I563172), .Q(I563559) );
nand I_32991 (I563576,I563559,I563223);
and I_32992 (I563593,I563401,I563576);
DFFARX1 I_32993  ( .D(I563593), .CLK(I2702), .RSTB(I563172), .Q(I563164) );
not I_32994 (I563624,I563559);
nor I_32995 (I563641,I563240,I563624);
and I_32996 (I563658,I563559,I563641);
or I_32997 (I563675,I563463,I563658);
DFFARX1 I_32998  ( .D(I563675), .CLK(I2702), .RSTB(I563172), .Q(I563149) );
nand I_32999 (I563146,I563559,I563305);
DFFARX1 I_33000  ( .D(I563559), .CLK(I2702), .RSTB(I563172), .Q(I563137) );
not I_33001 (I563767,I2709);
nand I_33002 (I563784,I78184,I78196);
and I_33003 (I563801,I563784,I78205);
DFFARX1 I_33004  ( .D(I563801), .CLK(I2702), .RSTB(I563767), .Q(I563818) );
nor I_33005 (I563835,I78199,I78196);
nor I_33006 (I563852,I563835,I563818);
not I_33007 (I563750,I563835);
DFFARX1 I_33008  ( .D(I78193), .CLK(I2702), .RSTB(I563767), .Q(I563883) );
not I_33009 (I563900,I563883);
nor I_33010 (I563917,I563835,I563900);
nand I_33011 (I563753,I563883,I563852);
DFFARX1 I_33012  ( .D(I563883), .CLK(I2702), .RSTB(I563767), .Q(I563735) );
nand I_33013 (I563962,I78190,I78187);
and I_33014 (I563979,I563962,I78178);
DFFARX1 I_33015  ( .D(I563979), .CLK(I2702), .RSTB(I563767), .Q(I563996) );
nor I_33016 (I563756,I563996,I563818);
nand I_33017 (I563747,I563996,I563917);
DFFARX1 I_33018  ( .D(I78202), .CLK(I2702), .RSTB(I563767), .Q(I564041) );
and I_33019 (I564058,I564041,I78181);
DFFARX1 I_33020  ( .D(I564058), .CLK(I2702), .RSTB(I563767), .Q(I564075) );
not I_33021 (I563738,I564075);
nand I_33022 (I564106,I564058,I563996);
and I_33023 (I564123,I563818,I564106);
DFFARX1 I_33024  ( .D(I564123), .CLK(I2702), .RSTB(I563767), .Q(I563729) );
DFFARX1 I_33025  ( .D(I78175), .CLK(I2702), .RSTB(I563767), .Q(I564154) );
nand I_33026 (I564171,I564154,I563818);
and I_33027 (I564188,I563996,I564171);
DFFARX1 I_33028  ( .D(I564188), .CLK(I2702), .RSTB(I563767), .Q(I563759) );
not I_33029 (I564219,I564154);
nor I_33030 (I564236,I563835,I564219);
and I_33031 (I564253,I564154,I564236);
or I_33032 (I564270,I564058,I564253);
DFFARX1 I_33033  ( .D(I564270), .CLK(I2702), .RSTB(I563767), .Q(I563744) );
nand I_33034 (I563741,I564154,I563900);
DFFARX1 I_33035  ( .D(I564154), .CLK(I2702), .RSTB(I563767), .Q(I563732) );
not I_33036 (I564362,I2709);
nand I_33037 (I564379,I164094,I164106);
and I_33038 (I564396,I564379,I164085);
DFFARX1 I_33039  ( .D(I564396), .CLK(I2702), .RSTB(I564362), .Q(I564413) );
nor I_33040 (I564430,I164076,I164106);
nor I_33041 (I564447,I564430,I564413);
not I_33042 (I564345,I564430);
DFFARX1 I_33043  ( .D(I164088), .CLK(I2702), .RSTB(I564362), .Q(I564478) );
not I_33044 (I564495,I564478);
nor I_33045 (I564512,I564430,I564495);
nand I_33046 (I564348,I564478,I564447);
DFFARX1 I_33047  ( .D(I564478), .CLK(I2702), .RSTB(I564362), .Q(I564330) );
nand I_33048 (I564557,I164103,I164091);
and I_33049 (I564574,I564557,I164079);
DFFARX1 I_33050  ( .D(I564574), .CLK(I2702), .RSTB(I564362), .Q(I564591) );
nor I_33051 (I564351,I564591,I564413);
nand I_33052 (I564342,I564591,I564512);
DFFARX1 I_33053  ( .D(I164097), .CLK(I2702), .RSTB(I564362), .Q(I564636) );
and I_33054 (I564653,I564636,I164082);
DFFARX1 I_33055  ( .D(I564653), .CLK(I2702), .RSTB(I564362), .Q(I564670) );
not I_33056 (I564333,I564670);
nand I_33057 (I564701,I564653,I564591);
and I_33058 (I564718,I564413,I564701);
DFFARX1 I_33059  ( .D(I564718), .CLK(I2702), .RSTB(I564362), .Q(I564324) );
DFFARX1 I_33060  ( .D(I164100), .CLK(I2702), .RSTB(I564362), .Q(I564749) );
nand I_33061 (I564766,I564749,I564413);
and I_33062 (I564783,I564591,I564766);
DFFARX1 I_33063  ( .D(I564783), .CLK(I2702), .RSTB(I564362), .Q(I564354) );
not I_33064 (I564814,I564749);
nor I_33065 (I564831,I564430,I564814);
and I_33066 (I564848,I564749,I564831);
or I_33067 (I564865,I564653,I564848);
DFFARX1 I_33068  ( .D(I564865), .CLK(I2702), .RSTB(I564362), .Q(I564339) );
nand I_33069 (I564336,I564749,I564495);
DFFARX1 I_33070  ( .D(I564749), .CLK(I2702), .RSTB(I564362), .Q(I564327) );
not I_33071 (I564957,I2709);
nand I_33072 (I564974,I91104,I91116);
and I_33073 (I564991,I564974,I91125);
DFFARX1 I_33074  ( .D(I564991), .CLK(I2702), .RSTB(I564957), .Q(I565008) );
nor I_33075 (I565025,I91119,I91116);
nor I_33076 (I565042,I565025,I565008);
not I_33077 (I564940,I565025);
DFFARX1 I_33078  ( .D(I91113), .CLK(I2702), .RSTB(I564957), .Q(I565073) );
not I_33079 (I565090,I565073);
nor I_33080 (I565107,I565025,I565090);
nand I_33081 (I564943,I565073,I565042);
DFFARX1 I_33082  ( .D(I565073), .CLK(I2702), .RSTB(I564957), .Q(I564925) );
nand I_33083 (I565152,I91110,I91107);
and I_33084 (I565169,I565152,I91098);
DFFARX1 I_33085  ( .D(I565169), .CLK(I2702), .RSTB(I564957), .Q(I565186) );
nor I_33086 (I564946,I565186,I565008);
nand I_33087 (I564937,I565186,I565107);
DFFARX1 I_33088  ( .D(I91122), .CLK(I2702), .RSTB(I564957), .Q(I565231) );
and I_33089 (I565248,I565231,I91101);
DFFARX1 I_33090  ( .D(I565248), .CLK(I2702), .RSTB(I564957), .Q(I565265) );
not I_33091 (I564928,I565265);
nand I_33092 (I565296,I565248,I565186);
and I_33093 (I565313,I565008,I565296);
DFFARX1 I_33094  ( .D(I565313), .CLK(I2702), .RSTB(I564957), .Q(I564919) );
DFFARX1 I_33095  ( .D(I91095), .CLK(I2702), .RSTB(I564957), .Q(I565344) );
nand I_33096 (I565361,I565344,I565008);
and I_33097 (I565378,I565186,I565361);
DFFARX1 I_33098  ( .D(I565378), .CLK(I2702), .RSTB(I564957), .Q(I564949) );
not I_33099 (I565409,I565344);
nor I_33100 (I565426,I565025,I565409);
and I_33101 (I565443,I565344,I565426);
or I_33102 (I565460,I565248,I565443);
DFFARX1 I_33103  ( .D(I565460), .CLK(I2702), .RSTB(I564957), .Q(I564934) );
nand I_33104 (I564931,I565344,I565090);
DFFARX1 I_33105  ( .D(I565344), .CLK(I2702), .RSTB(I564957), .Q(I564922) );
not I_33106 (I565552,I2709);
nand I_33107 (I565569,I138262,I138274);
and I_33108 (I565586,I565569,I138283);
DFFARX1 I_33109  ( .D(I565586), .CLK(I2702), .RSTB(I565552), .Q(I565603) );
nor I_33110 (I565620,I138277,I138274);
nor I_33111 (I565637,I565620,I565603);
not I_33112 (I565535,I565620);
DFFARX1 I_33113  ( .D(I138271), .CLK(I2702), .RSTB(I565552), .Q(I565668) );
not I_33114 (I565685,I565668);
nor I_33115 (I565702,I565620,I565685);
nand I_33116 (I565538,I565668,I565637);
DFFARX1 I_33117  ( .D(I565668), .CLK(I2702), .RSTB(I565552), .Q(I565520) );
nand I_33118 (I565747,I138268,I138265);
and I_33119 (I565764,I565747,I138256);
DFFARX1 I_33120  ( .D(I565764), .CLK(I2702), .RSTB(I565552), .Q(I565781) );
nor I_33121 (I565541,I565781,I565603);
nand I_33122 (I565532,I565781,I565702);
DFFARX1 I_33123  ( .D(I138280), .CLK(I2702), .RSTB(I565552), .Q(I565826) );
and I_33124 (I565843,I565826,I138259);
DFFARX1 I_33125  ( .D(I565843), .CLK(I2702), .RSTB(I565552), .Q(I565860) );
not I_33126 (I565523,I565860);
nand I_33127 (I565891,I565843,I565781);
and I_33128 (I565908,I565603,I565891);
DFFARX1 I_33129  ( .D(I565908), .CLK(I2702), .RSTB(I565552), .Q(I565514) );
DFFARX1 I_33130  ( .D(I138253), .CLK(I2702), .RSTB(I565552), .Q(I565939) );
nand I_33131 (I565956,I565939,I565603);
and I_33132 (I565973,I565781,I565956);
DFFARX1 I_33133  ( .D(I565973), .CLK(I2702), .RSTB(I565552), .Q(I565544) );
not I_33134 (I566004,I565939);
nor I_33135 (I566021,I565620,I566004);
and I_33136 (I566038,I565939,I566021);
or I_33137 (I566055,I565843,I566038);
DFFARX1 I_33138  ( .D(I566055), .CLK(I2702), .RSTB(I565552), .Q(I565529) );
nand I_33139 (I565526,I565939,I565685);
DFFARX1 I_33140  ( .D(I565939), .CLK(I2702), .RSTB(I565552), .Q(I565517) );
not I_33141 (I566147,I2709);
nand I_33142 (I566164,I652691,I652682);
and I_33143 (I566181,I566164,I652700);
DFFARX1 I_33144  ( .D(I566181), .CLK(I2702), .RSTB(I566147), .Q(I566198) );
nor I_33145 (I566215,I652697,I652682);
nor I_33146 (I566232,I566215,I566198);
not I_33147 (I566130,I566215);
DFFARX1 I_33148  ( .D(I652679), .CLK(I2702), .RSTB(I566147), .Q(I566263) );
not I_33149 (I566280,I566263);
nor I_33150 (I566297,I566215,I566280);
nand I_33151 (I566133,I566263,I566232);
DFFARX1 I_33152  ( .D(I566263), .CLK(I2702), .RSTB(I566147), .Q(I566115) );
nand I_33153 (I566342,I652688,I652703);
and I_33154 (I566359,I566342,I652694);
DFFARX1 I_33155  ( .D(I566359), .CLK(I2702), .RSTB(I566147), .Q(I566376) );
nor I_33156 (I566136,I566376,I566198);
nand I_33157 (I566127,I566376,I566297);
DFFARX1 I_33158  ( .D(I652676), .CLK(I2702), .RSTB(I566147), .Q(I566421) );
and I_33159 (I566438,I566421,I652685);
DFFARX1 I_33160  ( .D(I566438), .CLK(I2702), .RSTB(I566147), .Q(I566455) );
not I_33161 (I566118,I566455);
nand I_33162 (I566486,I566438,I566376);
and I_33163 (I566503,I566198,I566486);
DFFARX1 I_33164  ( .D(I566503), .CLK(I2702), .RSTB(I566147), .Q(I566109) );
DFFARX1 I_33165  ( .D(I652673), .CLK(I2702), .RSTB(I566147), .Q(I566534) );
nand I_33166 (I566551,I566534,I566198);
and I_33167 (I566568,I566376,I566551);
DFFARX1 I_33168  ( .D(I566568), .CLK(I2702), .RSTB(I566147), .Q(I566139) );
not I_33169 (I566599,I566534);
nor I_33170 (I566616,I566215,I566599);
and I_33171 (I566633,I566534,I566616);
or I_33172 (I566650,I566438,I566633);
DFFARX1 I_33173  ( .D(I566650), .CLK(I2702), .RSTB(I566147), .Q(I566124) );
nand I_33174 (I566121,I566534,I566280);
DFFARX1 I_33175  ( .D(I566534), .CLK(I2702), .RSTB(I566147), .Q(I566112) );
not I_33176 (I566742,I2709);
nand I_33177 (I566759,I601229,I601220);
and I_33178 (I566776,I566759,I601238);
DFFARX1 I_33179  ( .D(I566776), .CLK(I2702), .RSTB(I566742), .Q(I566793) );
nor I_33180 (I566810,I601217,I601220);
nor I_33181 (I566827,I566810,I566793);
not I_33182 (I566725,I566810);
DFFARX1 I_33183  ( .D(I601226), .CLK(I2702), .RSTB(I566742), .Q(I566858) );
not I_33184 (I566875,I566858);
nor I_33185 (I566892,I566810,I566875);
nand I_33186 (I566728,I566858,I566827);
DFFARX1 I_33187  ( .D(I566858), .CLK(I2702), .RSTB(I566742), .Q(I566710) );
nand I_33188 (I566937,I601241,I601223);
and I_33189 (I566954,I566937,I601244);
DFFARX1 I_33190  ( .D(I566954), .CLK(I2702), .RSTB(I566742), .Q(I566971) );
nor I_33191 (I566731,I566971,I566793);
nand I_33192 (I566722,I566971,I566892);
DFFARX1 I_33193  ( .D(I601232), .CLK(I2702), .RSTB(I566742), .Q(I567016) );
and I_33194 (I567033,I567016,I601214);
DFFARX1 I_33195  ( .D(I567033), .CLK(I2702), .RSTB(I566742), .Q(I567050) );
not I_33196 (I566713,I567050);
nand I_33197 (I567081,I567033,I566971);
and I_33198 (I567098,I566793,I567081);
DFFARX1 I_33199  ( .D(I567098), .CLK(I2702), .RSTB(I566742), .Q(I566704) );
DFFARX1 I_33200  ( .D(I601235), .CLK(I2702), .RSTB(I566742), .Q(I567129) );
nand I_33201 (I567146,I567129,I566793);
and I_33202 (I567163,I566971,I567146);
DFFARX1 I_33203  ( .D(I567163), .CLK(I2702), .RSTB(I566742), .Q(I566734) );
not I_33204 (I567194,I567129);
nor I_33205 (I567211,I566810,I567194);
and I_33206 (I567228,I567129,I567211);
or I_33207 (I567245,I567033,I567228);
DFFARX1 I_33208  ( .D(I567245), .CLK(I2702), .RSTB(I566742), .Q(I566719) );
nand I_33209 (I566716,I567129,I566875);
DFFARX1 I_33210  ( .D(I567129), .CLK(I2702), .RSTB(I566742), .Q(I566707) );
not I_33211 (I567337,I2709);
nand I_33212 (I567354,I291390,I291396);
and I_33213 (I567371,I567354,I291378);
DFFARX1 I_33214  ( .D(I567371), .CLK(I2702), .RSTB(I567337), .Q(I567388) );
nor I_33215 (I567405,I291372,I291396);
nor I_33216 (I567422,I567405,I567388);
not I_33217 (I567320,I567405);
DFFARX1 I_33218  ( .D(I291402), .CLK(I2702), .RSTB(I567337), .Q(I567453) );
not I_33219 (I567470,I567453);
nor I_33220 (I567487,I567405,I567470);
nand I_33221 (I567323,I567453,I567422);
DFFARX1 I_33222  ( .D(I567453), .CLK(I2702), .RSTB(I567337), .Q(I567305) );
nand I_33223 (I567532,I291393,I291384);
and I_33224 (I567549,I567532,I291387);
DFFARX1 I_33225  ( .D(I567549), .CLK(I2702), .RSTB(I567337), .Q(I567566) );
nor I_33226 (I567326,I567566,I567388);
nand I_33227 (I567317,I567566,I567487);
DFFARX1 I_33228  ( .D(I291399), .CLK(I2702), .RSTB(I567337), .Q(I567611) );
and I_33229 (I567628,I567611,I291375);
DFFARX1 I_33230  ( .D(I567628), .CLK(I2702), .RSTB(I567337), .Q(I567645) );
not I_33231 (I567308,I567645);
nand I_33232 (I567676,I567628,I567566);
and I_33233 (I567693,I567388,I567676);
DFFARX1 I_33234  ( .D(I567693), .CLK(I2702), .RSTB(I567337), .Q(I567299) );
DFFARX1 I_33235  ( .D(I291381), .CLK(I2702), .RSTB(I567337), .Q(I567724) );
nand I_33236 (I567741,I567724,I567388);
and I_33237 (I567758,I567566,I567741);
DFFARX1 I_33238  ( .D(I567758), .CLK(I2702), .RSTB(I567337), .Q(I567329) );
not I_33239 (I567789,I567724);
nor I_33240 (I567806,I567405,I567789);
and I_33241 (I567823,I567724,I567806);
or I_33242 (I567840,I567628,I567823);
DFFARX1 I_33243  ( .D(I567840), .CLK(I2702), .RSTB(I567337), .Q(I567314) );
nand I_33244 (I567311,I567724,I567470);
DFFARX1 I_33245  ( .D(I567724), .CLK(I2702), .RSTB(I567337), .Q(I567302) );
not I_33246 (I567932,I2709);
nand I_33247 (I567949,I656465,I656456);
and I_33248 (I567966,I567949,I656474);
DFFARX1 I_33249  ( .D(I567966), .CLK(I2702), .RSTB(I567932), .Q(I567983) );
nor I_33250 (I568000,I656471,I656456);
nor I_33251 (I568017,I568000,I567983);
not I_33252 (I567915,I568000);
DFFARX1 I_33253  ( .D(I656453), .CLK(I2702), .RSTB(I567932), .Q(I568048) );
not I_33254 (I568065,I568048);
nor I_33255 (I568082,I568000,I568065);
nand I_33256 (I567918,I568048,I568017);
DFFARX1 I_33257  ( .D(I568048), .CLK(I2702), .RSTB(I567932), .Q(I567900) );
nand I_33258 (I568127,I656462,I656477);
and I_33259 (I568144,I568127,I656468);
DFFARX1 I_33260  ( .D(I568144), .CLK(I2702), .RSTB(I567932), .Q(I568161) );
nor I_33261 (I567921,I568161,I567983);
nand I_33262 (I567912,I568161,I568082);
DFFARX1 I_33263  ( .D(I656450), .CLK(I2702), .RSTB(I567932), .Q(I568206) );
and I_33264 (I568223,I568206,I656459);
DFFARX1 I_33265  ( .D(I568223), .CLK(I2702), .RSTB(I567932), .Q(I568240) );
not I_33266 (I567903,I568240);
nand I_33267 (I568271,I568223,I568161);
and I_33268 (I568288,I567983,I568271);
DFFARX1 I_33269  ( .D(I568288), .CLK(I2702), .RSTB(I567932), .Q(I567894) );
DFFARX1 I_33270  ( .D(I656447), .CLK(I2702), .RSTB(I567932), .Q(I568319) );
nand I_33271 (I568336,I568319,I567983);
and I_33272 (I568353,I568161,I568336);
DFFARX1 I_33273  ( .D(I568353), .CLK(I2702), .RSTB(I567932), .Q(I567924) );
not I_33274 (I568384,I568319);
nor I_33275 (I568401,I568000,I568384);
and I_33276 (I568418,I568319,I568401);
or I_33277 (I568435,I568223,I568418);
DFFARX1 I_33278  ( .D(I568435), .CLK(I2702), .RSTB(I567932), .Q(I567909) );
nand I_33279 (I567906,I568319,I568065);
DFFARX1 I_33280  ( .D(I568319), .CLK(I2702), .RSTB(I567932), .Q(I567897) );
not I_33281 (I568527,I2709);
nand I_33282 (I568544,I607179,I607170);
and I_33283 (I568561,I568544,I607188);
DFFARX1 I_33284  ( .D(I568561), .CLK(I2702), .RSTB(I568527), .Q(I568578) );
nor I_33285 (I568595,I607167,I607170);
nor I_33286 (I568612,I568595,I568578);
not I_33287 (I568510,I568595);
DFFARX1 I_33288  ( .D(I607176), .CLK(I2702), .RSTB(I568527), .Q(I568643) );
not I_33289 (I568660,I568643);
nor I_33290 (I568677,I568595,I568660);
nand I_33291 (I568513,I568643,I568612);
DFFARX1 I_33292  ( .D(I568643), .CLK(I2702), .RSTB(I568527), .Q(I568495) );
nand I_33293 (I568722,I607191,I607173);
and I_33294 (I568739,I568722,I607194);
DFFARX1 I_33295  ( .D(I568739), .CLK(I2702), .RSTB(I568527), .Q(I568756) );
nor I_33296 (I568516,I568756,I568578);
nand I_33297 (I568507,I568756,I568677);
DFFARX1 I_33298  ( .D(I607182), .CLK(I2702), .RSTB(I568527), .Q(I568801) );
and I_33299 (I568818,I568801,I607164);
DFFARX1 I_33300  ( .D(I568818), .CLK(I2702), .RSTB(I568527), .Q(I568835) );
not I_33301 (I568498,I568835);
nand I_33302 (I568866,I568818,I568756);
and I_33303 (I568883,I568578,I568866);
DFFARX1 I_33304  ( .D(I568883), .CLK(I2702), .RSTB(I568527), .Q(I568489) );
DFFARX1 I_33305  ( .D(I607185), .CLK(I2702), .RSTB(I568527), .Q(I568914) );
nand I_33306 (I568931,I568914,I568578);
and I_33307 (I568948,I568756,I568931);
DFFARX1 I_33308  ( .D(I568948), .CLK(I2702), .RSTB(I568527), .Q(I568519) );
not I_33309 (I568979,I568914);
nor I_33310 (I568996,I568595,I568979);
and I_33311 (I569013,I568914,I568996);
or I_33312 (I569030,I568818,I569013);
DFFARX1 I_33313  ( .D(I569030), .CLK(I2702), .RSTB(I568527), .Q(I568504) );
nand I_33314 (I568501,I568914,I568660);
DFFARX1 I_33315  ( .D(I568914), .CLK(I2702), .RSTB(I568527), .Q(I568492) );
not I_33316 (I569122,I2709);
nand I_33317 (I569139,I12252,I12258);
and I_33318 (I569156,I569139,I12255);
DFFARX1 I_33319  ( .D(I569156), .CLK(I2702), .RSTB(I569122), .Q(I569173) );
nor I_33320 (I569190,I12279,I12258);
nor I_33321 (I569207,I569190,I569173);
not I_33322 (I569105,I569190);
DFFARX1 I_33323  ( .D(I12270), .CLK(I2702), .RSTB(I569122), .Q(I569238) );
not I_33324 (I569255,I569238);
nor I_33325 (I569272,I569190,I569255);
nand I_33326 (I569108,I569238,I569207);
DFFARX1 I_33327  ( .D(I569238), .CLK(I2702), .RSTB(I569122), .Q(I569090) );
nand I_33328 (I569317,I12273,I12276);
and I_33329 (I569334,I569317,I12249);
DFFARX1 I_33330  ( .D(I569334), .CLK(I2702), .RSTB(I569122), .Q(I569351) );
nor I_33331 (I569111,I569351,I569173);
nand I_33332 (I569102,I569351,I569272);
DFFARX1 I_33333  ( .D(I12267), .CLK(I2702), .RSTB(I569122), .Q(I569396) );
and I_33334 (I569413,I569396,I12261);
DFFARX1 I_33335  ( .D(I569413), .CLK(I2702), .RSTB(I569122), .Q(I569430) );
not I_33336 (I569093,I569430);
nand I_33337 (I569461,I569413,I569351);
and I_33338 (I569478,I569173,I569461);
DFFARX1 I_33339  ( .D(I569478), .CLK(I2702), .RSTB(I569122), .Q(I569084) );
DFFARX1 I_33340  ( .D(I12264), .CLK(I2702), .RSTB(I569122), .Q(I569509) );
nand I_33341 (I569526,I569509,I569173);
and I_33342 (I569543,I569351,I569526);
DFFARX1 I_33343  ( .D(I569543), .CLK(I2702), .RSTB(I569122), .Q(I569114) );
not I_33344 (I569574,I569509);
nor I_33345 (I569591,I569190,I569574);
and I_33346 (I569608,I569509,I569591);
or I_33347 (I569625,I569413,I569608);
DFFARX1 I_33348  ( .D(I569625), .CLK(I2702), .RSTB(I569122), .Q(I569099) );
nand I_33349 (I569096,I569509,I569255);
DFFARX1 I_33350  ( .D(I569509), .CLK(I2702), .RSTB(I569122), .Q(I569087) );
not I_33351 (I569717,I2709);
nand I_33352 (I569734,I39180,I39186);
and I_33353 (I569751,I569734,I39183);
DFFARX1 I_33354  ( .D(I569751), .CLK(I2702), .RSTB(I569717), .Q(I569768) );
nor I_33355 (I569785,I39207,I39186);
nor I_33356 (I569802,I569785,I569768);
not I_33357 (I569700,I569785);
DFFARX1 I_33358  ( .D(I39198), .CLK(I2702), .RSTB(I569717), .Q(I569833) );
not I_33359 (I569850,I569833);
nor I_33360 (I569867,I569785,I569850);
nand I_33361 (I569703,I569833,I569802);
DFFARX1 I_33362  ( .D(I569833), .CLK(I2702), .RSTB(I569717), .Q(I569685) );
nand I_33363 (I569912,I39201,I39204);
and I_33364 (I569929,I569912,I39177);
DFFARX1 I_33365  ( .D(I569929), .CLK(I2702), .RSTB(I569717), .Q(I569946) );
nor I_33366 (I569706,I569946,I569768);
nand I_33367 (I569697,I569946,I569867);
DFFARX1 I_33368  ( .D(I39195), .CLK(I2702), .RSTB(I569717), .Q(I569991) );
and I_33369 (I570008,I569991,I39189);
DFFARX1 I_33370  ( .D(I570008), .CLK(I2702), .RSTB(I569717), .Q(I570025) );
not I_33371 (I569688,I570025);
nand I_33372 (I570056,I570008,I569946);
and I_33373 (I570073,I569768,I570056);
DFFARX1 I_33374  ( .D(I570073), .CLK(I2702), .RSTB(I569717), .Q(I569679) );
DFFARX1 I_33375  ( .D(I39192), .CLK(I2702), .RSTB(I569717), .Q(I570104) );
nand I_33376 (I570121,I570104,I569768);
and I_33377 (I570138,I569946,I570121);
DFFARX1 I_33378  ( .D(I570138), .CLK(I2702), .RSTB(I569717), .Q(I569709) );
not I_33379 (I570169,I570104);
nor I_33380 (I570186,I569785,I570169);
and I_33381 (I570203,I570104,I570186);
or I_33382 (I570220,I570008,I570203);
DFFARX1 I_33383  ( .D(I570220), .CLK(I2702), .RSTB(I569717), .Q(I569694) );
nand I_33384 (I569691,I570104,I569850);
DFFARX1 I_33385  ( .D(I570104), .CLK(I2702), .RSTB(I569717), .Q(I569682) );
not I_33386 (I570312,I2709);
nand I_33387 (I570329,I366751,I366763);
and I_33388 (I570346,I570329,I366745);
DFFARX1 I_33389  ( .D(I570346), .CLK(I2702), .RSTB(I570312), .Q(I570363) );
nor I_33390 (I570380,I366757,I366763);
nor I_33391 (I570397,I570380,I570363);
not I_33392 (I570295,I570380);
DFFARX1 I_33393  ( .D(I366742), .CLK(I2702), .RSTB(I570312), .Q(I570428) );
not I_33394 (I570445,I570428);
nor I_33395 (I570462,I570380,I570445);
nand I_33396 (I570298,I570428,I570397);
DFFARX1 I_33397  ( .D(I570428), .CLK(I2702), .RSTB(I570312), .Q(I570280) );
nand I_33398 (I570507,I366733,I366748);
and I_33399 (I570524,I570507,I366739);
DFFARX1 I_33400  ( .D(I570524), .CLK(I2702), .RSTB(I570312), .Q(I570541) );
nor I_33401 (I570301,I570541,I570363);
nand I_33402 (I570292,I570541,I570462);
DFFARX1 I_33403  ( .D(I366760), .CLK(I2702), .RSTB(I570312), .Q(I570586) );
and I_33404 (I570603,I570586,I366754);
DFFARX1 I_33405  ( .D(I570603), .CLK(I2702), .RSTB(I570312), .Q(I570620) );
not I_33406 (I570283,I570620);
nand I_33407 (I570651,I570603,I570541);
and I_33408 (I570668,I570363,I570651);
DFFARX1 I_33409  ( .D(I570668), .CLK(I2702), .RSTB(I570312), .Q(I570274) );
DFFARX1 I_33410  ( .D(I366736), .CLK(I2702), .RSTB(I570312), .Q(I570699) );
nand I_33411 (I570716,I570699,I570363);
and I_33412 (I570733,I570541,I570716);
DFFARX1 I_33413  ( .D(I570733), .CLK(I2702), .RSTB(I570312), .Q(I570304) );
not I_33414 (I570764,I570699);
nor I_33415 (I570781,I570380,I570764);
and I_33416 (I570798,I570699,I570781);
or I_33417 (I570815,I570603,I570798);
DFFARX1 I_33418  ( .D(I570815), .CLK(I2702), .RSTB(I570312), .Q(I570289) );
nand I_33419 (I570286,I570699,I570445);
DFFARX1 I_33420  ( .D(I570699), .CLK(I2702), .RSTB(I570312), .Q(I570277) );
not I_33421 (I570907,I2709);
nand I_33422 (I570924,I715228,I715234);
and I_33423 (I570941,I570924,I715225);
DFFARX1 I_33424  ( .D(I570941), .CLK(I2702), .RSTB(I570907), .Q(I570958) );
nor I_33425 (I570975,I715237,I715234);
nor I_33426 (I570992,I570975,I570958);
not I_33427 (I570890,I570975);
DFFARX1 I_33428  ( .D(I715216), .CLK(I2702), .RSTB(I570907), .Q(I571023) );
not I_33429 (I571040,I571023);
nor I_33430 (I571057,I570975,I571040);
nand I_33431 (I570893,I571023,I570992);
DFFARX1 I_33432  ( .D(I571023), .CLK(I2702), .RSTB(I570907), .Q(I570875) );
nand I_33433 (I571102,I715240,I715222);
and I_33434 (I571119,I571102,I715231);
DFFARX1 I_33435  ( .D(I571119), .CLK(I2702), .RSTB(I570907), .Q(I571136) );
nor I_33436 (I570896,I571136,I570958);
nand I_33437 (I570887,I571136,I571057);
DFFARX1 I_33438  ( .D(I715246), .CLK(I2702), .RSTB(I570907), .Q(I571181) );
and I_33439 (I571198,I571181,I715219);
DFFARX1 I_33440  ( .D(I571198), .CLK(I2702), .RSTB(I570907), .Q(I571215) );
not I_33441 (I570878,I571215);
nand I_33442 (I571246,I571198,I571136);
and I_33443 (I571263,I570958,I571246);
DFFARX1 I_33444  ( .D(I571263), .CLK(I2702), .RSTB(I570907), .Q(I570869) );
DFFARX1 I_33445  ( .D(I715243), .CLK(I2702), .RSTB(I570907), .Q(I571294) );
nand I_33446 (I571311,I571294,I570958);
and I_33447 (I571328,I571136,I571311);
DFFARX1 I_33448  ( .D(I571328), .CLK(I2702), .RSTB(I570907), .Q(I570899) );
not I_33449 (I571359,I571294);
nor I_33450 (I571376,I570975,I571359);
and I_33451 (I571393,I571294,I571376);
or I_33452 (I571410,I571198,I571393);
DFFARX1 I_33453  ( .D(I571410), .CLK(I2702), .RSTB(I570907), .Q(I570884) );
nand I_33454 (I570881,I571294,I571040);
DFFARX1 I_33455  ( .D(I571294), .CLK(I2702), .RSTB(I570907), .Q(I570872) );
not I_33456 (I571502,I2709);
nand I_33457 (I571519,I466822,I466825);
and I_33458 (I571536,I571519,I466819);
DFFARX1 I_33459  ( .D(I571536), .CLK(I2702), .RSTB(I571502), .Q(I571553) );
nor I_33460 (I571570,I466816,I466825);
nor I_33461 (I571587,I571570,I571553);
not I_33462 (I571485,I571570);
DFFARX1 I_33463  ( .D(I466798), .CLK(I2702), .RSTB(I571502), .Q(I571618) );
not I_33464 (I571635,I571618);
nor I_33465 (I571652,I571570,I571635);
nand I_33466 (I571488,I571618,I571587);
DFFARX1 I_33467  ( .D(I571618), .CLK(I2702), .RSTB(I571502), .Q(I571470) );
nand I_33468 (I571697,I466807,I466804);
and I_33469 (I571714,I571697,I466813);
DFFARX1 I_33470  ( .D(I571714), .CLK(I2702), .RSTB(I571502), .Q(I571731) );
nor I_33471 (I571491,I571731,I571553);
nand I_33472 (I571482,I571731,I571652);
DFFARX1 I_33473  ( .D(I466795), .CLK(I2702), .RSTB(I571502), .Q(I571776) );
and I_33474 (I571793,I571776,I466810);
DFFARX1 I_33475  ( .D(I571793), .CLK(I2702), .RSTB(I571502), .Q(I571810) );
not I_33476 (I571473,I571810);
nand I_33477 (I571841,I571793,I571731);
and I_33478 (I571858,I571553,I571841);
DFFARX1 I_33479  ( .D(I571858), .CLK(I2702), .RSTB(I571502), .Q(I571464) );
DFFARX1 I_33480  ( .D(I466801), .CLK(I2702), .RSTB(I571502), .Q(I571889) );
nand I_33481 (I571906,I571889,I571553);
and I_33482 (I571923,I571731,I571906);
DFFARX1 I_33483  ( .D(I571923), .CLK(I2702), .RSTB(I571502), .Q(I571494) );
not I_33484 (I571954,I571889);
nor I_33485 (I571971,I571570,I571954);
and I_33486 (I571988,I571889,I571971);
or I_33487 (I572005,I571793,I571988);
DFFARX1 I_33488  ( .D(I572005), .CLK(I2702), .RSTB(I571502), .Q(I571479) );
nand I_33489 (I571476,I571889,I571635);
DFFARX1 I_33490  ( .D(I571889), .CLK(I2702), .RSTB(I571502), .Q(I571467) );
not I_33491 (I572097,I2709);
nand I_33492 (I572114,I697310,I697316);
and I_33493 (I572131,I572114,I697307);
DFFARX1 I_33494  ( .D(I572131), .CLK(I2702), .RSTB(I572097), .Q(I572148) );
nor I_33495 (I572165,I697319,I697316);
nor I_33496 (I572182,I572165,I572148);
not I_33497 (I572080,I572165);
DFFARX1 I_33498  ( .D(I697298), .CLK(I2702), .RSTB(I572097), .Q(I572213) );
not I_33499 (I572230,I572213);
nor I_33500 (I572247,I572165,I572230);
nand I_33501 (I572083,I572213,I572182);
DFFARX1 I_33502  ( .D(I572213), .CLK(I2702), .RSTB(I572097), .Q(I572065) );
nand I_33503 (I572292,I697322,I697304);
and I_33504 (I572309,I572292,I697313);
DFFARX1 I_33505  ( .D(I572309), .CLK(I2702), .RSTB(I572097), .Q(I572326) );
nor I_33506 (I572086,I572326,I572148);
nand I_33507 (I572077,I572326,I572247);
DFFARX1 I_33508  ( .D(I697328), .CLK(I2702), .RSTB(I572097), .Q(I572371) );
and I_33509 (I572388,I572371,I697301);
DFFARX1 I_33510  ( .D(I572388), .CLK(I2702), .RSTB(I572097), .Q(I572405) );
not I_33511 (I572068,I572405);
nand I_33512 (I572436,I572388,I572326);
and I_33513 (I572453,I572148,I572436);
DFFARX1 I_33514  ( .D(I572453), .CLK(I2702), .RSTB(I572097), .Q(I572059) );
DFFARX1 I_33515  ( .D(I697325), .CLK(I2702), .RSTB(I572097), .Q(I572484) );
nand I_33516 (I572501,I572484,I572148);
and I_33517 (I572518,I572326,I572501);
DFFARX1 I_33518  ( .D(I572518), .CLK(I2702), .RSTB(I572097), .Q(I572089) );
not I_33519 (I572549,I572484);
nor I_33520 (I572566,I572165,I572549);
and I_33521 (I572583,I572484,I572566);
or I_33522 (I572600,I572388,I572583);
DFFARX1 I_33523  ( .D(I572600), .CLK(I2702), .RSTB(I572097), .Q(I572074) );
nand I_33524 (I572071,I572484,I572230);
DFFARX1 I_33525  ( .D(I572484), .CLK(I2702), .RSTB(I572097), .Q(I572062) );
not I_33526 (I572692,I2709);
nand I_33527 (I572709,I45351,I45357);
and I_33528 (I572726,I572709,I45354);
DFFARX1 I_33529  ( .D(I572726), .CLK(I2702), .RSTB(I572692), .Q(I572743) );
nor I_33530 (I572760,I45378,I45357);
nor I_33531 (I572777,I572760,I572743);
not I_33532 (I572675,I572760);
DFFARX1 I_33533  ( .D(I45369), .CLK(I2702), .RSTB(I572692), .Q(I572808) );
not I_33534 (I572825,I572808);
nor I_33535 (I572842,I572760,I572825);
nand I_33536 (I572678,I572808,I572777);
DFFARX1 I_33537  ( .D(I572808), .CLK(I2702), .RSTB(I572692), .Q(I572660) );
nand I_33538 (I572887,I45372,I45375);
and I_33539 (I572904,I572887,I45348);
DFFARX1 I_33540  ( .D(I572904), .CLK(I2702), .RSTB(I572692), .Q(I572921) );
nor I_33541 (I572681,I572921,I572743);
nand I_33542 (I572672,I572921,I572842);
DFFARX1 I_33543  ( .D(I45366), .CLK(I2702), .RSTB(I572692), .Q(I572966) );
and I_33544 (I572983,I572966,I45360);
DFFARX1 I_33545  ( .D(I572983), .CLK(I2702), .RSTB(I572692), .Q(I573000) );
not I_33546 (I572663,I573000);
nand I_33547 (I573031,I572983,I572921);
and I_33548 (I573048,I572743,I573031);
DFFARX1 I_33549  ( .D(I573048), .CLK(I2702), .RSTB(I572692), .Q(I572654) );
DFFARX1 I_33550  ( .D(I45363), .CLK(I2702), .RSTB(I572692), .Q(I573079) );
nand I_33551 (I573096,I573079,I572743);
and I_33552 (I573113,I572921,I573096);
DFFARX1 I_33553  ( .D(I573113), .CLK(I2702), .RSTB(I572692), .Q(I572684) );
not I_33554 (I573144,I573079);
nor I_33555 (I573161,I572760,I573144);
and I_33556 (I573178,I573079,I573161);
or I_33557 (I573195,I572983,I573178);
DFFARX1 I_33558  ( .D(I573195), .CLK(I2702), .RSTB(I572692), .Q(I572669) );
nand I_33559 (I572666,I573079,I572825);
DFFARX1 I_33560  ( .D(I573079), .CLK(I2702), .RSTB(I572692), .Q(I572657) );
not I_33561 (I573287,I2709);
nand I_33562 (I573304,I441968,I441971);
and I_33563 (I573321,I573304,I441965);
DFFARX1 I_33564  ( .D(I573321), .CLK(I2702), .RSTB(I573287), .Q(I573338) );
nor I_33565 (I573355,I441962,I441971);
nor I_33566 (I573372,I573355,I573338);
not I_33567 (I573270,I573355);
DFFARX1 I_33568  ( .D(I441944), .CLK(I2702), .RSTB(I573287), .Q(I573403) );
not I_33569 (I573420,I573403);
nor I_33570 (I573437,I573355,I573420);
nand I_33571 (I573273,I573403,I573372);
DFFARX1 I_33572  ( .D(I573403), .CLK(I2702), .RSTB(I573287), .Q(I573255) );
nand I_33573 (I573482,I441953,I441950);
and I_33574 (I573499,I573482,I441959);
DFFARX1 I_33575  ( .D(I573499), .CLK(I2702), .RSTB(I573287), .Q(I573516) );
nor I_33576 (I573276,I573516,I573338);
nand I_33577 (I573267,I573516,I573437);
DFFARX1 I_33578  ( .D(I441941), .CLK(I2702), .RSTB(I573287), .Q(I573561) );
and I_33579 (I573578,I573561,I441956);
DFFARX1 I_33580  ( .D(I573578), .CLK(I2702), .RSTB(I573287), .Q(I573595) );
not I_33581 (I573258,I573595);
nand I_33582 (I573626,I573578,I573516);
and I_33583 (I573643,I573338,I573626);
DFFARX1 I_33584  ( .D(I573643), .CLK(I2702), .RSTB(I573287), .Q(I573249) );
DFFARX1 I_33585  ( .D(I441947), .CLK(I2702), .RSTB(I573287), .Q(I573674) );
nand I_33586 (I573691,I573674,I573338);
and I_33587 (I573708,I573516,I573691);
DFFARX1 I_33588  ( .D(I573708), .CLK(I2702), .RSTB(I573287), .Q(I573279) );
not I_33589 (I573739,I573674);
nor I_33590 (I573756,I573355,I573739);
and I_33591 (I573773,I573674,I573756);
or I_33592 (I573790,I573578,I573773);
DFFARX1 I_33593  ( .D(I573790), .CLK(I2702), .RSTB(I573287), .Q(I573264) );
nand I_33594 (I573261,I573674,I573420);
DFFARX1 I_33595  ( .D(I573674), .CLK(I2702), .RSTB(I573287), .Q(I573252) );
not I_33596 (I573882,I2709);
nand I_33597 (I573899,I284097,I284103);
and I_33598 (I573916,I573899,I284085);
DFFARX1 I_33599  ( .D(I573916), .CLK(I2702), .RSTB(I573882), .Q(I573933) );
nor I_33600 (I573950,I284079,I284103);
nor I_33601 (I573967,I573950,I573933);
not I_33602 (I573865,I573950);
DFFARX1 I_33603  ( .D(I284109), .CLK(I2702), .RSTB(I573882), .Q(I573998) );
not I_33604 (I574015,I573998);
nor I_33605 (I574032,I573950,I574015);
nand I_33606 (I573868,I573998,I573967);
DFFARX1 I_33607  ( .D(I573998), .CLK(I2702), .RSTB(I573882), .Q(I573850) );
nand I_33608 (I574077,I284100,I284091);
and I_33609 (I574094,I574077,I284094);
DFFARX1 I_33610  ( .D(I574094), .CLK(I2702), .RSTB(I573882), .Q(I574111) );
nor I_33611 (I573871,I574111,I573933);
nand I_33612 (I573862,I574111,I574032);
DFFARX1 I_33613  ( .D(I284106), .CLK(I2702), .RSTB(I573882), .Q(I574156) );
and I_33614 (I574173,I574156,I284082);
DFFARX1 I_33615  ( .D(I574173), .CLK(I2702), .RSTB(I573882), .Q(I574190) );
not I_33616 (I573853,I574190);
nand I_33617 (I574221,I574173,I574111);
and I_33618 (I574238,I573933,I574221);
DFFARX1 I_33619  ( .D(I574238), .CLK(I2702), .RSTB(I573882), .Q(I573844) );
DFFARX1 I_33620  ( .D(I284088), .CLK(I2702), .RSTB(I573882), .Q(I574269) );
nand I_33621 (I574286,I574269,I573933);
and I_33622 (I574303,I574111,I574286);
DFFARX1 I_33623  ( .D(I574303), .CLK(I2702), .RSTB(I573882), .Q(I573874) );
not I_33624 (I574334,I574269);
nor I_33625 (I574351,I573950,I574334);
and I_33626 (I574368,I574269,I574351);
or I_33627 (I574385,I574173,I574368);
DFFARX1 I_33628  ( .D(I574385), .CLK(I2702), .RSTB(I573882), .Q(I573859) );
nand I_33629 (I573856,I574269,I574015);
DFFARX1 I_33630  ( .D(I574269), .CLK(I2702), .RSTB(I573882), .Q(I573847) );
not I_33631 (I574477,I2709);
nand I_33632 (I574494,I465088,I465091);
and I_33633 (I574511,I574494,I465085);
DFFARX1 I_33634  ( .D(I574511), .CLK(I2702), .RSTB(I574477), .Q(I574528) );
nor I_33635 (I574545,I465082,I465091);
nor I_33636 (I574562,I574545,I574528);
not I_33637 (I574460,I574545);
DFFARX1 I_33638  ( .D(I465064), .CLK(I2702), .RSTB(I574477), .Q(I574593) );
not I_33639 (I574610,I574593);
nor I_33640 (I574627,I574545,I574610);
nand I_33641 (I574463,I574593,I574562);
DFFARX1 I_33642  ( .D(I574593), .CLK(I2702), .RSTB(I574477), .Q(I574445) );
nand I_33643 (I574672,I465073,I465070);
and I_33644 (I574689,I574672,I465079);
DFFARX1 I_33645  ( .D(I574689), .CLK(I2702), .RSTB(I574477), .Q(I574706) );
nor I_33646 (I574466,I574706,I574528);
nand I_33647 (I574457,I574706,I574627);
DFFARX1 I_33648  ( .D(I465061), .CLK(I2702), .RSTB(I574477), .Q(I574751) );
and I_33649 (I574768,I574751,I465076);
DFFARX1 I_33650  ( .D(I574768), .CLK(I2702), .RSTB(I574477), .Q(I574785) );
not I_33651 (I574448,I574785);
nand I_33652 (I574816,I574768,I574706);
and I_33653 (I574833,I574528,I574816);
DFFARX1 I_33654  ( .D(I574833), .CLK(I2702), .RSTB(I574477), .Q(I574439) );
DFFARX1 I_33655  ( .D(I465067), .CLK(I2702), .RSTB(I574477), .Q(I574864) );
nand I_33656 (I574881,I574864,I574528);
and I_33657 (I574898,I574706,I574881);
DFFARX1 I_33658  ( .D(I574898), .CLK(I2702), .RSTB(I574477), .Q(I574469) );
not I_33659 (I574929,I574864);
nor I_33660 (I574946,I574545,I574929);
and I_33661 (I574963,I574864,I574946);
or I_33662 (I574980,I574768,I574963);
DFFARX1 I_33663  ( .D(I574980), .CLK(I2702), .RSTB(I574477), .Q(I574454) );
nand I_33664 (I574451,I574864,I574610);
DFFARX1 I_33665  ( .D(I574864), .CLK(I2702), .RSTB(I574477), .Q(I574442) );
not I_33666 (I575072,I2709);
nand I_33667 (I575089,I480694,I480697);
and I_33668 (I575106,I575089,I480691);
DFFARX1 I_33669  ( .D(I575106), .CLK(I2702), .RSTB(I575072), .Q(I575123) );
nor I_33670 (I575140,I480688,I480697);
nor I_33671 (I575157,I575140,I575123);
not I_33672 (I575055,I575140);
DFFARX1 I_33673  ( .D(I480670), .CLK(I2702), .RSTB(I575072), .Q(I575188) );
not I_33674 (I575205,I575188);
nor I_33675 (I575222,I575140,I575205);
nand I_33676 (I575058,I575188,I575157);
DFFARX1 I_33677  ( .D(I575188), .CLK(I2702), .RSTB(I575072), .Q(I575040) );
nand I_33678 (I575267,I480679,I480676);
and I_33679 (I575284,I575267,I480685);
DFFARX1 I_33680  ( .D(I575284), .CLK(I2702), .RSTB(I575072), .Q(I575301) );
nor I_33681 (I575061,I575301,I575123);
nand I_33682 (I575052,I575301,I575222);
DFFARX1 I_33683  ( .D(I480667), .CLK(I2702), .RSTB(I575072), .Q(I575346) );
and I_33684 (I575363,I575346,I480682);
DFFARX1 I_33685  ( .D(I575363), .CLK(I2702), .RSTB(I575072), .Q(I575380) );
not I_33686 (I575043,I575380);
nand I_33687 (I575411,I575363,I575301);
and I_33688 (I575428,I575123,I575411);
DFFARX1 I_33689  ( .D(I575428), .CLK(I2702), .RSTB(I575072), .Q(I575034) );
DFFARX1 I_33690  ( .D(I480673), .CLK(I2702), .RSTB(I575072), .Q(I575459) );
nand I_33691 (I575476,I575459,I575123);
and I_33692 (I575493,I575301,I575476);
DFFARX1 I_33693  ( .D(I575493), .CLK(I2702), .RSTB(I575072), .Q(I575064) );
not I_33694 (I575524,I575459);
nor I_33695 (I575541,I575140,I575524);
and I_33696 (I575558,I575459,I575541);
or I_33697 (I575575,I575363,I575558);
DFFARX1 I_33698  ( .D(I575575), .CLK(I2702), .RSTB(I575072), .Q(I575049) );
nand I_33699 (I575046,I575459,I575205);
DFFARX1 I_33700  ( .D(I575459), .CLK(I2702), .RSTB(I575072), .Q(I575037) );
not I_33701 (I575667,I2709);
nand I_33702 (I575684,I356415,I356427);
and I_33703 (I575701,I575684,I356409);
DFFARX1 I_33704  ( .D(I575701), .CLK(I2702), .RSTB(I575667), .Q(I575718) );
nor I_33705 (I575735,I356421,I356427);
nor I_33706 (I575752,I575735,I575718);
not I_33707 (I575650,I575735);
DFFARX1 I_33708  ( .D(I356406), .CLK(I2702), .RSTB(I575667), .Q(I575783) );
not I_33709 (I575800,I575783);
nor I_33710 (I575817,I575735,I575800);
nand I_33711 (I575653,I575783,I575752);
DFFARX1 I_33712  ( .D(I575783), .CLK(I2702), .RSTB(I575667), .Q(I575635) );
nand I_33713 (I575862,I356397,I356412);
and I_33714 (I575879,I575862,I356403);
DFFARX1 I_33715  ( .D(I575879), .CLK(I2702), .RSTB(I575667), .Q(I575896) );
nor I_33716 (I575656,I575896,I575718);
nand I_33717 (I575647,I575896,I575817);
DFFARX1 I_33718  ( .D(I356424), .CLK(I2702), .RSTB(I575667), .Q(I575941) );
and I_33719 (I575958,I575941,I356418);
DFFARX1 I_33720  ( .D(I575958), .CLK(I2702), .RSTB(I575667), .Q(I575975) );
not I_33721 (I575638,I575975);
nand I_33722 (I576006,I575958,I575896);
and I_33723 (I576023,I575718,I576006);
DFFARX1 I_33724  ( .D(I576023), .CLK(I2702), .RSTB(I575667), .Q(I575629) );
DFFARX1 I_33725  ( .D(I356400), .CLK(I2702), .RSTB(I575667), .Q(I576054) );
nand I_33726 (I576071,I576054,I575718);
and I_33727 (I576088,I575896,I576071);
DFFARX1 I_33728  ( .D(I576088), .CLK(I2702), .RSTB(I575667), .Q(I575659) );
not I_33729 (I576119,I576054);
nor I_33730 (I576136,I575735,I576119);
and I_33731 (I576153,I576054,I576136);
or I_33732 (I576170,I575958,I576153);
DFFARX1 I_33733  ( .D(I576170), .CLK(I2702), .RSTB(I575667), .Q(I575644) );
nand I_33734 (I575641,I576054,I575800);
DFFARX1 I_33735  ( .D(I576054), .CLK(I2702), .RSTB(I575667), .Q(I575632) );
not I_33736 (I576262,I2709);
nand I_33737 (I576279,I369335,I369347);
and I_33738 (I576296,I576279,I369329);
DFFARX1 I_33739  ( .D(I576296), .CLK(I2702), .RSTB(I576262), .Q(I576313) );
nor I_33740 (I576330,I369341,I369347);
nor I_33741 (I576347,I576330,I576313);
not I_33742 (I576245,I576330);
DFFARX1 I_33743  ( .D(I369326), .CLK(I2702), .RSTB(I576262), .Q(I576378) );
not I_33744 (I576395,I576378);
nor I_33745 (I576412,I576330,I576395);
nand I_33746 (I576248,I576378,I576347);
DFFARX1 I_33747  ( .D(I576378), .CLK(I2702), .RSTB(I576262), .Q(I576230) );
nand I_33748 (I576457,I369317,I369332);
and I_33749 (I576474,I576457,I369323);
DFFARX1 I_33750  ( .D(I576474), .CLK(I2702), .RSTB(I576262), .Q(I576491) );
nor I_33751 (I576251,I576491,I576313);
nand I_33752 (I576242,I576491,I576412);
DFFARX1 I_33753  ( .D(I369344), .CLK(I2702), .RSTB(I576262), .Q(I576536) );
and I_33754 (I576553,I576536,I369338);
DFFARX1 I_33755  ( .D(I576553), .CLK(I2702), .RSTB(I576262), .Q(I576570) );
not I_33756 (I576233,I576570);
nand I_33757 (I576601,I576553,I576491);
and I_33758 (I576618,I576313,I576601);
DFFARX1 I_33759  ( .D(I576618), .CLK(I2702), .RSTB(I576262), .Q(I576224) );
DFFARX1 I_33760  ( .D(I369320), .CLK(I2702), .RSTB(I576262), .Q(I576649) );
nand I_33761 (I576666,I576649,I576313);
and I_33762 (I576683,I576491,I576666);
DFFARX1 I_33763  ( .D(I576683), .CLK(I2702), .RSTB(I576262), .Q(I576254) );
not I_33764 (I576714,I576649);
nor I_33765 (I576731,I576330,I576714);
and I_33766 (I576748,I576649,I576731);
or I_33767 (I576765,I576553,I576748);
DFFARX1 I_33768  ( .D(I576765), .CLK(I2702), .RSTB(I576262), .Q(I576239) );
nand I_33769 (I576236,I576649,I576395);
DFFARX1 I_33770  ( .D(I576649), .CLK(I2702), .RSTB(I576262), .Q(I576227) );
not I_33771 (I576857,I2709);
nand I_33772 (I576874,I88538,I88514);
and I_33773 (I576891,I576874,I88523);
DFFARX1 I_33774  ( .D(I576891), .CLK(I2702), .RSTB(I576857), .Q(I576908) );
nor I_33775 (I576925,I88517,I88514);
DFFARX1 I_33776  ( .D(I88532), .CLK(I2702), .RSTB(I576857), .Q(I576942) );
nand I_33777 (I576959,I576942,I576925);
DFFARX1 I_33778  ( .D(I576942), .CLK(I2702), .RSTB(I576857), .Q(I576828) );
nand I_33779 (I576990,I88526,I88541);
and I_33780 (I577007,I576990,I88520);
DFFARX1 I_33781  ( .D(I577007), .CLK(I2702), .RSTB(I576857), .Q(I577024) );
not I_33782 (I577041,I577024);
nor I_33783 (I577058,I576908,I577041);
and I_33784 (I577075,I576925,I577058);
and I_33785 (I577092,I577024,I576959);
DFFARX1 I_33786  ( .D(I577092), .CLK(I2702), .RSTB(I576857), .Q(I576825) );
DFFARX1 I_33787  ( .D(I577024), .CLK(I2702), .RSTB(I576857), .Q(I576819) );
DFFARX1 I_33788  ( .D(I88511), .CLK(I2702), .RSTB(I576857), .Q(I577137) );
and I_33789 (I577154,I577137,I88529);
nand I_33790 (I577171,I577154,I577024);
nor I_33791 (I576846,I577154,I576925);
not I_33792 (I577202,I577154);
nor I_33793 (I577219,I576908,I577202);
nand I_33794 (I576837,I576942,I577219);
nand I_33795 (I576831,I577024,I577202);
or I_33796 (I577264,I577154,I577075);
DFFARX1 I_33797  ( .D(I577264), .CLK(I2702), .RSTB(I576857), .Q(I576834) );
DFFARX1 I_33798  ( .D(I88535), .CLK(I2702), .RSTB(I576857), .Q(I577295) );
and I_33799 (I577312,I577295,I577171);
DFFARX1 I_33800  ( .D(I577312), .CLK(I2702), .RSTB(I576857), .Q(I576849) );
nor I_33801 (I577343,I577295,I576908);
nand I_33802 (I576843,I577154,I577343);
not I_33803 (I576840,I577295);
DFFARX1 I_33804  ( .D(I577295), .CLK(I2702), .RSTB(I576857), .Q(I577388) );
and I_33805 (I576822,I577295,I577388);
not I_33806 (I577452,I2709);
nand I_33807 (I577469,I359645,I359657);
and I_33808 (I577486,I577469,I359648);
DFFARX1 I_33809  ( .D(I577486), .CLK(I2702), .RSTB(I577452), .Q(I577503) );
nor I_33810 (I577520,I359642,I359657);
DFFARX1 I_33811  ( .D(I359633), .CLK(I2702), .RSTB(I577452), .Q(I577537) );
nand I_33812 (I577554,I577537,I577520);
DFFARX1 I_33813  ( .D(I577537), .CLK(I2702), .RSTB(I577452), .Q(I577423) );
nand I_33814 (I577585,I359639,I359630);
and I_33815 (I577602,I577585,I359636);
DFFARX1 I_33816  ( .D(I577602), .CLK(I2702), .RSTB(I577452), .Q(I577619) );
not I_33817 (I577636,I577619);
nor I_33818 (I577653,I577503,I577636);
and I_33819 (I577670,I577520,I577653);
and I_33820 (I577687,I577619,I577554);
DFFARX1 I_33821  ( .D(I577687), .CLK(I2702), .RSTB(I577452), .Q(I577420) );
DFFARX1 I_33822  ( .D(I577619), .CLK(I2702), .RSTB(I577452), .Q(I577414) );
DFFARX1 I_33823  ( .D(I359651), .CLK(I2702), .RSTB(I577452), .Q(I577732) );
and I_33824 (I577749,I577732,I359627);
nand I_33825 (I577766,I577749,I577619);
nor I_33826 (I577441,I577749,I577520);
not I_33827 (I577797,I577749);
nor I_33828 (I577814,I577503,I577797);
nand I_33829 (I577432,I577537,I577814);
nand I_33830 (I577426,I577619,I577797);
or I_33831 (I577859,I577749,I577670);
DFFARX1 I_33832  ( .D(I577859), .CLK(I2702), .RSTB(I577452), .Q(I577429) );
DFFARX1 I_33833  ( .D(I359654), .CLK(I2702), .RSTB(I577452), .Q(I577890) );
and I_33834 (I577907,I577890,I577766);
DFFARX1 I_33835  ( .D(I577907), .CLK(I2702), .RSTB(I577452), .Q(I577444) );
nor I_33836 (I577938,I577890,I577503);
nand I_33837 (I577438,I577749,I577938);
not I_33838 (I577435,I577890);
DFFARX1 I_33839  ( .D(I577890), .CLK(I2702), .RSTB(I577452), .Q(I577983) );
and I_33840 (I577417,I577890,I577983);
not I_33841 (I578047,I2709);
nand I_33842 (I578064,I208238,I208223);
and I_33843 (I578081,I578064,I208235);
DFFARX1 I_33844  ( .D(I578081), .CLK(I2702), .RSTB(I578047), .Q(I578098) );
nor I_33845 (I578115,I208226,I208223);
DFFARX1 I_33846  ( .D(I208217), .CLK(I2702), .RSTB(I578047), .Q(I578132) );
nand I_33847 (I578149,I578132,I578115);
DFFARX1 I_33848  ( .D(I578132), .CLK(I2702), .RSTB(I578047), .Q(I578018) );
nand I_33849 (I578180,I208208,I208232);
and I_33850 (I578197,I578180,I208211);
DFFARX1 I_33851  ( .D(I578197), .CLK(I2702), .RSTB(I578047), .Q(I578214) );
not I_33852 (I578231,I578214);
nor I_33853 (I578248,I578098,I578231);
and I_33854 (I578265,I578115,I578248);
and I_33855 (I578282,I578214,I578149);
DFFARX1 I_33856  ( .D(I578282), .CLK(I2702), .RSTB(I578047), .Q(I578015) );
DFFARX1 I_33857  ( .D(I578214), .CLK(I2702), .RSTB(I578047), .Q(I578009) );
DFFARX1 I_33858  ( .D(I208229), .CLK(I2702), .RSTB(I578047), .Q(I578327) );
and I_33859 (I578344,I578327,I208214);
nand I_33860 (I578361,I578344,I578214);
nor I_33861 (I578036,I578344,I578115);
not I_33862 (I578392,I578344);
nor I_33863 (I578409,I578098,I578392);
nand I_33864 (I578027,I578132,I578409);
nand I_33865 (I578021,I578214,I578392);
or I_33866 (I578454,I578344,I578265);
DFFARX1 I_33867  ( .D(I578454), .CLK(I2702), .RSTB(I578047), .Q(I578024) );
DFFARX1 I_33868  ( .D(I208220), .CLK(I2702), .RSTB(I578047), .Q(I578485) );
and I_33869 (I578502,I578485,I578361);
DFFARX1 I_33870  ( .D(I578502), .CLK(I2702), .RSTB(I578047), .Q(I578039) );
nor I_33871 (I578533,I578485,I578098);
nand I_33872 (I578033,I578344,I578533);
not I_33873 (I578030,I578485);
DFFARX1 I_33874  ( .D(I578485), .CLK(I2702), .RSTB(I578047), .Q(I578578) );
and I_33875 (I578012,I578485,I578578);
not I_33876 (I578642,I2709);
nand I_33877 (I578659,I273501,I273471);
and I_33878 (I578676,I578659,I273489);
DFFARX1 I_33879  ( .D(I578676), .CLK(I2702), .RSTB(I578642), .Q(I578693) );
nor I_33880 (I578710,I273483,I273471);
DFFARX1 I_33881  ( .D(I273480), .CLK(I2702), .RSTB(I578642), .Q(I578727) );
nand I_33882 (I578744,I578727,I578710);
DFFARX1 I_33883  ( .D(I578727), .CLK(I2702), .RSTB(I578642), .Q(I578613) );
nand I_33884 (I578775,I273474,I273477);
and I_33885 (I578792,I578775,I273495);
DFFARX1 I_33886  ( .D(I578792), .CLK(I2702), .RSTB(I578642), .Q(I578809) );
not I_33887 (I578826,I578809);
nor I_33888 (I578843,I578693,I578826);
and I_33889 (I578860,I578710,I578843);
and I_33890 (I578877,I578809,I578744);
DFFARX1 I_33891  ( .D(I578877), .CLK(I2702), .RSTB(I578642), .Q(I578610) );
DFFARX1 I_33892  ( .D(I578809), .CLK(I2702), .RSTB(I578642), .Q(I578604) );
DFFARX1 I_33893  ( .D(I273498), .CLK(I2702), .RSTB(I578642), .Q(I578922) );
and I_33894 (I578939,I578922,I273492);
nand I_33895 (I578956,I578939,I578809);
nor I_33896 (I578631,I578939,I578710);
not I_33897 (I578987,I578939);
nor I_33898 (I579004,I578693,I578987);
nand I_33899 (I578622,I578727,I579004);
nand I_33900 (I578616,I578809,I578987);
or I_33901 (I579049,I578939,I578860);
DFFARX1 I_33902  ( .D(I579049), .CLK(I2702), .RSTB(I578642), .Q(I578619) );
DFFARX1 I_33903  ( .D(I273486), .CLK(I2702), .RSTB(I578642), .Q(I579080) );
and I_33904 (I579097,I579080,I578956);
DFFARX1 I_33905  ( .D(I579097), .CLK(I2702), .RSTB(I578642), .Q(I578634) );
nor I_33906 (I579128,I579080,I578693);
nand I_33907 (I578628,I578939,I579128);
not I_33908 (I578625,I579080);
DFFARX1 I_33909  ( .D(I579080), .CLK(I2702), .RSTB(I578642), .Q(I579173) );
and I_33910 (I578607,I579080,I579173);
not I_33911 (I579237,I2709);
nand I_33912 (I579254,I391945,I391957);
and I_33913 (I579271,I579254,I391948);
DFFARX1 I_33914  ( .D(I579271), .CLK(I2702), .RSTB(I579237), .Q(I579288) );
nor I_33915 (I579305,I391942,I391957);
DFFARX1 I_33916  ( .D(I391933), .CLK(I2702), .RSTB(I579237), .Q(I579322) );
nand I_33917 (I579339,I579322,I579305);
DFFARX1 I_33918  ( .D(I579322), .CLK(I2702), .RSTB(I579237), .Q(I579208) );
nand I_33919 (I579370,I391939,I391930);
and I_33920 (I579387,I579370,I391936);
DFFARX1 I_33921  ( .D(I579387), .CLK(I2702), .RSTB(I579237), .Q(I579404) );
not I_33922 (I579421,I579404);
nor I_33923 (I579438,I579288,I579421);
and I_33924 (I579455,I579305,I579438);
and I_33925 (I579472,I579404,I579339);
DFFARX1 I_33926  ( .D(I579472), .CLK(I2702), .RSTB(I579237), .Q(I579205) );
DFFARX1 I_33927  ( .D(I579404), .CLK(I2702), .RSTB(I579237), .Q(I579199) );
DFFARX1 I_33928  ( .D(I391951), .CLK(I2702), .RSTB(I579237), .Q(I579517) );
and I_33929 (I579534,I579517,I391927);
nand I_33930 (I579551,I579534,I579404);
nor I_33931 (I579226,I579534,I579305);
not I_33932 (I579582,I579534);
nor I_33933 (I579599,I579288,I579582);
nand I_33934 (I579217,I579322,I579599);
nand I_33935 (I579211,I579404,I579582);
or I_33936 (I579644,I579534,I579455);
DFFARX1 I_33937  ( .D(I579644), .CLK(I2702), .RSTB(I579237), .Q(I579214) );
DFFARX1 I_33938  ( .D(I391954), .CLK(I2702), .RSTB(I579237), .Q(I579675) );
and I_33939 (I579692,I579675,I579551);
DFFARX1 I_33940  ( .D(I579692), .CLK(I2702), .RSTB(I579237), .Q(I579229) );
nor I_33941 (I579723,I579675,I579288);
nand I_33942 (I579223,I579534,I579723);
not I_33943 (I579220,I579675);
DFFARX1 I_33944  ( .D(I579675), .CLK(I2702), .RSTB(I579237), .Q(I579768) );
and I_33945 (I579202,I579675,I579768);
not I_33946 (I579832,I2709);
nand I_33947 (I579849,I214783,I214768);
and I_33948 (I579866,I579849,I214780);
DFFARX1 I_33949  ( .D(I579866), .CLK(I2702), .RSTB(I579832), .Q(I579883) );
nor I_33950 (I579900,I214771,I214768);
DFFARX1 I_33951  ( .D(I214762), .CLK(I2702), .RSTB(I579832), .Q(I579917) );
nand I_33952 (I579934,I579917,I579900);
DFFARX1 I_33953  ( .D(I579917), .CLK(I2702), .RSTB(I579832), .Q(I579803) );
nand I_33954 (I579965,I214753,I214777);
and I_33955 (I579982,I579965,I214756);
DFFARX1 I_33956  ( .D(I579982), .CLK(I2702), .RSTB(I579832), .Q(I579999) );
not I_33957 (I580016,I579999);
nor I_33958 (I580033,I579883,I580016);
and I_33959 (I580050,I579900,I580033);
and I_33960 (I580067,I579999,I579934);
DFFARX1 I_33961  ( .D(I580067), .CLK(I2702), .RSTB(I579832), .Q(I579800) );
DFFARX1 I_33962  ( .D(I579999), .CLK(I2702), .RSTB(I579832), .Q(I579794) );
DFFARX1 I_33963  ( .D(I214774), .CLK(I2702), .RSTB(I579832), .Q(I580112) );
and I_33964 (I580129,I580112,I214759);
nand I_33965 (I580146,I580129,I579999);
nor I_33966 (I579821,I580129,I579900);
not I_33967 (I580177,I580129);
nor I_33968 (I580194,I579883,I580177);
nand I_33969 (I579812,I579917,I580194);
nand I_33970 (I579806,I579999,I580177);
or I_33971 (I580239,I580129,I580050);
DFFARX1 I_33972  ( .D(I580239), .CLK(I2702), .RSTB(I579832), .Q(I579809) );
DFFARX1 I_33973  ( .D(I214765), .CLK(I2702), .RSTB(I579832), .Q(I580270) );
and I_33974 (I580287,I580270,I580146);
DFFARX1 I_33975  ( .D(I580287), .CLK(I2702), .RSTB(I579832), .Q(I579824) );
nor I_33976 (I580318,I580270,I579883);
nand I_33977 (I579818,I580129,I580318);
not I_33978 (I579815,I580270);
DFFARX1 I_33979  ( .D(I580270), .CLK(I2702), .RSTB(I579832), .Q(I580363) );
and I_33980 (I579797,I580270,I580363);
not I_33981 (I580427,I2709);
nand I_33982 (I580444,I195903,I195924);
and I_33983 (I580461,I580444,I195909);
DFFARX1 I_33984  ( .D(I580461), .CLK(I2702), .RSTB(I580427), .Q(I580478) );
nor I_33985 (I580495,I195927,I195924);
DFFARX1 I_33986  ( .D(I195930), .CLK(I2702), .RSTB(I580427), .Q(I580512) );
nand I_33987 (I580529,I580512,I580495);
DFFARX1 I_33988  ( .D(I580512), .CLK(I2702), .RSTB(I580427), .Q(I580398) );
nand I_33989 (I580560,I195900,I195912);
and I_33990 (I580577,I580560,I195921);
DFFARX1 I_33991  ( .D(I580577), .CLK(I2702), .RSTB(I580427), .Q(I580594) );
not I_33992 (I580611,I580594);
nor I_33993 (I580628,I580478,I580611);
and I_33994 (I580645,I580495,I580628);
and I_33995 (I580662,I580594,I580529);
DFFARX1 I_33996  ( .D(I580662), .CLK(I2702), .RSTB(I580427), .Q(I580395) );
DFFARX1 I_33997  ( .D(I580594), .CLK(I2702), .RSTB(I580427), .Q(I580389) );
DFFARX1 I_33998  ( .D(I195915), .CLK(I2702), .RSTB(I580427), .Q(I580707) );
and I_33999 (I580724,I580707,I195918);
nand I_34000 (I580741,I580724,I580594);
nor I_34001 (I580416,I580724,I580495);
not I_34002 (I580772,I580724);
nor I_34003 (I580789,I580478,I580772);
nand I_34004 (I580407,I580512,I580789);
nand I_34005 (I580401,I580594,I580772);
or I_34006 (I580834,I580724,I580645);
DFFARX1 I_34007  ( .D(I580834), .CLK(I2702), .RSTB(I580427), .Q(I580404) );
DFFARX1 I_34008  ( .D(I195906), .CLK(I2702), .RSTB(I580427), .Q(I580865) );
and I_34009 (I580882,I580865,I580741);
DFFARX1 I_34010  ( .D(I580882), .CLK(I2702), .RSTB(I580427), .Q(I580419) );
nor I_34011 (I580913,I580865,I580478);
nand I_34012 (I580413,I580724,I580913);
not I_34013 (I580410,I580865);
DFFARX1 I_34014  ( .D(I580865), .CLK(I2702), .RSTB(I580427), .Q(I580958) );
and I_34015 (I580392,I580865,I580958);
not I_34016 (I581022,I2709);
nand I_34017 (I581039,I379671,I379683);
and I_34018 (I581056,I581039,I379674);
DFFARX1 I_34019  ( .D(I581056), .CLK(I2702), .RSTB(I581022), .Q(I581073) );
nor I_34020 (I581090,I379668,I379683);
DFFARX1 I_34021  ( .D(I379659), .CLK(I2702), .RSTB(I581022), .Q(I581107) );
nand I_34022 (I581124,I581107,I581090);
DFFARX1 I_34023  ( .D(I581107), .CLK(I2702), .RSTB(I581022), .Q(I580993) );
nand I_34024 (I581155,I379665,I379656);
and I_34025 (I581172,I581155,I379662);
DFFARX1 I_34026  ( .D(I581172), .CLK(I2702), .RSTB(I581022), .Q(I581189) );
not I_34027 (I581206,I581189);
nor I_34028 (I581223,I581073,I581206);
and I_34029 (I581240,I581090,I581223);
and I_34030 (I581257,I581189,I581124);
DFFARX1 I_34031  ( .D(I581257), .CLK(I2702), .RSTB(I581022), .Q(I580990) );
DFFARX1 I_34032  ( .D(I581189), .CLK(I2702), .RSTB(I581022), .Q(I580984) );
DFFARX1 I_34033  ( .D(I379677), .CLK(I2702), .RSTB(I581022), .Q(I581302) );
and I_34034 (I581319,I581302,I379653);
nand I_34035 (I581336,I581319,I581189);
nor I_34036 (I581011,I581319,I581090);
not I_34037 (I581367,I581319);
nor I_34038 (I581384,I581073,I581367);
nand I_34039 (I581002,I581107,I581384);
nand I_34040 (I580996,I581189,I581367);
or I_34041 (I581429,I581319,I581240);
DFFARX1 I_34042  ( .D(I581429), .CLK(I2702), .RSTB(I581022), .Q(I580999) );
DFFARX1 I_34043  ( .D(I379680), .CLK(I2702), .RSTB(I581022), .Q(I581460) );
and I_34044 (I581477,I581460,I581336);
DFFARX1 I_34045  ( .D(I581477), .CLK(I2702), .RSTB(I581022), .Q(I581014) );
nor I_34046 (I581508,I581460,I581073);
nand I_34047 (I581008,I581319,I581508);
not I_34048 (I581005,I581460);
DFFARX1 I_34049  ( .D(I581460), .CLK(I2702), .RSTB(I581022), .Q(I581553) );
and I_34050 (I580987,I581460,I581553);
not I_34051 (I581617,I2709);
nand I_34052 (I581634,I355123,I355135);
and I_34053 (I581651,I581634,I355126);
DFFARX1 I_34054  ( .D(I581651), .CLK(I2702), .RSTB(I581617), .Q(I581668) );
nor I_34055 (I581685,I355120,I355135);
DFFARX1 I_34056  ( .D(I355111), .CLK(I2702), .RSTB(I581617), .Q(I581702) );
nand I_34057 (I581719,I581702,I581685);
DFFARX1 I_34058  ( .D(I581702), .CLK(I2702), .RSTB(I581617), .Q(I581588) );
nand I_34059 (I581750,I355117,I355108);
and I_34060 (I581767,I581750,I355114);
DFFARX1 I_34061  ( .D(I581767), .CLK(I2702), .RSTB(I581617), .Q(I581784) );
not I_34062 (I581801,I581784);
nor I_34063 (I581818,I581668,I581801);
and I_34064 (I581835,I581685,I581818);
and I_34065 (I581852,I581784,I581719);
DFFARX1 I_34066  ( .D(I581852), .CLK(I2702), .RSTB(I581617), .Q(I581585) );
DFFARX1 I_34067  ( .D(I581784), .CLK(I2702), .RSTB(I581617), .Q(I581579) );
DFFARX1 I_34068  ( .D(I355129), .CLK(I2702), .RSTB(I581617), .Q(I581897) );
and I_34069 (I581914,I581897,I355105);
nand I_34070 (I581931,I581914,I581784);
nor I_34071 (I581606,I581914,I581685);
not I_34072 (I581962,I581914);
nor I_34073 (I581979,I581668,I581962);
nand I_34074 (I581597,I581702,I581979);
nand I_34075 (I581591,I581784,I581962);
or I_34076 (I582024,I581914,I581835);
DFFARX1 I_34077  ( .D(I582024), .CLK(I2702), .RSTB(I581617), .Q(I581594) );
DFFARX1 I_34078  ( .D(I355132), .CLK(I2702), .RSTB(I581617), .Q(I582055) );
and I_34079 (I582072,I582055,I581931);
DFFARX1 I_34080  ( .D(I582072), .CLK(I2702), .RSTB(I581617), .Q(I581609) );
nor I_34081 (I582103,I582055,I581668);
nand I_34082 (I581603,I581914,I582103);
not I_34083 (I581600,I582055);
DFFARX1 I_34084  ( .D(I582055), .CLK(I2702), .RSTB(I581617), .Q(I582148) );
and I_34085 (I581582,I582055,I582148);
not I_34086 (I582212,I2709);
nand I_34087 (I582229,I408095,I408107);
and I_34088 (I582246,I582229,I408098);
DFFARX1 I_34089  ( .D(I582246), .CLK(I2702), .RSTB(I582212), .Q(I582263) );
nor I_34090 (I582280,I408092,I408107);
DFFARX1 I_34091  ( .D(I408083), .CLK(I2702), .RSTB(I582212), .Q(I582297) );
nand I_34092 (I582314,I582297,I582280);
DFFARX1 I_34093  ( .D(I582297), .CLK(I2702), .RSTB(I582212), .Q(I582183) );
nand I_34094 (I582345,I408089,I408080);
and I_34095 (I582362,I582345,I408086);
DFFARX1 I_34096  ( .D(I582362), .CLK(I2702), .RSTB(I582212), .Q(I582379) );
not I_34097 (I582396,I582379);
nor I_34098 (I582413,I582263,I582396);
and I_34099 (I582430,I582280,I582413);
and I_34100 (I582447,I582379,I582314);
DFFARX1 I_34101  ( .D(I582447), .CLK(I2702), .RSTB(I582212), .Q(I582180) );
DFFARX1 I_34102  ( .D(I582379), .CLK(I2702), .RSTB(I582212), .Q(I582174) );
DFFARX1 I_34103  ( .D(I408101), .CLK(I2702), .RSTB(I582212), .Q(I582492) );
and I_34104 (I582509,I582492,I408077);
nand I_34105 (I582526,I582509,I582379);
nor I_34106 (I582201,I582509,I582280);
not I_34107 (I582557,I582509);
nor I_34108 (I582574,I582263,I582557);
nand I_34109 (I582192,I582297,I582574);
nand I_34110 (I582186,I582379,I582557);
or I_34111 (I582619,I582509,I582430);
DFFARX1 I_34112  ( .D(I582619), .CLK(I2702), .RSTB(I582212), .Q(I582189) );
DFFARX1 I_34113  ( .D(I408104), .CLK(I2702), .RSTB(I582212), .Q(I582650) );
and I_34114 (I582667,I582650,I582526);
DFFARX1 I_34115  ( .D(I582667), .CLK(I2702), .RSTB(I582212), .Q(I582204) );
nor I_34116 (I582698,I582650,I582263);
nand I_34117 (I582198,I582509,I582698);
not I_34118 (I582195,I582650);
DFFARX1 I_34119  ( .D(I582650), .CLK(I2702), .RSTB(I582212), .Q(I582743) );
and I_34120 (I582177,I582650,I582743);
not I_34121 (I582807,I2709);
nand I_34122 (I582824,I517929,I517914);
and I_34123 (I582841,I582824,I517920);
DFFARX1 I_34124  ( .D(I582841), .CLK(I2702), .RSTB(I582807), .Q(I582858) );
nor I_34125 (I582875,I517923,I517914);
DFFARX1 I_34126  ( .D(I517935), .CLK(I2702), .RSTB(I582807), .Q(I582892) );
nand I_34127 (I582909,I582892,I582875);
DFFARX1 I_34128  ( .D(I582892), .CLK(I2702), .RSTB(I582807), .Q(I582778) );
nand I_34129 (I582940,I517926,I517917);
and I_34130 (I582957,I582940,I517944);
DFFARX1 I_34131  ( .D(I582957), .CLK(I2702), .RSTB(I582807), .Q(I582974) );
not I_34132 (I582991,I582974);
nor I_34133 (I583008,I582858,I582991);
and I_34134 (I583025,I582875,I583008);
and I_34135 (I583042,I582974,I582909);
DFFARX1 I_34136  ( .D(I583042), .CLK(I2702), .RSTB(I582807), .Q(I582775) );
DFFARX1 I_34137  ( .D(I582974), .CLK(I2702), .RSTB(I582807), .Q(I582769) );
DFFARX1 I_34138  ( .D(I517932), .CLK(I2702), .RSTB(I582807), .Q(I583087) );
and I_34139 (I583104,I583087,I517938);
nand I_34140 (I583121,I583104,I582974);
nor I_34141 (I582796,I583104,I582875);
not I_34142 (I583152,I583104);
nor I_34143 (I583169,I582858,I583152);
nand I_34144 (I582787,I582892,I583169);
nand I_34145 (I582781,I582974,I583152);
or I_34146 (I583214,I583104,I583025);
DFFARX1 I_34147  ( .D(I583214), .CLK(I2702), .RSTB(I582807), .Q(I582784) );
DFFARX1 I_34148  ( .D(I517941), .CLK(I2702), .RSTB(I582807), .Q(I583245) );
and I_34149 (I583262,I583245,I583121);
DFFARX1 I_34150  ( .D(I583262), .CLK(I2702), .RSTB(I582807), .Q(I582799) );
nor I_34151 (I583293,I583245,I582858);
nand I_34152 (I582793,I583104,I583293);
not I_34153 (I582790,I583245);
DFFARX1 I_34154  ( .D(I583245), .CLK(I2702), .RSTB(I582807), .Q(I583338) );
and I_34155 (I582772,I583245,I583338);
not I_34156 (I583402,I2709);
nand I_34157 (I583419,I237366,I237363);
and I_34158 (I583436,I583419,I237390);
DFFARX1 I_34159  ( .D(I583436), .CLK(I2702), .RSTB(I583402), .Q(I583453) );
nor I_34160 (I583470,I237393,I237363);
DFFARX1 I_34161  ( .D(I237381), .CLK(I2702), .RSTB(I583402), .Q(I583487) );
nand I_34162 (I583504,I583487,I583470);
DFFARX1 I_34163  ( .D(I583487), .CLK(I2702), .RSTB(I583402), .Q(I583373) );
nand I_34164 (I583535,I237387,I237372);
and I_34165 (I583552,I583535,I237378);
DFFARX1 I_34166  ( .D(I583552), .CLK(I2702), .RSTB(I583402), .Q(I583569) );
not I_34167 (I583586,I583569);
nor I_34168 (I583603,I583453,I583586);
and I_34169 (I583620,I583470,I583603);
and I_34170 (I583637,I583569,I583504);
DFFARX1 I_34171  ( .D(I583637), .CLK(I2702), .RSTB(I583402), .Q(I583370) );
DFFARX1 I_34172  ( .D(I583569), .CLK(I2702), .RSTB(I583402), .Q(I583364) );
DFFARX1 I_34173  ( .D(I237369), .CLK(I2702), .RSTB(I583402), .Q(I583682) );
and I_34174 (I583699,I583682,I237375);
nand I_34175 (I583716,I583699,I583569);
nor I_34176 (I583391,I583699,I583470);
not I_34177 (I583747,I583699);
nor I_34178 (I583764,I583453,I583747);
nand I_34179 (I583382,I583487,I583764);
nand I_34180 (I583376,I583569,I583747);
or I_34181 (I583809,I583699,I583620);
DFFARX1 I_34182  ( .D(I583809), .CLK(I2702), .RSTB(I583402), .Q(I583379) );
DFFARX1 I_34183  ( .D(I237384), .CLK(I2702), .RSTB(I583402), .Q(I583840) );
and I_34184 (I583857,I583840,I583716);
DFFARX1 I_34185  ( .D(I583857), .CLK(I2702), .RSTB(I583402), .Q(I583394) );
nor I_34186 (I583888,I583840,I583453);
nand I_34187 (I583388,I583699,I583888);
not I_34188 (I583385,I583840);
DFFARX1 I_34189  ( .D(I583840), .CLK(I2702), .RSTB(I583402), .Q(I583933) );
and I_34190 (I583367,I583840,I583933);
not I_34191 (I583997,I2709);
nand I_34192 (I584014,I371919,I371931);
and I_34193 (I584031,I584014,I371922);
DFFARX1 I_34194  ( .D(I584031), .CLK(I2702), .RSTB(I583997), .Q(I584048) );
nor I_34195 (I584065,I371916,I371931);
DFFARX1 I_34196  ( .D(I371907), .CLK(I2702), .RSTB(I583997), .Q(I584082) );
nand I_34197 (I584099,I584082,I584065);
DFFARX1 I_34198  ( .D(I584082), .CLK(I2702), .RSTB(I583997), .Q(I583968) );
nand I_34199 (I584130,I371913,I371904);
and I_34200 (I584147,I584130,I371910);
DFFARX1 I_34201  ( .D(I584147), .CLK(I2702), .RSTB(I583997), .Q(I584164) );
not I_34202 (I584181,I584164);
nor I_34203 (I584198,I584048,I584181);
and I_34204 (I584215,I584065,I584198);
and I_34205 (I584232,I584164,I584099);
DFFARX1 I_34206  ( .D(I584232), .CLK(I2702), .RSTB(I583997), .Q(I583965) );
DFFARX1 I_34207  ( .D(I584164), .CLK(I2702), .RSTB(I583997), .Q(I583959) );
DFFARX1 I_34208  ( .D(I371925), .CLK(I2702), .RSTB(I583997), .Q(I584277) );
and I_34209 (I584294,I584277,I371901);
nand I_34210 (I584311,I584294,I584164);
nor I_34211 (I583986,I584294,I584065);
not I_34212 (I584342,I584294);
nor I_34213 (I584359,I584048,I584342);
nand I_34214 (I583977,I584082,I584359);
nand I_34215 (I583971,I584164,I584342);
or I_34216 (I584404,I584294,I584215);
DFFARX1 I_34217  ( .D(I584404), .CLK(I2702), .RSTB(I583997), .Q(I583974) );
DFFARX1 I_34218  ( .D(I371928), .CLK(I2702), .RSTB(I583997), .Q(I584435) );
and I_34219 (I584452,I584435,I584311);
DFFARX1 I_34220  ( .D(I584452), .CLK(I2702), .RSTB(I583997), .Q(I583989) );
nor I_34221 (I584483,I584435,I584048);
nand I_34222 (I583983,I584294,I584483);
not I_34223 (I583980,I584435);
DFFARX1 I_34224  ( .D(I584435), .CLK(I2702), .RSTB(I583997), .Q(I584528) );
and I_34225 (I583962,I584435,I584528);
not I_34226 (I584592,I2709);
nand I_34227 (I584609,I12813,I12828);
and I_34228 (I584626,I584609,I12834);
DFFARX1 I_34229  ( .D(I584626), .CLK(I2702), .RSTB(I584592), .Q(I584643) );
nor I_34230 (I584660,I12822,I12828);
DFFARX1 I_34231  ( .D(I12810), .CLK(I2702), .RSTB(I584592), .Q(I584677) );
nand I_34232 (I584694,I584677,I584660);
DFFARX1 I_34233  ( .D(I584677), .CLK(I2702), .RSTB(I584592), .Q(I584563) );
nand I_34234 (I584725,I12816,I12819);
and I_34235 (I584742,I584725,I12825);
DFFARX1 I_34236  ( .D(I584742), .CLK(I2702), .RSTB(I584592), .Q(I584759) );
not I_34237 (I584776,I584759);
nor I_34238 (I584793,I584643,I584776);
and I_34239 (I584810,I584660,I584793);
and I_34240 (I584827,I584759,I584694);
DFFARX1 I_34241  ( .D(I584827), .CLK(I2702), .RSTB(I584592), .Q(I584560) );
DFFARX1 I_34242  ( .D(I584759), .CLK(I2702), .RSTB(I584592), .Q(I584554) );
DFFARX1 I_34243  ( .D(I12831), .CLK(I2702), .RSTB(I584592), .Q(I584872) );
and I_34244 (I584889,I584872,I12840);
nand I_34245 (I584906,I584889,I584759);
nor I_34246 (I584581,I584889,I584660);
not I_34247 (I584937,I584889);
nor I_34248 (I584954,I584643,I584937);
nand I_34249 (I584572,I584677,I584954);
nand I_34250 (I584566,I584759,I584937);
or I_34251 (I584999,I584889,I584810);
DFFARX1 I_34252  ( .D(I584999), .CLK(I2702), .RSTB(I584592), .Q(I584569) );
DFFARX1 I_34253  ( .D(I12837), .CLK(I2702), .RSTB(I584592), .Q(I585030) );
and I_34254 (I585047,I585030,I584906);
DFFARX1 I_34255  ( .D(I585047), .CLK(I2702), .RSTB(I584592), .Q(I584584) );
nor I_34256 (I585078,I585030,I584643);
nand I_34257 (I584578,I584889,I585078);
not I_34258 (I584575,I585030);
DFFARX1 I_34259  ( .D(I585030), .CLK(I2702), .RSTB(I584592), .Q(I585123) );
and I_34260 (I584557,I585030,I585123);
not I_34261 (I585187,I2709);
nand I_34262 (I585204,I254274,I254244);
and I_34263 (I585221,I585204,I254262);
DFFARX1 I_34264  ( .D(I585221), .CLK(I2702), .RSTB(I585187), .Q(I585238) );
nor I_34265 (I585255,I254256,I254244);
DFFARX1 I_34266  ( .D(I254253), .CLK(I2702), .RSTB(I585187), .Q(I585272) );
nand I_34267 (I585289,I585272,I585255);
DFFARX1 I_34268  ( .D(I585272), .CLK(I2702), .RSTB(I585187), .Q(I585158) );
nand I_34269 (I585320,I254247,I254250);
and I_34270 (I585337,I585320,I254268);
DFFARX1 I_34271  ( .D(I585337), .CLK(I2702), .RSTB(I585187), .Q(I585354) );
not I_34272 (I585371,I585354);
nor I_34273 (I585388,I585238,I585371);
and I_34274 (I585405,I585255,I585388);
and I_34275 (I585422,I585354,I585289);
DFFARX1 I_34276  ( .D(I585422), .CLK(I2702), .RSTB(I585187), .Q(I585155) );
DFFARX1 I_34277  ( .D(I585354), .CLK(I2702), .RSTB(I585187), .Q(I585149) );
DFFARX1 I_34278  ( .D(I254271), .CLK(I2702), .RSTB(I585187), .Q(I585467) );
and I_34279 (I585484,I585467,I254265);
nand I_34280 (I585501,I585484,I585354);
nor I_34281 (I585176,I585484,I585255);
not I_34282 (I585532,I585484);
nor I_34283 (I585549,I585238,I585532);
nand I_34284 (I585167,I585272,I585549);
nand I_34285 (I585161,I585354,I585532);
or I_34286 (I585594,I585484,I585405);
DFFARX1 I_34287  ( .D(I585594), .CLK(I2702), .RSTB(I585187), .Q(I585164) );
DFFARX1 I_34288  ( .D(I254259), .CLK(I2702), .RSTB(I585187), .Q(I585625) );
and I_34289 (I585642,I585625,I585501);
DFFARX1 I_34290  ( .D(I585642), .CLK(I2702), .RSTB(I585187), .Q(I585179) );
nor I_34291 (I585673,I585625,I585238);
nand I_34292 (I585173,I585484,I585673);
not I_34293 (I585170,I585625);
DFFARX1 I_34294  ( .D(I585625), .CLK(I2702), .RSTB(I585187), .Q(I585718) );
and I_34295 (I585152,I585625,I585718);
not I_34296 (I585782,I2709);
nand I_34297 (I585799,I102750,I102726);
and I_34298 (I585816,I585799,I102735);
DFFARX1 I_34299  ( .D(I585816), .CLK(I2702), .RSTB(I585782), .Q(I585833) );
nor I_34300 (I585850,I102729,I102726);
DFFARX1 I_34301  ( .D(I102744), .CLK(I2702), .RSTB(I585782), .Q(I585867) );
nand I_34302 (I585884,I585867,I585850);
DFFARX1 I_34303  ( .D(I585867), .CLK(I2702), .RSTB(I585782), .Q(I585753) );
nand I_34304 (I585915,I102738,I102753);
and I_34305 (I585932,I585915,I102732);
DFFARX1 I_34306  ( .D(I585932), .CLK(I2702), .RSTB(I585782), .Q(I585949) );
not I_34307 (I585966,I585949);
nor I_34308 (I585983,I585833,I585966);
and I_34309 (I586000,I585850,I585983);
and I_34310 (I586017,I585949,I585884);
DFFARX1 I_34311  ( .D(I586017), .CLK(I2702), .RSTB(I585782), .Q(I585750) );
DFFARX1 I_34312  ( .D(I585949), .CLK(I2702), .RSTB(I585782), .Q(I585744) );
DFFARX1 I_34313  ( .D(I102723), .CLK(I2702), .RSTB(I585782), .Q(I586062) );
and I_34314 (I586079,I586062,I102741);
nand I_34315 (I586096,I586079,I585949);
nor I_34316 (I585771,I586079,I585850);
not I_34317 (I586127,I586079);
nor I_34318 (I586144,I585833,I586127);
nand I_34319 (I585762,I585867,I586144);
nand I_34320 (I585756,I585949,I586127);
or I_34321 (I586189,I586079,I586000);
DFFARX1 I_34322  ( .D(I586189), .CLK(I2702), .RSTB(I585782), .Q(I585759) );
DFFARX1 I_34323  ( .D(I102747), .CLK(I2702), .RSTB(I585782), .Q(I586220) );
and I_34324 (I586237,I586220,I586096);
DFFARX1 I_34325  ( .D(I586237), .CLK(I2702), .RSTB(I585782), .Q(I585774) );
nor I_34326 (I586268,I586220,I585833);
nand I_34327 (I585768,I586079,I586268);
not I_34328 (I585765,I586220);
DFFARX1 I_34329  ( .D(I586220), .CLK(I2702), .RSTB(I585782), .Q(I586313) );
and I_34330 (I585747,I586220,I586313);
not I_34331 (I586377,I2709);
nand I_34332 (I586394,I446577,I446592);
and I_34333 (I586411,I586394,I446589);
DFFARX1 I_34334  ( .D(I586411), .CLK(I2702), .RSTB(I586377), .Q(I586428) );
nor I_34335 (I586445,I446565,I446592);
DFFARX1 I_34336  ( .D(I446583), .CLK(I2702), .RSTB(I586377), .Q(I586462) );
nand I_34337 (I586479,I586462,I586445);
DFFARX1 I_34338  ( .D(I586462), .CLK(I2702), .RSTB(I586377), .Q(I586348) );
nand I_34339 (I586510,I446586,I446574);
and I_34340 (I586527,I586510,I446580);
DFFARX1 I_34341  ( .D(I586527), .CLK(I2702), .RSTB(I586377), .Q(I586544) );
not I_34342 (I586561,I586544);
nor I_34343 (I586578,I586428,I586561);
and I_34344 (I586595,I586445,I586578);
and I_34345 (I586612,I586544,I586479);
DFFARX1 I_34346  ( .D(I586612), .CLK(I2702), .RSTB(I586377), .Q(I586345) );
DFFARX1 I_34347  ( .D(I586544), .CLK(I2702), .RSTB(I586377), .Q(I586339) );
DFFARX1 I_34348  ( .D(I446571), .CLK(I2702), .RSTB(I586377), .Q(I586657) );
and I_34349 (I586674,I586657,I446595);
nand I_34350 (I586691,I586674,I586544);
nor I_34351 (I586366,I586674,I586445);
not I_34352 (I586722,I586674);
nor I_34353 (I586739,I586428,I586722);
nand I_34354 (I586357,I586462,I586739);
nand I_34355 (I586351,I586544,I586722);
or I_34356 (I586784,I586674,I586595);
DFFARX1 I_34357  ( .D(I586784), .CLK(I2702), .RSTB(I586377), .Q(I586354) );
DFFARX1 I_34358  ( .D(I446568), .CLK(I2702), .RSTB(I586377), .Q(I586815) );
and I_34359 (I586832,I586815,I586691);
DFFARX1 I_34360  ( .D(I586832), .CLK(I2702), .RSTB(I586377), .Q(I586369) );
nor I_34361 (I586863,I586815,I586428);
nand I_34362 (I586363,I586674,I586863);
not I_34363 (I586360,I586815);
DFFARX1 I_34364  ( .D(I586815), .CLK(I2702), .RSTB(I586377), .Q(I586908) );
and I_34365 (I586342,I586815,I586908);
not I_34366 (I586972,I2709);
nand I_34367 (I586989,I226088,I226073);
and I_34368 (I587006,I586989,I226085);
DFFARX1 I_34369  ( .D(I587006), .CLK(I2702), .RSTB(I586972), .Q(I587023) );
nor I_34370 (I587040,I226076,I226073);
DFFARX1 I_34371  ( .D(I226067), .CLK(I2702), .RSTB(I586972), .Q(I587057) );
nand I_34372 (I587074,I587057,I587040);
DFFARX1 I_34373  ( .D(I587057), .CLK(I2702), .RSTB(I586972), .Q(I586943) );
nand I_34374 (I587105,I226058,I226082);
and I_34375 (I587122,I587105,I226061);
DFFARX1 I_34376  ( .D(I587122), .CLK(I2702), .RSTB(I586972), .Q(I587139) );
not I_34377 (I587156,I587139);
nor I_34378 (I587173,I587023,I587156);
and I_34379 (I587190,I587040,I587173);
and I_34380 (I587207,I587139,I587074);
DFFARX1 I_34381  ( .D(I587207), .CLK(I2702), .RSTB(I586972), .Q(I586940) );
DFFARX1 I_34382  ( .D(I587139), .CLK(I2702), .RSTB(I586972), .Q(I586934) );
DFFARX1 I_34383  ( .D(I226079), .CLK(I2702), .RSTB(I586972), .Q(I587252) );
and I_34384 (I587269,I587252,I226064);
nand I_34385 (I587286,I587269,I587139);
nor I_34386 (I586961,I587269,I587040);
not I_34387 (I587317,I587269);
nor I_34388 (I587334,I587023,I587317);
nand I_34389 (I586952,I587057,I587334);
nand I_34390 (I586946,I587139,I587317);
or I_34391 (I587379,I587269,I587190);
DFFARX1 I_34392  ( .D(I587379), .CLK(I2702), .RSTB(I586972), .Q(I586949) );
DFFARX1 I_34393  ( .D(I226070), .CLK(I2702), .RSTB(I586972), .Q(I587410) );
and I_34394 (I587427,I587410,I587286);
DFFARX1 I_34395  ( .D(I587427), .CLK(I2702), .RSTB(I586972), .Q(I586964) );
nor I_34396 (I587458,I587410,I587023);
nand I_34397 (I586958,I587269,I587458);
not I_34398 (I586955,I587410);
DFFARX1 I_34399  ( .D(I587410), .CLK(I2702), .RSTB(I586972), .Q(I587503) );
and I_34400 (I586937,I587410,I587503);
not I_34401 (I587567,I2709);
nand I_34402 (I587584,I481257,I481272);
and I_34403 (I587601,I587584,I481269);
DFFARX1 I_34404  ( .D(I587601), .CLK(I2702), .RSTB(I587567), .Q(I587618) );
nor I_34405 (I587635,I481245,I481272);
DFFARX1 I_34406  ( .D(I481263), .CLK(I2702), .RSTB(I587567), .Q(I587652) );
nand I_34407 (I587669,I587652,I587635);
DFFARX1 I_34408  ( .D(I587652), .CLK(I2702), .RSTB(I587567), .Q(I587538) );
nand I_34409 (I587700,I481266,I481254);
and I_34410 (I587717,I587700,I481260);
DFFARX1 I_34411  ( .D(I587717), .CLK(I2702), .RSTB(I587567), .Q(I587734) );
not I_34412 (I587751,I587734);
nor I_34413 (I587768,I587618,I587751);
and I_34414 (I587785,I587635,I587768);
and I_34415 (I587802,I587734,I587669);
DFFARX1 I_34416  ( .D(I587802), .CLK(I2702), .RSTB(I587567), .Q(I587535) );
DFFARX1 I_34417  ( .D(I587734), .CLK(I2702), .RSTB(I587567), .Q(I587529) );
DFFARX1 I_34418  ( .D(I481251), .CLK(I2702), .RSTB(I587567), .Q(I587847) );
and I_34419 (I587864,I587847,I481275);
nand I_34420 (I587881,I587864,I587734);
nor I_34421 (I587556,I587864,I587635);
not I_34422 (I587912,I587864);
nor I_34423 (I587929,I587618,I587912);
nand I_34424 (I587547,I587652,I587929);
nand I_34425 (I587541,I587734,I587912);
or I_34426 (I587974,I587864,I587785);
DFFARX1 I_34427  ( .D(I587974), .CLK(I2702), .RSTB(I587567), .Q(I587544) );
DFFARX1 I_34428  ( .D(I481248), .CLK(I2702), .RSTB(I587567), .Q(I588005) );
and I_34429 (I588022,I588005,I587881);
DFFARX1 I_34430  ( .D(I588022), .CLK(I2702), .RSTB(I587567), .Q(I587559) );
nor I_34431 (I588053,I588005,I587618);
nand I_34432 (I587553,I587864,I588053);
not I_34433 (I587550,I588005);
DFFARX1 I_34434  ( .D(I588005), .CLK(I2702), .RSTB(I587567), .Q(I588098) );
and I_34435 (I587532,I588005,I588098);
not I_34436 (I588162,I2709);
nand I_34437 (I588179,I262230,I262200);
and I_34438 (I588196,I588179,I262218);
DFFARX1 I_34439  ( .D(I588196), .CLK(I2702), .RSTB(I588162), .Q(I588213) );
nor I_34440 (I588230,I262212,I262200);
DFFARX1 I_34441  ( .D(I262209), .CLK(I2702), .RSTB(I588162), .Q(I588247) );
nand I_34442 (I588264,I588247,I588230);
DFFARX1 I_34443  ( .D(I588247), .CLK(I2702), .RSTB(I588162), .Q(I588133) );
nand I_34444 (I588295,I262203,I262206);
and I_34445 (I588312,I588295,I262224);
DFFARX1 I_34446  ( .D(I588312), .CLK(I2702), .RSTB(I588162), .Q(I588329) );
not I_34447 (I588346,I588329);
nor I_34448 (I588363,I588213,I588346);
and I_34449 (I588380,I588230,I588363);
and I_34450 (I588397,I588329,I588264);
DFFARX1 I_34451  ( .D(I588397), .CLK(I2702), .RSTB(I588162), .Q(I588130) );
DFFARX1 I_34452  ( .D(I588329), .CLK(I2702), .RSTB(I588162), .Q(I588124) );
DFFARX1 I_34453  ( .D(I262227), .CLK(I2702), .RSTB(I588162), .Q(I588442) );
and I_34454 (I588459,I588442,I262221);
nand I_34455 (I588476,I588459,I588329);
nor I_34456 (I588151,I588459,I588230);
not I_34457 (I588507,I588459);
nor I_34458 (I588524,I588213,I588507);
nand I_34459 (I588142,I588247,I588524);
nand I_34460 (I588136,I588329,I588507);
or I_34461 (I588569,I588459,I588380);
DFFARX1 I_34462  ( .D(I588569), .CLK(I2702), .RSTB(I588162), .Q(I588139) );
DFFARX1 I_34463  ( .D(I262215), .CLK(I2702), .RSTB(I588162), .Q(I588600) );
and I_34464 (I588617,I588600,I588476);
DFFARX1 I_34465  ( .D(I588617), .CLK(I2702), .RSTB(I588162), .Q(I588154) );
nor I_34466 (I588648,I588600,I588213);
nand I_34467 (I588148,I588459,I588648);
not I_34468 (I588145,I588600);
DFFARX1 I_34469  ( .D(I588600), .CLK(I2702), .RSTB(I588162), .Q(I588693) );
and I_34470 (I588127,I588600,I588693);
not I_34471 (I588757,I2709);
nand I_34472 (I588774,I701344,I701347);
and I_34473 (I588791,I588774,I701356);
DFFARX1 I_34474  ( .D(I588791), .CLK(I2702), .RSTB(I588757), .Q(I588808) );
nor I_34475 (I588825,I701350,I701347);
DFFARX1 I_34476  ( .D(I701371), .CLK(I2702), .RSTB(I588757), .Q(I588842) );
nand I_34477 (I588859,I588842,I588825);
DFFARX1 I_34478  ( .D(I588842), .CLK(I2702), .RSTB(I588757), .Q(I588728) );
nand I_34479 (I588890,I701368,I701374);
and I_34480 (I588907,I588890,I701359);
DFFARX1 I_34481  ( .D(I588907), .CLK(I2702), .RSTB(I588757), .Q(I588924) );
not I_34482 (I588941,I588924);
nor I_34483 (I588958,I588808,I588941);
and I_34484 (I588975,I588825,I588958);
and I_34485 (I588992,I588924,I588859);
DFFARX1 I_34486  ( .D(I588992), .CLK(I2702), .RSTB(I588757), .Q(I588725) );
DFFARX1 I_34487  ( .D(I588924), .CLK(I2702), .RSTB(I588757), .Q(I588719) );
DFFARX1 I_34488  ( .D(I701362), .CLK(I2702), .RSTB(I588757), .Q(I589037) );
and I_34489 (I589054,I589037,I701365);
nand I_34490 (I589071,I589054,I588924);
nor I_34491 (I588746,I589054,I588825);
not I_34492 (I589102,I589054);
nor I_34493 (I589119,I588808,I589102);
nand I_34494 (I588737,I588842,I589119);
nand I_34495 (I588731,I588924,I589102);
or I_34496 (I589164,I589054,I588975);
DFFARX1 I_34497  ( .D(I589164), .CLK(I2702), .RSTB(I588757), .Q(I588734) );
DFFARX1 I_34498  ( .D(I701353), .CLK(I2702), .RSTB(I588757), .Q(I589195) );
and I_34499 (I589212,I589195,I589071);
DFFARX1 I_34500  ( .D(I589212), .CLK(I2702), .RSTB(I588757), .Q(I588749) );
nor I_34501 (I589243,I589195,I588808);
nand I_34502 (I588743,I589054,I589243);
not I_34503 (I588740,I589195);
DFFARX1 I_34504  ( .D(I589195), .CLK(I2702), .RSTB(I588757), .Q(I589288) );
and I_34505 (I588722,I589195,I589288);
not I_34506 (I589352,I2709);
nand I_34507 (I589369,I285435,I285405);
and I_34508 (I589386,I589369,I285423);
DFFARX1 I_34509  ( .D(I589386), .CLK(I2702), .RSTB(I589352), .Q(I589403) );
nor I_34510 (I589420,I285417,I285405);
DFFARX1 I_34511  ( .D(I285414), .CLK(I2702), .RSTB(I589352), .Q(I589437) );
nand I_34512 (I589454,I589437,I589420);
DFFARX1 I_34513  ( .D(I589437), .CLK(I2702), .RSTB(I589352), .Q(I589323) );
nand I_34514 (I589485,I285408,I285411);
and I_34515 (I589502,I589485,I285429);
DFFARX1 I_34516  ( .D(I589502), .CLK(I2702), .RSTB(I589352), .Q(I589519) );
not I_34517 (I589536,I589519);
nor I_34518 (I589553,I589403,I589536);
and I_34519 (I589570,I589420,I589553);
and I_34520 (I589587,I589519,I589454);
DFFARX1 I_34521  ( .D(I589587), .CLK(I2702), .RSTB(I589352), .Q(I589320) );
DFFARX1 I_34522  ( .D(I589519), .CLK(I2702), .RSTB(I589352), .Q(I589314) );
DFFARX1 I_34523  ( .D(I285432), .CLK(I2702), .RSTB(I589352), .Q(I589632) );
and I_34524 (I589649,I589632,I285426);
nand I_34525 (I589666,I589649,I589519);
nor I_34526 (I589341,I589649,I589420);
not I_34527 (I589697,I589649);
nor I_34528 (I589714,I589403,I589697);
nand I_34529 (I589332,I589437,I589714);
nand I_34530 (I589326,I589519,I589697);
or I_34531 (I589759,I589649,I589570);
DFFARX1 I_34532  ( .D(I589759), .CLK(I2702), .RSTB(I589352), .Q(I589329) );
DFFARX1 I_34533  ( .D(I285420), .CLK(I2702), .RSTB(I589352), .Q(I589790) );
and I_34534 (I589807,I589790,I589666);
DFFARX1 I_34535  ( .D(I589807), .CLK(I2702), .RSTB(I589352), .Q(I589344) );
nor I_34536 (I589838,I589790,I589403);
nand I_34537 (I589338,I589649,I589838);
not I_34538 (I589335,I589790);
DFFARX1 I_34539  ( .D(I589790), .CLK(I2702), .RSTB(I589352), .Q(I589883) );
and I_34540 (I589317,I589790,I589883);
not I_34541 (I589947,I2709);
nand I_34542 (I589964,I286761,I286731);
and I_34543 (I589981,I589964,I286749);
DFFARX1 I_34544  ( .D(I589981), .CLK(I2702), .RSTB(I589947), .Q(I589998) );
nor I_34545 (I590015,I286743,I286731);
DFFARX1 I_34546  ( .D(I286740), .CLK(I2702), .RSTB(I589947), .Q(I590032) );
nand I_34547 (I590049,I590032,I590015);
DFFARX1 I_34548  ( .D(I590032), .CLK(I2702), .RSTB(I589947), .Q(I589918) );
nand I_34549 (I590080,I286734,I286737);
and I_34550 (I590097,I590080,I286755);
DFFARX1 I_34551  ( .D(I590097), .CLK(I2702), .RSTB(I589947), .Q(I590114) );
not I_34552 (I590131,I590114);
nor I_34553 (I590148,I589998,I590131);
and I_34554 (I590165,I590015,I590148);
and I_34555 (I590182,I590114,I590049);
DFFARX1 I_34556  ( .D(I590182), .CLK(I2702), .RSTB(I589947), .Q(I589915) );
DFFARX1 I_34557  ( .D(I590114), .CLK(I2702), .RSTB(I589947), .Q(I589909) );
DFFARX1 I_34558  ( .D(I286758), .CLK(I2702), .RSTB(I589947), .Q(I590227) );
and I_34559 (I590244,I590227,I286752);
nand I_34560 (I590261,I590244,I590114);
nor I_34561 (I589936,I590244,I590015);
not I_34562 (I590292,I590244);
nor I_34563 (I590309,I589998,I590292);
nand I_34564 (I589927,I590032,I590309);
nand I_34565 (I589921,I590114,I590292);
or I_34566 (I590354,I590244,I590165);
DFFARX1 I_34567  ( .D(I590354), .CLK(I2702), .RSTB(I589947), .Q(I589924) );
DFFARX1 I_34568  ( .D(I286746), .CLK(I2702), .RSTB(I589947), .Q(I590385) );
and I_34569 (I590402,I590385,I590261);
DFFARX1 I_34570  ( .D(I590402), .CLK(I2702), .RSTB(I589947), .Q(I589939) );
nor I_34571 (I590433,I590385,I589998);
nand I_34572 (I589933,I590244,I590433);
not I_34573 (I589930,I590385);
DFFARX1 I_34574  ( .D(I590385), .CLK(I2702), .RSTB(I589947), .Q(I590478) );
and I_34575 (I589912,I590385,I590478);
not I_34576 (I590542,I2709);
nand I_34577 (I590559,I67220,I67196);
and I_34578 (I590576,I590559,I67205);
DFFARX1 I_34579  ( .D(I590576), .CLK(I2702), .RSTB(I590542), .Q(I590593) );
nor I_34580 (I590610,I67199,I67196);
DFFARX1 I_34581  ( .D(I67214), .CLK(I2702), .RSTB(I590542), .Q(I590627) );
nand I_34582 (I590644,I590627,I590610);
DFFARX1 I_34583  ( .D(I590627), .CLK(I2702), .RSTB(I590542), .Q(I590513) );
nand I_34584 (I590675,I67208,I67223);
and I_34585 (I590692,I590675,I67202);
DFFARX1 I_34586  ( .D(I590692), .CLK(I2702), .RSTB(I590542), .Q(I590709) );
not I_34587 (I590726,I590709);
nor I_34588 (I590743,I590593,I590726);
and I_34589 (I590760,I590610,I590743);
and I_34590 (I590777,I590709,I590644);
DFFARX1 I_34591  ( .D(I590777), .CLK(I2702), .RSTB(I590542), .Q(I590510) );
DFFARX1 I_34592  ( .D(I590709), .CLK(I2702), .RSTB(I590542), .Q(I590504) );
DFFARX1 I_34593  ( .D(I67193), .CLK(I2702), .RSTB(I590542), .Q(I590822) );
and I_34594 (I590839,I590822,I67211);
nand I_34595 (I590856,I590839,I590709);
nor I_34596 (I590531,I590839,I590610);
not I_34597 (I590887,I590839);
nor I_34598 (I590904,I590593,I590887);
nand I_34599 (I590522,I590627,I590904);
nand I_34600 (I590516,I590709,I590887);
or I_34601 (I590949,I590839,I590760);
DFFARX1 I_34602  ( .D(I590949), .CLK(I2702), .RSTB(I590542), .Q(I590519) );
DFFARX1 I_34603  ( .D(I67217), .CLK(I2702), .RSTB(I590542), .Q(I590980) );
and I_34604 (I590997,I590980,I590856);
DFFARX1 I_34605  ( .D(I590997), .CLK(I2702), .RSTB(I590542), .Q(I590534) );
nor I_34606 (I591028,I590980,I590593);
nand I_34607 (I590528,I590839,I591028);
not I_34608 (I590525,I590980);
DFFARX1 I_34609  ( .D(I590980), .CLK(I2702), .RSTB(I590542), .Q(I591073) );
and I_34610 (I590507,I590980,I591073);
not I_34611 (I591137,I2709);
nand I_34612 (I591154,I127944,I127920);
and I_34613 (I591171,I591154,I127929);
DFFARX1 I_34614  ( .D(I591171), .CLK(I2702), .RSTB(I591137), .Q(I591188) );
nor I_34615 (I591205,I127923,I127920);
DFFARX1 I_34616  ( .D(I127938), .CLK(I2702), .RSTB(I591137), .Q(I591222) );
nand I_34617 (I591239,I591222,I591205);
DFFARX1 I_34618  ( .D(I591222), .CLK(I2702), .RSTB(I591137), .Q(I591108) );
nand I_34619 (I591270,I127932,I127947);
and I_34620 (I591287,I591270,I127926);
DFFARX1 I_34621  ( .D(I591287), .CLK(I2702), .RSTB(I591137), .Q(I591304) );
not I_34622 (I591321,I591304);
nor I_34623 (I591338,I591188,I591321);
and I_34624 (I591355,I591205,I591338);
and I_34625 (I591372,I591304,I591239);
DFFARX1 I_34626  ( .D(I591372), .CLK(I2702), .RSTB(I591137), .Q(I591105) );
DFFARX1 I_34627  ( .D(I591304), .CLK(I2702), .RSTB(I591137), .Q(I591099) );
DFFARX1 I_34628  ( .D(I127917), .CLK(I2702), .RSTB(I591137), .Q(I591417) );
and I_34629 (I591434,I591417,I127935);
nand I_34630 (I591451,I591434,I591304);
nor I_34631 (I591126,I591434,I591205);
not I_34632 (I591482,I591434);
nor I_34633 (I591499,I591188,I591482);
nand I_34634 (I591117,I591222,I591499);
nand I_34635 (I591111,I591304,I591482);
or I_34636 (I591544,I591434,I591355);
DFFARX1 I_34637  ( .D(I591544), .CLK(I2702), .RSTB(I591137), .Q(I591114) );
DFFARX1 I_34638  ( .D(I127941), .CLK(I2702), .RSTB(I591137), .Q(I591575) );
and I_34639 (I591592,I591575,I591451);
DFFARX1 I_34640  ( .D(I591592), .CLK(I2702), .RSTB(I591137), .Q(I591129) );
nor I_34641 (I591623,I591575,I591188);
nand I_34642 (I591123,I591434,I591623);
not I_34643 (I591120,I591575);
DFFARX1 I_34644  ( .D(I591575), .CLK(I2702), .RSTB(I591137), .Q(I591668) );
and I_34645 (I591102,I591575,I591668);
not I_34646 (I591732,I2709);
nand I_34647 (I591749,I224898,I224883);
and I_34648 (I591766,I591749,I224895);
DFFARX1 I_34649  ( .D(I591766), .CLK(I2702), .RSTB(I591732), .Q(I591783) );
nor I_34650 (I591800,I224886,I224883);
DFFARX1 I_34651  ( .D(I224877), .CLK(I2702), .RSTB(I591732), .Q(I591817) );
nand I_34652 (I591834,I591817,I591800);
DFFARX1 I_34653  ( .D(I591817), .CLK(I2702), .RSTB(I591732), .Q(I591703) );
nand I_34654 (I591865,I224868,I224892);
and I_34655 (I591882,I591865,I224871);
DFFARX1 I_34656  ( .D(I591882), .CLK(I2702), .RSTB(I591732), .Q(I591899) );
not I_34657 (I591916,I591899);
nor I_34658 (I591933,I591783,I591916);
and I_34659 (I591950,I591800,I591933);
and I_34660 (I591967,I591899,I591834);
DFFARX1 I_34661  ( .D(I591967), .CLK(I2702), .RSTB(I591732), .Q(I591700) );
DFFARX1 I_34662  ( .D(I591899), .CLK(I2702), .RSTB(I591732), .Q(I591694) );
DFFARX1 I_34663  ( .D(I224889), .CLK(I2702), .RSTB(I591732), .Q(I592012) );
and I_34664 (I592029,I592012,I224874);
nand I_34665 (I592046,I592029,I591899);
nor I_34666 (I591721,I592029,I591800);
not I_34667 (I592077,I592029);
nor I_34668 (I592094,I591783,I592077);
nand I_34669 (I591712,I591817,I592094);
nand I_34670 (I591706,I591899,I592077);
or I_34671 (I592139,I592029,I591950);
DFFARX1 I_34672  ( .D(I592139), .CLK(I2702), .RSTB(I591732), .Q(I591709) );
DFFARX1 I_34673  ( .D(I224880), .CLK(I2702), .RSTB(I591732), .Q(I592170) );
and I_34674 (I592187,I592170,I592046);
DFFARX1 I_34675  ( .D(I592187), .CLK(I2702), .RSTB(I591732), .Q(I591724) );
nor I_34676 (I592218,I592170,I591783);
nand I_34677 (I591718,I592029,I592218);
not I_34678 (I591715,I592170);
DFFARX1 I_34679  ( .D(I592170), .CLK(I2702), .RSTB(I591732), .Q(I592263) );
and I_34680 (I591697,I592170,I592263);
not I_34681 (I592327,I2709);
nand I_34682 (I592344,I293391,I293361);
and I_34683 (I592361,I592344,I293379);
DFFARX1 I_34684  ( .D(I592361), .CLK(I2702), .RSTB(I592327), .Q(I592378) );
nor I_34685 (I592395,I293373,I293361);
DFFARX1 I_34686  ( .D(I293370), .CLK(I2702), .RSTB(I592327), .Q(I592412) );
nand I_34687 (I592429,I592412,I592395);
DFFARX1 I_34688  ( .D(I592412), .CLK(I2702), .RSTB(I592327), .Q(I592298) );
nand I_34689 (I592460,I293364,I293367);
and I_34690 (I592477,I592460,I293385);
DFFARX1 I_34691  ( .D(I592477), .CLK(I2702), .RSTB(I592327), .Q(I592494) );
not I_34692 (I592511,I592494);
nor I_34693 (I592528,I592378,I592511);
and I_34694 (I592545,I592395,I592528);
and I_34695 (I592562,I592494,I592429);
DFFARX1 I_34696  ( .D(I592562), .CLK(I2702), .RSTB(I592327), .Q(I592295) );
DFFARX1 I_34697  ( .D(I592494), .CLK(I2702), .RSTB(I592327), .Q(I592289) );
DFFARX1 I_34698  ( .D(I293388), .CLK(I2702), .RSTB(I592327), .Q(I592607) );
and I_34699 (I592624,I592607,I293382);
nand I_34700 (I592641,I592624,I592494);
nor I_34701 (I592316,I592624,I592395);
not I_34702 (I592672,I592624);
nor I_34703 (I592689,I592378,I592672);
nand I_34704 (I592307,I592412,I592689);
nand I_34705 (I592301,I592494,I592672);
or I_34706 (I592734,I592624,I592545);
DFFARX1 I_34707  ( .D(I592734), .CLK(I2702), .RSTB(I592327), .Q(I592304) );
DFFARX1 I_34708  ( .D(I293376), .CLK(I2702), .RSTB(I592327), .Q(I592765) );
and I_34709 (I592782,I592765,I592641);
DFFARX1 I_34710  ( .D(I592782), .CLK(I2702), .RSTB(I592327), .Q(I592319) );
nor I_34711 (I592813,I592765,I592378);
nand I_34712 (I592313,I592624,I592813);
not I_34713 (I592310,I592765);
DFFARX1 I_34714  ( .D(I592765), .CLK(I2702), .RSTB(I592327), .Q(I592858) );
and I_34715 (I592292,I592765,I592858);
not I_34716 (I592922,I2709);
nand I_34717 (I592939,I330519,I330489);
and I_34718 (I592956,I592939,I330507);
DFFARX1 I_34719  ( .D(I592956), .CLK(I2702), .RSTB(I592922), .Q(I592973) );
nor I_34720 (I592990,I330501,I330489);
DFFARX1 I_34721  ( .D(I330498), .CLK(I2702), .RSTB(I592922), .Q(I593007) );
nand I_34722 (I593024,I593007,I592990);
DFFARX1 I_34723  ( .D(I593007), .CLK(I2702), .RSTB(I592922), .Q(I592893) );
nand I_34724 (I593055,I330492,I330495);
and I_34725 (I593072,I593055,I330513);
DFFARX1 I_34726  ( .D(I593072), .CLK(I2702), .RSTB(I592922), .Q(I593089) );
not I_34727 (I593106,I593089);
nor I_34728 (I593123,I592973,I593106);
and I_34729 (I593140,I592990,I593123);
and I_34730 (I593157,I593089,I593024);
DFFARX1 I_34731  ( .D(I593157), .CLK(I2702), .RSTB(I592922), .Q(I592890) );
DFFARX1 I_34732  ( .D(I593089), .CLK(I2702), .RSTB(I592922), .Q(I592884) );
DFFARX1 I_34733  ( .D(I330516), .CLK(I2702), .RSTB(I592922), .Q(I593202) );
and I_34734 (I593219,I593202,I330510);
nand I_34735 (I593236,I593219,I593089);
nor I_34736 (I592911,I593219,I592990);
not I_34737 (I593267,I593219);
nor I_34738 (I593284,I592973,I593267);
nand I_34739 (I592902,I593007,I593284);
nand I_34740 (I592896,I593089,I593267);
or I_34741 (I593329,I593219,I593140);
DFFARX1 I_34742  ( .D(I593329), .CLK(I2702), .RSTB(I592922), .Q(I592899) );
DFFARX1 I_34743  ( .D(I330504), .CLK(I2702), .RSTB(I592922), .Q(I593360) );
and I_34744 (I593377,I593360,I593236);
DFFARX1 I_34745  ( .D(I593377), .CLK(I2702), .RSTB(I592922), .Q(I592914) );
nor I_34746 (I593408,I593360,I592973);
nand I_34747 (I592908,I593219,I593408);
not I_34748 (I592905,I593360);
DFFARX1 I_34749  ( .D(I593360), .CLK(I2702), .RSTB(I592922), .Q(I593453) );
and I_34750 (I592887,I593360,I593453);
not I_34751 (I593517,I2709);
nand I_34752 (I593534,I685411,I685399);
and I_34753 (I593551,I593534,I685384);
DFFARX1 I_34754  ( .D(I593551), .CLK(I2702), .RSTB(I593517), .Q(I593568) );
nor I_34755 (I593585,I685396,I685399);
DFFARX1 I_34756  ( .D(I685408), .CLK(I2702), .RSTB(I593517), .Q(I593602) );
nand I_34757 (I593619,I593602,I593585);
DFFARX1 I_34758  ( .D(I593602), .CLK(I2702), .RSTB(I593517), .Q(I593488) );
nand I_34759 (I593650,I685381,I685405);
and I_34760 (I593667,I593650,I685390);
DFFARX1 I_34761  ( .D(I593667), .CLK(I2702), .RSTB(I593517), .Q(I593684) );
not I_34762 (I593701,I593684);
nor I_34763 (I593718,I593568,I593701);
and I_34764 (I593735,I593585,I593718);
and I_34765 (I593752,I593684,I593619);
DFFARX1 I_34766  ( .D(I593752), .CLK(I2702), .RSTB(I593517), .Q(I593485) );
DFFARX1 I_34767  ( .D(I593684), .CLK(I2702), .RSTB(I593517), .Q(I593479) );
DFFARX1 I_34768  ( .D(I685393), .CLK(I2702), .RSTB(I593517), .Q(I593797) );
and I_34769 (I593814,I593797,I685402);
nand I_34770 (I593831,I593814,I593684);
nor I_34771 (I593506,I593814,I593585);
not I_34772 (I593862,I593814);
nor I_34773 (I593879,I593568,I593862);
nand I_34774 (I593497,I593602,I593879);
nand I_34775 (I593491,I593684,I593862);
or I_34776 (I593924,I593814,I593735);
DFFARX1 I_34777  ( .D(I593924), .CLK(I2702), .RSTB(I593517), .Q(I593494) );
DFFARX1 I_34778  ( .D(I685387), .CLK(I2702), .RSTB(I593517), .Q(I593955) );
and I_34779 (I593972,I593955,I593831);
DFFARX1 I_34780  ( .D(I593972), .CLK(I2702), .RSTB(I593517), .Q(I593509) );
nor I_34781 (I594003,I593955,I593568);
nand I_34782 (I593503,I593814,I594003);
not I_34783 (I593500,I593955);
DFFARX1 I_34784  ( .D(I593955), .CLK(I2702), .RSTB(I593517), .Q(I594048) );
and I_34785 (I593482,I593955,I594048);
not I_34786 (I594112,I2709);
nand I_34787 (I594129,I178002,I178023);
and I_34788 (I594146,I594129,I178008);
DFFARX1 I_34789  ( .D(I594146), .CLK(I2702), .RSTB(I594112), .Q(I594163) );
nor I_34790 (I594180,I178026,I178023);
DFFARX1 I_34791  ( .D(I178029), .CLK(I2702), .RSTB(I594112), .Q(I594197) );
nand I_34792 (I594214,I594197,I594180);
DFFARX1 I_34793  ( .D(I594197), .CLK(I2702), .RSTB(I594112), .Q(I594083) );
nand I_34794 (I594245,I177999,I178011);
and I_34795 (I594262,I594245,I178020);
DFFARX1 I_34796  ( .D(I594262), .CLK(I2702), .RSTB(I594112), .Q(I594279) );
not I_34797 (I594296,I594279);
nor I_34798 (I594313,I594163,I594296);
and I_34799 (I594330,I594180,I594313);
and I_34800 (I594347,I594279,I594214);
DFFARX1 I_34801  ( .D(I594347), .CLK(I2702), .RSTB(I594112), .Q(I594080) );
DFFARX1 I_34802  ( .D(I594279), .CLK(I2702), .RSTB(I594112), .Q(I594074) );
DFFARX1 I_34803  ( .D(I178014), .CLK(I2702), .RSTB(I594112), .Q(I594392) );
and I_34804 (I594409,I594392,I178017);
nand I_34805 (I594426,I594409,I594279);
nor I_34806 (I594101,I594409,I594180);
not I_34807 (I594457,I594409);
nor I_34808 (I594474,I594163,I594457);
nand I_34809 (I594092,I594197,I594474);
nand I_34810 (I594086,I594279,I594457);
or I_34811 (I594519,I594409,I594330);
DFFARX1 I_34812  ( .D(I594519), .CLK(I2702), .RSTB(I594112), .Q(I594089) );
DFFARX1 I_34813  ( .D(I178005), .CLK(I2702), .RSTB(I594112), .Q(I594550) );
and I_34814 (I594567,I594550,I594426);
DFFARX1 I_34815  ( .D(I594567), .CLK(I2702), .RSTB(I594112), .Q(I594104) );
nor I_34816 (I594598,I594550,I594163);
nand I_34817 (I594098,I594409,I594598);
not I_34818 (I594095,I594550);
DFFARX1 I_34819  ( .D(I594550), .CLK(I2702), .RSTB(I594112), .Q(I594643) );
and I_34820 (I594077,I594550,I594643);
not I_34821 (I594707,I2709);
nand I_34822 (I594724,I726776,I726779);
and I_34823 (I594741,I594724,I726788);
DFFARX1 I_34824  ( .D(I594741), .CLK(I2702), .RSTB(I594707), .Q(I594758) );
nor I_34825 (I594775,I726782,I726779);
DFFARX1 I_34826  ( .D(I726803), .CLK(I2702), .RSTB(I594707), .Q(I594792) );
nand I_34827 (I594809,I594792,I594775);
DFFARX1 I_34828  ( .D(I594792), .CLK(I2702), .RSTB(I594707), .Q(I594678) );
nand I_34829 (I594840,I726800,I726806);
and I_34830 (I594857,I594840,I726791);
DFFARX1 I_34831  ( .D(I594857), .CLK(I2702), .RSTB(I594707), .Q(I594874) );
not I_34832 (I594891,I594874);
nor I_34833 (I594908,I594758,I594891);
and I_34834 (I594925,I594775,I594908);
and I_34835 (I594942,I594874,I594809);
DFFARX1 I_34836  ( .D(I594942), .CLK(I2702), .RSTB(I594707), .Q(I594675) );
DFFARX1 I_34837  ( .D(I594874), .CLK(I2702), .RSTB(I594707), .Q(I594669) );
DFFARX1 I_34838  ( .D(I726794), .CLK(I2702), .RSTB(I594707), .Q(I594987) );
and I_34839 (I595004,I594987,I726797);
nand I_34840 (I595021,I595004,I594874);
nor I_34841 (I594696,I595004,I594775);
not I_34842 (I595052,I595004);
nor I_34843 (I595069,I594758,I595052);
nand I_34844 (I594687,I594792,I595069);
nand I_34845 (I594681,I594874,I595052);
or I_34846 (I595114,I595004,I594925);
DFFARX1 I_34847  ( .D(I595114), .CLK(I2702), .RSTB(I594707), .Q(I594684) );
DFFARX1 I_34848  ( .D(I726785), .CLK(I2702), .RSTB(I594707), .Q(I595145) );
and I_34849 (I595162,I595145,I595021);
DFFARX1 I_34850  ( .D(I595162), .CLK(I2702), .RSTB(I594707), .Q(I594699) );
nor I_34851 (I595193,I595145,I594758);
nand I_34852 (I594693,I595004,I595193);
not I_34853 (I594690,I595145);
DFFARX1 I_34854  ( .D(I595145), .CLK(I2702), .RSTB(I594707), .Q(I595238) );
and I_34855 (I594672,I595145,I595238);
not I_34856 (I595302,I2709);
nand I_34857 (I595319,I237961,I237958);
and I_34858 (I595336,I595319,I237985);
DFFARX1 I_34859  ( .D(I595336), .CLK(I2702), .RSTB(I595302), .Q(I595353) );
nor I_34860 (I595370,I237988,I237958);
DFFARX1 I_34861  ( .D(I237976), .CLK(I2702), .RSTB(I595302), .Q(I595387) );
nand I_34862 (I595404,I595387,I595370);
DFFARX1 I_34863  ( .D(I595387), .CLK(I2702), .RSTB(I595302), .Q(I595273) );
nand I_34864 (I595435,I237982,I237967);
and I_34865 (I595452,I595435,I237973);
DFFARX1 I_34866  ( .D(I595452), .CLK(I2702), .RSTB(I595302), .Q(I595469) );
not I_34867 (I595486,I595469);
nor I_34868 (I595503,I595353,I595486);
and I_34869 (I595520,I595370,I595503);
and I_34870 (I595537,I595469,I595404);
DFFARX1 I_34871  ( .D(I595537), .CLK(I2702), .RSTB(I595302), .Q(I595270) );
DFFARX1 I_34872  ( .D(I595469), .CLK(I2702), .RSTB(I595302), .Q(I595264) );
DFFARX1 I_34873  ( .D(I237964), .CLK(I2702), .RSTB(I595302), .Q(I595582) );
and I_34874 (I595599,I595582,I237970);
nand I_34875 (I595616,I595599,I595469);
nor I_34876 (I595291,I595599,I595370);
not I_34877 (I595647,I595599);
nor I_34878 (I595664,I595353,I595647);
nand I_34879 (I595282,I595387,I595664);
nand I_34880 (I595276,I595469,I595647);
or I_34881 (I595709,I595599,I595520);
DFFARX1 I_34882  ( .D(I595709), .CLK(I2702), .RSTB(I595302), .Q(I595279) );
DFFARX1 I_34883  ( .D(I237979), .CLK(I2702), .RSTB(I595302), .Q(I595740) );
and I_34884 (I595757,I595740,I595616);
DFFARX1 I_34885  ( .D(I595757), .CLK(I2702), .RSTB(I595302), .Q(I595294) );
nor I_34886 (I595788,I595740,I595353);
nand I_34887 (I595288,I595599,I595788);
not I_34888 (I595285,I595740);
DFFARX1 I_34889  ( .D(I595740), .CLK(I2702), .RSTB(I595302), .Q(I595833) );
and I_34890 (I595267,I595740,I595833);
not I_34891 (I595897,I2709);
nand I_34892 (I595914,I341557,I341569);
and I_34893 (I595931,I595914,I341560);
DFFARX1 I_34894  ( .D(I595931), .CLK(I2702), .RSTB(I595897), .Q(I595948) );
nor I_34895 (I595965,I341554,I341569);
DFFARX1 I_34896  ( .D(I341545), .CLK(I2702), .RSTB(I595897), .Q(I595982) );
nand I_34897 (I595999,I595982,I595965);
DFFARX1 I_34898  ( .D(I595982), .CLK(I2702), .RSTB(I595897), .Q(I595868) );
nand I_34899 (I596030,I341551,I341542);
and I_34900 (I596047,I596030,I341548);
DFFARX1 I_34901  ( .D(I596047), .CLK(I2702), .RSTB(I595897), .Q(I596064) );
not I_34902 (I596081,I596064);
nor I_34903 (I596098,I595948,I596081);
and I_34904 (I596115,I595965,I596098);
and I_34905 (I596132,I596064,I595999);
DFFARX1 I_34906  ( .D(I596132), .CLK(I2702), .RSTB(I595897), .Q(I595865) );
DFFARX1 I_34907  ( .D(I596064), .CLK(I2702), .RSTB(I595897), .Q(I595859) );
DFFARX1 I_34908  ( .D(I341563), .CLK(I2702), .RSTB(I595897), .Q(I596177) );
and I_34909 (I596194,I596177,I341539);
nand I_34910 (I596211,I596194,I596064);
nor I_34911 (I595886,I596194,I595965);
not I_34912 (I596242,I596194);
nor I_34913 (I596259,I595948,I596242);
nand I_34914 (I595877,I595982,I596259);
nand I_34915 (I595871,I596064,I596242);
or I_34916 (I596304,I596194,I596115);
DFFARX1 I_34917  ( .D(I596304), .CLK(I2702), .RSTB(I595897), .Q(I595874) );
DFFARX1 I_34918  ( .D(I341566), .CLK(I2702), .RSTB(I595897), .Q(I596335) );
and I_34919 (I596352,I596335,I596211);
DFFARX1 I_34920  ( .D(I596352), .CLK(I2702), .RSTB(I595897), .Q(I595889) );
nor I_34921 (I596383,I596335,I595948);
nand I_34922 (I595883,I596194,I596383);
not I_34923 (I595880,I596335);
DFFARX1 I_34924  ( .D(I596335), .CLK(I2702), .RSTB(I595897), .Q(I596428) );
and I_34925 (I595862,I596335,I596428);
not I_34926 (I596492,I2709);
nand I_34927 (I596509,I300021,I299991);
and I_34928 (I596526,I596509,I300009);
DFFARX1 I_34929  ( .D(I596526), .CLK(I2702), .RSTB(I596492), .Q(I596543) );
nor I_34930 (I596560,I300003,I299991);
DFFARX1 I_34931  ( .D(I300000), .CLK(I2702), .RSTB(I596492), .Q(I596577) );
nand I_34932 (I596594,I596577,I596560);
DFFARX1 I_34933  ( .D(I596577), .CLK(I2702), .RSTB(I596492), .Q(I596463) );
nand I_34934 (I596625,I299994,I299997);
and I_34935 (I596642,I596625,I300015);
DFFARX1 I_34936  ( .D(I596642), .CLK(I2702), .RSTB(I596492), .Q(I596659) );
not I_34937 (I596676,I596659);
nor I_34938 (I596693,I596543,I596676);
and I_34939 (I596710,I596560,I596693);
and I_34940 (I596727,I596659,I596594);
DFFARX1 I_34941  ( .D(I596727), .CLK(I2702), .RSTB(I596492), .Q(I596460) );
DFFARX1 I_34942  ( .D(I596659), .CLK(I2702), .RSTB(I596492), .Q(I596454) );
DFFARX1 I_34943  ( .D(I300018), .CLK(I2702), .RSTB(I596492), .Q(I596772) );
and I_34944 (I596789,I596772,I300012);
nand I_34945 (I596806,I596789,I596659);
nor I_34946 (I596481,I596789,I596560);
not I_34947 (I596837,I596789);
nor I_34948 (I596854,I596543,I596837);
nand I_34949 (I596472,I596577,I596854);
nand I_34950 (I596466,I596659,I596837);
or I_34951 (I596899,I596789,I596710);
DFFARX1 I_34952  ( .D(I596899), .CLK(I2702), .RSTB(I596492), .Q(I596469) );
DFFARX1 I_34953  ( .D(I300006), .CLK(I2702), .RSTB(I596492), .Q(I596930) );
and I_34954 (I596947,I596930,I596806);
DFFARX1 I_34955  ( .D(I596947), .CLK(I2702), .RSTB(I596492), .Q(I596484) );
nor I_34956 (I596978,I596930,I596543);
nand I_34957 (I596478,I596789,I596978);
not I_34958 (I596475,I596930);
DFFARX1 I_34959  ( .D(I596930), .CLK(I2702), .RSTB(I596492), .Q(I597023) );
and I_34960 (I596457,I596930,I597023);
not I_34961 (I597087,I2709);
nand I_34962 (I597104,I235581,I235578);
and I_34963 (I597121,I597104,I235605);
DFFARX1 I_34964  ( .D(I597121), .CLK(I2702), .RSTB(I597087), .Q(I597138) );
nor I_34965 (I597155,I235608,I235578);
DFFARX1 I_34966  ( .D(I235596), .CLK(I2702), .RSTB(I597087), .Q(I597172) );
nand I_34967 (I597189,I597172,I597155);
DFFARX1 I_34968  ( .D(I597172), .CLK(I2702), .RSTB(I597087), .Q(I597058) );
nand I_34969 (I597220,I235602,I235587);
and I_34970 (I597237,I597220,I235593);
DFFARX1 I_34971  ( .D(I597237), .CLK(I2702), .RSTB(I597087), .Q(I597254) );
not I_34972 (I597271,I597254);
nor I_34973 (I597288,I597138,I597271);
and I_34974 (I597305,I597155,I597288);
and I_34975 (I597322,I597254,I597189);
DFFARX1 I_34976  ( .D(I597322), .CLK(I2702), .RSTB(I597087), .Q(I597055) );
DFFARX1 I_34977  ( .D(I597254), .CLK(I2702), .RSTB(I597087), .Q(I597049) );
DFFARX1 I_34978  ( .D(I235584), .CLK(I2702), .RSTB(I597087), .Q(I597367) );
and I_34979 (I597384,I597367,I235590);
nand I_34980 (I597401,I597384,I597254);
nor I_34981 (I597076,I597384,I597155);
not I_34982 (I597432,I597384);
nor I_34983 (I597449,I597138,I597432);
nand I_34984 (I597067,I597172,I597449);
nand I_34985 (I597061,I597254,I597432);
or I_34986 (I597494,I597384,I597305);
DFFARX1 I_34987  ( .D(I597494), .CLK(I2702), .RSTB(I597087), .Q(I597064) );
DFFARX1 I_34988  ( .D(I235599), .CLK(I2702), .RSTB(I597087), .Q(I597525) );
and I_34989 (I597542,I597525,I597401);
DFFARX1 I_34990  ( .D(I597542), .CLK(I2702), .RSTB(I597087), .Q(I597079) );
nor I_34991 (I597573,I597525,I597138);
nand I_34992 (I597073,I597384,I597573);
not I_34993 (I597070,I597525);
DFFARX1 I_34994  ( .D(I597525), .CLK(I2702), .RSTB(I597087), .Q(I597618) );
and I_34995 (I597052,I597525,I597618);
not I_34996 (I597682,I2709);
nand I_34997 (I597699,I710014,I710017);
and I_34998 (I597716,I597699,I710026);
DFFARX1 I_34999  ( .D(I597716), .CLK(I2702), .RSTB(I597682), .Q(I597733) );
nor I_35000 (I597750,I710020,I710017);
DFFARX1 I_35001  ( .D(I710041), .CLK(I2702), .RSTB(I597682), .Q(I597767) );
nand I_35002 (I597784,I597767,I597750);
DFFARX1 I_35003  ( .D(I597767), .CLK(I2702), .RSTB(I597682), .Q(I597653) );
nand I_35004 (I597815,I710038,I710044);
and I_35005 (I597832,I597815,I710029);
DFFARX1 I_35006  ( .D(I597832), .CLK(I2702), .RSTB(I597682), .Q(I597849) );
not I_35007 (I597866,I597849);
nor I_35008 (I597883,I597733,I597866);
and I_35009 (I597900,I597750,I597883);
and I_35010 (I597917,I597849,I597784);
DFFARX1 I_35011  ( .D(I597917), .CLK(I2702), .RSTB(I597682), .Q(I597650) );
DFFARX1 I_35012  ( .D(I597849), .CLK(I2702), .RSTB(I597682), .Q(I597644) );
DFFARX1 I_35013  ( .D(I710032), .CLK(I2702), .RSTB(I597682), .Q(I597962) );
and I_35014 (I597979,I597962,I710035);
nand I_35015 (I597996,I597979,I597849);
nor I_35016 (I597671,I597979,I597750);
not I_35017 (I598027,I597979);
nor I_35018 (I598044,I597733,I598027);
nand I_35019 (I597662,I597767,I598044);
nand I_35020 (I597656,I597849,I598027);
or I_35021 (I598089,I597979,I597900);
DFFARX1 I_35022  ( .D(I598089), .CLK(I2702), .RSTB(I597682), .Q(I597659) );
DFFARX1 I_35023  ( .D(I710023), .CLK(I2702), .RSTB(I597682), .Q(I598120) );
and I_35024 (I598137,I598120,I597996);
DFFARX1 I_35025  ( .D(I598137), .CLK(I2702), .RSTB(I597682), .Q(I597674) );
nor I_35026 (I598168,I598120,I597733);
nand I_35027 (I597668,I597979,I598168);
not I_35028 (I597665,I598120);
DFFARX1 I_35029  ( .D(I598120), .CLK(I2702), .RSTB(I597682), .Q(I598213) );
and I_35030 (I597647,I598120,I598213);
not I_35031 (I598277,I2709);
nand I_35032 (I598294,I536969,I536954);
and I_35033 (I598311,I598294,I536960);
DFFARX1 I_35034  ( .D(I598311), .CLK(I2702), .RSTB(I598277), .Q(I598328) );
nor I_35035 (I598345,I536963,I536954);
DFFARX1 I_35036  ( .D(I536975), .CLK(I2702), .RSTB(I598277), .Q(I598362) );
nand I_35037 (I598379,I598362,I598345);
DFFARX1 I_35038  ( .D(I598362), .CLK(I2702), .RSTB(I598277), .Q(I598248) );
nand I_35039 (I598410,I536966,I536957);
and I_35040 (I598427,I598410,I536984);
DFFARX1 I_35041  ( .D(I598427), .CLK(I2702), .RSTB(I598277), .Q(I598444) );
not I_35042 (I598461,I598444);
nor I_35043 (I598478,I598328,I598461);
and I_35044 (I598495,I598345,I598478);
and I_35045 (I598512,I598444,I598379);
DFFARX1 I_35046  ( .D(I598512), .CLK(I2702), .RSTB(I598277), .Q(I598245) );
DFFARX1 I_35047  ( .D(I598444), .CLK(I2702), .RSTB(I598277), .Q(I598239) );
DFFARX1 I_35048  ( .D(I536972), .CLK(I2702), .RSTB(I598277), .Q(I598557) );
and I_35049 (I598574,I598557,I536978);
nand I_35050 (I598591,I598574,I598444);
nor I_35051 (I598266,I598574,I598345);
not I_35052 (I598622,I598574);
nor I_35053 (I598639,I598328,I598622);
nand I_35054 (I598257,I598362,I598639);
nand I_35055 (I598251,I598444,I598622);
or I_35056 (I598684,I598574,I598495);
DFFARX1 I_35057  ( .D(I598684), .CLK(I2702), .RSTB(I598277), .Q(I598254) );
DFFARX1 I_35058  ( .D(I536981), .CLK(I2702), .RSTB(I598277), .Q(I598715) );
and I_35059 (I598732,I598715,I598591);
DFFARX1 I_35060  ( .D(I598732), .CLK(I2702), .RSTB(I598277), .Q(I598269) );
nor I_35061 (I598763,I598715,I598328);
nand I_35062 (I598263,I598574,I598763);
not I_35063 (I598260,I598715);
DFFARX1 I_35064  ( .D(I598715), .CLK(I2702), .RSTB(I598277), .Q(I598808) );
and I_35065 (I598242,I598715,I598808);
not I_35066 (I598872,I2709);
nand I_35067 (I598889,I263556,I263526);
and I_35068 (I598906,I598889,I263544);
DFFARX1 I_35069  ( .D(I598906), .CLK(I2702), .RSTB(I598872), .Q(I598923) );
nor I_35070 (I598940,I263538,I263526);
DFFARX1 I_35071  ( .D(I263535), .CLK(I2702), .RSTB(I598872), .Q(I598957) );
nand I_35072 (I598974,I598957,I598940);
DFFARX1 I_35073  ( .D(I598957), .CLK(I2702), .RSTB(I598872), .Q(I598843) );
nand I_35074 (I599005,I263529,I263532);
and I_35075 (I599022,I599005,I263550);
DFFARX1 I_35076  ( .D(I599022), .CLK(I2702), .RSTB(I598872), .Q(I599039) );
not I_35077 (I599056,I599039);
nor I_35078 (I599073,I598923,I599056);
and I_35079 (I599090,I598940,I599073);
and I_35080 (I599107,I599039,I598974);
DFFARX1 I_35081  ( .D(I599107), .CLK(I2702), .RSTB(I598872), .Q(I598840) );
DFFARX1 I_35082  ( .D(I599039), .CLK(I2702), .RSTB(I598872), .Q(I598834) );
DFFARX1 I_35083  ( .D(I263553), .CLK(I2702), .RSTB(I598872), .Q(I599152) );
and I_35084 (I599169,I599152,I263547);
nand I_35085 (I599186,I599169,I599039);
nor I_35086 (I598861,I599169,I598940);
not I_35087 (I599217,I599169);
nor I_35088 (I599234,I598923,I599217);
nand I_35089 (I598852,I598957,I599234);
nand I_35090 (I598846,I599039,I599217);
or I_35091 (I599279,I599169,I599090);
DFFARX1 I_35092  ( .D(I599279), .CLK(I2702), .RSTB(I598872), .Q(I598849) );
DFFARX1 I_35093  ( .D(I263541), .CLK(I2702), .RSTB(I598872), .Q(I599310) );
and I_35094 (I599327,I599310,I599186);
DFFARX1 I_35095  ( .D(I599327), .CLK(I2702), .RSTB(I598872), .Q(I598864) );
nor I_35096 (I599358,I599310,I598923);
nand I_35097 (I598858,I599169,I599358);
not I_35098 (I598855,I599310);
DFFARX1 I_35099  ( .D(I599310), .CLK(I2702), .RSTB(I598872), .Q(I599403) );
and I_35100 (I598837,I599310,I599403);
not I_35101 (I599467,I2709);
nand I_35102 (I599484,I631317,I631305);
and I_35103 (I599501,I599484,I631290);
DFFARX1 I_35104  ( .D(I599501), .CLK(I2702), .RSTB(I599467), .Q(I599518) );
nor I_35105 (I599535,I631302,I631305);
DFFARX1 I_35106  ( .D(I631314), .CLK(I2702), .RSTB(I599467), .Q(I599552) );
nand I_35107 (I599569,I599552,I599535);
DFFARX1 I_35108  ( .D(I599552), .CLK(I2702), .RSTB(I599467), .Q(I599438) );
nand I_35109 (I599600,I631287,I631311);
and I_35110 (I599617,I599600,I631296);
DFFARX1 I_35111  ( .D(I599617), .CLK(I2702), .RSTB(I599467), .Q(I599634) );
not I_35112 (I599651,I599634);
nor I_35113 (I599668,I599518,I599651);
and I_35114 (I599685,I599535,I599668);
and I_35115 (I599702,I599634,I599569);
DFFARX1 I_35116  ( .D(I599702), .CLK(I2702), .RSTB(I599467), .Q(I599435) );
DFFARX1 I_35117  ( .D(I599634), .CLK(I2702), .RSTB(I599467), .Q(I599429) );
DFFARX1 I_35118  ( .D(I631299), .CLK(I2702), .RSTB(I599467), .Q(I599747) );
and I_35119 (I599764,I599747,I631308);
nand I_35120 (I599781,I599764,I599634);
nor I_35121 (I599456,I599764,I599535);
not I_35122 (I599812,I599764);
nor I_35123 (I599829,I599518,I599812);
nand I_35124 (I599447,I599552,I599829);
nand I_35125 (I599441,I599634,I599812);
or I_35126 (I599874,I599764,I599685);
DFFARX1 I_35127  ( .D(I599874), .CLK(I2702), .RSTB(I599467), .Q(I599444) );
DFFARX1 I_35128  ( .D(I631293), .CLK(I2702), .RSTB(I599467), .Q(I599905) );
and I_35129 (I599922,I599905,I599781);
DFFARX1 I_35130  ( .D(I599922), .CLK(I2702), .RSTB(I599467), .Q(I599459) );
nor I_35131 (I599953,I599905,I599518);
nand I_35132 (I599453,I599764,I599953);
not I_35133 (I599450,I599905);
DFFARX1 I_35134  ( .D(I599905), .CLK(I2702), .RSTB(I599467), .Q(I599998) );
and I_35135 (I599432,I599905,I599998);
not I_35136 (I600062,I2709);
nand I_35137 (I600079,I724464,I724467);
and I_35138 (I600096,I600079,I724476);
DFFARX1 I_35139  ( .D(I600096), .CLK(I2702), .RSTB(I600062), .Q(I600113) );
nor I_35140 (I600130,I724470,I724467);
DFFARX1 I_35141  ( .D(I724491), .CLK(I2702), .RSTB(I600062), .Q(I600147) );
nand I_35142 (I600164,I600147,I600130);
DFFARX1 I_35143  ( .D(I600147), .CLK(I2702), .RSTB(I600062), .Q(I600033) );
nand I_35144 (I600195,I724488,I724494);
and I_35145 (I600212,I600195,I724479);
DFFARX1 I_35146  ( .D(I600212), .CLK(I2702), .RSTB(I600062), .Q(I600229) );
not I_35147 (I600246,I600229);
nor I_35148 (I600263,I600113,I600246);
and I_35149 (I600280,I600130,I600263);
and I_35150 (I600297,I600229,I600164);
DFFARX1 I_35151  ( .D(I600297), .CLK(I2702), .RSTB(I600062), .Q(I600030) );
DFFARX1 I_35152  ( .D(I600229), .CLK(I2702), .RSTB(I600062), .Q(I600024) );
DFFARX1 I_35153  ( .D(I724482), .CLK(I2702), .RSTB(I600062), .Q(I600342) );
and I_35154 (I600359,I600342,I724485);
nand I_35155 (I600376,I600359,I600229);
nor I_35156 (I600051,I600359,I600130);
not I_35157 (I600407,I600359);
nor I_35158 (I600424,I600113,I600407);
nand I_35159 (I600042,I600147,I600424);
nand I_35160 (I600036,I600229,I600407);
or I_35161 (I600469,I600359,I600280);
DFFARX1 I_35162  ( .D(I600469), .CLK(I2702), .RSTB(I600062), .Q(I600039) );
DFFARX1 I_35163  ( .D(I724473), .CLK(I2702), .RSTB(I600062), .Q(I600500) );
and I_35164 (I600517,I600500,I600376);
DFFARX1 I_35165  ( .D(I600517), .CLK(I2702), .RSTB(I600062), .Q(I600054) );
nor I_35166 (I600548,I600500,I600113);
nand I_35167 (I600048,I600359,I600548);
not I_35168 (I600045,I600500);
DFFARX1 I_35169  ( .D(I600500), .CLK(I2702), .RSTB(I600062), .Q(I600593) );
and I_35170 (I600027,I600500,I600593);
not I_35171 (I600657,I2709);
nand I_35172 (I600674,I23472,I23487);
and I_35173 (I600691,I600674,I23493);
DFFARX1 I_35174  ( .D(I600691), .CLK(I2702), .RSTB(I600657), .Q(I600708) );
nor I_35175 (I600725,I23481,I23487);
DFFARX1 I_35176  ( .D(I23469), .CLK(I2702), .RSTB(I600657), .Q(I600742) );
nand I_35177 (I600759,I600742,I600725);
DFFARX1 I_35178  ( .D(I600742), .CLK(I2702), .RSTB(I600657), .Q(I600628) );
nand I_35179 (I600790,I23475,I23478);
and I_35180 (I600807,I600790,I23484);
DFFARX1 I_35181  ( .D(I600807), .CLK(I2702), .RSTB(I600657), .Q(I600824) );
not I_35182 (I600841,I600824);
nor I_35183 (I600858,I600708,I600841);
and I_35184 (I600875,I600725,I600858);
and I_35185 (I600892,I600824,I600759);
DFFARX1 I_35186  ( .D(I600892), .CLK(I2702), .RSTB(I600657), .Q(I600625) );
DFFARX1 I_35187  ( .D(I600824), .CLK(I2702), .RSTB(I600657), .Q(I600619) );
DFFARX1 I_35188  ( .D(I23490), .CLK(I2702), .RSTB(I600657), .Q(I600937) );
and I_35189 (I600954,I600937,I23499);
nand I_35190 (I600971,I600954,I600824);
nor I_35191 (I600646,I600954,I600725);
not I_35192 (I601002,I600954);
nor I_35193 (I601019,I600708,I601002);
nand I_35194 (I600637,I600742,I601019);
nand I_35195 (I600631,I600824,I601002);
or I_35196 (I601064,I600954,I600875);
DFFARX1 I_35197  ( .D(I601064), .CLK(I2702), .RSTB(I600657), .Q(I600634) );
DFFARX1 I_35198  ( .D(I23496), .CLK(I2702), .RSTB(I600657), .Q(I601095) );
and I_35199 (I601112,I601095,I600971);
DFFARX1 I_35200  ( .D(I601112), .CLK(I2702), .RSTB(I600657), .Q(I600649) );
nor I_35201 (I601143,I601095,I600708);
nand I_35202 (I600643,I600954,I601143);
not I_35203 (I600640,I601095);
DFFARX1 I_35204  ( .D(I601095), .CLK(I2702), .RSTB(I600657), .Q(I601188) );
and I_35205 (I600622,I601095,I601188);
not I_35206 (I601252,I2709);
nand I_35207 (I601269,I686669,I686657);
and I_35208 (I601286,I601269,I686642);
DFFARX1 I_35209  ( .D(I601286), .CLK(I2702), .RSTB(I601252), .Q(I601303) );
nor I_35210 (I601320,I686654,I686657);
DFFARX1 I_35211  ( .D(I686666), .CLK(I2702), .RSTB(I601252), .Q(I601337) );
nand I_35212 (I601354,I601337,I601320);
DFFARX1 I_35213  ( .D(I601337), .CLK(I2702), .RSTB(I601252), .Q(I601223) );
nand I_35214 (I601385,I686639,I686663);
and I_35215 (I601402,I601385,I686648);
DFFARX1 I_35216  ( .D(I601402), .CLK(I2702), .RSTB(I601252), .Q(I601419) );
not I_35217 (I601436,I601419);
nor I_35218 (I601453,I601303,I601436);
and I_35219 (I601470,I601320,I601453);
and I_35220 (I601487,I601419,I601354);
DFFARX1 I_35221  ( .D(I601487), .CLK(I2702), .RSTB(I601252), .Q(I601220) );
DFFARX1 I_35222  ( .D(I601419), .CLK(I2702), .RSTB(I601252), .Q(I601214) );
DFFARX1 I_35223  ( .D(I686651), .CLK(I2702), .RSTB(I601252), .Q(I601532) );
and I_35224 (I601549,I601532,I686660);
nand I_35225 (I601566,I601549,I601419);
nor I_35226 (I601241,I601549,I601320);
not I_35227 (I601597,I601549);
nor I_35228 (I601614,I601303,I601597);
nand I_35229 (I601232,I601337,I601614);
nand I_35230 (I601226,I601419,I601597);
or I_35231 (I601659,I601549,I601470);
DFFARX1 I_35232  ( .D(I601659), .CLK(I2702), .RSTB(I601252), .Q(I601229) );
DFFARX1 I_35233  ( .D(I686645), .CLK(I2702), .RSTB(I601252), .Q(I601690) );
and I_35234 (I601707,I601690,I601566);
DFFARX1 I_35235  ( .D(I601707), .CLK(I2702), .RSTB(I601252), .Q(I601244) );
nor I_35236 (I601738,I601690,I601303);
nand I_35237 (I601238,I601549,I601738);
not I_35238 (I601235,I601690);
DFFARX1 I_35239  ( .D(I601690), .CLK(I2702), .RSTB(I601252), .Q(I601783) );
and I_35240 (I601217,I601690,I601783);
not I_35241 (I601847,I2709);
nand I_35242 (I601864,I276816,I276786);
and I_35243 (I601881,I601864,I276804);
DFFARX1 I_35244  ( .D(I601881), .CLK(I2702), .RSTB(I601847), .Q(I601898) );
nor I_35245 (I601915,I276798,I276786);
DFFARX1 I_35246  ( .D(I276795), .CLK(I2702), .RSTB(I601847), .Q(I601932) );
nand I_35247 (I601949,I601932,I601915);
DFFARX1 I_35248  ( .D(I601932), .CLK(I2702), .RSTB(I601847), .Q(I601818) );
nand I_35249 (I601980,I276789,I276792);
and I_35250 (I601997,I601980,I276810);
DFFARX1 I_35251  ( .D(I601997), .CLK(I2702), .RSTB(I601847), .Q(I602014) );
not I_35252 (I602031,I602014);
nor I_35253 (I602048,I601898,I602031);
and I_35254 (I602065,I601915,I602048);
and I_35255 (I602082,I602014,I601949);
DFFARX1 I_35256  ( .D(I602082), .CLK(I2702), .RSTB(I601847), .Q(I601815) );
DFFARX1 I_35257  ( .D(I602014), .CLK(I2702), .RSTB(I601847), .Q(I601809) );
DFFARX1 I_35258  ( .D(I276813), .CLK(I2702), .RSTB(I601847), .Q(I602127) );
and I_35259 (I602144,I602127,I276807);
nand I_35260 (I602161,I602144,I602014);
nor I_35261 (I601836,I602144,I601915);
not I_35262 (I602192,I602144);
nor I_35263 (I602209,I601898,I602192);
nand I_35264 (I601827,I601932,I602209);
nand I_35265 (I601821,I602014,I602192);
or I_35266 (I602254,I602144,I602065);
DFFARX1 I_35267  ( .D(I602254), .CLK(I2702), .RSTB(I601847), .Q(I601824) );
DFFARX1 I_35268  ( .D(I276801), .CLK(I2702), .RSTB(I601847), .Q(I602285) );
and I_35269 (I602302,I602285,I602161);
DFFARX1 I_35270  ( .D(I602302), .CLK(I2702), .RSTB(I601847), .Q(I601839) );
nor I_35271 (I602333,I602285,I601898);
nand I_35272 (I601833,I602144,I602333);
not I_35273 (I601830,I602285);
DFFARX1 I_35274  ( .D(I602285), .CLK(I2702), .RSTB(I601847), .Q(I602378) );
and I_35275 (I601812,I602285,I602378);
not I_35276 (I602442,I2709);
nand I_35277 (I602459,I260904,I260874);
and I_35278 (I602476,I602459,I260892);
DFFARX1 I_35279  ( .D(I602476), .CLK(I2702), .RSTB(I602442), .Q(I602493) );
nor I_35280 (I602510,I260886,I260874);
DFFARX1 I_35281  ( .D(I260883), .CLK(I2702), .RSTB(I602442), .Q(I602527) );
nand I_35282 (I602544,I602527,I602510);
DFFARX1 I_35283  ( .D(I602527), .CLK(I2702), .RSTB(I602442), .Q(I602413) );
nand I_35284 (I602575,I260877,I260880);
and I_35285 (I602592,I602575,I260898);
DFFARX1 I_35286  ( .D(I602592), .CLK(I2702), .RSTB(I602442), .Q(I602609) );
not I_35287 (I602626,I602609);
nor I_35288 (I602643,I602493,I602626);
and I_35289 (I602660,I602510,I602643);
and I_35290 (I602677,I602609,I602544);
DFFARX1 I_35291  ( .D(I602677), .CLK(I2702), .RSTB(I602442), .Q(I602410) );
DFFARX1 I_35292  ( .D(I602609), .CLK(I2702), .RSTB(I602442), .Q(I602404) );
DFFARX1 I_35293  ( .D(I260901), .CLK(I2702), .RSTB(I602442), .Q(I602722) );
and I_35294 (I602739,I602722,I260895);
nand I_35295 (I602756,I602739,I602609);
nor I_35296 (I602431,I602739,I602510);
not I_35297 (I602787,I602739);
nor I_35298 (I602804,I602493,I602787);
nand I_35299 (I602422,I602527,I602804);
nand I_35300 (I602416,I602609,I602787);
or I_35301 (I602849,I602739,I602660);
DFFARX1 I_35302  ( .D(I602849), .CLK(I2702), .RSTB(I602442), .Q(I602419) );
DFFARX1 I_35303  ( .D(I260889), .CLK(I2702), .RSTB(I602442), .Q(I602880) );
and I_35304 (I602897,I602880,I602756);
DFFARX1 I_35305  ( .D(I602897), .CLK(I2702), .RSTB(I602442), .Q(I602434) );
nor I_35306 (I602928,I602880,I602493);
nand I_35307 (I602428,I602739,I602928);
not I_35308 (I602425,I602880);
DFFARX1 I_35309  ( .D(I602880), .CLK(I2702), .RSTB(I602442), .Q(I602973) );
and I_35310 (I602407,I602880,I602973);
not I_35311 (I603037,I2709);
nand I_35312 (I603054,I485303,I485318);
and I_35313 (I603071,I603054,I485315);
DFFARX1 I_35314  ( .D(I603071), .CLK(I2702), .RSTB(I603037), .Q(I603088) );
nor I_35315 (I603105,I485291,I485318);
DFFARX1 I_35316  ( .D(I485309), .CLK(I2702), .RSTB(I603037), .Q(I603122) );
nand I_35317 (I603139,I603122,I603105);
DFFARX1 I_35318  ( .D(I603122), .CLK(I2702), .RSTB(I603037), .Q(I603008) );
nand I_35319 (I603170,I485312,I485300);
and I_35320 (I603187,I603170,I485306);
DFFARX1 I_35321  ( .D(I603187), .CLK(I2702), .RSTB(I603037), .Q(I603204) );
not I_35322 (I603221,I603204);
nor I_35323 (I603238,I603088,I603221);
and I_35324 (I603255,I603105,I603238);
and I_35325 (I603272,I603204,I603139);
DFFARX1 I_35326  ( .D(I603272), .CLK(I2702), .RSTB(I603037), .Q(I603005) );
DFFARX1 I_35327  ( .D(I603204), .CLK(I2702), .RSTB(I603037), .Q(I602999) );
DFFARX1 I_35328  ( .D(I485297), .CLK(I2702), .RSTB(I603037), .Q(I603317) );
and I_35329 (I603334,I603317,I485321);
nand I_35330 (I603351,I603334,I603204);
nor I_35331 (I603026,I603334,I603105);
not I_35332 (I603382,I603334);
nor I_35333 (I603399,I603088,I603382);
nand I_35334 (I603017,I603122,I603399);
nand I_35335 (I603011,I603204,I603382);
or I_35336 (I603444,I603334,I603255);
DFFARX1 I_35337  ( .D(I603444), .CLK(I2702), .RSTB(I603037), .Q(I603014) );
DFFARX1 I_35338  ( .D(I485294), .CLK(I2702), .RSTB(I603037), .Q(I603475) );
and I_35339 (I603492,I603475,I603351);
DFFARX1 I_35340  ( .D(I603492), .CLK(I2702), .RSTB(I603037), .Q(I603029) );
nor I_35341 (I603523,I603475,I603088);
nand I_35342 (I603023,I603334,I603523);
not I_35343 (I603020,I603475);
DFFARX1 I_35344  ( .D(I603475), .CLK(I2702), .RSTB(I603037), .Q(I603568) );
and I_35345 (I603002,I603475,I603568);
not I_35346 (I603632,I2709);
nand I_35347 (I603649,I506029,I506014);
and I_35348 (I603666,I603649,I506020);
DFFARX1 I_35349  ( .D(I603666), .CLK(I2702), .RSTB(I603632), .Q(I603683) );
nor I_35350 (I603700,I506023,I506014);
DFFARX1 I_35351  ( .D(I506035), .CLK(I2702), .RSTB(I603632), .Q(I603717) );
nand I_35352 (I603734,I603717,I603700);
DFFARX1 I_35353  ( .D(I603717), .CLK(I2702), .RSTB(I603632), .Q(I603603) );
nand I_35354 (I603765,I506026,I506017);
and I_35355 (I603782,I603765,I506044);
DFFARX1 I_35356  ( .D(I603782), .CLK(I2702), .RSTB(I603632), .Q(I603799) );
not I_35357 (I603816,I603799);
nor I_35358 (I603833,I603683,I603816);
and I_35359 (I603850,I603700,I603833);
and I_35360 (I603867,I603799,I603734);
DFFARX1 I_35361  ( .D(I603867), .CLK(I2702), .RSTB(I603632), .Q(I603600) );
DFFARX1 I_35362  ( .D(I603799), .CLK(I2702), .RSTB(I603632), .Q(I603594) );
DFFARX1 I_35363  ( .D(I506032), .CLK(I2702), .RSTB(I603632), .Q(I603912) );
and I_35364 (I603929,I603912,I506038);
nand I_35365 (I603946,I603929,I603799);
nor I_35366 (I603621,I603929,I603700);
not I_35367 (I603977,I603929);
nor I_35368 (I603994,I603683,I603977);
nand I_35369 (I603612,I603717,I603994);
nand I_35370 (I603606,I603799,I603977);
or I_35371 (I604039,I603929,I603850);
DFFARX1 I_35372  ( .D(I604039), .CLK(I2702), .RSTB(I603632), .Q(I603609) );
DFFARX1 I_35373  ( .D(I506041), .CLK(I2702), .RSTB(I603632), .Q(I604070) );
and I_35374 (I604087,I604070,I603946);
DFFARX1 I_35375  ( .D(I604087), .CLK(I2702), .RSTB(I603632), .Q(I603624) );
nor I_35376 (I604118,I604070,I603683);
nand I_35377 (I603618,I603929,I604118);
not I_35378 (I603615,I604070);
DFFARX1 I_35379  ( .D(I604070), .CLK(I2702), .RSTB(I603632), .Q(I604163) );
and I_35380 (I603597,I604070,I604163);
not I_35381 (I604227,I2709);
nand I_35382 (I604244,I637607,I637595);
and I_35383 (I604261,I604244,I637580);
DFFARX1 I_35384  ( .D(I604261), .CLK(I2702), .RSTB(I604227), .Q(I604278) );
nor I_35385 (I604295,I637592,I637595);
DFFARX1 I_35386  ( .D(I637604), .CLK(I2702), .RSTB(I604227), .Q(I604312) );
nand I_35387 (I604329,I604312,I604295);
DFFARX1 I_35388  ( .D(I604312), .CLK(I2702), .RSTB(I604227), .Q(I604198) );
nand I_35389 (I604360,I637577,I637601);
and I_35390 (I604377,I604360,I637586);
DFFARX1 I_35391  ( .D(I604377), .CLK(I2702), .RSTB(I604227), .Q(I604394) );
not I_35392 (I604411,I604394);
nor I_35393 (I604428,I604278,I604411);
and I_35394 (I604445,I604295,I604428);
and I_35395 (I604462,I604394,I604329);
DFFARX1 I_35396  ( .D(I604462), .CLK(I2702), .RSTB(I604227), .Q(I604195) );
DFFARX1 I_35397  ( .D(I604394), .CLK(I2702), .RSTB(I604227), .Q(I604189) );
DFFARX1 I_35398  ( .D(I637589), .CLK(I2702), .RSTB(I604227), .Q(I604507) );
and I_35399 (I604524,I604507,I637598);
nand I_35400 (I604541,I604524,I604394);
nor I_35401 (I604216,I604524,I604295);
not I_35402 (I604572,I604524);
nor I_35403 (I604589,I604278,I604572);
nand I_35404 (I604207,I604312,I604589);
nand I_35405 (I604201,I604394,I604572);
or I_35406 (I604634,I604524,I604445);
DFFARX1 I_35407  ( .D(I604634), .CLK(I2702), .RSTB(I604227), .Q(I604204) );
DFFARX1 I_35408  ( .D(I637583), .CLK(I2702), .RSTB(I604227), .Q(I604665) );
and I_35409 (I604682,I604665,I604541);
DFFARX1 I_35410  ( .D(I604682), .CLK(I2702), .RSTB(I604227), .Q(I604219) );
nor I_35411 (I604713,I604665,I604278);
nand I_35412 (I604213,I604524,I604713);
not I_35413 (I604210,I604665);
DFFARX1 I_35414  ( .D(I604665), .CLK(I2702), .RSTB(I604227), .Q(I604758) );
and I_35415 (I604192,I604665,I604758);
not I_35416 (I604822,I2709);
nand I_35417 (I604839,I532209,I532194);
and I_35418 (I604856,I604839,I532200);
DFFARX1 I_35419  ( .D(I604856), .CLK(I2702), .RSTB(I604822), .Q(I604873) );
nor I_35420 (I604890,I532203,I532194);
DFFARX1 I_35421  ( .D(I532215), .CLK(I2702), .RSTB(I604822), .Q(I604907) );
nand I_35422 (I604924,I604907,I604890);
DFFARX1 I_35423  ( .D(I604907), .CLK(I2702), .RSTB(I604822), .Q(I604793) );
nand I_35424 (I604955,I532206,I532197);
and I_35425 (I604972,I604955,I532224);
DFFARX1 I_35426  ( .D(I604972), .CLK(I2702), .RSTB(I604822), .Q(I604989) );
not I_35427 (I605006,I604989);
nor I_35428 (I605023,I604873,I605006);
and I_35429 (I605040,I604890,I605023);
and I_35430 (I605057,I604989,I604924);
DFFARX1 I_35431  ( .D(I605057), .CLK(I2702), .RSTB(I604822), .Q(I604790) );
DFFARX1 I_35432  ( .D(I604989), .CLK(I2702), .RSTB(I604822), .Q(I604784) );
DFFARX1 I_35433  ( .D(I532212), .CLK(I2702), .RSTB(I604822), .Q(I605102) );
and I_35434 (I605119,I605102,I532218);
nand I_35435 (I605136,I605119,I604989);
nor I_35436 (I604811,I605119,I604890);
not I_35437 (I605167,I605119);
nor I_35438 (I605184,I604873,I605167);
nand I_35439 (I604802,I604907,I605184);
nand I_35440 (I604796,I604989,I605167);
or I_35441 (I605229,I605119,I605040);
DFFARX1 I_35442  ( .D(I605229), .CLK(I2702), .RSTB(I604822), .Q(I604799) );
DFFARX1 I_35443  ( .D(I532221), .CLK(I2702), .RSTB(I604822), .Q(I605260) );
and I_35444 (I605277,I605260,I605136);
DFFARX1 I_35445  ( .D(I605277), .CLK(I2702), .RSTB(I604822), .Q(I604814) );
nor I_35446 (I605308,I605260,I604873);
nand I_35447 (I604808,I605119,I605308);
not I_35448 (I604805,I605260);
DFFARX1 I_35449  ( .D(I605260), .CLK(I2702), .RSTB(I604822), .Q(I605353) );
and I_35450 (I604787,I605260,I605353);
not I_35451 (I605417,I2709);
nand I_35452 (I605434,I655848,I655836);
and I_35453 (I605451,I605434,I655821);
DFFARX1 I_35454  ( .D(I605451), .CLK(I2702), .RSTB(I605417), .Q(I605468) );
nor I_35455 (I605485,I655833,I655836);
DFFARX1 I_35456  ( .D(I655845), .CLK(I2702), .RSTB(I605417), .Q(I605502) );
nand I_35457 (I605519,I605502,I605485);
DFFARX1 I_35458  ( .D(I605502), .CLK(I2702), .RSTB(I605417), .Q(I605388) );
nand I_35459 (I605550,I655818,I655842);
and I_35460 (I605567,I605550,I655827);
DFFARX1 I_35461  ( .D(I605567), .CLK(I2702), .RSTB(I605417), .Q(I605584) );
not I_35462 (I605601,I605584);
nor I_35463 (I605618,I605468,I605601);
and I_35464 (I605635,I605485,I605618);
and I_35465 (I605652,I605584,I605519);
DFFARX1 I_35466  ( .D(I605652), .CLK(I2702), .RSTB(I605417), .Q(I605385) );
DFFARX1 I_35467  ( .D(I605584), .CLK(I2702), .RSTB(I605417), .Q(I605379) );
DFFARX1 I_35468  ( .D(I655830), .CLK(I2702), .RSTB(I605417), .Q(I605697) );
and I_35469 (I605714,I605697,I655839);
nand I_35470 (I605731,I605714,I605584);
nor I_35471 (I605406,I605714,I605485);
not I_35472 (I605762,I605714);
nor I_35473 (I605779,I605468,I605762);
nand I_35474 (I605397,I605502,I605779);
nand I_35475 (I605391,I605584,I605762);
or I_35476 (I605824,I605714,I605635);
DFFARX1 I_35477  ( .D(I605824), .CLK(I2702), .RSTB(I605417), .Q(I605394) );
DFFARX1 I_35478  ( .D(I655824), .CLK(I2702), .RSTB(I605417), .Q(I605855) );
and I_35479 (I605872,I605855,I605731);
DFFARX1 I_35480  ( .D(I605872), .CLK(I2702), .RSTB(I605417), .Q(I605409) );
nor I_35481 (I605903,I605855,I605468);
nand I_35482 (I605403,I605714,I605903);
not I_35483 (I605400,I605855);
DFFARX1 I_35484  ( .D(I605855), .CLK(I2702), .RSTB(I605417), .Q(I605948) );
and I_35485 (I605382,I605855,I605948);
not I_35486 (I606012,I2709);
nand I_35487 (I606029,I563744,I563729);
and I_35488 (I606046,I606029,I563735);
DFFARX1 I_35489  ( .D(I606046), .CLK(I2702), .RSTB(I606012), .Q(I606063) );
nor I_35490 (I606080,I563738,I563729);
DFFARX1 I_35491  ( .D(I563750), .CLK(I2702), .RSTB(I606012), .Q(I606097) );
nand I_35492 (I606114,I606097,I606080);
DFFARX1 I_35493  ( .D(I606097), .CLK(I2702), .RSTB(I606012), .Q(I605983) );
nand I_35494 (I606145,I563741,I563732);
and I_35495 (I606162,I606145,I563759);
DFFARX1 I_35496  ( .D(I606162), .CLK(I2702), .RSTB(I606012), .Q(I606179) );
not I_35497 (I606196,I606179);
nor I_35498 (I606213,I606063,I606196);
and I_35499 (I606230,I606080,I606213);
and I_35500 (I606247,I606179,I606114);
DFFARX1 I_35501  ( .D(I606247), .CLK(I2702), .RSTB(I606012), .Q(I605980) );
DFFARX1 I_35502  ( .D(I606179), .CLK(I2702), .RSTB(I606012), .Q(I605974) );
DFFARX1 I_35503  ( .D(I563747), .CLK(I2702), .RSTB(I606012), .Q(I606292) );
and I_35504 (I606309,I606292,I563753);
nand I_35505 (I606326,I606309,I606179);
nor I_35506 (I606001,I606309,I606080);
not I_35507 (I606357,I606309);
nor I_35508 (I606374,I606063,I606357);
nand I_35509 (I605992,I606097,I606374);
nand I_35510 (I605986,I606179,I606357);
or I_35511 (I606419,I606309,I606230);
DFFARX1 I_35512  ( .D(I606419), .CLK(I2702), .RSTB(I606012), .Q(I605989) );
DFFARX1 I_35513  ( .D(I563756), .CLK(I2702), .RSTB(I606012), .Q(I606450) );
and I_35514 (I606467,I606450,I606326);
DFFARX1 I_35515  ( .D(I606467), .CLK(I2702), .RSTB(I606012), .Q(I606004) );
nor I_35516 (I606498,I606450,I606063);
nand I_35517 (I605998,I606309,I606498);
not I_35518 (I605995,I606450);
DFFARX1 I_35519  ( .D(I606450), .CLK(I2702), .RSTB(I606012), .Q(I606543) );
and I_35520 (I605977,I606450,I606543);
not I_35521 (I606607,I2709);
nand I_35522 (I606624,I526854,I526839);
and I_35523 (I606641,I606624,I526845);
DFFARX1 I_35524  ( .D(I606641), .CLK(I2702), .RSTB(I606607), .Q(I606658) );
nor I_35525 (I606675,I526848,I526839);
DFFARX1 I_35526  ( .D(I526860), .CLK(I2702), .RSTB(I606607), .Q(I606692) );
nand I_35527 (I606709,I606692,I606675);
DFFARX1 I_35528  ( .D(I606692), .CLK(I2702), .RSTB(I606607), .Q(I606578) );
nand I_35529 (I606740,I526851,I526842);
and I_35530 (I606757,I606740,I526869);
DFFARX1 I_35531  ( .D(I606757), .CLK(I2702), .RSTB(I606607), .Q(I606774) );
not I_35532 (I606791,I606774);
nor I_35533 (I606808,I606658,I606791);
and I_35534 (I606825,I606675,I606808);
and I_35535 (I606842,I606774,I606709);
DFFARX1 I_35536  ( .D(I606842), .CLK(I2702), .RSTB(I606607), .Q(I606575) );
DFFARX1 I_35537  ( .D(I606774), .CLK(I2702), .RSTB(I606607), .Q(I606569) );
DFFARX1 I_35538  ( .D(I526857), .CLK(I2702), .RSTB(I606607), .Q(I606887) );
and I_35539 (I606904,I606887,I526863);
nand I_35540 (I606921,I606904,I606774);
nor I_35541 (I606596,I606904,I606675);
not I_35542 (I606952,I606904);
nor I_35543 (I606969,I606658,I606952);
nand I_35544 (I606587,I606692,I606969);
nand I_35545 (I606581,I606774,I606952);
or I_35546 (I607014,I606904,I606825);
DFFARX1 I_35547  ( .D(I607014), .CLK(I2702), .RSTB(I606607), .Q(I606584) );
DFFARX1 I_35548  ( .D(I526866), .CLK(I2702), .RSTB(I606607), .Q(I607045) );
and I_35549 (I607062,I607045,I606921);
DFFARX1 I_35550  ( .D(I607062), .CLK(I2702), .RSTB(I606607), .Q(I606599) );
nor I_35551 (I607093,I607045,I606658);
nand I_35552 (I606593,I606904,I607093);
not I_35553 (I606590,I607045);
DFFARX1 I_35554  ( .D(I607045), .CLK(I2702), .RSTB(I606607), .Q(I607138) );
and I_35555 (I606572,I607045,I607138);
not I_35556 (I607202,I2709);
nand I_35557 (I607219,I58822,I58798);
and I_35558 (I607236,I607219,I58807);
DFFARX1 I_35559  ( .D(I607236), .CLK(I2702), .RSTB(I607202), .Q(I607253) );
nor I_35560 (I607270,I58801,I58798);
DFFARX1 I_35561  ( .D(I58816), .CLK(I2702), .RSTB(I607202), .Q(I607287) );
nand I_35562 (I607304,I607287,I607270);
DFFARX1 I_35563  ( .D(I607287), .CLK(I2702), .RSTB(I607202), .Q(I607173) );
nand I_35564 (I607335,I58810,I58825);
and I_35565 (I607352,I607335,I58804);
DFFARX1 I_35566  ( .D(I607352), .CLK(I2702), .RSTB(I607202), .Q(I607369) );
not I_35567 (I607386,I607369);
nor I_35568 (I607403,I607253,I607386);
and I_35569 (I607420,I607270,I607403);
and I_35570 (I607437,I607369,I607304);
DFFARX1 I_35571  ( .D(I607437), .CLK(I2702), .RSTB(I607202), .Q(I607170) );
DFFARX1 I_35572  ( .D(I607369), .CLK(I2702), .RSTB(I607202), .Q(I607164) );
DFFARX1 I_35573  ( .D(I58795), .CLK(I2702), .RSTB(I607202), .Q(I607482) );
and I_35574 (I607499,I607482,I58813);
nand I_35575 (I607516,I607499,I607369);
nor I_35576 (I607191,I607499,I607270);
not I_35577 (I607547,I607499);
nor I_35578 (I607564,I607253,I607547);
nand I_35579 (I607182,I607287,I607564);
nand I_35580 (I607176,I607369,I607547);
or I_35581 (I607609,I607499,I607420);
DFFARX1 I_35582  ( .D(I607609), .CLK(I2702), .RSTB(I607202), .Q(I607179) );
DFFARX1 I_35583  ( .D(I58819), .CLK(I2702), .RSTB(I607202), .Q(I607640) );
and I_35584 (I607657,I607640,I607516);
DFFARX1 I_35585  ( .D(I607657), .CLK(I2702), .RSTB(I607202), .Q(I607194) );
nor I_35586 (I607688,I607640,I607253);
nand I_35587 (I607188,I607499,I607688);
not I_35588 (I607185,I607640);
DFFARX1 I_35589  ( .D(I607640), .CLK(I2702), .RSTB(I607202), .Q(I607733) );
and I_35590 (I607167,I607640,I607733);
not I_35591 (I607797,I2709);
nand I_35592 (I607814,I571479,I571464);
and I_35593 (I607831,I607814,I571470);
DFFARX1 I_35594  ( .D(I607831), .CLK(I2702), .RSTB(I607797), .Q(I607848) );
nor I_35595 (I607865,I571473,I571464);
DFFARX1 I_35596  ( .D(I571485), .CLK(I2702), .RSTB(I607797), .Q(I607882) );
nand I_35597 (I607899,I607882,I607865);
DFFARX1 I_35598  ( .D(I607882), .CLK(I2702), .RSTB(I607797), .Q(I607768) );
nand I_35599 (I607930,I571476,I571467);
and I_35600 (I607947,I607930,I571494);
DFFARX1 I_35601  ( .D(I607947), .CLK(I2702), .RSTB(I607797), .Q(I607964) );
not I_35602 (I607981,I607964);
nor I_35603 (I607998,I607848,I607981);
and I_35604 (I608015,I607865,I607998);
and I_35605 (I608032,I607964,I607899);
DFFARX1 I_35606  ( .D(I608032), .CLK(I2702), .RSTB(I607797), .Q(I607765) );
DFFARX1 I_35607  ( .D(I607964), .CLK(I2702), .RSTB(I607797), .Q(I607759) );
DFFARX1 I_35608  ( .D(I571482), .CLK(I2702), .RSTB(I607797), .Q(I608077) );
and I_35609 (I608094,I608077,I571488);
nand I_35610 (I608111,I608094,I607964);
nor I_35611 (I607786,I608094,I607865);
not I_35612 (I608142,I608094);
nor I_35613 (I608159,I607848,I608142);
nand I_35614 (I607777,I607882,I608159);
nand I_35615 (I607771,I607964,I608142);
or I_35616 (I608204,I608094,I608015);
DFFARX1 I_35617  ( .D(I608204), .CLK(I2702), .RSTB(I607797), .Q(I607774) );
DFFARX1 I_35618  ( .D(I571491), .CLK(I2702), .RSTB(I607797), .Q(I608235) );
and I_35619 (I608252,I608235,I608111);
DFFARX1 I_35620  ( .D(I608252), .CLK(I2702), .RSTB(I607797), .Q(I607789) );
nor I_35621 (I608283,I608235,I607848);
nand I_35622 (I607783,I608094,I608283);
not I_35623 (I607780,I608235);
DFFARX1 I_35624  ( .D(I608235), .CLK(I2702), .RSTB(I607797), .Q(I608328) );
and I_35625 (I607762,I608235,I608328);
not I_35626 (I608392,I2709);
nand I_35627 (I608409,I229631,I229628);
and I_35628 (I608426,I608409,I229655);
DFFARX1 I_35629  ( .D(I608426), .CLK(I2702), .RSTB(I608392), .Q(I608443) );
nor I_35630 (I608460,I229658,I229628);
DFFARX1 I_35631  ( .D(I229646), .CLK(I2702), .RSTB(I608392), .Q(I608477) );
nand I_35632 (I608494,I608477,I608460);
DFFARX1 I_35633  ( .D(I608477), .CLK(I2702), .RSTB(I608392), .Q(I608363) );
nand I_35634 (I608525,I229652,I229637);
and I_35635 (I608542,I608525,I229643);
DFFARX1 I_35636  ( .D(I608542), .CLK(I2702), .RSTB(I608392), .Q(I608559) );
not I_35637 (I608576,I608559);
nor I_35638 (I608593,I608443,I608576);
and I_35639 (I608610,I608460,I608593);
and I_35640 (I608627,I608559,I608494);
DFFARX1 I_35641  ( .D(I608627), .CLK(I2702), .RSTB(I608392), .Q(I608360) );
DFFARX1 I_35642  ( .D(I608559), .CLK(I2702), .RSTB(I608392), .Q(I608354) );
DFFARX1 I_35643  ( .D(I229634), .CLK(I2702), .RSTB(I608392), .Q(I608672) );
and I_35644 (I608689,I608672,I229640);
nand I_35645 (I608706,I608689,I608559);
nor I_35646 (I608381,I608689,I608460);
not I_35647 (I608737,I608689);
nor I_35648 (I608754,I608443,I608737);
nand I_35649 (I608372,I608477,I608754);
nand I_35650 (I608366,I608559,I608737);
or I_35651 (I608799,I608689,I608610);
DFFARX1 I_35652  ( .D(I608799), .CLK(I2702), .RSTB(I608392), .Q(I608369) );
DFFARX1 I_35653  ( .D(I229649), .CLK(I2702), .RSTB(I608392), .Q(I608830) );
and I_35654 (I608847,I608830,I608706);
DFFARX1 I_35655  ( .D(I608847), .CLK(I2702), .RSTB(I608392), .Q(I608384) );
nor I_35656 (I608878,I608830,I608443);
nand I_35657 (I608378,I608689,I608878);
not I_35658 (I608375,I608830);
DFFARX1 I_35659  ( .D(I608830), .CLK(I2702), .RSTB(I608392), .Q(I608923) );
and I_35660 (I608357,I608830,I608923);
not I_35661 (I608987,I2709);
nand I_35662 (I609004,I294054,I294024);
and I_35663 (I609021,I609004,I294042);
DFFARX1 I_35664  ( .D(I609021), .CLK(I2702), .RSTB(I608987), .Q(I609038) );
nor I_35665 (I609055,I294036,I294024);
DFFARX1 I_35666  ( .D(I294033), .CLK(I2702), .RSTB(I608987), .Q(I609072) );
nand I_35667 (I609089,I609072,I609055);
DFFARX1 I_35668  ( .D(I609072), .CLK(I2702), .RSTB(I608987), .Q(I608958) );
nand I_35669 (I609120,I294027,I294030);
and I_35670 (I609137,I609120,I294048);
DFFARX1 I_35671  ( .D(I609137), .CLK(I2702), .RSTB(I608987), .Q(I609154) );
not I_35672 (I609171,I609154);
nor I_35673 (I609188,I609038,I609171);
and I_35674 (I609205,I609055,I609188);
and I_35675 (I609222,I609154,I609089);
DFFARX1 I_35676  ( .D(I609222), .CLK(I2702), .RSTB(I608987), .Q(I608955) );
DFFARX1 I_35677  ( .D(I609154), .CLK(I2702), .RSTB(I608987), .Q(I608949) );
DFFARX1 I_35678  ( .D(I294051), .CLK(I2702), .RSTB(I608987), .Q(I609267) );
and I_35679 (I609284,I609267,I294045);
nand I_35680 (I609301,I609284,I609154);
nor I_35681 (I608976,I609284,I609055);
not I_35682 (I609332,I609284);
nor I_35683 (I609349,I609038,I609332);
nand I_35684 (I608967,I609072,I609349);
nand I_35685 (I608961,I609154,I609332);
or I_35686 (I609394,I609284,I609205);
DFFARX1 I_35687  ( .D(I609394), .CLK(I2702), .RSTB(I608987), .Q(I608964) );
DFFARX1 I_35688  ( .D(I294039), .CLK(I2702), .RSTB(I608987), .Q(I609425) );
and I_35689 (I609442,I609425,I609301);
DFFARX1 I_35690  ( .D(I609442), .CLK(I2702), .RSTB(I608987), .Q(I608979) );
nor I_35691 (I609473,I609425,I609038);
nand I_35692 (I608973,I609284,I609473);
not I_35693 (I608970,I609425);
DFFARX1 I_35694  ( .D(I609425), .CLK(I2702), .RSTB(I608987), .Q(I609518) );
and I_35695 (I608952,I609425,I609518);
not I_35696 (I609582,I2709);
nand I_35697 (I609599,I541729,I541714);
and I_35698 (I609616,I609599,I541720);
DFFARX1 I_35699  ( .D(I609616), .CLK(I2702), .RSTB(I609582), .Q(I609633) );
nor I_35700 (I609650,I541723,I541714);
DFFARX1 I_35701  ( .D(I541735), .CLK(I2702), .RSTB(I609582), .Q(I609667) );
nand I_35702 (I609684,I609667,I609650);
DFFARX1 I_35703  ( .D(I609667), .CLK(I2702), .RSTB(I609582), .Q(I609553) );
nand I_35704 (I609715,I541726,I541717);
and I_35705 (I609732,I609715,I541744);
DFFARX1 I_35706  ( .D(I609732), .CLK(I2702), .RSTB(I609582), .Q(I609749) );
not I_35707 (I609766,I609749);
nor I_35708 (I609783,I609633,I609766);
and I_35709 (I609800,I609650,I609783);
and I_35710 (I609817,I609749,I609684);
DFFARX1 I_35711  ( .D(I609817), .CLK(I2702), .RSTB(I609582), .Q(I609550) );
DFFARX1 I_35712  ( .D(I609749), .CLK(I2702), .RSTB(I609582), .Q(I609544) );
DFFARX1 I_35713  ( .D(I541732), .CLK(I2702), .RSTB(I609582), .Q(I609862) );
and I_35714 (I609879,I609862,I541738);
nand I_35715 (I609896,I609879,I609749);
nor I_35716 (I609571,I609879,I609650);
not I_35717 (I609927,I609879);
nor I_35718 (I609944,I609633,I609927);
nand I_35719 (I609562,I609667,I609944);
nand I_35720 (I609556,I609749,I609927);
or I_35721 (I609989,I609879,I609800);
DFFARX1 I_35722  ( .D(I609989), .CLK(I2702), .RSTB(I609582), .Q(I609559) );
DFFARX1 I_35723  ( .D(I541741), .CLK(I2702), .RSTB(I609582), .Q(I610020) );
and I_35724 (I610037,I610020,I609896);
DFFARX1 I_35725  ( .D(I610037), .CLK(I2702), .RSTB(I609582), .Q(I609574) );
nor I_35726 (I610068,I610020,I609633);
nand I_35727 (I609568,I609879,I610068);
not I_35728 (I609565,I610020);
DFFARX1 I_35729  ( .D(I610020), .CLK(I2702), .RSTB(I609582), .Q(I610113) );
and I_35730 (I609547,I610020,I610113);
not I_35731 (I610177,I2709);
nand I_35732 (I610194,I677863,I677851);
and I_35733 (I610211,I610194,I677836);
DFFARX1 I_35734  ( .D(I610211), .CLK(I2702), .RSTB(I610177), .Q(I610228) );
nor I_35735 (I610245,I677848,I677851);
DFFARX1 I_35736  ( .D(I677860), .CLK(I2702), .RSTB(I610177), .Q(I610262) );
nand I_35737 (I610279,I610262,I610245);
DFFARX1 I_35738  ( .D(I610262), .CLK(I2702), .RSTB(I610177), .Q(I610148) );
nand I_35739 (I610310,I677833,I677857);
and I_35740 (I610327,I610310,I677842);
DFFARX1 I_35741  ( .D(I610327), .CLK(I2702), .RSTB(I610177), .Q(I610344) );
not I_35742 (I610361,I610344);
nor I_35743 (I610378,I610228,I610361);
and I_35744 (I610395,I610245,I610378);
and I_35745 (I610412,I610344,I610279);
DFFARX1 I_35746  ( .D(I610412), .CLK(I2702), .RSTB(I610177), .Q(I610145) );
DFFARX1 I_35747  ( .D(I610344), .CLK(I2702), .RSTB(I610177), .Q(I610139) );
DFFARX1 I_35748  ( .D(I677845), .CLK(I2702), .RSTB(I610177), .Q(I610457) );
and I_35749 (I610474,I610457,I677854);
nand I_35750 (I610491,I610474,I610344);
nor I_35751 (I610166,I610474,I610245);
not I_35752 (I610522,I610474);
nor I_35753 (I610539,I610228,I610522);
nand I_35754 (I610157,I610262,I610539);
nand I_35755 (I610151,I610344,I610522);
or I_35756 (I610584,I610474,I610395);
DFFARX1 I_35757  ( .D(I610584), .CLK(I2702), .RSTB(I610177), .Q(I610154) );
DFFARX1 I_35758  ( .D(I677839), .CLK(I2702), .RSTB(I610177), .Q(I610615) );
and I_35759 (I610632,I610615,I610491);
DFFARX1 I_35760  ( .D(I610632), .CLK(I2702), .RSTB(I610177), .Q(I610169) );
nor I_35761 (I610663,I610615,I610228);
nand I_35762 (I610163,I610474,I610663);
not I_35763 (I610160,I610615);
DFFARX1 I_35764  ( .D(I610615), .CLK(I2702), .RSTB(I610177), .Q(I610708) );
and I_35765 (I610142,I610615,I610708);
not I_35766 (I610772,I2709);
nand I_35767 (I610789,I226683,I226668);
and I_35768 (I610806,I610789,I226680);
DFFARX1 I_35769  ( .D(I610806), .CLK(I2702), .RSTB(I610772), .Q(I610823) );
nor I_35770 (I610840,I226671,I226668);
DFFARX1 I_35771  ( .D(I226662), .CLK(I2702), .RSTB(I610772), .Q(I610857) );
nand I_35772 (I610874,I610857,I610840);
DFFARX1 I_35773  ( .D(I610857), .CLK(I2702), .RSTB(I610772), .Q(I610743) );
nand I_35774 (I610905,I226653,I226677);
and I_35775 (I610922,I610905,I226656);
DFFARX1 I_35776  ( .D(I610922), .CLK(I2702), .RSTB(I610772), .Q(I610939) );
not I_35777 (I610956,I610939);
nor I_35778 (I610973,I610823,I610956);
and I_35779 (I610990,I610840,I610973);
and I_35780 (I611007,I610939,I610874);
DFFARX1 I_35781  ( .D(I611007), .CLK(I2702), .RSTB(I610772), .Q(I610740) );
DFFARX1 I_35782  ( .D(I610939), .CLK(I2702), .RSTB(I610772), .Q(I610734) );
DFFARX1 I_35783  ( .D(I226674), .CLK(I2702), .RSTB(I610772), .Q(I611052) );
and I_35784 (I611069,I611052,I226659);
nand I_35785 (I611086,I611069,I610939);
nor I_35786 (I610761,I611069,I610840);
not I_35787 (I611117,I611069);
nor I_35788 (I611134,I610823,I611117);
nand I_35789 (I610752,I610857,I611134);
nand I_35790 (I610746,I610939,I611117);
or I_35791 (I611179,I611069,I610990);
DFFARX1 I_35792  ( .D(I611179), .CLK(I2702), .RSTB(I610772), .Q(I610749) );
DFFARX1 I_35793  ( .D(I226665), .CLK(I2702), .RSTB(I610772), .Q(I611210) );
and I_35794 (I611227,I611210,I611086);
DFFARX1 I_35795  ( .D(I611227), .CLK(I2702), .RSTB(I610772), .Q(I610764) );
nor I_35796 (I611258,I611210,I610823);
nand I_35797 (I610758,I611069,I611258);
not I_35798 (I610755,I611210);
DFFARX1 I_35799  ( .D(I611210), .CLK(I2702), .RSTB(I610772), .Q(I611303) );
and I_35800 (I610737,I611210,I611303);
not I_35801 (I611367,I2709);
nand I_35802 (I611384,I182643,I182664);
and I_35803 (I611401,I611384,I182649);
DFFARX1 I_35804  ( .D(I611401), .CLK(I2702), .RSTB(I611367), .Q(I611418) );
nor I_35805 (I611435,I182667,I182664);
DFFARX1 I_35806  ( .D(I182670), .CLK(I2702), .RSTB(I611367), .Q(I611452) );
nand I_35807 (I611469,I611452,I611435);
DFFARX1 I_35808  ( .D(I611452), .CLK(I2702), .RSTB(I611367), .Q(I611338) );
nand I_35809 (I611500,I182640,I182652);
and I_35810 (I611517,I611500,I182661);
DFFARX1 I_35811  ( .D(I611517), .CLK(I2702), .RSTB(I611367), .Q(I611534) );
not I_35812 (I611551,I611534);
nor I_35813 (I611568,I611418,I611551);
and I_35814 (I611585,I611435,I611568);
and I_35815 (I611602,I611534,I611469);
DFFARX1 I_35816  ( .D(I611602), .CLK(I2702), .RSTB(I611367), .Q(I611335) );
DFFARX1 I_35817  ( .D(I611534), .CLK(I2702), .RSTB(I611367), .Q(I611329) );
DFFARX1 I_35818  ( .D(I182655), .CLK(I2702), .RSTB(I611367), .Q(I611647) );
and I_35819 (I611664,I611647,I182658);
nand I_35820 (I611681,I611664,I611534);
nor I_35821 (I611356,I611664,I611435);
not I_35822 (I611712,I611664);
nor I_35823 (I611729,I611418,I611712);
nand I_35824 (I611347,I611452,I611729);
nand I_35825 (I611341,I611534,I611712);
or I_35826 (I611774,I611664,I611585);
DFFARX1 I_35827  ( .D(I611774), .CLK(I2702), .RSTB(I611367), .Q(I611344) );
DFFARX1 I_35828  ( .D(I182646), .CLK(I2702), .RSTB(I611367), .Q(I611805) );
and I_35829 (I611822,I611805,I611681);
DFFARX1 I_35830  ( .D(I611822), .CLK(I2702), .RSTB(I611367), .Q(I611359) );
nor I_35831 (I611853,I611805,I611418);
nand I_35832 (I611353,I611664,I611853);
not I_35833 (I611350,I611805);
DFFARX1 I_35834  ( .D(I611805), .CLK(I2702), .RSTB(I611367), .Q(I611898) );
and I_35835 (I611332,I611805,I611898);
not I_35836 (I611962,I2709);
nand I_35837 (I611979,I122776,I122752);
and I_35838 (I611996,I611979,I122761);
DFFARX1 I_35839  ( .D(I611996), .CLK(I2702), .RSTB(I611962), .Q(I612013) );
nor I_35840 (I612030,I122755,I122752);
DFFARX1 I_35841  ( .D(I122770), .CLK(I2702), .RSTB(I611962), .Q(I612047) );
nand I_35842 (I612064,I612047,I612030);
DFFARX1 I_35843  ( .D(I612047), .CLK(I2702), .RSTB(I611962), .Q(I611933) );
nand I_35844 (I612095,I122764,I122779);
and I_35845 (I612112,I612095,I122758);
DFFARX1 I_35846  ( .D(I612112), .CLK(I2702), .RSTB(I611962), .Q(I612129) );
not I_35847 (I612146,I612129);
nor I_35848 (I612163,I612013,I612146);
and I_35849 (I612180,I612030,I612163);
and I_35850 (I612197,I612129,I612064);
DFFARX1 I_35851  ( .D(I612197), .CLK(I2702), .RSTB(I611962), .Q(I611930) );
DFFARX1 I_35852  ( .D(I612129), .CLK(I2702), .RSTB(I611962), .Q(I611924) );
DFFARX1 I_35853  ( .D(I122749), .CLK(I2702), .RSTB(I611962), .Q(I612242) );
and I_35854 (I612259,I612242,I122767);
nand I_35855 (I612276,I612259,I612129);
nor I_35856 (I611951,I612259,I612030);
not I_35857 (I612307,I612259);
nor I_35858 (I612324,I612013,I612307);
nand I_35859 (I611942,I612047,I612324);
nand I_35860 (I611936,I612129,I612307);
or I_35861 (I612369,I612259,I612180);
DFFARX1 I_35862  ( .D(I612369), .CLK(I2702), .RSTB(I611962), .Q(I611939) );
DFFARX1 I_35863  ( .D(I122773), .CLK(I2702), .RSTB(I611962), .Q(I612400) );
and I_35864 (I612417,I612400,I612276);
DFFARX1 I_35865  ( .D(I612417), .CLK(I2702), .RSTB(I611962), .Q(I611954) );
nor I_35866 (I612448,I612400,I612013);
nand I_35867 (I611948,I612259,I612448);
not I_35868 (I611945,I612400);
DFFARX1 I_35869  ( .D(I612400), .CLK(I2702), .RSTB(I611962), .Q(I612493) );
and I_35870 (I611927,I612400,I612493);
not I_35871 (I612557,I2709);
nand I_35872 (I612574,I200503,I200488);
and I_35873 (I612591,I612574,I200500);
DFFARX1 I_35874  ( .D(I612591), .CLK(I2702), .RSTB(I612557), .Q(I612608) );
nor I_35875 (I612625,I200491,I200488);
DFFARX1 I_35876  ( .D(I200482), .CLK(I2702), .RSTB(I612557), .Q(I612642) );
nand I_35877 (I612659,I612642,I612625);
DFFARX1 I_35878  ( .D(I612642), .CLK(I2702), .RSTB(I612557), .Q(I612528) );
nand I_35879 (I612690,I200473,I200497);
and I_35880 (I612707,I612690,I200476);
DFFARX1 I_35881  ( .D(I612707), .CLK(I2702), .RSTB(I612557), .Q(I612724) );
not I_35882 (I612741,I612724);
nor I_35883 (I612758,I612608,I612741);
and I_35884 (I612775,I612625,I612758);
and I_35885 (I612792,I612724,I612659);
DFFARX1 I_35886  ( .D(I612792), .CLK(I2702), .RSTB(I612557), .Q(I612525) );
DFFARX1 I_35887  ( .D(I612724), .CLK(I2702), .RSTB(I612557), .Q(I612519) );
DFFARX1 I_35888  ( .D(I200494), .CLK(I2702), .RSTB(I612557), .Q(I612837) );
and I_35889 (I612854,I612837,I200479);
nand I_35890 (I612871,I612854,I612724);
nor I_35891 (I612546,I612854,I612625);
not I_35892 (I612902,I612854);
nor I_35893 (I612919,I612608,I612902);
nand I_35894 (I612537,I612642,I612919);
nand I_35895 (I612531,I612724,I612902);
or I_35896 (I612964,I612854,I612775);
DFFARX1 I_35897  ( .D(I612964), .CLK(I2702), .RSTB(I612557), .Q(I612534) );
DFFARX1 I_35898  ( .D(I200485), .CLK(I2702), .RSTB(I612557), .Q(I612995) );
and I_35899 (I613012,I612995,I612871);
DFFARX1 I_35900  ( .D(I613012), .CLK(I2702), .RSTB(I612557), .Q(I612549) );
nor I_35901 (I613043,I612995,I612608);
nand I_35902 (I612543,I612854,I613043);
not I_35903 (I612540,I612995);
DFFARX1 I_35904  ( .D(I612995), .CLK(I2702), .RSTB(I612557), .Q(I613088) );
and I_35905 (I612522,I612995,I613088);
not I_35906 (I613152,I2709);
nand I_35907 (I613169,I461605,I461620);
and I_35908 (I613186,I613169,I461617);
DFFARX1 I_35909  ( .D(I613186), .CLK(I2702), .RSTB(I613152), .Q(I613203) );
nor I_35910 (I613220,I461593,I461620);
DFFARX1 I_35911  ( .D(I461611), .CLK(I2702), .RSTB(I613152), .Q(I613237) );
nand I_35912 (I613254,I613237,I613220);
DFFARX1 I_35913  ( .D(I613237), .CLK(I2702), .RSTB(I613152), .Q(I613123) );
nand I_35914 (I613285,I461614,I461602);
and I_35915 (I613302,I613285,I461608);
DFFARX1 I_35916  ( .D(I613302), .CLK(I2702), .RSTB(I613152), .Q(I613319) );
not I_35917 (I613336,I613319);
nor I_35918 (I613353,I613203,I613336);
and I_35919 (I613370,I613220,I613353);
and I_35920 (I613387,I613319,I613254);
DFFARX1 I_35921  ( .D(I613387), .CLK(I2702), .RSTB(I613152), .Q(I613120) );
DFFARX1 I_35922  ( .D(I613319), .CLK(I2702), .RSTB(I613152), .Q(I613114) );
DFFARX1 I_35923  ( .D(I461599), .CLK(I2702), .RSTB(I613152), .Q(I613432) );
and I_35924 (I613449,I613432,I461623);
nand I_35925 (I613466,I613449,I613319);
nor I_35926 (I613141,I613449,I613220);
not I_35927 (I613497,I613449);
nor I_35928 (I613514,I613203,I613497);
nand I_35929 (I613132,I613237,I613514);
nand I_35930 (I613126,I613319,I613497);
or I_35931 (I613559,I613449,I613370);
DFFARX1 I_35932  ( .D(I613559), .CLK(I2702), .RSTB(I613152), .Q(I613129) );
DFFARX1 I_35933  ( .D(I461596), .CLK(I2702), .RSTB(I613152), .Q(I613590) );
and I_35934 (I613607,I613590,I613466);
DFFARX1 I_35935  ( .D(I613607), .CLK(I2702), .RSTB(I613152), .Q(I613144) );
nor I_35936 (I613638,I613590,I613203);
nand I_35937 (I613138,I613449,I613638);
not I_35938 (I613135,I613590);
DFFARX1 I_35939  ( .D(I613590), .CLK(I2702), .RSTB(I613152), .Q(I613683) );
and I_35940 (I613117,I613590,I613683);
not I_35941 (I613747,I2709);
nand I_35942 (I613764,I29082,I29097);
and I_35943 (I613781,I613764,I29103);
DFFARX1 I_35944  ( .D(I613781), .CLK(I2702), .RSTB(I613747), .Q(I613798) );
nor I_35945 (I613815,I29091,I29097);
DFFARX1 I_35946  ( .D(I29079), .CLK(I2702), .RSTB(I613747), .Q(I613832) );
nand I_35947 (I613849,I613832,I613815);
DFFARX1 I_35948  ( .D(I613832), .CLK(I2702), .RSTB(I613747), .Q(I613718) );
nand I_35949 (I613880,I29085,I29088);
and I_35950 (I613897,I613880,I29094);
DFFARX1 I_35951  ( .D(I613897), .CLK(I2702), .RSTB(I613747), .Q(I613914) );
not I_35952 (I613931,I613914);
nor I_35953 (I613948,I613798,I613931);
and I_35954 (I613965,I613815,I613948);
and I_35955 (I613982,I613914,I613849);
DFFARX1 I_35956  ( .D(I613982), .CLK(I2702), .RSTB(I613747), .Q(I613715) );
DFFARX1 I_35957  ( .D(I613914), .CLK(I2702), .RSTB(I613747), .Q(I613709) );
DFFARX1 I_35958  ( .D(I29100), .CLK(I2702), .RSTB(I613747), .Q(I614027) );
and I_35959 (I614044,I614027,I29109);
nand I_35960 (I614061,I614044,I613914);
nor I_35961 (I613736,I614044,I613815);
not I_35962 (I614092,I614044);
nor I_35963 (I614109,I613798,I614092);
nand I_35964 (I613727,I613832,I614109);
nand I_35965 (I613721,I613914,I614092);
or I_35966 (I614154,I614044,I613965);
DFFARX1 I_35967  ( .D(I614154), .CLK(I2702), .RSTB(I613747), .Q(I613724) );
DFFARX1 I_35968  ( .D(I29106), .CLK(I2702), .RSTB(I613747), .Q(I614185) );
and I_35969 (I614202,I614185,I614061);
DFFARX1 I_35970  ( .D(I614202), .CLK(I2702), .RSTB(I613747), .Q(I613739) );
nor I_35971 (I614233,I614185,I613798);
nand I_35972 (I613733,I614044,I614233);
not I_35973 (I613730,I614185);
DFFARX1 I_35974  ( .D(I614185), .CLK(I2702), .RSTB(I613747), .Q(I614278) );
and I_35975 (I613712,I614185,I614278);
not I_35976 (I614342,I2709);
not I_35977 (I614359,I278130);
nor I_35978 (I614376,I278136,I278115);
nand I_35979 (I614393,I614376,I278121);
nor I_35980 (I614410,I614359,I278136);
nand I_35981 (I614427,I614410,I278127);
not I_35982 (I614444,I278136);
not I_35983 (I614461,I614444);
not I_35984 (I614478,I278124);
nor I_35985 (I614495,I614478,I278142);
and I_35986 (I614512,I614495,I278133);
or I_35987 (I614529,I614512,I278112);
DFFARX1 I_35988  ( .D(I614529), .CLK(I2702), .RSTB(I614342), .Q(I614546) );
nand I_35989 (I614563,I614359,I278124);
or I_35990 (I614331,I614563,I614546);
not I_35991 (I614594,I614563);
nor I_35992 (I614611,I614546,I614594);
and I_35993 (I614628,I614444,I614611);
nand I_35994 (I614304,I614563,I614461);
DFFARX1 I_35995  ( .D(I278139), .CLK(I2702), .RSTB(I614342), .Q(I614659) );
or I_35996 (I614325,I614659,I614546);
nor I_35997 (I614690,I614659,I614427);
nor I_35998 (I614707,I614659,I614461);
nand I_35999 (I614310,I614393,I614707);
or I_36000 (I614738,I614659,I614628);
DFFARX1 I_36001  ( .D(I614738), .CLK(I2702), .RSTB(I614342), .Q(I614307) );
not I_36002 (I614313,I614659);
DFFARX1 I_36003  ( .D(I278118), .CLK(I2702), .RSTB(I614342), .Q(I614783) );
not I_36004 (I614800,I614783);
nor I_36005 (I614817,I614800,I614393);
DFFARX1 I_36006  ( .D(I614817), .CLK(I2702), .RSTB(I614342), .Q(I614319) );
nor I_36007 (I614334,I614659,I614800);
nor I_36008 (I614322,I614800,I614563);
not I_36009 (I614876,I614800);
and I_36010 (I614893,I614427,I614876);
nor I_36011 (I614328,I614563,I614893);
nand I_36012 (I614316,I614800,I614690);
not I_36013 (I614971,I2709);
not I_36014 (I614988,I539935);
nor I_36015 (I615005,I539953,I539932);
nand I_36016 (I615022,I615005,I539956);
nor I_36017 (I615039,I614988,I539953);
nand I_36018 (I615056,I615039,I539950);
not I_36019 (I615073,I539953);
not I_36020 (I615090,I615073);
not I_36021 (I615107,I539941);
nor I_36022 (I615124,I615107,I539929);
and I_36023 (I615141,I615124,I539947);
or I_36024 (I615158,I615141,I539959);
DFFARX1 I_36025  ( .D(I615158), .CLK(I2702), .RSTB(I614971), .Q(I615175) );
nand I_36026 (I615192,I614988,I539941);
or I_36027 (I614960,I615192,I615175);
not I_36028 (I615223,I615192);
nor I_36029 (I615240,I615175,I615223);
and I_36030 (I615257,I615073,I615240);
nand I_36031 (I614933,I615192,I615090);
DFFARX1 I_36032  ( .D(I539938), .CLK(I2702), .RSTB(I614971), .Q(I615288) );
or I_36033 (I614954,I615288,I615175);
nor I_36034 (I615319,I615288,I615056);
nor I_36035 (I615336,I615288,I615090);
nand I_36036 (I614939,I615022,I615336);
or I_36037 (I615367,I615288,I615257);
DFFARX1 I_36038  ( .D(I615367), .CLK(I2702), .RSTB(I614971), .Q(I614936) );
not I_36039 (I614942,I615288);
DFFARX1 I_36040  ( .D(I539944), .CLK(I2702), .RSTB(I614971), .Q(I615412) );
not I_36041 (I615429,I615412);
nor I_36042 (I615446,I615429,I615022);
DFFARX1 I_36043  ( .D(I615446), .CLK(I2702), .RSTB(I614971), .Q(I614948) );
nor I_36044 (I614963,I615288,I615429);
nor I_36045 (I614951,I615429,I615192);
not I_36046 (I615505,I615429);
and I_36047 (I615522,I615056,I615505);
nor I_36048 (I614957,I615192,I615522);
nand I_36049 (I614945,I615429,I615319);
not I_36050 (I615600,I2709);
not I_36051 (I615617,I194586);
nor I_36052 (I615634,I194577,I194601);
nand I_36053 (I615651,I615634,I194604);
nor I_36054 (I615668,I615617,I194577);
nand I_36055 (I615685,I615668,I194595);
not I_36056 (I615702,I194577);
not I_36057 (I615719,I615702);
not I_36058 (I615736,I194589);
nor I_36059 (I615753,I615736,I194583);
and I_36060 (I615770,I615753,I194592);
or I_36061 (I615787,I615770,I194580);
DFFARX1 I_36062  ( .D(I615787), .CLK(I2702), .RSTB(I615600), .Q(I615804) );
nand I_36063 (I615821,I615617,I194589);
or I_36064 (I615589,I615821,I615804);
not I_36065 (I615852,I615821);
nor I_36066 (I615869,I615804,I615852);
and I_36067 (I615886,I615702,I615869);
nand I_36068 (I615562,I615821,I615719);
DFFARX1 I_36069  ( .D(I194574), .CLK(I2702), .RSTB(I615600), .Q(I615917) );
or I_36070 (I615583,I615917,I615804);
nor I_36071 (I615948,I615917,I615685);
nor I_36072 (I615965,I615917,I615719);
nand I_36073 (I615568,I615651,I615965);
or I_36074 (I615996,I615917,I615886);
DFFARX1 I_36075  ( .D(I615996), .CLK(I2702), .RSTB(I615600), .Q(I615565) );
not I_36076 (I615571,I615917);
DFFARX1 I_36077  ( .D(I194598), .CLK(I2702), .RSTB(I615600), .Q(I616041) );
not I_36078 (I616058,I616041);
nor I_36079 (I616075,I616058,I615651);
DFFARX1 I_36080  ( .D(I616075), .CLK(I2702), .RSTB(I615600), .Q(I615577) );
nor I_36081 (I615592,I615917,I616058);
nor I_36082 (I615580,I616058,I615821);
not I_36083 (I616134,I616058);
and I_36084 (I616151,I615685,I616134);
nor I_36085 (I615586,I615821,I616151);
nand I_36086 (I615574,I616058,I615948);
not I_36087 (I616229,I2709);
not I_36088 (I616246,I307965);
nor I_36089 (I616263,I307971,I307950);
nand I_36090 (I616280,I616263,I307956);
nor I_36091 (I616297,I616246,I307971);
nand I_36092 (I616314,I616297,I307962);
not I_36093 (I616331,I307971);
not I_36094 (I616348,I616331);
not I_36095 (I616365,I307959);
nor I_36096 (I616382,I616365,I307977);
and I_36097 (I616399,I616382,I307968);
or I_36098 (I616416,I616399,I307947);
DFFARX1 I_36099  ( .D(I616416), .CLK(I2702), .RSTB(I616229), .Q(I616433) );
nand I_36100 (I616450,I616246,I307959);
or I_36101 (I616218,I616450,I616433);
not I_36102 (I616481,I616450);
nor I_36103 (I616498,I616433,I616481);
and I_36104 (I616515,I616331,I616498);
nand I_36105 (I616191,I616450,I616348);
DFFARX1 I_36106  ( .D(I307974), .CLK(I2702), .RSTB(I616229), .Q(I616546) );
or I_36107 (I616212,I616546,I616433);
nor I_36108 (I616577,I616546,I616314);
nor I_36109 (I616594,I616546,I616348);
nand I_36110 (I616197,I616280,I616594);
or I_36111 (I616625,I616546,I616515);
DFFARX1 I_36112  ( .D(I616625), .CLK(I2702), .RSTB(I616229), .Q(I616194) );
not I_36113 (I616200,I616546);
DFFARX1 I_36114  ( .D(I307953), .CLK(I2702), .RSTB(I616229), .Q(I616670) );
not I_36115 (I616687,I616670);
nor I_36116 (I616704,I616687,I616280);
DFFARX1 I_36117  ( .D(I616704), .CLK(I2702), .RSTB(I616229), .Q(I616206) );
nor I_36118 (I616221,I616546,I616687);
nor I_36119 (I616209,I616687,I616450);
not I_36120 (I616763,I616687);
and I_36121 (I616780,I616314,I616763);
nor I_36122 (I616215,I616450,I616780);
nand I_36123 (I616203,I616687,I616577);
not I_36124 (I616858,I2709);
not I_36125 (I616875,I274152);
nor I_36126 (I616892,I274158,I274137);
nand I_36127 (I616909,I616892,I274143);
nor I_36128 (I616926,I616875,I274158);
nand I_36129 (I616943,I616926,I274149);
not I_36130 (I616960,I274158);
not I_36131 (I616977,I616960);
not I_36132 (I616994,I274146);
nor I_36133 (I617011,I616994,I274164);
and I_36134 (I617028,I617011,I274155);
or I_36135 (I617045,I617028,I274134);
DFFARX1 I_36136  ( .D(I617045), .CLK(I2702), .RSTB(I616858), .Q(I617062) );
nand I_36137 (I617079,I616875,I274146);
or I_36138 (I616847,I617079,I617062);
not I_36139 (I617110,I617079);
nor I_36140 (I617127,I617062,I617110);
and I_36141 (I617144,I616960,I617127);
nand I_36142 (I616820,I617079,I616977);
DFFARX1 I_36143  ( .D(I274161), .CLK(I2702), .RSTB(I616858), .Q(I617175) );
or I_36144 (I616841,I617175,I617062);
nor I_36145 (I617206,I617175,I616943);
nor I_36146 (I617223,I617175,I616977);
nand I_36147 (I616826,I616909,I617223);
or I_36148 (I617254,I617175,I617144);
DFFARX1 I_36149  ( .D(I617254), .CLK(I2702), .RSTB(I616858), .Q(I616823) );
not I_36150 (I616829,I617175);
DFFARX1 I_36151  ( .D(I274140), .CLK(I2702), .RSTB(I616858), .Q(I617299) );
not I_36152 (I617316,I617299);
nor I_36153 (I617333,I617316,I616909);
DFFARX1 I_36154  ( .D(I617333), .CLK(I2702), .RSTB(I616858), .Q(I616835) );
nor I_36155 (I616850,I617175,I617316);
nor I_36156 (I616838,I617316,I617079);
not I_36157 (I617392,I617316);
and I_36158 (I617409,I616943,I617392);
nor I_36159 (I616844,I617079,I617409);
nand I_36160 (I616832,I617316,I617206);
not I_36161 (I617487,I2709);
not I_36162 (I617504,I51695);
nor I_36163 (I617521,I51713,I51692);
nand I_36164 (I617538,I617521,I51710);
nor I_36165 (I617555,I617504,I51713);
nand I_36166 (I617572,I617555,I51704);
not I_36167 (I617589,I51713);
not I_36168 (I617606,I617589);
not I_36169 (I617623,I51707);
nor I_36170 (I617640,I617623,I51701);
and I_36171 (I617657,I617640,I51698);
or I_36172 (I617674,I617657,I51689);
DFFARX1 I_36173  ( .D(I617674), .CLK(I2702), .RSTB(I617487), .Q(I617691) );
nand I_36174 (I617708,I617504,I51707);
or I_36175 (I617476,I617708,I617691);
not I_36176 (I617739,I617708);
nor I_36177 (I617756,I617691,I617739);
and I_36178 (I617773,I617589,I617756);
nand I_36179 (I617449,I617708,I617606);
DFFARX1 I_36180  ( .D(I51719), .CLK(I2702), .RSTB(I617487), .Q(I617804) );
or I_36181 (I617470,I617804,I617691);
nor I_36182 (I617835,I617804,I617572);
nor I_36183 (I617852,I617804,I617606);
nand I_36184 (I617455,I617538,I617852);
or I_36185 (I617883,I617804,I617773);
DFFARX1 I_36186  ( .D(I617883), .CLK(I2702), .RSTB(I617487), .Q(I617452) );
not I_36187 (I617458,I617804);
DFFARX1 I_36188  ( .D(I51716), .CLK(I2702), .RSTB(I617487), .Q(I617928) );
not I_36189 (I617945,I617928);
nor I_36190 (I617962,I617945,I617538);
DFFARX1 I_36191  ( .D(I617962), .CLK(I2702), .RSTB(I617487), .Q(I617464) );
nor I_36192 (I617479,I617804,I617945);
nor I_36193 (I617467,I617945,I617708);
not I_36194 (I618021,I617945);
and I_36195 (I618038,I617572,I618021);
nor I_36196 (I617473,I617708,I618038);
nand I_36197 (I617461,I617945,I617835);
not I_36198 (I618116,I2709);
not I_36199 (I618133,I210618);
nor I_36200 (I618150,I210594,I210609);
nand I_36201 (I618167,I618150,I210591);
nor I_36202 (I618184,I618133,I210594);
nand I_36203 (I618201,I618184,I210606);
not I_36204 (I618218,I210594);
not I_36205 (I618235,I618218);
not I_36206 (I618252,I210597);
nor I_36207 (I618269,I618252,I210612);
and I_36208 (I618286,I618269,I210603);
or I_36209 (I618303,I618286,I210588);
DFFARX1 I_36210  ( .D(I618303), .CLK(I2702), .RSTB(I618116), .Q(I618320) );
nand I_36211 (I618337,I618133,I210597);
or I_36212 (I618105,I618337,I618320);
not I_36213 (I618368,I618337);
nor I_36214 (I618385,I618320,I618368);
and I_36215 (I618402,I618218,I618385);
nand I_36216 (I618078,I618337,I618235);
DFFARX1 I_36217  ( .D(I210600), .CLK(I2702), .RSTB(I618116), .Q(I618433) );
or I_36218 (I618099,I618433,I618320);
nor I_36219 (I618464,I618433,I618201);
nor I_36220 (I618481,I618433,I618235);
nand I_36221 (I618084,I618167,I618481);
or I_36222 (I618512,I618433,I618402);
DFFARX1 I_36223  ( .D(I618512), .CLK(I2702), .RSTB(I618116), .Q(I618081) );
not I_36224 (I618087,I618433);
DFFARX1 I_36225  ( .D(I210615), .CLK(I2702), .RSTB(I618116), .Q(I618557) );
not I_36226 (I618574,I618557);
nor I_36227 (I618591,I618574,I618167);
DFFARX1 I_36228  ( .D(I618591), .CLK(I2702), .RSTB(I618116), .Q(I618093) );
nor I_36229 (I618108,I618433,I618574);
nor I_36230 (I618096,I618574,I618337);
not I_36231 (I618650,I618574);
and I_36232 (I618667,I618201,I618650);
nor I_36233 (I618102,I618337,I618667);
nand I_36234 (I618090,I618574,I618464);
not I_36235 (I618745,I2709);
not I_36236 (I618762,I574445);
nor I_36237 (I618779,I574463,I574442);
nand I_36238 (I618796,I618779,I574466);
nor I_36239 (I618813,I618762,I574463);
nand I_36240 (I618830,I618813,I574460);
not I_36241 (I618847,I574463);
not I_36242 (I618864,I618847);
not I_36243 (I618881,I574451);
nor I_36244 (I618898,I618881,I574439);
and I_36245 (I618915,I618898,I574457);
or I_36246 (I618932,I618915,I574469);
DFFARX1 I_36247  ( .D(I618932), .CLK(I2702), .RSTB(I618745), .Q(I618949) );
nand I_36248 (I618966,I618762,I574451);
or I_36249 (I618734,I618966,I618949);
not I_36250 (I618997,I618966);
nor I_36251 (I619014,I618949,I618997);
and I_36252 (I619031,I618847,I619014);
nand I_36253 (I618707,I618966,I618864);
DFFARX1 I_36254  ( .D(I574448), .CLK(I2702), .RSTB(I618745), .Q(I619062) );
or I_36255 (I618728,I619062,I618949);
nor I_36256 (I619093,I619062,I618830);
nor I_36257 (I619110,I619062,I618864);
nand I_36258 (I618713,I618796,I619110);
or I_36259 (I619141,I619062,I619031);
DFFARX1 I_36260  ( .D(I619141), .CLK(I2702), .RSTB(I618745), .Q(I618710) );
not I_36261 (I618716,I619062);
DFFARX1 I_36262  ( .D(I574454), .CLK(I2702), .RSTB(I618745), .Q(I619186) );
not I_36263 (I619203,I619186);
nor I_36264 (I619220,I619203,I618796);
DFFARX1 I_36265  ( .D(I619220), .CLK(I2702), .RSTB(I618745), .Q(I618722) );
nor I_36266 (I618737,I619062,I619203);
nor I_36267 (I618725,I619203,I618966);
not I_36268 (I619279,I619203);
and I_36269 (I619296,I618830,I619279);
nor I_36270 (I618731,I618966,I619296);
nand I_36271 (I618719,I619203,I619093);
not I_36272 (I619374,I2709);
not I_36273 (I619391,I722158);
nor I_36274 (I619408,I722182,I722167);
nand I_36275 (I619425,I619408,I722152);
nor I_36276 (I619442,I619391,I722182);
nand I_36277 (I619459,I619442,I722179);
not I_36278 (I619476,I722182);
not I_36279 (I619493,I619476);
not I_36280 (I619510,I722161);
nor I_36281 (I619527,I619510,I722155);
and I_36282 (I619544,I619527,I722176);
or I_36283 (I619561,I619544,I722164);
DFFARX1 I_36284  ( .D(I619561), .CLK(I2702), .RSTB(I619374), .Q(I619578) );
nand I_36285 (I619595,I619391,I722161);
or I_36286 (I619363,I619595,I619578);
not I_36287 (I619626,I619595);
nor I_36288 (I619643,I619578,I619626);
and I_36289 (I619660,I619476,I619643);
nand I_36290 (I619336,I619595,I619493);
DFFARX1 I_36291  ( .D(I722173), .CLK(I2702), .RSTB(I619374), .Q(I619691) );
or I_36292 (I619357,I619691,I619578);
nor I_36293 (I619722,I619691,I619459);
nor I_36294 (I619739,I619691,I619493);
nand I_36295 (I619342,I619425,I619739);
or I_36296 (I619770,I619691,I619660);
DFFARX1 I_36297  ( .D(I619770), .CLK(I2702), .RSTB(I619374), .Q(I619339) );
not I_36298 (I619345,I619691);
DFFARX1 I_36299  ( .D(I722170), .CLK(I2702), .RSTB(I619374), .Q(I619815) );
not I_36300 (I619832,I619815);
nor I_36301 (I619849,I619832,I619425);
DFFARX1 I_36302  ( .D(I619849), .CLK(I2702), .RSTB(I619374), .Q(I619351) );
nor I_36303 (I619366,I619691,I619832);
nor I_36304 (I619354,I619832,I619595);
not I_36305 (I619908,I619832);
and I_36306 (I619925,I619459,I619908);
nor I_36307 (I619360,I619595,I619925);
nand I_36308 (I619348,I619832,I619722);
not I_36309 (I620003,I2709);
not I_36310 (I620020,I575635);
nor I_36311 (I620037,I575653,I575632);
nand I_36312 (I620054,I620037,I575656);
nor I_36313 (I620071,I620020,I575653);
nand I_36314 (I620088,I620071,I575650);
not I_36315 (I620105,I575653);
not I_36316 (I620122,I620105);
not I_36317 (I620139,I575641);
nor I_36318 (I620156,I620139,I575629);
and I_36319 (I620173,I620156,I575647);
or I_36320 (I620190,I620173,I575659);
DFFARX1 I_36321  ( .D(I620190), .CLK(I2702), .RSTB(I620003), .Q(I620207) );
nand I_36322 (I620224,I620020,I575641);
or I_36323 (I619992,I620224,I620207);
not I_36324 (I620255,I620224);
nor I_36325 (I620272,I620207,I620255);
and I_36326 (I620289,I620105,I620272);
nand I_36327 (I619965,I620224,I620122);
DFFARX1 I_36328  ( .D(I575638), .CLK(I2702), .RSTB(I620003), .Q(I620320) );
or I_36329 (I619986,I620320,I620207);
nor I_36330 (I620351,I620320,I620088);
nor I_36331 (I620368,I620320,I620122);
nand I_36332 (I619971,I620054,I620368);
or I_36333 (I620399,I620320,I620289);
DFFARX1 I_36334  ( .D(I620399), .CLK(I2702), .RSTB(I620003), .Q(I619968) );
not I_36335 (I619974,I620320);
DFFARX1 I_36336  ( .D(I575644), .CLK(I2702), .RSTB(I620003), .Q(I620444) );
not I_36337 (I620461,I620444);
nor I_36338 (I620478,I620461,I620054);
DFFARX1 I_36339  ( .D(I620478), .CLK(I2702), .RSTB(I620003), .Q(I619980) );
nor I_36340 (I619995,I620320,I620461);
nor I_36341 (I619983,I620461,I620224);
not I_36342 (I620537,I620461);
and I_36343 (I620554,I620088,I620537);
nor I_36344 (I619989,I620224,I620554);
nand I_36345 (I619977,I620461,I620351);
not I_36346 (I620632,I2709);
not I_36347 (I620649,I542315);
nor I_36348 (I620666,I542333,I542312);
nand I_36349 (I620683,I620666,I542336);
nor I_36350 (I620700,I620649,I542333);
nand I_36351 (I620717,I620700,I542330);
not I_36352 (I620734,I542333);
not I_36353 (I620751,I620734);
not I_36354 (I620768,I542321);
nor I_36355 (I620785,I620768,I542309);
and I_36356 (I620802,I620785,I542327);
or I_36357 (I620819,I620802,I542339);
DFFARX1 I_36358  ( .D(I620819), .CLK(I2702), .RSTB(I620632), .Q(I620836) );
nand I_36359 (I620853,I620649,I542321);
or I_36360 (I620621,I620853,I620836);
not I_36361 (I620884,I620853);
nor I_36362 (I620901,I620836,I620884);
and I_36363 (I620918,I620734,I620901);
nand I_36364 (I620594,I620853,I620751);
DFFARX1 I_36365  ( .D(I542318), .CLK(I2702), .RSTB(I620632), .Q(I620949) );
or I_36366 (I620615,I620949,I620836);
nor I_36367 (I620980,I620949,I620717);
nor I_36368 (I620997,I620949,I620751);
nand I_36369 (I620600,I620683,I620997);
or I_36370 (I621028,I620949,I620918);
DFFARX1 I_36371  ( .D(I621028), .CLK(I2702), .RSTB(I620632), .Q(I620597) );
not I_36372 (I620603,I620949);
DFFARX1 I_36373  ( .D(I542324), .CLK(I2702), .RSTB(I620632), .Q(I621073) );
not I_36374 (I621090,I621073);
nor I_36375 (I621107,I621090,I620683);
DFFARX1 I_36376  ( .D(I621107), .CLK(I2702), .RSTB(I620632), .Q(I620609) );
nor I_36377 (I620624,I620949,I621090);
nor I_36378 (I620612,I621090,I620853);
not I_36379 (I621166,I621090);
and I_36380 (I621183,I620717,I621166);
nor I_36381 (I620618,I620853,I621183);
nand I_36382 (I620606,I621090,I620980);
not I_36383 (I621261,I2709);
not I_36384 (I621278,I561950);
nor I_36385 (I621295,I561968,I561947);
nand I_36386 (I621312,I621295,I561971);
nor I_36387 (I621329,I621278,I561968);
nand I_36388 (I621346,I621329,I561965);
not I_36389 (I621363,I561968);
not I_36390 (I621380,I621363);
not I_36391 (I621397,I561956);
nor I_36392 (I621414,I621397,I561944);
and I_36393 (I621431,I621414,I561962);
or I_36394 (I621448,I621431,I561974);
DFFARX1 I_36395  ( .D(I621448), .CLK(I2702), .RSTB(I621261), .Q(I621465) );
nand I_36396 (I621482,I621278,I561956);
or I_36397 (I621250,I621482,I621465);
not I_36398 (I621513,I621482);
nor I_36399 (I621530,I621465,I621513);
and I_36400 (I621547,I621363,I621530);
nand I_36401 (I621223,I621482,I621380);
DFFARX1 I_36402  ( .D(I561953), .CLK(I2702), .RSTB(I621261), .Q(I621578) );
or I_36403 (I621244,I621578,I621465);
nor I_36404 (I621609,I621578,I621346);
nor I_36405 (I621626,I621578,I621380);
nand I_36406 (I621229,I621312,I621626);
or I_36407 (I621657,I621578,I621547);
DFFARX1 I_36408  ( .D(I621657), .CLK(I2702), .RSTB(I621261), .Q(I621226) );
not I_36409 (I621232,I621578);
DFFARX1 I_36410  ( .D(I561959), .CLK(I2702), .RSTB(I621261), .Q(I621702) );
not I_36411 (I621719,I621702);
nor I_36412 (I621736,I621719,I621312);
DFFARX1 I_36413  ( .D(I621736), .CLK(I2702), .RSTB(I621261), .Q(I621238) );
nor I_36414 (I621253,I621578,I621719);
nor I_36415 (I621241,I621719,I621482);
not I_36416 (I621795,I621719);
and I_36417 (I621812,I621346,I621795);
nor I_36418 (I621247,I621482,I621812);
nand I_36419 (I621235,I621719,I621609);
not I_36420 (I621890,I2709);
not I_36421 (I621907,I113711);
nor I_36422 (I621924,I113729,I113708);
nand I_36423 (I621941,I621924,I113726);
nor I_36424 (I621958,I621907,I113729);
nand I_36425 (I621975,I621958,I113720);
not I_36426 (I621992,I113729);
not I_36427 (I622009,I621992);
not I_36428 (I622026,I113723);
nor I_36429 (I622043,I622026,I113717);
and I_36430 (I622060,I622043,I113714);
or I_36431 (I622077,I622060,I113705);
DFFARX1 I_36432  ( .D(I622077), .CLK(I2702), .RSTB(I621890), .Q(I622094) );
nand I_36433 (I622111,I621907,I113723);
or I_36434 (I621879,I622111,I622094);
not I_36435 (I622142,I622111);
nor I_36436 (I622159,I622094,I622142);
and I_36437 (I622176,I621992,I622159);
nand I_36438 (I621852,I622111,I622009);
DFFARX1 I_36439  ( .D(I113735), .CLK(I2702), .RSTB(I621890), .Q(I622207) );
or I_36440 (I621873,I622207,I622094);
nor I_36441 (I622238,I622207,I621975);
nor I_36442 (I622255,I622207,I622009);
nand I_36443 (I621858,I621941,I622255);
or I_36444 (I622286,I622207,I622176);
DFFARX1 I_36445  ( .D(I622286), .CLK(I2702), .RSTB(I621890), .Q(I621855) );
not I_36446 (I621861,I622207);
DFFARX1 I_36447  ( .D(I113732), .CLK(I2702), .RSTB(I621890), .Q(I622331) );
not I_36448 (I622348,I622331);
nor I_36449 (I622365,I622348,I621941);
DFFARX1 I_36450  ( .D(I622365), .CLK(I2702), .RSTB(I621890), .Q(I621867) );
nor I_36451 (I621882,I622207,I622348);
nor I_36452 (I621870,I622348,I622111);
not I_36453 (I622424,I622348);
and I_36454 (I622441,I621975,I622424);
nor I_36455 (I621876,I622111,I622441);
nand I_36456 (I621864,I622348,I622238);
not I_36457 (I622519,I2709);
not I_36458 (I622536,I442549);
nor I_36459 (I622553,I442522,I442540);
nand I_36460 (I622570,I622553,I442525);
nor I_36461 (I622587,I622536,I442522);
nand I_36462 (I622604,I622587,I442543);
not I_36463 (I622621,I442522);
not I_36464 (I622638,I622621);
not I_36465 (I622655,I442519);
nor I_36466 (I622672,I622655,I442546);
and I_36467 (I622689,I622672,I442537);
or I_36468 (I622706,I622689,I442528);
DFFARX1 I_36469  ( .D(I622706), .CLK(I2702), .RSTB(I622519), .Q(I622723) );
nand I_36470 (I622740,I622536,I442519);
or I_36471 (I622508,I622740,I622723);
not I_36472 (I622771,I622740);
nor I_36473 (I622788,I622723,I622771);
and I_36474 (I622805,I622621,I622788);
nand I_36475 (I622481,I622740,I622638);
DFFARX1 I_36476  ( .D(I442531), .CLK(I2702), .RSTB(I622519), .Q(I622836) );
or I_36477 (I622502,I622836,I622723);
nor I_36478 (I622867,I622836,I622604);
nor I_36479 (I622884,I622836,I622638);
nand I_36480 (I622487,I622570,I622884);
or I_36481 (I622915,I622836,I622805);
DFFARX1 I_36482  ( .D(I622915), .CLK(I2702), .RSTB(I622519), .Q(I622484) );
not I_36483 (I622490,I622836);
DFFARX1 I_36484  ( .D(I442534), .CLK(I2702), .RSTB(I622519), .Q(I622960) );
not I_36485 (I622977,I622960);
nor I_36486 (I622994,I622977,I622570);
DFFARX1 I_36487  ( .D(I622994), .CLK(I2702), .RSTB(I622519), .Q(I622496) );
nor I_36488 (I622511,I622836,I622977);
nor I_36489 (I622499,I622977,I622740);
not I_36490 (I623053,I622977);
and I_36491 (I623070,I622604,I623053);
nor I_36492 (I622505,I622740,I623070);
nand I_36493 (I622493,I622977,I622867);
not I_36494 (I623148,I2709);
not I_36495 (I623165,I111773);
nor I_36496 (I623182,I111791,I111770);
nand I_36497 (I623199,I623182,I111788);
nor I_36498 (I623216,I623165,I111791);
nand I_36499 (I623233,I623216,I111782);
not I_36500 (I623250,I111791);
not I_36501 (I623267,I623250);
not I_36502 (I623284,I111785);
nor I_36503 (I623301,I623284,I111779);
and I_36504 (I623318,I623301,I111776);
or I_36505 (I623335,I623318,I111767);
DFFARX1 I_36506  ( .D(I623335), .CLK(I2702), .RSTB(I623148), .Q(I623352) );
nand I_36507 (I623369,I623165,I111785);
or I_36508 (I623137,I623369,I623352);
not I_36509 (I623400,I623369);
nor I_36510 (I623417,I623352,I623400);
and I_36511 (I623434,I623250,I623417);
nand I_36512 (I623110,I623369,I623267);
DFFARX1 I_36513  ( .D(I111797), .CLK(I2702), .RSTB(I623148), .Q(I623465) );
or I_36514 (I623131,I623465,I623352);
nor I_36515 (I623496,I623465,I623233);
nor I_36516 (I623513,I623465,I623267);
nand I_36517 (I623116,I623199,I623513);
or I_36518 (I623544,I623465,I623434);
DFFARX1 I_36519  ( .D(I623544), .CLK(I2702), .RSTB(I623148), .Q(I623113) );
not I_36520 (I623119,I623465);
DFFARX1 I_36521  ( .D(I111794), .CLK(I2702), .RSTB(I623148), .Q(I623589) );
not I_36522 (I623606,I623589);
nor I_36523 (I623623,I623606,I623199);
DFFARX1 I_36524  ( .D(I623623), .CLK(I2702), .RSTB(I623148), .Q(I623125) );
nor I_36525 (I623140,I623465,I623606);
nor I_36526 (I623128,I623606,I623369);
not I_36527 (I623682,I623606);
and I_36528 (I623699,I623233,I623682);
nor I_36529 (I623134,I623369,I623699);
nand I_36530 (I623122,I623606,I623496);
not I_36531 (I623777,I2709);
not I_36532 (I623794,I103375);
nor I_36533 (I623811,I103393,I103372);
nand I_36534 (I623828,I623811,I103390);
nor I_36535 (I623845,I623794,I103393);
nand I_36536 (I623862,I623845,I103384);
not I_36537 (I623879,I103393);
not I_36538 (I623896,I623879);
not I_36539 (I623913,I103387);
nor I_36540 (I623930,I623913,I103381);
and I_36541 (I623947,I623930,I103378);
or I_36542 (I623964,I623947,I103369);
DFFARX1 I_36543  ( .D(I623964), .CLK(I2702), .RSTB(I623777), .Q(I623981) );
nand I_36544 (I623998,I623794,I103387);
or I_36545 (I623766,I623998,I623981);
not I_36546 (I624029,I623998);
nor I_36547 (I624046,I623981,I624029);
and I_36548 (I624063,I623879,I624046);
nand I_36549 (I623739,I623998,I623896);
DFFARX1 I_36550  ( .D(I103399), .CLK(I2702), .RSTB(I623777), .Q(I624094) );
or I_36551 (I623760,I624094,I623981);
nor I_36552 (I624125,I624094,I623862);
nor I_36553 (I624142,I624094,I623896);
nand I_36554 (I623745,I623828,I624142);
or I_36555 (I624173,I624094,I624063);
DFFARX1 I_36556  ( .D(I624173), .CLK(I2702), .RSTB(I623777), .Q(I623742) );
not I_36557 (I623748,I624094);
DFFARX1 I_36558  ( .D(I103396), .CLK(I2702), .RSTB(I623777), .Q(I624218) );
not I_36559 (I624235,I624218);
nor I_36560 (I624252,I624235,I623828);
DFFARX1 I_36561  ( .D(I624252), .CLK(I2702), .RSTB(I623777), .Q(I623754) );
nor I_36562 (I623769,I624094,I624235);
nor I_36563 (I623757,I624235,I623998);
not I_36564 (I624311,I624235);
and I_36565 (I624328,I623862,I624311);
nor I_36566 (I623763,I623998,I624328);
nand I_36567 (I623751,I624235,I624125);
not I_36568 (I624406,I2709);
not I_36569 (I624423,I233823);
nor I_36570 (I624440,I233793,I233796);
nand I_36571 (I624457,I624440,I233814);
nor I_36572 (I624474,I624423,I233793);
nand I_36573 (I624491,I624474,I233820);
not I_36574 (I624508,I233793);
not I_36575 (I624525,I624508);
not I_36576 (I624542,I233817);
nor I_36577 (I624559,I624542,I233802);
and I_36578 (I624576,I624559,I233811);
or I_36579 (I624593,I624576,I233808);
DFFARX1 I_36580  ( .D(I624593), .CLK(I2702), .RSTB(I624406), .Q(I624610) );
nand I_36581 (I624627,I624423,I233817);
or I_36582 (I624395,I624627,I624610);
not I_36583 (I624658,I624627);
nor I_36584 (I624675,I624610,I624658);
and I_36585 (I624692,I624508,I624675);
nand I_36586 (I624368,I624627,I624525);
DFFARX1 I_36587  ( .D(I233799), .CLK(I2702), .RSTB(I624406), .Q(I624723) );
or I_36588 (I624389,I624723,I624610);
nor I_36589 (I624754,I624723,I624491);
nor I_36590 (I624771,I624723,I624525);
nand I_36591 (I624374,I624457,I624771);
or I_36592 (I624802,I624723,I624692);
DFFARX1 I_36593  ( .D(I624802), .CLK(I2702), .RSTB(I624406), .Q(I624371) );
not I_36594 (I624377,I624723);
DFFARX1 I_36595  ( .D(I233805), .CLK(I2702), .RSTB(I624406), .Q(I624847) );
not I_36596 (I624864,I624847);
nor I_36597 (I624881,I624864,I624457);
DFFARX1 I_36598  ( .D(I624881), .CLK(I2702), .RSTB(I624406), .Q(I624383) );
nor I_36599 (I624398,I624723,I624864);
nor I_36600 (I624386,I624864,I624627);
not I_36601 (I624940,I624864);
and I_36602 (I624957,I624491,I624940);
nor I_36603 (I624392,I624627,I624957);
nand I_36604 (I624380,I624864,I624754);
not I_36605 (I625035,I2709);
not I_36606 (I625052,I46473);
nor I_36607 (I625069,I46476,I46485);
nand I_36608 (I625086,I625069,I46500);
nor I_36609 (I625103,I625052,I46476);
nand I_36610 (I625120,I625103,I46479);
not I_36611 (I625137,I46476);
not I_36612 (I625154,I625137);
not I_36613 (I625171,I46470);
nor I_36614 (I625188,I625171,I46494);
and I_36615 (I625205,I625188,I46482);
or I_36616 (I625222,I625205,I46488);
DFFARX1 I_36617  ( .D(I625222), .CLK(I2702), .RSTB(I625035), .Q(I625239) );
nand I_36618 (I625256,I625052,I46470);
or I_36619 (I625024,I625256,I625239);
not I_36620 (I625287,I625256);
nor I_36621 (I625304,I625239,I625287);
and I_36622 (I625321,I625137,I625304);
nand I_36623 (I624997,I625256,I625154);
DFFARX1 I_36624  ( .D(I46491), .CLK(I2702), .RSTB(I625035), .Q(I625352) );
or I_36625 (I625018,I625352,I625239);
nor I_36626 (I625383,I625352,I625120);
nor I_36627 (I625400,I625352,I625154);
nand I_36628 (I625003,I625086,I625400);
or I_36629 (I625431,I625352,I625321);
DFFARX1 I_36630  ( .D(I625431), .CLK(I2702), .RSTB(I625035), .Q(I625000) );
not I_36631 (I625006,I625352);
DFFARX1 I_36632  ( .D(I46497), .CLK(I2702), .RSTB(I625035), .Q(I625476) );
not I_36633 (I625493,I625476);
nor I_36634 (I625510,I625493,I625086);
DFFARX1 I_36635  ( .D(I625510), .CLK(I2702), .RSTB(I625035), .Q(I625012) );
nor I_36636 (I625027,I625352,I625493);
nor I_36637 (I625015,I625493,I625256);
not I_36638 (I625569,I625493);
and I_36639 (I625586,I625120,I625569);
nor I_36640 (I625021,I625256,I625586);
nand I_36641 (I625009,I625493,I625383);
not I_36642 (I625664,I2709);
not I_36643 (I625681,I450063);
nor I_36644 (I625698,I450036,I450054);
nand I_36645 (I625715,I625698,I450039);
nor I_36646 (I625732,I625681,I450036);
nand I_36647 (I625749,I625732,I450057);
not I_36648 (I625766,I450036);
not I_36649 (I625783,I625766);
not I_36650 (I625800,I450033);
nor I_36651 (I625817,I625800,I450060);
and I_36652 (I625834,I625817,I450051);
or I_36653 (I625851,I625834,I450042);
DFFARX1 I_36654  ( .D(I625851), .CLK(I2702), .RSTB(I625664), .Q(I625868) );
nand I_36655 (I625885,I625681,I450033);
or I_36656 (I625653,I625885,I625868);
not I_36657 (I625916,I625885);
nor I_36658 (I625933,I625868,I625916);
and I_36659 (I625950,I625766,I625933);
nand I_36660 (I625626,I625885,I625783);
DFFARX1 I_36661  ( .D(I450045), .CLK(I2702), .RSTB(I625664), .Q(I625981) );
or I_36662 (I625647,I625981,I625868);
nor I_36663 (I626012,I625981,I625749);
nor I_36664 (I626029,I625981,I625783);
nand I_36665 (I625632,I625715,I626029);
or I_36666 (I626060,I625981,I625950);
DFFARX1 I_36667  ( .D(I626060), .CLK(I2702), .RSTB(I625664), .Q(I625629) );
not I_36668 (I625635,I625981);
DFFARX1 I_36669  ( .D(I450048), .CLK(I2702), .RSTB(I625664), .Q(I626105) );
not I_36670 (I626122,I626105);
nor I_36671 (I626139,I626122,I625715);
DFFARX1 I_36672  ( .D(I626139), .CLK(I2702), .RSTB(I625664), .Q(I625641) );
nor I_36673 (I625656,I625981,I626122);
nor I_36674 (I625644,I626122,I625885);
not I_36675 (I626198,I626122);
and I_36676 (I626215,I625749,I626198);
nor I_36677 (I625650,I625885,I626215);
nand I_36678 (I625638,I626122,I626012);
not I_36679 (I626293,I2709);
not I_36680 (I626310,I393883);
nor I_36681 (I626327,I393892,I393895);
nand I_36682 (I626344,I626327,I393880);
nor I_36683 (I626361,I626310,I393892);
nand I_36684 (I626378,I626361,I393877);
not I_36685 (I626395,I393892);
not I_36686 (I626412,I626395);
not I_36687 (I626429,I393865);
nor I_36688 (I626446,I626429,I393871);
and I_36689 (I626463,I626446,I393868);
or I_36690 (I626480,I626463,I393889);
DFFARX1 I_36691  ( .D(I626480), .CLK(I2702), .RSTB(I626293), .Q(I626497) );
nand I_36692 (I626514,I626310,I393865);
or I_36693 (I626282,I626514,I626497);
not I_36694 (I626545,I626514);
nor I_36695 (I626562,I626497,I626545);
and I_36696 (I626579,I626395,I626562);
nand I_36697 (I626255,I626514,I626412);
DFFARX1 I_36698  ( .D(I393874), .CLK(I2702), .RSTB(I626293), .Q(I626610) );
or I_36699 (I626276,I626610,I626497);
nor I_36700 (I626641,I626610,I626378);
nor I_36701 (I626658,I626610,I626412);
nand I_36702 (I626261,I626344,I626658);
or I_36703 (I626689,I626610,I626579);
DFFARX1 I_36704  ( .D(I626689), .CLK(I2702), .RSTB(I626293), .Q(I626258) );
not I_36705 (I626264,I626610);
DFFARX1 I_36706  ( .D(I393886), .CLK(I2702), .RSTB(I626293), .Q(I626734) );
not I_36707 (I626751,I626734);
nor I_36708 (I626768,I626751,I626344);
DFFARX1 I_36709  ( .D(I626768), .CLK(I2702), .RSTB(I626293), .Q(I626270) );
nor I_36710 (I626285,I626610,I626751);
nor I_36711 (I626273,I626751,I626514);
not I_36712 (I626827,I626751);
and I_36713 (I626844,I626378,I626827);
nor I_36714 (I626279,I626514,I626844);
nand I_36715 (I626267,I626751,I626641);
not I_36716 (I626922,I2709);
not I_36717 (I626939,I711176);
nor I_36718 (I626956,I711200,I711185);
nand I_36719 (I626973,I626956,I711170);
nor I_36720 (I626990,I626939,I711200);
nand I_36721 (I627007,I626990,I711197);
not I_36722 (I627024,I711200);
not I_36723 (I627041,I627024);
not I_36724 (I627058,I711179);
nor I_36725 (I627075,I627058,I711173);
and I_36726 (I627092,I627075,I711194);
or I_36727 (I627109,I627092,I711182);
DFFARX1 I_36728  ( .D(I627109), .CLK(I2702), .RSTB(I626922), .Q(I627126) );
nand I_36729 (I627143,I626939,I711179);
or I_36730 (I626911,I627143,I627126);
not I_36731 (I627174,I627143);
nor I_36732 (I627191,I627126,I627174);
and I_36733 (I627208,I627024,I627191);
nand I_36734 (I626884,I627143,I627041);
DFFARX1 I_36735  ( .D(I711191), .CLK(I2702), .RSTB(I626922), .Q(I627239) );
or I_36736 (I626905,I627239,I627126);
nor I_36737 (I627270,I627239,I627007);
nor I_36738 (I627287,I627239,I627041);
nand I_36739 (I626890,I626973,I627287);
or I_36740 (I627318,I627239,I627208);
DFFARX1 I_36741  ( .D(I627318), .CLK(I2702), .RSTB(I626922), .Q(I626887) );
not I_36742 (I626893,I627239);
DFFARX1 I_36743  ( .D(I711188), .CLK(I2702), .RSTB(I626922), .Q(I627363) );
not I_36744 (I627380,I627363);
nor I_36745 (I627397,I627380,I626973);
DFFARX1 I_36746  ( .D(I627397), .CLK(I2702), .RSTB(I626922), .Q(I626899) );
nor I_36747 (I626914,I627239,I627380);
nor I_36748 (I626902,I627380,I627143);
not I_36749 (I627456,I627380);
and I_36750 (I627473,I627007,I627456);
nor I_36751 (I626908,I627143,I627473);
nand I_36752 (I626896,I627380,I627270);
not I_36753 (I627551,I2709);
not I_36754 (I627568,I47034);
nor I_36755 (I627585,I47037,I47046);
nand I_36756 (I627602,I627585,I47061);
nor I_36757 (I627619,I627568,I47037);
nand I_36758 (I627636,I627619,I47040);
not I_36759 (I627653,I47037);
not I_36760 (I627670,I627653);
not I_36761 (I627687,I47031);
nor I_36762 (I627704,I627687,I47055);
and I_36763 (I627721,I627704,I47043);
or I_36764 (I627738,I627721,I47049);
DFFARX1 I_36765  ( .D(I627738), .CLK(I2702), .RSTB(I627551), .Q(I627755) );
nand I_36766 (I627772,I627568,I47031);
or I_36767 (I627540,I627772,I627755);
not I_36768 (I627803,I627772);
nor I_36769 (I627820,I627755,I627803);
and I_36770 (I627837,I627653,I627820);
nand I_36771 (I627513,I627772,I627670);
DFFARX1 I_36772  ( .D(I47052), .CLK(I2702), .RSTB(I627551), .Q(I627868) );
or I_36773 (I627534,I627868,I627755);
nor I_36774 (I627899,I627868,I627636);
nor I_36775 (I627916,I627868,I627670);
nand I_36776 (I627519,I627602,I627916);
or I_36777 (I627947,I627868,I627837);
DFFARX1 I_36778  ( .D(I627947), .CLK(I2702), .RSTB(I627551), .Q(I627516) );
not I_36779 (I627522,I627868);
DFFARX1 I_36780  ( .D(I47058), .CLK(I2702), .RSTB(I627551), .Q(I627992) );
not I_36781 (I628009,I627992);
nor I_36782 (I628026,I628009,I627602);
DFFARX1 I_36783  ( .D(I628026), .CLK(I2702), .RSTB(I627551), .Q(I627528) );
nor I_36784 (I627543,I627868,I628009);
nor I_36785 (I627531,I628009,I627772);
not I_36786 (I628085,I628009);
and I_36787 (I628102,I627636,I628085);
nor I_36788 (I627537,I627772,I628102);
nand I_36789 (I627525,I628009,I627899);
not I_36790 (I628180,I2709);
not I_36791 (I628197,I553025);
nor I_36792 (I628214,I553043,I553022);
nand I_36793 (I628231,I628214,I553046);
nor I_36794 (I628248,I628197,I553043);
nand I_36795 (I628265,I628248,I553040);
not I_36796 (I628282,I553043);
not I_36797 (I628299,I628282);
not I_36798 (I628316,I553031);
nor I_36799 (I628333,I628316,I553019);
and I_36800 (I628350,I628333,I553037);
or I_36801 (I628367,I628350,I553049);
DFFARX1 I_36802  ( .D(I628367), .CLK(I2702), .RSTB(I628180), .Q(I628384) );
nand I_36803 (I628401,I628197,I553031);
or I_36804 (I628169,I628401,I628384);
not I_36805 (I628432,I628401);
nor I_36806 (I628449,I628384,I628432);
and I_36807 (I628466,I628282,I628449);
nand I_36808 (I628142,I628401,I628299);
DFFARX1 I_36809  ( .D(I553028), .CLK(I2702), .RSTB(I628180), .Q(I628497) );
or I_36810 (I628163,I628497,I628384);
nor I_36811 (I628528,I628497,I628265);
nor I_36812 (I628545,I628497,I628299);
nand I_36813 (I628148,I628231,I628545);
or I_36814 (I628576,I628497,I628466);
DFFARX1 I_36815  ( .D(I628576), .CLK(I2702), .RSTB(I628180), .Q(I628145) );
not I_36816 (I628151,I628497);
DFFARX1 I_36817  ( .D(I553034), .CLK(I2702), .RSTB(I628180), .Q(I628621) );
not I_36818 (I628638,I628621);
nor I_36819 (I628655,I628638,I628231);
DFFARX1 I_36820  ( .D(I628655), .CLK(I2702), .RSTB(I628180), .Q(I628157) );
nor I_36821 (I628172,I628497,I628638);
nor I_36822 (I628160,I628638,I628401);
not I_36823 (I628714,I628638);
and I_36824 (I628731,I628265,I628714);
nor I_36825 (I628166,I628401,I628731);
nand I_36826 (I628154,I628638,I628528);
not I_36827 (I628809,I2709);
not I_36828 (I628826,I63323);
nor I_36829 (I628843,I63341,I63320);
nand I_36830 (I628860,I628843,I63338);
nor I_36831 (I628877,I628826,I63341);
nand I_36832 (I628894,I628877,I63332);
not I_36833 (I628911,I63341);
not I_36834 (I628928,I628911);
not I_36835 (I628945,I63335);
nor I_36836 (I628962,I628945,I63329);
and I_36837 (I628979,I628962,I63326);
or I_36838 (I628996,I628979,I63317);
DFFARX1 I_36839  ( .D(I628996), .CLK(I2702), .RSTB(I628809), .Q(I629013) );
nand I_36840 (I629030,I628826,I63335);
or I_36841 (I628798,I629030,I629013);
not I_36842 (I629061,I629030);
nor I_36843 (I629078,I629013,I629061);
and I_36844 (I629095,I628911,I629078);
nand I_36845 (I628771,I629030,I628928);
DFFARX1 I_36846  ( .D(I63347), .CLK(I2702), .RSTB(I628809), .Q(I629126) );
or I_36847 (I628792,I629126,I629013);
nor I_36848 (I629157,I629126,I628894);
nor I_36849 (I629174,I629126,I628928);
nand I_36850 (I628777,I628860,I629174);
or I_36851 (I629205,I629126,I629095);
DFFARX1 I_36852  ( .D(I629205), .CLK(I2702), .RSTB(I628809), .Q(I628774) );
not I_36853 (I628780,I629126);
DFFARX1 I_36854  ( .D(I63344), .CLK(I2702), .RSTB(I628809), .Q(I629250) );
not I_36855 (I629267,I629250);
nor I_36856 (I629284,I629267,I628860);
DFFARX1 I_36857  ( .D(I629284), .CLK(I2702), .RSTB(I628809), .Q(I628786) );
nor I_36858 (I628801,I629126,I629267);
nor I_36859 (I628789,I629267,I629030);
not I_36860 (I629343,I629267);
and I_36861 (I629360,I628894,I629343);
nor I_36862 (I628795,I629030,I629360);
nand I_36863 (I628783,I629267,I629157);
not I_36864 (I629438,I2709);
not I_36865 (I629455,I152817);
nor I_36866 (I629472,I152808,I152832);
nand I_36867 (I629489,I629472,I152835);
nor I_36868 (I629506,I629455,I152808);
nand I_36869 (I629523,I629506,I152826);
not I_36870 (I629540,I152808);
not I_36871 (I629557,I629540);
not I_36872 (I629574,I152820);
nor I_36873 (I629591,I629574,I152814);
and I_36874 (I629608,I629591,I152823);
or I_36875 (I629625,I629608,I152811);
DFFARX1 I_36876  ( .D(I629625), .CLK(I2702), .RSTB(I629438), .Q(I629642) );
nand I_36877 (I629659,I629455,I152820);
or I_36878 (I629427,I629659,I629642);
not I_36879 (I629690,I629659);
nor I_36880 (I629707,I629642,I629690);
and I_36881 (I629724,I629540,I629707);
nand I_36882 (I629400,I629659,I629557);
DFFARX1 I_36883  ( .D(I152805), .CLK(I2702), .RSTB(I629438), .Q(I629755) );
or I_36884 (I629421,I629755,I629642);
nor I_36885 (I629786,I629755,I629523);
nor I_36886 (I629803,I629755,I629557);
nand I_36887 (I629406,I629489,I629803);
or I_36888 (I629834,I629755,I629724);
DFFARX1 I_36889  ( .D(I629834), .CLK(I2702), .RSTB(I629438), .Q(I629403) );
not I_36890 (I629409,I629755);
DFFARX1 I_36891  ( .D(I152829), .CLK(I2702), .RSTB(I629438), .Q(I629879) );
not I_36892 (I629896,I629879);
nor I_36893 (I629913,I629896,I629489);
DFFARX1 I_36894  ( .D(I629913), .CLK(I2702), .RSTB(I629438), .Q(I629415) );
nor I_36895 (I629430,I629755,I629896);
nor I_36896 (I629418,I629896,I629659);
not I_36897 (I629972,I629896);
and I_36898 (I629989,I629523,I629972);
nor I_36899 (I629424,I629659,I629989);
nand I_36900 (I629412,I629896,I629786);
not I_36901 (I630067,I2709);
not I_36902 (I630084,I411325);
nor I_36903 (I630101,I411334,I411337);
nand I_36904 (I630118,I630101,I411322);
nor I_36905 (I630135,I630084,I411334);
nand I_36906 (I630152,I630135,I411319);
not I_36907 (I630169,I411334);
not I_36908 (I630186,I630169);
not I_36909 (I630203,I411307);
nor I_36910 (I630220,I630203,I411313);
and I_36911 (I630237,I630220,I411310);
or I_36912 (I630254,I630237,I411331);
DFFARX1 I_36913  ( .D(I630254), .CLK(I2702), .RSTB(I630067), .Q(I630271) );
nand I_36914 (I630288,I630084,I411307);
or I_36915 (I630056,I630288,I630271);
not I_36916 (I630319,I630288);
nor I_36917 (I630336,I630271,I630319);
and I_36918 (I630353,I630169,I630336);
nand I_36919 (I630029,I630288,I630186);
DFFARX1 I_36920  ( .D(I411316), .CLK(I2702), .RSTB(I630067), .Q(I630384) );
or I_36921 (I630050,I630384,I630271);
nor I_36922 (I630415,I630384,I630152);
nor I_36923 (I630432,I630384,I630186);
nand I_36924 (I630035,I630118,I630432);
or I_36925 (I630463,I630384,I630353);
DFFARX1 I_36926  ( .D(I630463), .CLK(I2702), .RSTB(I630067), .Q(I630032) );
not I_36927 (I630038,I630384);
DFFARX1 I_36928  ( .D(I411328), .CLK(I2702), .RSTB(I630067), .Q(I630508) );
not I_36929 (I630525,I630508);
nor I_36930 (I630542,I630525,I630118);
DFFARX1 I_36931  ( .D(I630542), .CLK(I2702), .RSTB(I630067), .Q(I630044) );
nor I_36932 (I630059,I630384,I630525);
nor I_36933 (I630047,I630525,I630288);
not I_36934 (I630601,I630525);
and I_36935 (I630618,I630152,I630601);
nor I_36936 (I630053,I630288,I630618);
nand I_36937 (I630041,I630525,I630415);
not I_36938 (I630696,I2709);
not I_36939 (I630713,I256251);
nor I_36940 (I630730,I256257,I256236);
nand I_36941 (I630747,I630730,I256242);
nor I_36942 (I630764,I630713,I256257);
nand I_36943 (I630781,I630764,I256248);
not I_36944 (I630798,I256257);
not I_36945 (I630815,I630798);
not I_36946 (I630832,I256245);
nor I_36947 (I630849,I630832,I256263);
and I_36948 (I630866,I630849,I256254);
or I_36949 (I630883,I630866,I256233);
DFFARX1 I_36950  ( .D(I630883), .CLK(I2702), .RSTB(I630696), .Q(I630900) );
nand I_36951 (I630917,I630713,I256245);
or I_36952 (I630685,I630917,I630900);
not I_36953 (I630948,I630917);
nor I_36954 (I630965,I630900,I630948);
and I_36955 (I630982,I630798,I630965);
nand I_36956 (I630658,I630917,I630815);
DFFARX1 I_36957  ( .D(I256260), .CLK(I2702), .RSTB(I630696), .Q(I631013) );
or I_36958 (I630679,I631013,I630900);
nor I_36959 (I631044,I631013,I630781);
nor I_36960 (I631061,I631013,I630815);
nand I_36961 (I630664,I630747,I631061);
or I_36962 (I631092,I631013,I630982);
DFFARX1 I_36963  ( .D(I631092), .CLK(I2702), .RSTB(I630696), .Q(I630661) );
not I_36964 (I630667,I631013);
DFFARX1 I_36965  ( .D(I256239), .CLK(I2702), .RSTB(I630696), .Q(I631137) );
not I_36966 (I631154,I631137);
nor I_36967 (I631171,I631154,I630747);
DFFARX1 I_36968  ( .D(I631171), .CLK(I2702), .RSTB(I630696), .Q(I630673) );
nor I_36969 (I630688,I631013,I631154);
nor I_36970 (I630676,I631154,I630917);
not I_36971 (I631230,I631154);
and I_36972 (I631247,I630781,I631230);
nor I_36973 (I630682,I630917,I631247);
nand I_36974 (I630670,I631154,I631044);
not I_36975 (I631325,I2709);
not I_36976 (I631342,I600033);
nor I_36977 (I631359,I600036,I600045);
nand I_36978 (I631376,I631359,I600030);
nor I_36979 (I631393,I631342,I600036);
nand I_36980 (I631410,I631393,I600039);
not I_36981 (I631427,I600036);
not I_36982 (I631444,I631427);
not I_36983 (I631461,I600054);
nor I_36984 (I631478,I631461,I600042);
and I_36985 (I631495,I631478,I600027);
or I_36986 (I631512,I631495,I600024);
DFFARX1 I_36987  ( .D(I631512), .CLK(I2702), .RSTB(I631325), .Q(I631529) );
nand I_36988 (I631546,I631342,I600054);
or I_36989 (I631314,I631546,I631529);
not I_36990 (I631577,I631546);
nor I_36991 (I631594,I631529,I631577);
and I_36992 (I631611,I631427,I631594);
nand I_36993 (I631287,I631546,I631444);
DFFARX1 I_36994  ( .D(I600048), .CLK(I2702), .RSTB(I631325), .Q(I631642) );
or I_36995 (I631308,I631642,I631529);
nor I_36996 (I631673,I631642,I631410);
nor I_36997 (I631690,I631642,I631444);
nand I_36998 (I631293,I631376,I631690);
or I_36999 (I631721,I631642,I631611);
DFFARX1 I_37000  ( .D(I631721), .CLK(I2702), .RSTB(I631325), .Q(I631290) );
not I_37001 (I631296,I631642);
DFFARX1 I_37002  ( .D(I600051), .CLK(I2702), .RSTB(I631325), .Q(I631766) );
not I_37003 (I631783,I631766);
nor I_37004 (I631800,I631783,I631376);
DFFARX1 I_37005  ( .D(I631800), .CLK(I2702), .RSTB(I631325), .Q(I631302) );
nor I_37006 (I631317,I631642,I631783);
nor I_37007 (I631305,I631783,I631546);
not I_37008 (I631859,I631783);
and I_37009 (I631876,I631410,I631859);
nor I_37010 (I631311,I631546,I631876);
nand I_37011 (I631299,I631783,I631673);
not I_37012 (I631954,I2709);
not I_37013 (I631971,I603008);
nor I_37014 (I631988,I603011,I603020);
nand I_37015 (I632005,I631988,I603005);
nor I_37016 (I632022,I631971,I603011);
nand I_37017 (I632039,I632022,I603014);
not I_37018 (I632056,I603011);
not I_37019 (I632073,I632056);
not I_37020 (I632090,I603029);
nor I_37021 (I632107,I632090,I603017);
and I_37022 (I632124,I632107,I603002);
or I_37023 (I632141,I632124,I602999);
DFFARX1 I_37024  ( .D(I632141), .CLK(I2702), .RSTB(I631954), .Q(I632158) );
nand I_37025 (I632175,I631971,I603029);
or I_37026 (I631943,I632175,I632158);
not I_37027 (I632206,I632175);
nor I_37028 (I632223,I632158,I632206);
and I_37029 (I632240,I632056,I632223);
nand I_37030 (I631916,I632175,I632073);
DFFARX1 I_37031  ( .D(I603023), .CLK(I2702), .RSTB(I631954), .Q(I632271) );
or I_37032 (I631937,I632271,I632158);
nor I_37033 (I632302,I632271,I632039);
nor I_37034 (I632319,I632271,I632073);
nand I_37035 (I631922,I632005,I632319);
or I_37036 (I632350,I632271,I632240);
DFFARX1 I_37037  ( .D(I632350), .CLK(I2702), .RSTB(I631954), .Q(I631919) );
not I_37038 (I631925,I632271);
DFFARX1 I_37039  ( .D(I603026), .CLK(I2702), .RSTB(I631954), .Q(I632395) );
not I_37040 (I632412,I632395);
nor I_37041 (I632429,I632412,I632005);
DFFARX1 I_37042  ( .D(I632429), .CLK(I2702), .RSTB(I631954), .Q(I631931) );
nor I_37043 (I631946,I632271,I632412);
nor I_37044 (I631934,I632412,I632175);
not I_37045 (I632488,I632412);
and I_37046 (I632505,I632039,I632488);
nor I_37047 (I631940,I632175,I632505);
nand I_37048 (I631928,I632412,I632302);
not I_37049 (I632583,I2709);
not I_37050 (I632600,I1551);
nor I_37051 (I632617,I2687,I2503);
nand I_37052 (I632634,I632617,I1911);
nor I_37053 (I632651,I632600,I2687);
nand I_37054 (I632668,I632651,I2591);
not I_37055 (I632685,I2687);
not I_37056 (I632702,I632685);
not I_37057 (I632719,I1295);
nor I_37058 (I632736,I632719,I2103);
and I_37059 (I632753,I632736,I1871);
or I_37060 (I632770,I632753,I1783);
DFFARX1 I_37061  ( .D(I632770), .CLK(I2702), .RSTB(I632583), .Q(I632787) );
nand I_37062 (I632804,I632600,I1295);
or I_37063 (I632572,I632804,I632787);
not I_37064 (I632835,I632804);
nor I_37065 (I632852,I632787,I632835);
and I_37066 (I632869,I632685,I632852);
nand I_37067 (I632545,I632804,I632702);
DFFARX1 I_37068  ( .D(I1647), .CLK(I2702), .RSTB(I632583), .Q(I632900) );
or I_37069 (I632566,I632900,I632787);
nor I_37070 (I632931,I632900,I632668);
nor I_37071 (I632948,I632900,I632702);
nand I_37072 (I632551,I632634,I632948);
or I_37073 (I632979,I632900,I632869);
DFFARX1 I_37074  ( .D(I632979), .CLK(I2702), .RSTB(I632583), .Q(I632548) );
not I_37075 (I632554,I632900);
DFFARX1 I_37076  ( .D(I2407), .CLK(I2702), .RSTB(I632583), .Q(I633024) );
not I_37077 (I633041,I633024);
nor I_37078 (I633058,I633041,I632634);
DFFARX1 I_37079  ( .D(I633058), .CLK(I2702), .RSTB(I632583), .Q(I632560) );
nor I_37080 (I632575,I632900,I633041);
nor I_37081 (I632563,I633041,I632804);
not I_37082 (I633117,I633041);
and I_37083 (I633134,I632668,I633117);
nor I_37084 (I632569,I632804,I633134);
nand I_37085 (I632557,I633041,I632931);
not I_37086 (I633212,I2709);
not I_37087 (I633229,I94331);
nor I_37088 (I633246,I94349,I94328);
nand I_37089 (I633263,I633246,I94346);
nor I_37090 (I633280,I633229,I94349);
nand I_37091 (I633297,I633280,I94340);
not I_37092 (I633314,I94349);
not I_37093 (I633331,I633314);
not I_37094 (I633348,I94343);
nor I_37095 (I633365,I633348,I94337);
and I_37096 (I633382,I633365,I94334);
or I_37097 (I633399,I633382,I94325);
DFFARX1 I_37098  ( .D(I633399), .CLK(I2702), .RSTB(I633212), .Q(I633416) );
nand I_37099 (I633433,I633229,I94343);
or I_37100 (I633201,I633433,I633416);
not I_37101 (I633464,I633433);
nor I_37102 (I633481,I633416,I633464);
and I_37103 (I633498,I633314,I633481);
nand I_37104 (I633174,I633433,I633331);
DFFARX1 I_37105  ( .D(I94355), .CLK(I2702), .RSTB(I633212), .Q(I633529) );
or I_37106 (I633195,I633529,I633416);
nor I_37107 (I633560,I633529,I633297);
nor I_37108 (I633577,I633529,I633331);
nand I_37109 (I633180,I633263,I633577);
or I_37110 (I633608,I633529,I633498);
DFFARX1 I_37111  ( .D(I633608), .CLK(I2702), .RSTB(I633212), .Q(I633177) );
not I_37112 (I633183,I633529);
DFFARX1 I_37113  ( .D(I94352), .CLK(I2702), .RSTB(I633212), .Q(I633653) );
not I_37114 (I633670,I633653);
nor I_37115 (I633687,I633670,I633263);
DFFARX1 I_37116  ( .D(I633687), .CLK(I2702), .RSTB(I633212), .Q(I633189) );
nor I_37117 (I633204,I633529,I633670);
nor I_37118 (I633192,I633670,I633433);
not I_37119 (I633746,I633670);
and I_37120 (I633763,I633297,I633746);
nor I_37121 (I633198,I633433,I633763);
nand I_37122 (I633186,I633670,I633560);
not I_37123 (I633841,I2709);
not I_37124 (I633858,I351893);
nor I_37125 (I633875,I351902,I351905);
nand I_37126 (I633892,I633875,I351890);
nor I_37127 (I633909,I633858,I351902);
nand I_37128 (I633926,I633909,I351887);
not I_37129 (I633943,I351902);
not I_37130 (I633960,I633943);
not I_37131 (I633977,I351875);
nor I_37132 (I633994,I633977,I351881);
and I_37133 (I634011,I633994,I351878);
or I_37134 (I634028,I634011,I351899);
DFFARX1 I_37135  ( .D(I634028), .CLK(I2702), .RSTB(I633841), .Q(I634045) );
nand I_37136 (I634062,I633858,I351875);
or I_37137 (I633830,I634062,I634045);
not I_37138 (I634093,I634062);
nor I_37139 (I634110,I634045,I634093);
and I_37140 (I634127,I633943,I634110);
nand I_37141 (I633803,I634062,I633960);
DFFARX1 I_37142  ( .D(I351884), .CLK(I2702), .RSTB(I633841), .Q(I634158) );
or I_37143 (I633824,I634158,I634045);
nor I_37144 (I634189,I634158,I633926);
nor I_37145 (I634206,I634158,I633960);
nand I_37146 (I633809,I633892,I634206);
or I_37147 (I634237,I634158,I634127);
DFFARX1 I_37148  ( .D(I634237), .CLK(I2702), .RSTB(I633841), .Q(I633806) );
not I_37149 (I633812,I634158);
DFFARX1 I_37150  ( .D(I351896), .CLK(I2702), .RSTB(I633841), .Q(I634282) );
not I_37151 (I634299,I634282);
nor I_37152 (I634316,I634299,I633892);
DFFARX1 I_37153  ( .D(I634316), .CLK(I2702), .RSTB(I633841), .Q(I633818) );
nor I_37154 (I633833,I634158,I634299);
nor I_37155 (I633821,I634299,I634062);
not I_37156 (I634375,I634299);
and I_37157 (I634392,I633926,I634375);
nor I_37158 (I633827,I634062,I634392);
nand I_37159 (I633815,I634299,I634189);
not I_37160 (I634470,I2709);
not I_37161 (I634487,I220733);
nor I_37162 (I634504,I220709,I220724);
nand I_37163 (I634521,I634504,I220706);
nor I_37164 (I634538,I634487,I220709);
nand I_37165 (I634555,I634538,I220721);
not I_37166 (I634572,I220709);
not I_37167 (I634589,I634572);
not I_37168 (I634606,I220712);
nor I_37169 (I634623,I634606,I220727);
and I_37170 (I634640,I634623,I220718);
or I_37171 (I634657,I634640,I220703);
DFFARX1 I_37172  ( .D(I634657), .CLK(I2702), .RSTB(I634470), .Q(I634674) );
nand I_37173 (I634691,I634487,I220712);
or I_37174 (I634459,I634691,I634674);
not I_37175 (I634722,I634691);
nor I_37176 (I634739,I634674,I634722);
and I_37177 (I634756,I634572,I634739);
nand I_37178 (I634432,I634691,I634589);
DFFARX1 I_37179  ( .D(I220715), .CLK(I2702), .RSTB(I634470), .Q(I634787) );
or I_37180 (I634453,I634787,I634674);
nor I_37181 (I634818,I634787,I634555);
nor I_37182 (I634835,I634787,I634589);
nand I_37183 (I634438,I634521,I634835);
or I_37184 (I634866,I634787,I634756);
DFFARX1 I_37185  ( .D(I634866), .CLK(I2702), .RSTB(I634470), .Q(I634435) );
not I_37186 (I634441,I634787);
DFFARX1 I_37187  ( .D(I220730), .CLK(I2702), .RSTB(I634470), .Q(I634911) );
not I_37188 (I634928,I634911);
nor I_37189 (I634945,I634928,I634521);
DFFARX1 I_37190  ( .D(I634945), .CLK(I2702), .RSTB(I634470), .Q(I634447) );
nor I_37191 (I634462,I634787,I634928);
nor I_37192 (I634450,I634928,I634691);
not I_37193 (I635004,I634928);
and I_37194 (I635021,I634555,I635004);
nor I_37195 (I634456,I634691,I635021);
nand I_37196 (I634444,I634928,I634818);
not I_37197 (I635099,I2709);
not I_37198 (I635116,I437347);
nor I_37199 (I635133,I437320,I437338);
nand I_37200 (I635150,I635133,I437323);
nor I_37201 (I635167,I635116,I437320);
nand I_37202 (I635184,I635167,I437341);
not I_37203 (I635201,I437320);
not I_37204 (I635218,I635201);
not I_37205 (I635235,I437317);
nor I_37206 (I635252,I635235,I437344);
and I_37207 (I635269,I635252,I437335);
or I_37208 (I635286,I635269,I437326);
DFFARX1 I_37209  ( .D(I635286), .CLK(I2702), .RSTB(I635099), .Q(I635303) );
nand I_37210 (I635320,I635116,I437317);
or I_37211 (I635088,I635320,I635303);
not I_37212 (I635351,I635320);
nor I_37213 (I635368,I635303,I635351);
and I_37214 (I635385,I635201,I635368);
nand I_37215 (I635061,I635320,I635218);
DFFARX1 I_37216  ( .D(I437329), .CLK(I2702), .RSTB(I635099), .Q(I635416) );
or I_37217 (I635082,I635416,I635303);
nor I_37218 (I635447,I635416,I635184);
nor I_37219 (I635464,I635416,I635218);
nand I_37220 (I635067,I635150,I635464);
or I_37221 (I635495,I635416,I635385);
DFFARX1 I_37222  ( .D(I635495), .CLK(I2702), .RSTB(I635099), .Q(I635064) );
not I_37223 (I635070,I635416);
DFFARX1 I_37224  ( .D(I437332), .CLK(I2702), .RSTB(I635099), .Q(I635540) );
not I_37225 (I635557,I635540);
nor I_37226 (I635574,I635557,I635150);
DFFARX1 I_37227  ( .D(I635574), .CLK(I2702), .RSTB(I635099), .Q(I635076) );
nor I_37228 (I635091,I635416,I635557);
nor I_37229 (I635079,I635557,I635320);
not I_37230 (I635633,I635557);
and I_37231 (I635650,I635184,I635633);
nor I_37232 (I635085,I635320,I635650);
nand I_37233 (I635073,I635557,I635447);
not I_37234 (I635728,I2709);
not I_37235 (I635745,I150828);
nor I_37236 (I635762,I150819,I150843);
nand I_37237 (I635779,I635762,I150846);
nor I_37238 (I635796,I635745,I150819);
nand I_37239 (I635813,I635796,I150837);
not I_37240 (I635830,I150819);
not I_37241 (I635847,I635830);
not I_37242 (I635864,I150831);
nor I_37243 (I635881,I635864,I150825);
and I_37244 (I635898,I635881,I150834);
or I_37245 (I635915,I635898,I150822);
DFFARX1 I_37246  ( .D(I635915), .CLK(I2702), .RSTB(I635728), .Q(I635932) );
nand I_37247 (I635949,I635745,I150831);
or I_37248 (I635717,I635949,I635932);
not I_37249 (I635980,I635949);
nor I_37250 (I635997,I635932,I635980);
and I_37251 (I636014,I635830,I635997);
nand I_37252 (I635690,I635949,I635847);
DFFARX1 I_37253  ( .D(I150816), .CLK(I2702), .RSTB(I635728), .Q(I636045) );
or I_37254 (I635711,I636045,I635932);
nor I_37255 (I636076,I636045,I635813);
nor I_37256 (I636093,I636045,I635847);
nand I_37257 (I635696,I635779,I636093);
or I_37258 (I636124,I636045,I636014);
DFFARX1 I_37259  ( .D(I636124), .CLK(I2702), .RSTB(I635728), .Q(I635693) );
not I_37260 (I635699,I636045);
DFFARX1 I_37261  ( .D(I150840), .CLK(I2702), .RSTB(I635728), .Q(I636169) );
not I_37262 (I636186,I636169);
nor I_37263 (I636203,I636186,I635779);
DFFARX1 I_37264  ( .D(I636203), .CLK(I2702), .RSTB(I635728), .Q(I635705) );
nor I_37265 (I635720,I636045,I636186);
nor I_37266 (I635708,I636186,I635949);
not I_37267 (I636262,I636186);
and I_37268 (I636279,I635813,I636262);
nor I_37269 (I635714,I635949,I636279);
nand I_37270 (I635702,I636186,I636076);
not I_37271 (I636357,I2709);
not I_37272 (I636374,I529820);
nor I_37273 (I636391,I529838,I529817);
nand I_37274 (I636408,I636391,I529841);
nor I_37275 (I636425,I636374,I529838);
nand I_37276 (I636442,I636425,I529835);
not I_37277 (I636459,I529838);
not I_37278 (I636476,I636459);
not I_37279 (I636493,I529826);
nor I_37280 (I636510,I636493,I529814);
and I_37281 (I636527,I636510,I529832);
or I_37282 (I636544,I636527,I529844);
DFFARX1 I_37283  ( .D(I636544), .CLK(I2702), .RSTB(I636357), .Q(I636561) );
nand I_37284 (I636578,I636374,I529826);
or I_37285 (I636346,I636578,I636561);
not I_37286 (I636609,I636578);
nor I_37287 (I636626,I636561,I636609);
and I_37288 (I636643,I636459,I636626);
nand I_37289 (I636319,I636578,I636476);
DFFARX1 I_37290  ( .D(I529823), .CLK(I2702), .RSTB(I636357), .Q(I636674) );
or I_37291 (I636340,I636674,I636561);
nor I_37292 (I636705,I636674,I636442);
nor I_37293 (I636722,I636674,I636476);
nand I_37294 (I636325,I636408,I636722);
or I_37295 (I636753,I636674,I636643);
DFFARX1 I_37296  ( .D(I636753), .CLK(I2702), .RSTB(I636357), .Q(I636322) );
not I_37297 (I636328,I636674);
DFFARX1 I_37298  ( .D(I529829), .CLK(I2702), .RSTB(I636357), .Q(I636798) );
not I_37299 (I636815,I636798);
nor I_37300 (I636832,I636815,I636408);
DFFARX1 I_37301  ( .D(I636832), .CLK(I2702), .RSTB(I636357), .Q(I636334) );
nor I_37302 (I636349,I636674,I636815);
nor I_37303 (I636337,I636815,I636578);
not I_37304 (I636891,I636815);
and I_37305 (I636908,I636442,I636891);
nor I_37306 (I636343,I636578,I636908);
nand I_37307 (I636331,I636815,I636705);
not I_37308 (I636986,I2709);
not I_37309 (I637003,I260229);
nor I_37310 (I637020,I260235,I260214);
nand I_37311 (I637037,I637020,I260220);
nor I_37312 (I637054,I637003,I260235);
nand I_37313 (I637071,I637054,I260226);
not I_37314 (I637088,I260235);
not I_37315 (I637105,I637088);
not I_37316 (I637122,I260223);
nor I_37317 (I637139,I637122,I260241);
and I_37318 (I637156,I637139,I260232);
or I_37319 (I637173,I637156,I260211);
DFFARX1 I_37320  ( .D(I637173), .CLK(I2702), .RSTB(I636986), .Q(I637190) );
nand I_37321 (I637207,I637003,I260223);
or I_37322 (I636975,I637207,I637190);
not I_37323 (I637238,I637207);
nor I_37324 (I637255,I637190,I637238);
and I_37325 (I637272,I637088,I637255);
nand I_37326 (I636948,I637207,I637105);
DFFARX1 I_37327  ( .D(I260238), .CLK(I2702), .RSTB(I636986), .Q(I637303) );
or I_37328 (I636969,I637303,I637190);
nor I_37329 (I637334,I637303,I637071);
nor I_37330 (I637351,I637303,I637105);
nand I_37331 (I636954,I637037,I637351);
or I_37332 (I637382,I637303,I637272);
DFFARX1 I_37333  ( .D(I637382), .CLK(I2702), .RSTB(I636986), .Q(I636951) );
not I_37334 (I636957,I637303);
DFFARX1 I_37335  ( .D(I260217), .CLK(I2702), .RSTB(I636986), .Q(I637427) );
not I_37336 (I637444,I637427);
nor I_37337 (I637461,I637444,I637037);
DFFARX1 I_37338  ( .D(I637461), .CLK(I2702), .RSTB(I636986), .Q(I636963) );
nor I_37339 (I636978,I637303,I637444);
nor I_37340 (I636966,I637444,I637207);
not I_37341 (I637520,I637444);
and I_37342 (I637537,I637071,I637520);
nor I_37343 (I636972,I637207,I637537);
nand I_37344 (I636960,I637444,I637334);
not I_37345 (I637615,I2709);
not I_37346 (I637632,I21228);
nor I_37347 (I637649,I21231,I21240);
nand I_37348 (I637666,I637649,I21255);
nor I_37349 (I637683,I637632,I21231);
nand I_37350 (I637700,I637683,I21234);
not I_37351 (I637717,I21231);
not I_37352 (I637734,I637717);
not I_37353 (I637751,I21225);
nor I_37354 (I637768,I637751,I21249);
and I_37355 (I637785,I637768,I21237);
or I_37356 (I637802,I637785,I21243);
DFFARX1 I_37357  ( .D(I637802), .CLK(I2702), .RSTB(I637615), .Q(I637819) );
nand I_37358 (I637836,I637632,I21225);
or I_37359 (I637604,I637836,I637819);
not I_37360 (I637867,I637836);
nor I_37361 (I637884,I637819,I637867);
and I_37362 (I637901,I637717,I637884);
nand I_37363 (I637577,I637836,I637734);
DFFARX1 I_37364  ( .D(I21246), .CLK(I2702), .RSTB(I637615), .Q(I637932) );
or I_37365 (I637598,I637932,I637819);
nor I_37366 (I637963,I637932,I637700);
nor I_37367 (I637980,I637932,I637734);
nand I_37368 (I637583,I637666,I637980);
or I_37369 (I638011,I637932,I637901);
DFFARX1 I_37370  ( .D(I638011), .CLK(I2702), .RSTB(I637615), .Q(I637580) );
not I_37371 (I637586,I637932);
DFFARX1 I_37372  ( .D(I21252), .CLK(I2702), .RSTB(I637615), .Q(I638056) );
not I_37373 (I638073,I638056);
nor I_37374 (I638090,I638073,I637666);
DFFARX1 I_37375  ( .D(I638090), .CLK(I2702), .RSTB(I637615), .Q(I637592) );
nor I_37376 (I637607,I637932,I638073);
nor I_37377 (I637595,I638073,I637836);
not I_37378 (I638149,I638073);
and I_37379 (I638166,I637700,I638149);
nor I_37380 (I637601,I637836,I638166);
nand I_37381 (I637589,I638073,I637963);
not I_37382 (I638244,I2709);
not I_37383 (I638261,I138905);
nor I_37384 (I638278,I138923,I138902);
nand I_37385 (I638295,I638278,I138920);
nor I_37386 (I638312,I638261,I138923);
nand I_37387 (I638329,I638312,I138914);
not I_37388 (I638346,I138923);
not I_37389 (I638363,I638346);
not I_37390 (I638380,I138917);
nor I_37391 (I638397,I638380,I138911);
and I_37392 (I638414,I638397,I138908);
or I_37393 (I638431,I638414,I138899);
DFFARX1 I_37394  ( .D(I638431), .CLK(I2702), .RSTB(I638244), .Q(I638448) );
nand I_37395 (I638465,I638261,I138917);
or I_37396 (I638233,I638465,I638448);
not I_37397 (I638496,I638465);
nor I_37398 (I638513,I638448,I638496);
and I_37399 (I638530,I638346,I638513);
nand I_37400 (I638206,I638465,I638363);
DFFARX1 I_37401  ( .D(I138929), .CLK(I2702), .RSTB(I638244), .Q(I638561) );
or I_37402 (I638227,I638561,I638448);
nor I_37403 (I638592,I638561,I638329);
nor I_37404 (I638609,I638561,I638363);
nand I_37405 (I638212,I638295,I638609);
or I_37406 (I638640,I638561,I638530);
DFFARX1 I_37407  ( .D(I638640), .CLK(I2702), .RSTB(I638244), .Q(I638209) );
not I_37408 (I638215,I638561);
DFFARX1 I_37409  ( .D(I138926), .CLK(I2702), .RSTB(I638244), .Q(I638685) );
not I_37410 (I638702,I638685);
nor I_37411 (I638719,I638702,I638295);
DFFARX1 I_37412  ( .D(I638719), .CLK(I2702), .RSTB(I638244), .Q(I638221) );
nor I_37413 (I638236,I638561,I638702);
nor I_37414 (I638224,I638702,I638465);
not I_37415 (I638778,I638702);
and I_37416 (I638795,I638329,I638778);
nor I_37417 (I638230,I638465,I638795);
nand I_37418 (I638218,I638702,I638592);
not I_37419 (I638873,I2709);
not I_37420 (I638890,I349955);
nor I_37421 (I638907,I349964,I349967);
nand I_37422 (I638924,I638907,I349952);
nor I_37423 (I638941,I638890,I349964);
nand I_37424 (I638958,I638941,I349949);
not I_37425 (I638975,I349964);
not I_37426 (I638992,I638975);
not I_37427 (I639009,I349937);
nor I_37428 (I639026,I639009,I349943);
and I_37429 (I639043,I639026,I349940);
or I_37430 (I639060,I639043,I349961);
DFFARX1 I_37431  ( .D(I639060), .CLK(I2702), .RSTB(I638873), .Q(I639077) );
nand I_37432 (I639094,I638890,I349937);
or I_37433 (I638862,I639094,I639077);
not I_37434 (I639125,I639094);
nor I_37435 (I639142,I639077,I639125);
and I_37436 (I639159,I638975,I639142);
nand I_37437 (I638835,I639094,I638992);
DFFARX1 I_37438  ( .D(I349946), .CLK(I2702), .RSTB(I638873), .Q(I639190) );
or I_37439 (I638856,I639190,I639077);
nor I_37440 (I639221,I639190,I638958);
nor I_37441 (I639238,I639190,I638992);
nand I_37442 (I638841,I638924,I639238);
or I_37443 (I639269,I639190,I639159);
DFFARX1 I_37444  ( .D(I639269), .CLK(I2702), .RSTB(I638873), .Q(I638838) );
not I_37445 (I638844,I639190);
DFFARX1 I_37446  ( .D(I349958), .CLK(I2702), .RSTB(I638873), .Q(I639314) );
not I_37447 (I639331,I639314);
nor I_37448 (I639348,I639331,I638924);
DFFARX1 I_37449  ( .D(I639348), .CLK(I2702), .RSTB(I638873), .Q(I638850) );
nor I_37450 (I638865,I639190,I639331);
nor I_37451 (I638853,I639331,I639094);
not I_37452 (I639407,I639331);
and I_37453 (I639424,I638958,I639407);
nor I_37454 (I638859,I639094,I639424);
nand I_37455 (I638847,I639331,I639221);
not I_37456 (I639502,I2709);
not I_37457 (I639519,I443705);
nor I_37458 (I639536,I443678,I443696);
nand I_37459 (I639553,I639536,I443681);
nor I_37460 (I639570,I639519,I443678);
nand I_37461 (I639587,I639570,I443699);
not I_37462 (I639604,I443678);
not I_37463 (I639621,I639604);
not I_37464 (I639638,I443675);
nor I_37465 (I639655,I639638,I443702);
and I_37466 (I639672,I639655,I443693);
or I_37467 (I639689,I639672,I443684);
DFFARX1 I_37468  ( .D(I639689), .CLK(I2702), .RSTB(I639502), .Q(I639706) );
nand I_37469 (I639723,I639519,I443675);
or I_37470 (I639491,I639723,I639706);
not I_37471 (I639754,I639723);
nor I_37472 (I639771,I639706,I639754);
and I_37473 (I639788,I639604,I639771);
nand I_37474 (I639464,I639723,I639621);
DFFARX1 I_37475  ( .D(I443687), .CLK(I2702), .RSTB(I639502), .Q(I639819) );
or I_37476 (I639485,I639819,I639706);
nor I_37477 (I639850,I639819,I639587);
nor I_37478 (I639867,I639819,I639621);
nand I_37479 (I639470,I639553,I639867);
or I_37480 (I639898,I639819,I639788);
DFFARX1 I_37481  ( .D(I639898), .CLK(I2702), .RSTB(I639502), .Q(I639467) );
not I_37482 (I639473,I639819);
DFFARX1 I_37483  ( .D(I443690), .CLK(I2702), .RSTB(I639502), .Q(I639943) );
not I_37484 (I639960,I639943);
nor I_37485 (I639977,I639960,I639553);
DFFARX1 I_37486  ( .D(I639977), .CLK(I2702), .RSTB(I639502), .Q(I639479) );
nor I_37487 (I639494,I639819,I639960);
nor I_37488 (I639482,I639960,I639723);
not I_37489 (I640036,I639960);
and I_37490 (I640053,I639587,I640036);
nor I_37491 (I639488,I639723,I640053);
nand I_37492 (I639476,I639960,I639850);
not I_37493 (I640131,I2709);
not I_37494 (I640148,I383547);
nor I_37495 (I640165,I383556,I383559);
nand I_37496 (I640182,I640165,I383544);
nor I_37497 (I640199,I640148,I383556);
nand I_37498 (I640216,I640199,I383541);
not I_37499 (I640233,I383556);
not I_37500 (I640250,I640233);
not I_37501 (I640267,I383529);
nor I_37502 (I640284,I640267,I383535);
and I_37503 (I640301,I640284,I383532);
or I_37504 (I640318,I640301,I383553);
DFFARX1 I_37505  ( .D(I640318), .CLK(I2702), .RSTB(I640131), .Q(I640335) );
nand I_37506 (I640352,I640148,I383529);
or I_37507 (I640120,I640352,I640335);
not I_37508 (I640383,I640352);
nor I_37509 (I640400,I640335,I640383);
and I_37510 (I640417,I640233,I640400);
nand I_37511 (I640093,I640352,I640250);
DFFARX1 I_37512  ( .D(I383538), .CLK(I2702), .RSTB(I640131), .Q(I640448) );
or I_37513 (I640114,I640448,I640335);
nor I_37514 (I640479,I640448,I640216);
nor I_37515 (I640496,I640448,I640250);
nand I_37516 (I640099,I640182,I640496);
or I_37517 (I640527,I640448,I640417);
DFFARX1 I_37518  ( .D(I640527), .CLK(I2702), .RSTB(I640131), .Q(I640096) );
not I_37519 (I640102,I640448);
DFFARX1 I_37520  ( .D(I383550), .CLK(I2702), .RSTB(I640131), .Q(I640572) );
not I_37521 (I640589,I640572);
nor I_37522 (I640606,I640589,I640182);
DFFARX1 I_37523  ( .D(I640606), .CLK(I2702), .RSTB(I640131), .Q(I640108) );
nor I_37524 (I640123,I640448,I640589);
nor I_37525 (I640111,I640589,I640352);
not I_37526 (I640665,I640589);
and I_37527 (I640682,I640216,I640665);
nor I_37528 (I640117,I640352,I640682);
nand I_37529 (I640105,I640589,I640479);
not I_37530 (I640760,I2709);
not I_37531 (I640777,I531010);
nor I_37532 (I640794,I531028,I531007);
nand I_37533 (I640811,I640794,I531031);
nor I_37534 (I640828,I640777,I531028);
nand I_37535 (I640845,I640828,I531025);
not I_37536 (I640862,I531028);
not I_37537 (I640879,I640862);
not I_37538 (I640896,I531016);
nor I_37539 (I640913,I640896,I531004);
and I_37540 (I640930,I640913,I531022);
or I_37541 (I640947,I640930,I531034);
DFFARX1 I_37542  ( .D(I640947), .CLK(I2702), .RSTB(I640760), .Q(I640964) );
nand I_37543 (I640981,I640777,I531016);
or I_37544 (I640749,I640981,I640964);
not I_37545 (I641012,I640981);
nor I_37546 (I641029,I640964,I641012);
and I_37547 (I641046,I640862,I641029);
nand I_37548 (I640722,I640981,I640879);
DFFARX1 I_37549  ( .D(I531013), .CLK(I2702), .RSTB(I640760), .Q(I641077) );
or I_37550 (I640743,I641077,I640964);
nor I_37551 (I641108,I641077,I640845);
nor I_37552 (I641125,I641077,I640879);
nand I_37553 (I640728,I640811,I641125);
or I_37554 (I641156,I641077,I641046);
DFFARX1 I_37555  ( .D(I641156), .CLK(I2702), .RSTB(I640760), .Q(I640725) );
not I_37556 (I640731,I641077);
DFFARX1 I_37557  ( .D(I531019), .CLK(I2702), .RSTB(I640760), .Q(I641201) );
not I_37558 (I641218,I641201);
nor I_37559 (I641235,I641218,I640811);
DFFARX1 I_37560  ( .D(I641235), .CLK(I2702), .RSTB(I640760), .Q(I640737) );
nor I_37561 (I640752,I641077,I641218);
nor I_37562 (I640740,I641218,I640981);
not I_37563 (I641294,I641218);
and I_37564 (I641311,I640845,I641294);
nor I_37565 (I640746,I640981,I641311);
nand I_37566 (I640734,I641218,I641108);
not I_37567 (I641389,I2709);
not I_37568 (I641406,I706552);
nor I_37569 (I641423,I706576,I706561);
nand I_37570 (I641440,I641423,I706546);
nor I_37571 (I641457,I641406,I706576);
nand I_37572 (I641474,I641457,I706573);
not I_37573 (I641491,I706576);
not I_37574 (I641508,I641491);
not I_37575 (I641525,I706555);
nor I_37576 (I641542,I641525,I706549);
and I_37577 (I641559,I641542,I706570);
or I_37578 (I641576,I641559,I706558);
DFFARX1 I_37579  ( .D(I641576), .CLK(I2702), .RSTB(I641389), .Q(I641593) );
nand I_37580 (I641610,I641406,I706555);
or I_37581 (I641378,I641610,I641593);
not I_37582 (I641641,I641610);
nor I_37583 (I641658,I641593,I641641);
and I_37584 (I641675,I641491,I641658);
nand I_37585 (I641351,I641610,I641508);
DFFARX1 I_37586  ( .D(I706567), .CLK(I2702), .RSTB(I641389), .Q(I641706) );
or I_37587 (I641372,I641706,I641593);
nor I_37588 (I641737,I641706,I641474);
nor I_37589 (I641754,I641706,I641508);
nand I_37590 (I641357,I641440,I641754);
or I_37591 (I641785,I641706,I641675);
DFFARX1 I_37592  ( .D(I641785), .CLK(I2702), .RSTB(I641389), .Q(I641354) );
not I_37593 (I641360,I641706);
DFFARX1 I_37594  ( .D(I706564), .CLK(I2702), .RSTB(I641389), .Q(I641830) );
not I_37595 (I641847,I641830);
nor I_37596 (I641864,I641847,I641440);
DFFARX1 I_37597  ( .D(I641864), .CLK(I2702), .RSTB(I641389), .Q(I641366) );
nor I_37598 (I641381,I641706,I641847);
nor I_37599 (I641369,I641847,I641610);
not I_37600 (I641923,I641847);
and I_37601 (I641940,I641474,I641923);
nor I_37602 (I641375,I641610,I641940);
nand I_37603 (I641363,I641847,I641737);
not I_37604 (I642018,I2709);
not I_37605 (I642035,I37497);
nor I_37606 (I642052,I37500,I37509);
nand I_37607 (I642069,I642052,I37524);
nor I_37608 (I642086,I642035,I37500);
nand I_37609 (I642103,I642086,I37503);
not I_37610 (I642120,I37500);
not I_37611 (I642137,I642120);
not I_37612 (I642154,I37494);
nor I_37613 (I642171,I642154,I37518);
and I_37614 (I642188,I642171,I37506);
or I_37615 (I642205,I642188,I37512);
DFFARX1 I_37616  ( .D(I642205), .CLK(I2702), .RSTB(I642018), .Q(I642222) );
nand I_37617 (I642239,I642035,I37494);
or I_37618 (I642007,I642239,I642222);
not I_37619 (I642270,I642239);
nor I_37620 (I642287,I642222,I642270);
and I_37621 (I642304,I642120,I642287);
nand I_37622 (I641980,I642239,I642137);
DFFARX1 I_37623  ( .D(I37515), .CLK(I2702), .RSTB(I642018), .Q(I642335) );
or I_37624 (I642001,I642335,I642222);
nor I_37625 (I642366,I642335,I642103);
nor I_37626 (I642383,I642335,I642137);
nand I_37627 (I641986,I642069,I642383);
or I_37628 (I642414,I642335,I642304);
DFFARX1 I_37629  ( .D(I642414), .CLK(I2702), .RSTB(I642018), .Q(I641983) );
not I_37630 (I641989,I642335);
DFFARX1 I_37631  ( .D(I37521), .CLK(I2702), .RSTB(I642018), .Q(I642459) );
not I_37632 (I642476,I642459);
nor I_37633 (I642493,I642476,I642069);
DFFARX1 I_37634  ( .D(I642493), .CLK(I2702), .RSTB(I642018), .Q(I641995) );
nor I_37635 (I642010,I642335,I642476);
nor I_37636 (I641998,I642476,I642239);
not I_37637 (I642552,I642476);
and I_37638 (I642569,I642103,I642552);
nor I_37639 (I642004,I642239,I642569);
nand I_37640 (I641992,I642476,I642366);
not I_37641 (I642647,I2709);
not I_37642 (I642664,I696726);
nor I_37643 (I642681,I696750,I696735);
nand I_37644 (I642698,I642681,I696720);
nor I_37645 (I642715,I642664,I696750);
nand I_37646 (I642732,I642715,I696747);
not I_37647 (I642749,I696750);
not I_37648 (I642766,I642749);
not I_37649 (I642783,I696729);
nor I_37650 (I642800,I642783,I696723);
and I_37651 (I642817,I642800,I696744);
or I_37652 (I642834,I642817,I696732);
DFFARX1 I_37653  ( .D(I642834), .CLK(I2702), .RSTB(I642647), .Q(I642851) );
nand I_37654 (I642868,I642664,I696729);
or I_37655 (I642636,I642868,I642851);
not I_37656 (I642899,I642868);
nor I_37657 (I642916,I642851,I642899);
and I_37658 (I642933,I642749,I642916);
nand I_37659 (I642609,I642868,I642766);
DFFARX1 I_37660  ( .D(I696741), .CLK(I2702), .RSTB(I642647), .Q(I642964) );
or I_37661 (I642630,I642964,I642851);
nor I_37662 (I642995,I642964,I642732);
nor I_37663 (I643012,I642964,I642766);
nand I_37664 (I642615,I642698,I643012);
or I_37665 (I643043,I642964,I642933);
DFFARX1 I_37666  ( .D(I643043), .CLK(I2702), .RSTB(I642647), .Q(I642612) );
not I_37667 (I642618,I642964);
DFFARX1 I_37668  ( .D(I696738), .CLK(I2702), .RSTB(I642647), .Q(I643088) );
not I_37669 (I643105,I643088);
nor I_37670 (I643122,I643105,I642698);
DFFARX1 I_37671  ( .D(I643122), .CLK(I2702), .RSTB(I642647), .Q(I642624) );
nor I_37672 (I642639,I642964,I643105);
nor I_37673 (I642627,I643105,I642868);
not I_37674 (I643181,I643105);
and I_37675 (I643198,I642732,I643181);
nor I_37676 (I642633,I642868,I643198);
nand I_37677 (I642621,I643105,I642995);
not I_37678 (I643276,I2709);
not I_37679 (I643293,I470871);
nor I_37680 (I643310,I470844,I470862);
nand I_37681 (I643327,I643310,I470847);
nor I_37682 (I643344,I643293,I470844);
nand I_37683 (I643361,I643344,I470865);
not I_37684 (I643378,I470844);
not I_37685 (I643395,I643378);
not I_37686 (I643412,I470841);
nor I_37687 (I643429,I643412,I470868);
and I_37688 (I643446,I643429,I470859);
or I_37689 (I643463,I643446,I470850);
DFFARX1 I_37690  ( .D(I643463), .CLK(I2702), .RSTB(I643276), .Q(I643480) );
nand I_37691 (I643497,I643293,I470841);
or I_37692 (I643265,I643497,I643480);
not I_37693 (I643528,I643497);
nor I_37694 (I643545,I643480,I643528);
and I_37695 (I643562,I643378,I643545);
nand I_37696 (I643238,I643497,I643395);
DFFARX1 I_37697  ( .D(I470853), .CLK(I2702), .RSTB(I643276), .Q(I643593) );
or I_37698 (I643259,I643593,I643480);
nor I_37699 (I643624,I643593,I643361);
nor I_37700 (I643641,I643593,I643395);
nand I_37701 (I643244,I643327,I643641);
or I_37702 (I643672,I643593,I643562);
DFFARX1 I_37703  ( .D(I643672), .CLK(I2702), .RSTB(I643276), .Q(I643241) );
not I_37704 (I643247,I643593);
DFFARX1 I_37705  ( .D(I470856), .CLK(I2702), .RSTB(I643276), .Q(I643717) );
not I_37706 (I643734,I643717);
nor I_37707 (I643751,I643734,I643327);
DFFARX1 I_37708  ( .D(I643751), .CLK(I2702), .RSTB(I643276), .Q(I643253) );
nor I_37709 (I643268,I643593,I643734);
nor I_37710 (I643256,I643734,I643497);
not I_37711 (I643810,I643734);
and I_37712 (I643827,I643361,I643810);
nor I_37713 (I643262,I643497,I643827);
nand I_37714 (I643250,I643734,I643624);
not I_37715 (I643905,I2709);
not I_37716 (I643922,I302661);
nor I_37717 (I643939,I302667,I302646);
nand I_37718 (I643956,I643939,I302652);
nor I_37719 (I643973,I643922,I302667);
nand I_37720 (I643990,I643973,I302658);
not I_37721 (I644007,I302667);
not I_37722 (I644024,I644007);
not I_37723 (I644041,I302655);
nor I_37724 (I644058,I644041,I302673);
and I_37725 (I644075,I644058,I302664);
or I_37726 (I644092,I644075,I302643);
DFFARX1 I_37727  ( .D(I644092), .CLK(I2702), .RSTB(I643905), .Q(I644109) );
nand I_37728 (I644126,I643922,I302655);
or I_37729 (I643894,I644126,I644109);
not I_37730 (I644157,I644126);
nor I_37731 (I644174,I644109,I644157);
and I_37732 (I644191,I644007,I644174);
nand I_37733 (I643867,I644126,I644024);
DFFARX1 I_37734  ( .D(I302670), .CLK(I2702), .RSTB(I643905), .Q(I644222) );
or I_37735 (I643888,I644222,I644109);
nor I_37736 (I644253,I644222,I643990);
nor I_37737 (I644270,I644222,I644024);
nand I_37738 (I643873,I643956,I644270);
or I_37739 (I644301,I644222,I644191);
DFFARX1 I_37740  ( .D(I644301), .CLK(I2702), .RSTB(I643905), .Q(I643870) );
not I_37741 (I643876,I644222);
DFFARX1 I_37742  ( .D(I302649), .CLK(I2702), .RSTB(I643905), .Q(I644346) );
not I_37743 (I644363,I644346);
nor I_37744 (I644380,I644363,I643956);
DFFARX1 I_37745  ( .D(I644380), .CLK(I2702), .RSTB(I643905), .Q(I643882) );
nor I_37746 (I643897,I644222,I644363);
nor I_37747 (I643885,I644363,I644126);
not I_37748 (I644439,I644363);
and I_37749 (I644456,I643990,I644439);
nor I_37750 (I643891,I644126,I644456);
nand I_37751 (I643879,I644363,I644253);
not I_37752 (I644534,I2709);
not I_37753 (I644551,I171381);
nor I_37754 (I644568,I171372,I171396);
nand I_37755 (I644585,I644568,I171399);
nor I_37756 (I644602,I644551,I171372);
nand I_37757 (I644619,I644602,I171390);
not I_37758 (I644636,I171372);
not I_37759 (I644653,I644636);
not I_37760 (I644670,I171384);
nor I_37761 (I644687,I644670,I171378);
and I_37762 (I644704,I644687,I171387);
or I_37763 (I644721,I644704,I171375);
DFFARX1 I_37764  ( .D(I644721), .CLK(I2702), .RSTB(I644534), .Q(I644738) );
nand I_37765 (I644755,I644551,I171384);
or I_37766 (I644523,I644755,I644738);
not I_37767 (I644786,I644755);
nor I_37768 (I644803,I644738,I644786);
and I_37769 (I644820,I644636,I644803);
nand I_37770 (I644496,I644755,I644653);
DFFARX1 I_37771  ( .D(I171369), .CLK(I2702), .RSTB(I644534), .Q(I644851) );
or I_37772 (I644517,I644851,I644738);
nor I_37773 (I644882,I644851,I644619);
nor I_37774 (I644899,I644851,I644653);
nand I_37775 (I644502,I644585,I644899);
or I_37776 (I644930,I644851,I644820);
DFFARX1 I_37777  ( .D(I644930), .CLK(I2702), .RSTB(I644534), .Q(I644499) );
not I_37778 (I644505,I644851);
DFFARX1 I_37779  ( .D(I171393), .CLK(I2702), .RSTB(I644534), .Q(I644975) );
not I_37780 (I644992,I644975);
nor I_37781 (I645009,I644992,I644585);
DFFARX1 I_37782  ( .D(I645009), .CLK(I2702), .RSTB(I644534), .Q(I644511) );
nor I_37783 (I644526,I644851,I644992);
nor I_37784 (I644514,I644992,I644755);
not I_37785 (I645068,I644992);
and I_37786 (I645085,I644619,I645068);
nor I_37787 (I644520,I644755,I645085);
nand I_37788 (I644508,I644992,I644882);
not I_37789 (I645163,I2709);
not I_37790 (I645180,I337681);
nor I_37791 (I645197,I337690,I337693);
nand I_37792 (I645214,I645197,I337678);
nor I_37793 (I645231,I645180,I337690);
nand I_37794 (I645248,I645231,I337675);
not I_37795 (I645265,I337690);
not I_37796 (I645282,I645265);
not I_37797 (I645299,I337663);
nor I_37798 (I645316,I645299,I337669);
and I_37799 (I645333,I645316,I337666);
or I_37800 (I645350,I645333,I337687);
DFFARX1 I_37801  ( .D(I645350), .CLK(I2702), .RSTB(I645163), .Q(I645367) );
nand I_37802 (I645384,I645180,I337663);
or I_37803 (I645152,I645384,I645367);
not I_37804 (I645415,I645384);
nor I_37805 (I645432,I645367,I645415);
and I_37806 (I645449,I645265,I645432);
nand I_37807 (I645125,I645384,I645282);
DFFARX1 I_37808  ( .D(I337672), .CLK(I2702), .RSTB(I645163), .Q(I645480) );
or I_37809 (I645146,I645480,I645367);
nor I_37810 (I645511,I645480,I645248);
nor I_37811 (I645528,I645480,I645282);
nand I_37812 (I645131,I645214,I645528);
or I_37813 (I645559,I645480,I645449);
DFFARX1 I_37814  ( .D(I645559), .CLK(I2702), .RSTB(I645163), .Q(I645128) );
not I_37815 (I645134,I645480);
DFFARX1 I_37816  ( .D(I337684), .CLK(I2702), .RSTB(I645163), .Q(I645604) );
not I_37817 (I645621,I645604);
nor I_37818 (I645638,I645621,I645214);
DFFARX1 I_37819  ( .D(I645638), .CLK(I2702), .RSTB(I645163), .Q(I645140) );
nor I_37820 (I645155,I645480,I645621);
nor I_37821 (I645143,I645621,I645384);
not I_37822 (I645697,I645621);
and I_37823 (I645714,I645248,I645697);
nor I_37824 (I645149,I645384,I645714);
nand I_37825 (I645137,I645621,I645511);
not I_37826 (I645792,I2709);
not I_37827 (I645809,I2055);
nor I_37828 (I645826,I1287,I2167);
nand I_37829 (I645843,I645826,I2279);
nor I_37830 (I645860,I645809,I1287);
nand I_37831 (I645877,I645860,I2031);
not I_37832 (I645894,I1287);
not I_37833 (I645911,I645894);
not I_37834 (I645928,I2639);
nor I_37835 (I645945,I645928,I2215);
and I_37836 (I645962,I645945,I1575);
or I_37837 (I645979,I645962,I2303);
DFFARX1 I_37838  ( .D(I645979), .CLK(I2702), .RSTB(I645792), .Q(I645996) );
nand I_37839 (I646013,I645809,I2639);
or I_37840 (I645781,I646013,I645996);
not I_37841 (I646044,I646013);
nor I_37842 (I646061,I645996,I646044);
and I_37843 (I646078,I645894,I646061);
nand I_37844 (I645754,I646013,I645911);
DFFARX1 I_37845  ( .D(I2271), .CLK(I2702), .RSTB(I645792), .Q(I646109) );
or I_37846 (I645775,I646109,I645996);
nor I_37847 (I646140,I646109,I645877);
nor I_37848 (I646157,I646109,I645911);
nand I_37849 (I645760,I645843,I646157);
or I_37850 (I646188,I646109,I646078);
DFFARX1 I_37851  ( .D(I646188), .CLK(I2702), .RSTB(I645792), .Q(I645757) );
not I_37852 (I645763,I646109);
DFFARX1 I_37853  ( .D(I1263), .CLK(I2702), .RSTB(I645792), .Q(I646233) );
not I_37854 (I646250,I646233);
nor I_37855 (I646267,I646250,I645843);
DFFARX1 I_37856  ( .D(I646267), .CLK(I2702), .RSTB(I645792), .Q(I645769) );
nor I_37857 (I645784,I646109,I646250);
nor I_37858 (I645772,I646250,I646013);
not I_37859 (I646326,I646250);
and I_37860 (I646343,I645877,I646326);
nor I_37861 (I645778,I646013,I646343);
nand I_37862 (I645766,I646250,I646140);
not I_37863 (I646421,I2709);
not I_37864 (I646438,I110481);
nor I_37865 (I646455,I110499,I110478);
nand I_37866 (I646472,I646455,I110496);
nor I_37867 (I646489,I646438,I110499);
nand I_37868 (I646506,I646489,I110490);
not I_37869 (I646523,I110499);
not I_37870 (I646540,I646523);
not I_37871 (I646557,I110493);
nor I_37872 (I646574,I646557,I110487);
and I_37873 (I646591,I646574,I110484);
or I_37874 (I646608,I646591,I110475);
DFFARX1 I_37875  ( .D(I646608), .CLK(I2702), .RSTB(I646421), .Q(I646625) );
nand I_37876 (I646642,I646438,I110493);
or I_37877 (I646410,I646642,I646625);
not I_37878 (I646673,I646642);
nor I_37879 (I646690,I646625,I646673);
and I_37880 (I646707,I646523,I646690);
nand I_37881 (I646383,I646642,I646540);
DFFARX1 I_37882  ( .D(I110505), .CLK(I2702), .RSTB(I646421), .Q(I646738) );
or I_37883 (I646404,I646738,I646625);
nor I_37884 (I646769,I646738,I646506);
nor I_37885 (I646786,I646738,I646540);
nand I_37886 (I646389,I646472,I646786);
or I_37887 (I646817,I646738,I646707);
DFFARX1 I_37888  ( .D(I646817), .CLK(I2702), .RSTB(I646421), .Q(I646386) );
not I_37889 (I646392,I646738);
DFFARX1 I_37890  ( .D(I110502), .CLK(I2702), .RSTB(I646421), .Q(I646862) );
not I_37891 (I646879,I646862);
nor I_37892 (I646896,I646879,I646472);
DFFARX1 I_37893  ( .D(I646896), .CLK(I2702), .RSTB(I646421), .Q(I646398) );
nor I_37894 (I646413,I646738,I646879);
nor I_37895 (I646401,I646879,I646642);
not I_37896 (I646955,I646879);
and I_37897 (I646972,I646506,I646955);
nor I_37898 (I646407,I646642,I646972);
nand I_37899 (I646395,I646879,I646769);
not I_37900 (I647050,I2709);
not I_37901 (I647067,I202288);
nor I_37902 (I647084,I202264,I202279);
nand I_37903 (I647101,I647084,I202261);
nor I_37904 (I647118,I647067,I202264);
nand I_37905 (I647135,I647118,I202276);
not I_37906 (I647152,I202264);
not I_37907 (I647169,I647152);
not I_37908 (I647186,I202267);
nor I_37909 (I647203,I647186,I202282);
and I_37910 (I647220,I647203,I202273);
or I_37911 (I647237,I647220,I202258);
DFFARX1 I_37912  ( .D(I647237), .CLK(I2702), .RSTB(I647050), .Q(I647254) );
nand I_37913 (I647271,I647067,I202267);
or I_37914 (I647039,I647271,I647254);
not I_37915 (I647302,I647271);
nor I_37916 (I647319,I647254,I647302);
and I_37917 (I647336,I647152,I647319);
nand I_37918 (I647012,I647271,I647169);
DFFARX1 I_37919  ( .D(I202270), .CLK(I2702), .RSTB(I647050), .Q(I647367) );
or I_37920 (I647033,I647367,I647254);
nor I_37921 (I647398,I647367,I647135);
nor I_37922 (I647415,I647367,I647169);
nand I_37923 (I647018,I647101,I647415);
or I_37924 (I647446,I647367,I647336);
DFFARX1 I_37925  ( .D(I647446), .CLK(I2702), .RSTB(I647050), .Q(I647015) );
not I_37926 (I647021,I647367);
DFFARX1 I_37927  ( .D(I202285), .CLK(I2702), .RSTB(I647050), .Q(I647491) );
not I_37928 (I647508,I647491);
nor I_37929 (I647525,I647508,I647101);
DFFARX1 I_37930  ( .D(I647525), .CLK(I2702), .RSTB(I647050), .Q(I647027) );
nor I_37931 (I647042,I647367,I647508);
nor I_37932 (I647030,I647508,I647271);
not I_37933 (I647584,I647508);
and I_37934 (I647601,I647135,I647584);
nor I_37935 (I647036,I647271,I647601);
nand I_37936 (I647024,I647508,I647398);
not I_37937 (I647679,I2709);
not I_37938 (I647696,I481853);
nor I_37939 (I647713,I481826,I481844);
nand I_37940 (I647730,I647713,I481829);
nor I_37941 (I647747,I647696,I481826);
nand I_37942 (I647764,I647747,I481847);
not I_37943 (I647781,I481826);
not I_37944 (I647798,I647781);
not I_37945 (I647815,I481823);
nor I_37946 (I647832,I647815,I481850);
and I_37947 (I647849,I647832,I481841);
or I_37948 (I647866,I647849,I481832);
DFFARX1 I_37949  ( .D(I647866), .CLK(I2702), .RSTB(I647679), .Q(I647883) );
nand I_37950 (I647900,I647696,I481823);
or I_37951 (I647668,I647900,I647883);
not I_37952 (I647931,I647900);
nor I_37953 (I647948,I647883,I647931);
and I_37954 (I647965,I647781,I647948);
nand I_37955 (I647641,I647900,I647798);
DFFARX1 I_37956  ( .D(I481835), .CLK(I2702), .RSTB(I647679), .Q(I647996) );
or I_37957 (I647662,I647996,I647883);
nor I_37958 (I648027,I647996,I647764);
nor I_37959 (I648044,I647996,I647798);
nand I_37960 (I647647,I647730,I648044);
or I_37961 (I648075,I647996,I647965);
DFFARX1 I_37962  ( .D(I648075), .CLK(I2702), .RSTB(I647679), .Q(I647644) );
not I_37963 (I647650,I647996);
DFFARX1 I_37964  ( .D(I481838), .CLK(I2702), .RSTB(I647679), .Q(I648120) );
not I_37965 (I648137,I648120);
nor I_37966 (I648154,I648137,I647730);
DFFARX1 I_37967  ( .D(I648154), .CLK(I2702), .RSTB(I647679), .Q(I647656) );
nor I_37968 (I647671,I647996,I648137);
nor I_37969 (I647659,I648137,I647900);
not I_37970 (I648213,I648137);
and I_37971 (I648230,I647764,I648213);
nor I_37972 (I647665,I647900,I648230);
nand I_37973 (I647653,I648137,I648027);
not I_37974 (I648308,I2709);
not I_37975 (I648325,I218353);
nor I_37976 (I648342,I218329,I218344);
nand I_37977 (I648359,I648342,I218326);
nor I_37978 (I648376,I648325,I218329);
nand I_37979 (I648393,I648376,I218341);
not I_37980 (I648410,I218329);
not I_37981 (I648427,I648410);
not I_37982 (I648444,I218332);
nor I_37983 (I648461,I648444,I218347);
and I_37984 (I648478,I648461,I218338);
or I_37985 (I648495,I648478,I218323);
DFFARX1 I_37986  ( .D(I648495), .CLK(I2702), .RSTB(I648308), .Q(I648512) );
nand I_37987 (I648529,I648325,I218332);
or I_37988 (I648297,I648529,I648512);
not I_37989 (I648560,I648529);
nor I_37990 (I648577,I648512,I648560);
and I_37991 (I648594,I648410,I648577);
nand I_37992 (I648270,I648529,I648427);
DFFARX1 I_37993  ( .D(I218335), .CLK(I2702), .RSTB(I648308), .Q(I648625) );
or I_37994 (I648291,I648625,I648512);
nor I_37995 (I648656,I648625,I648393);
nor I_37996 (I648673,I648625,I648427);
nand I_37997 (I648276,I648359,I648673);
or I_37998 (I648704,I648625,I648594);
DFFARX1 I_37999  ( .D(I648704), .CLK(I2702), .RSTB(I648308), .Q(I648273) );
not I_38000 (I648279,I648625);
DFFARX1 I_38001  ( .D(I218350), .CLK(I2702), .RSTB(I648308), .Q(I648749) );
not I_38002 (I648766,I648749);
nor I_38003 (I648783,I648766,I648359);
DFFARX1 I_38004  ( .D(I648783), .CLK(I2702), .RSTB(I648308), .Q(I648285) );
nor I_38005 (I648300,I648625,I648766);
nor I_38006 (I648288,I648766,I648529);
not I_38007 (I648842,I648766);
and I_38008 (I648859,I648393,I648842);
nor I_38009 (I648294,I648529,I648859);
nand I_38010 (I648282,I648766,I648656);
not I_38011 (I648937,I2709);
not I_38012 (I648954,I239773);
nor I_38013 (I648971,I239743,I239746);
nand I_38014 (I648988,I648971,I239764);
nor I_38015 (I649005,I648954,I239743);
nand I_38016 (I649022,I649005,I239770);
not I_38017 (I649039,I239743);
not I_38018 (I649056,I649039);
not I_38019 (I649073,I239767);
nor I_38020 (I649090,I649073,I239752);
and I_38021 (I649107,I649090,I239761);
or I_38022 (I649124,I649107,I239758);
DFFARX1 I_38023  ( .D(I649124), .CLK(I2702), .RSTB(I648937), .Q(I649141) );
nand I_38024 (I649158,I648954,I239767);
or I_38025 (I648926,I649158,I649141);
not I_38026 (I649189,I649158);
nor I_38027 (I649206,I649141,I649189);
and I_38028 (I649223,I649039,I649206);
nand I_38029 (I648899,I649158,I649056);
DFFARX1 I_38030  ( .D(I239749), .CLK(I2702), .RSTB(I648937), .Q(I649254) );
or I_38031 (I648920,I649254,I649141);
nor I_38032 (I649285,I649254,I649022);
nor I_38033 (I649302,I649254,I649056);
nand I_38034 (I648905,I648988,I649302);
or I_38035 (I649333,I649254,I649223);
DFFARX1 I_38036  ( .D(I649333), .CLK(I2702), .RSTB(I648937), .Q(I648902) );
not I_38037 (I648908,I649254);
DFFARX1 I_38038  ( .D(I239755), .CLK(I2702), .RSTB(I648937), .Q(I649378) );
not I_38039 (I649395,I649378);
nor I_38040 (I649412,I649395,I648988);
DFFARX1 I_38041  ( .D(I649412), .CLK(I2702), .RSTB(I648937), .Q(I648914) );
nor I_38042 (I648929,I649254,I649395);
nor I_38043 (I648917,I649395,I649158);
not I_38044 (I649471,I649395);
and I_38045 (I649488,I649022,I649471);
nor I_38046 (I648923,I649158,I649488);
nand I_38047 (I648911,I649395,I649285);
not I_38048 (I649566,I2709);
not I_38049 (I649583,I489485);
nor I_38050 (I649600,I489476,I489503);
nand I_38051 (I649617,I649600,I489473);
nor I_38052 (I649634,I649583,I489476);
nand I_38053 (I649651,I649634,I489497);
not I_38054 (I649668,I489476);
not I_38055 (I649685,I649668);
not I_38056 (I649702,I489482);
nor I_38057 (I649719,I649702,I489500);
and I_38058 (I649736,I649719,I489491);
or I_38059 (I649753,I649736,I489488);
DFFARX1 I_38060  ( .D(I649753), .CLK(I2702), .RSTB(I649566), .Q(I649770) );
nand I_38061 (I649787,I649583,I489482);
or I_38062 (I649555,I649787,I649770);
not I_38063 (I649818,I649787);
nor I_38064 (I649835,I649770,I649818);
and I_38065 (I649852,I649668,I649835);
nand I_38066 (I649528,I649787,I649685);
DFFARX1 I_38067  ( .D(I489479), .CLK(I2702), .RSTB(I649566), .Q(I649883) );
or I_38068 (I649549,I649883,I649770);
nor I_38069 (I649914,I649883,I649651);
nor I_38070 (I649931,I649883,I649685);
nand I_38071 (I649534,I649617,I649931);
or I_38072 (I649962,I649883,I649852);
DFFARX1 I_38073  ( .D(I649962), .CLK(I2702), .RSTB(I649566), .Q(I649531) );
not I_38074 (I649537,I649883);
DFFARX1 I_38075  ( .D(I489494), .CLK(I2702), .RSTB(I649566), .Q(I650007) );
not I_38076 (I650024,I650007);
nor I_38077 (I650041,I650024,I649617);
DFFARX1 I_38078  ( .D(I650041), .CLK(I2702), .RSTB(I649566), .Q(I649543) );
nor I_38079 (I649558,I649883,I650024);
nor I_38080 (I649546,I650024,I649787);
not I_38081 (I650100,I650024);
and I_38082 (I650117,I649651,I650100);
nor I_38083 (I649552,I649787,I650117);
nand I_38084 (I649540,I650024,I649914);
not I_38085 (I650195,I2709);
not I_38086 (I650212,I723892);
nor I_38087 (I650229,I723916,I723901);
nand I_38088 (I650246,I650229,I723886);
nor I_38089 (I650263,I650212,I723916);
nand I_38090 (I650280,I650263,I723913);
not I_38091 (I650297,I723916);
not I_38092 (I650314,I650297);
not I_38093 (I650331,I723895);
nor I_38094 (I650348,I650331,I723889);
and I_38095 (I650365,I650348,I723910);
or I_38096 (I650382,I650365,I723898);
DFFARX1 I_38097  ( .D(I650382), .CLK(I2702), .RSTB(I650195), .Q(I650399) );
nand I_38098 (I650416,I650212,I723895);
or I_38099 (I650184,I650416,I650399);
not I_38100 (I650447,I650416);
nor I_38101 (I650464,I650399,I650447);
and I_38102 (I650481,I650297,I650464);
nand I_38103 (I650157,I650416,I650314);
DFFARX1 I_38104  ( .D(I723907), .CLK(I2702), .RSTB(I650195), .Q(I650512) );
or I_38105 (I650178,I650512,I650399);
nor I_38106 (I650543,I650512,I650280);
nor I_38107 (I650560,I650512,I650314);
nand I_38108 (I650163,I650246,I650560);
or I_38109 (I650591,I650512,I650481);
DFFARX1 I_38110  ( .D(I650591), .CLK(I2702), .RSTB(I650195), .Q(I650160) );
not I_38111 (I650166,I650512);
DFFARX1 I_38112  ( .D(I723904), .CLK(I2702), .RSTB(I650195), .Q(I650636) );
not I_38113 (I650653,I650636);
nor I_38114 (I650670,I650653,I650246);
DFFARX1 I_38115  ( .D(I650670), .CLK(I2702), .RSTB(I650195), .Q(I650172) );
nor I_38116 (I650187,I650512,I650653);
nor I_38117 (I650175,I650653,I650416);
not I_38118 (I650729,I650653);
and I_38119 (I650746,I650280,I650729);
nor I_38120 (I650181,I650416,I650746);
nand I_38121 (I650169,I650653,I650543);
not I_38122 (I650824,I2709);
not I_38123 (I650841,I114357);
nor I_38124 (I650858,I114375,I114354);
nand I_38125 (I650875,I650858,I114372);
nor I_38126 (I650892,I650841,I114375);
nand I_38127 (I650909,I650892,I114366);
not I_38128 (I650926,I114375);
not I_38129 (I650943,I650926);
not I_38130 (I650960,I114369);
nor I_38131 (I650977,I650960,I114363);
and I_38132 (I650994,I650977,I114360);
or I_38133 (I651011,I650994,I114351);
DFFARX1 I_38134  ( .D(I651011), .CLK(I2702), .RSTB(I650824), .Q(I651028) );
nand I_38135 (I651045,I650841,I114369);
or I_38136 (I650813,I651045,I651028);
not I_38137 (I651076,I651045);
nor I_38138 (I651093,I651028,I651076);
and I_38139 (I651110,I650926,I651093);
nand I_38140 (I650786,I651045,I650943);
DFFARX1 I_38141  ( .D(I114381), .CLK(I2702), .RSTB(I650824), .Q(I651141) );
or I_38142 (I650807,I651141,I651028);
nor I_38143 (I651172,I651141,I650909);
nor I_38144 (I651189,I651141,I650943);
nand I_38145 (I650792,I650875,I651189);
or I_38146 (I651220,I651141,I651110);
DFFARX1 I_38147  ( .D(I651220), .CLK(I2702), .RSTB(I650824), .Q(I650789) );
not I_38148 (I650795,I651141);
DFFARX1 I_38149  ( .D(I114378), .CLK(I2702), .RSTB(I650824), .Q(I651265) );
not I_38150 (I651282,I651265);
nor I_38151 (I651299,I651282,I650875);
DFFARX1 I_38152  ( .D(I651299), .CLK(I2702), .RSTB(I650824), .Q(I650801) );
nor I_38153 (I650816,I651141,I651282);
nor I_38154 (I650804,I651282,I651045);
not I_38155 (I651358,I651282);
and I_38156 (I651375,I650909,I651358);
nor I_38157 (I650810,I651045,I651375);
nand I_38158 (I650798,I651282,I651172);
not I_38159 (I651453,I2709);
not I_38160 (I651470,I578613);
nor I_38161 (I651487,I578616,I578625);
nand I_38162 (I651504,I651487,I578610);
nor I_38163 (I651521,I651470,I578616);
nand I_38164 (I651538,I651521,I578619);
not I_38165 (I651555,I578616);
not I_38166 (I651572,I651555);
not I_38167 (I651589,I578634);
nor I_38168 (I651606,I651589,I578622);
and I_38169 (I651623,I651606,I578607);
or I_38170 (I651640,I651623,I578604);
DFFARX1 I_38171  ( .D(I651640), .CLK(I2702), .RSTB(I651453), .Q(I651657) );
nand I_38172 (I651674,I651470,I578634);
or I_38173 (I651442,I651674,I651657);
not I_38174 (I651705,I651674);
nor I_38175 (I651722,I651657,I651705);
and I_38176 (I651739,I651555,I651722);
nand I_38177 (I651415,I651674,I651572);
DFFARX1 I_38178  ( .D(I578628), .CLK(I2702), .RSTB(I651453), .Q(I651770) );
or I_38179 (I651436,I651770,I651657);
nor I_38180 (I651801,I651770,I651538);
nor I_38181 (I651818,I651770,I651572);
nand I_38182 (I651421,I651504,I651818);
or I_38183 (I651849,I651770,I651739);
DFFARX1 I_38184  ( .D(I651849), .CLK(I2702), .RSTB(I651453), .Q(I651418) );
not I_38185 (I651424,I651770);
DFFARX1 I_38186  ( .D(I578631), .CLK(I2702), .RSTB(I651453), .Q(I651894) );
not I_38187 (I651911,I651894);
nor I_38188 (I651928,I651911,I651504);
DFFARX1 I_38189  ( .D(I651928), .CLK(I2702), .RSTB(I651453), .Q(I651430) );
nor I_38190 (I651445,I651770,I651911);
nor I_38191 (I651433,I651911,I651674);
not I_38192 (I651987,I651911);
and I_38193 (I652004,I651538,I651987);
nor I_38194 (I651439,I651674,I652004);
nand I_38195 (I651427,I651911,I651801);
not I_38196 (I652082,I2709);
not I_38197 (I652099,I56217);
nor I_38198 (I652116,I56235,I56214);
nand I_38199 (I652133,I652116,I56232);
nor I_38200 (I652150,I652099,I56235);
nand I_38201 (I652167,I652150,I56226);
not I_38202 (I652184,I56235);
not I_38203 (I652201,I652184);
not I_38204 (I652218,I56229);
nor I_38205 (I652235,I652218,I56223);
and I_38206 (I652252,I652235,I56220);
or I_38207 (I652269,I652252,I56211);
DFFARX1 I_38208  ( .D(I652269), .CLK(I2702), .RSTB(I652082), .Q(I652286) );
nand I_38209 (I652303,I652099,I56229);
or I_38210 (I652071,I652303,I652286);
not I_38211 (I652334,I652303);
nor I_38212 (I652351,I652286,I652334);
and I_38213 (I652368,I652184,I652351);
nand I_38214 (I652044,I652303,I652201);
DFFARX1 I_38215  ( .D(I56241), .CLK(I2702), .RSTB(I652082), .Q(I652399) );
or I_38216 (I652065,I652399,I652286);
nor I_38217 (I652430,I652399,I652167);
nor I_38218 (I652447,I652399,I652201);
nand I_38219 (I652050,I652133,I652447);
or I_38220 (I652478,I652399,I652368);
DFFARX1 I_38221  ( .D(I652478), .CLK(I2702), .RSTB(I652082), .Q(I652047) );
not I_38222 (I652053,I652399);
DFFARX1 I_38223  ( .D(I56238), .CLK(I2702), .RSTB(I652082), .Q(I652523) );
not I_38224 (I652540,I652523);
nor I_38225 (I652557,I652540,I652133);
DFFARX1 I_38226  ( .D(I652557), .CLK(I2702), .RSTB(I652082), .Q(I652059) );
nor I_38227 (I652074,I652399,I652540);
nor I_38228 (I652062,I652540,I652303);
not I_38229 (I652616,I652540);
and I_38230 (I652633,I652167,I652616);
nor I_38231 (I652068,I652303,I652633);
nand I_38232 (I652056,I652540,I652430);
not I_38233 (I652711,I2709);
not I_38234 (I652728,I613718);
nor I_38235 (I652745,I613721,I613730);
nand I_38236 (I652762,I652745,I613715);
nor I_38237 (I652779,I652728,I613721);
nand I_38238 (I652796,I652779,I613724);
not I_38239 (I652813,I613721);
not I_38240 (I652830,I652813);
not I_38241 (I652847,I613739);
nor I_38242 (I652864,I652847,I613727);
and I_38243 (I652881,I652864,I613712);
or I_38244 (I652898,I652881,I613709);
DFFARX1 I_38245  ( .D(I652898), .CLK(I2702), .RSTB(I652711), .Q(I652915) );
nand I_38246 (I652932,I652728,I613739);
or I_38247 (I652700,I652932,I652915);
not I_38248 (I652963,I652932);
nor I_38249 (I652980,I652915,I652963);
and I_38250 (I652997,I652813,I652980);
nand I_38251 (I652673,I652932,I652830);
DFFARX1 I_38252  ( .D(I613733), .CLK(I2702), .RSTB(I652711), .Q(I653028) );
or I_38253 (I652694,I653028,I652915);
nor I_38254 (I653059,I653028,I652796);
nor I_38255 (I653076,I653028,I652830);
nand I_38256 (I652679,I652762,I653076);
or I_38257 (I653107,I653028,I652997);
DFFARX1 I_38258  ( .D(I653107), .CLK(I2702), .RSTB(I652711), .Q(I652676) );
not I_38259 (I652682,I653028);
DFFARX1 I_38260  ( .D(I613736), .CLK(I2702), .RSTB(I652711), .Q(I653152) );
not I_38261 (I653169,I653152);
nor I_38262 (I653186,I653169,I652762);
DFFARX1 I_38263  ( .D(I653186), .CLK(I2702), .RSTB(I652711), .Q(I652688) );
nor I_38264 (I652703,I653028,I653169);
nor I_38265 (I652691,I653169,I652932);
not I_38266 (I653245,I653169);
and I_38267 (I653262,I652796,I653245);
nor I_38268 (I652697,I652932,I653262);
nand I_38269 (I652685,I653169,I653059);
not I_38270 (I653340,I2709);
not I_38271 (I653357,I85933);
nor I_38272 (I653374,I85951,I85930);
nand I_38273 (I653391,I653374,I85948);
nor I_38274 (I653408,I653357,I85951);
nand I_38275 (I653425,I653408,I85942);
not I_38276 (I653442,I85951);
not I_38277 (I653459,I653442);
not I_38278 (I653476,I85945);
nor I_38279 (I653493,I653476,I85939);
and I_38280 (I653510,I653493,I85936);
or I_38281 (I653527,I653510,I85927);
DFFARX1 I_38282  ( .D(I653527), .CLK(I2702), .RSTB(I653340), .Q(I653544) );
nand I_38283 (I653561,I653357,I85945);
or I_38284 (I653329,I653561,I653544);
not I_38285 (I653592,I653561);
nor I_38286 (I653609,I653544,I653592);
and I_38287 (I653626,I653442,I653609);
nand I_38288 (I653302,I653561,I653459);
DFFARX1 I_38289  ( .D(I85957), .CLK(I2702), .RSTB(I653340), .Q(I653657) );
or I_38290 (I653323,I653657,I653544);
nor I_38291 (I653688,I653657,I653425);
nor I_38292 (I653705,I653657,I653459);
nand I_38293 (I653308,I653391,I653705);
or I_38294 (I653736,I653657,I653626);
DFFARX1 I_38295  ( .D(I653736), .CLK(I2702), .RSTB(I653340), .Q(I653305) );
not I_38296 (I653311,I653657);
DFFARX1 I_38297  ( .D(I85954), .CLK(I2702), .RSTB(I653340), .Q(I653781) );
not I_38298 (I653798,I653781);
nor I_38299 (I653815,I653798,I653391);
DFFARX1 I_38300  ( .D(I653815), .CLK(I2702), .RSTB(I653340), .Q(I653317) );
nor I_38301 (I653332,I653657,I653798);
nor I_38302 (I653320,I653798,I653561);
not I_38303 (I653874,I653798);
and I_38304 (I653891,I653425,I653874);
nor I_38305 (I653326,I653561,I653891);
nand I_38306 (I653314,I653798,I653688);
not I_38307 (I653969,I2709);
not I_38308 (I653986,I29643);
nor I_38309 (I654003,I29646,I29655);
nand I_38310 (I654020,I654003,I29670);
nor I_38311 (I654037,I653986,I29646);
nand I_38312 (I654054,I654037,I29649);
not I_38313 (I654071,I29646);
not I_38314 (I654088,I654071);
not I_38315 (I654105,I29640);
nor I_38316 (I654122,I654105,I29664);
and I_38317 (I654139,I654122,I29652);
or I_38318 (I654156,I654139,I29658);
DFFARX1 I_38319  ( .D(I654156), .CLK(I2702), .RSTB(I653969), .Q(I654173) );
nand I_38320 (I654190,I653986,I29640);
or I_38321 (I653958,I654190,I654173);
not I_38322 (I654221,I654190);
nor I_38323 (I654238,I654173,I654221);
and I_38324 (I654255,I654071,I654238);
nand I_38325 (I653931,I654190,I654088);
DFFARX1 I_38326  ( .D(I29661), .CLK(I2702), .RSTB(I653969), .Q(I654286) );
or I_38327 (I653952,I654286,I654173);
nor I_38328 (I654317,I654286,I654054);
nor I_38329 (I654334,I654286,I654088);
nand I_38330 (I653937,I654020,I654334);
or I_38331 (I654365,I654286,I654255);
DFFARX1 I_38332  ( .D(I654365), .CLK(I2702), .RSTB(I653969), .Q(I653934) );
not I_38333 (I653940,I654286);
DFFARX1 I_38334  ( .D(I29667), .CLK(I2702), .RSTB(I653969), .Q(I654410) );
not I_38335 (I654427,I654410);
nor I_38336 (I654444,I654427,I654020);
DFFARX1 I_38337  ( .D(I654444), .CLK(I2702), .RSTB(I653969), .Q(I653946) );
nor I_38338 (I653961,I654286,I654427);
nor I_38339 (I653949,I654427,I654190);
not I_38340 (I654503,I654427);
and I_38341 (I654520,I654054,I654503);
nor I_38342 (I653955,I654190,I654520);
nand I_38343 (I653943,I654427,I654317);
not I_38344 (I654598,I2709);
not I_38345 (I654615,I533390);
nor I_38346 (I654632,I533408,I533387);
nand I_38347 (I654649,I654632,I533411);
nor I_38348 (I654666,I654615,I533408);
nand I_38349 (I654683,I654666,I533405);
not I_38350 (I654700,I533408);
not I_38351 (I654717,I654700);
not I_38352 (I654734,I533396);
nor I_38353 (I654751,I654734,I533384);
and I_38354 (I654768,I654751,I533402);
or I_38355 (I654785,I654768,I533414);
DFFARX1 I_38356  ( .D(I654785), .CLK(I2702), .RSTB(I654598), .Q(I654802) );
nand I_38357 (I654819,I654615,I533396);
or I_38358 (I654587,I654819,I654802);
not I_38359 (I654850,I654819);
nor I_38360 (I654867,I654802,I654850);
and I_38361 (I654884,I654700,I654867);
nand I_38362 (I654560,I654819,I654717);
DFFARX1 I_38363  ( .D(I533393), .CLK(I2702), .RSTB(I654598), .Q(I654915) );
or I_38364 (I654581,I654915,I654802);
nor I_38365 (I654946,I654915,I654683);
nor I_38366 (I654963,I654915,I654717);
nand I_38367 (I654566,I654649,I654963);
or I_38368 (I654994,I654915,I654884);
DFFARX1 I_38369  ( .D(I654994), .CLK(I2702), .RSTB(I654598), .Q(I654563) );
not I_38370 (I654569,I654915);
DFFARX1 I_38371  ( .D(I533399), .CLK(I2702), .RSTB(I654598), .Q(I655039) );
not I_38372 (I655056,I655039);
nor I_38373 (I655073,I655056,I654649);
DFFARX1 I_38374  ( .D(I655073), .CLK(I2702), .RSTB(I654598), .Q(I654575) );
nor I_38375 (I654590,I654915,I655056);
nor I_38376 (I654578,I655056,I654819);
not I_38377 (I655132,I655056);
and I_38378 (I655149,I654683,I655132);
nor I_38379 (I654584,I654819,I655149);
nand I_38380 (I654572,I655056,I654946);
not I_38381 (I655227,I2709);
not I_38382 (I655244,I170055);
nor I_38383 (I655261,I170046,I170070);
nand I_38384 (I655278,I655261,I170073);
nor I_38385 (I655295,I655244,I170046);
nand I_38386 (I655312,I655295,I170064);
not I_38387 (I655329,I170046);
not I_38388 (I655346,I655329);
not I_38389 (I655363,I170058);
nor I_38390 (I655380,I655363,I170052);
and I_38391 (I655397,I655380,I170061);
or I_38392 (I655414,I655397,I170049);
DFFARX1 I_38393  ( .D(I655414), .CLK(I2702), .RSTB(I655227), .Q(I655431) );
nand I_38394 (I655448,I655244,I170058);
or I_38395 (I655216,I655448,I655431);
not I_38396 (I655479,I655448);
nor I_38397 (I655496,I655431,I655479);
and I_38398 (I655513,I655329,I655496);
nand I_38399 (I655189,I655448,I655346);
DFFARX1 I_38400  ( .D(I170043), .CLK(I2702), .RSTB(I655227), .Q(I655544) );
or I_38401 (I655210,I655544,I655431);
nor I_38402 (I655575,I655544,I655312);
nor I_38403 (I655592,I655544,I655346);
nand I_38404 (I655195,I655278,I655592);
or I_38405 (I655623,I655544,I655513);
DFFARX1 I_38406  ( .D(I655623), .CLK(I2702), .RSTB(I655227), .Q(I655192) );
not I_38407 (I655198,I655544);
DFFARX1 I_38408  ( .D(I170067), .CLK(I2702), .RSTB(I655227), .Q(I655668) );
not I_38409 (I655685,I655668);
nor I_38410 (I655702,I655685,I655278);
DFFARX1 I_38411  ( .D(I655702), .CLK(I2702), .RSTB(I655227), .Q(I655204) );
nor I_38412 (I655219,I655544,I655685);
nor I_38413 (I655207,I655685,I655448);
not I_38414 (I655761,I655685);
and I_38415 (I655778,I655312,I655761);
nor I_38416 (I655213,I655448,I655778);
nand I_38417 (I655201,I655685,I655575);
not I_38418 (I655856,I2709);
not I_38419 (I655873,I165414);
nor I_38420 (I655890,I165405,I165429);
nand I_38421 (I655907,I655890,I165432);
nor I_38422 (I655924,I655873,I165405);
nand I_38423 (I655941,I655924,I165423);
not I_38424 (I655958,I165405);
not I_38425 (I655975,I655958);
not I_38426 (I655992,I165417);
nor I_38427 (I656009,I655992,I165411);
and I_38428 (I656026,I656009,I165420);
or I_38429 (I656043,I656026,I165408);
DFFARX1 I_38430  ( .D(I656043), .CLK(I2702), .RSTB(I655856), .Q(I656060) );
nand I_38431 (I656077,I655873,I165417);
or I_38432 (I655845,I656077,I656060);
not I_38433 (I656108,I656077);
nor I_38434 (I656125,I656060,I656108);
and I_38435 (I656142,I655958,I656125);
nand I_38436 (I655818,I656077,I655975);
DFFARX1 I_38437  ( .D(I165402), .CLK(I2702), .RSTB(I655856), .Q(I656173) );
or I_38438 (I655839,I656173,I656060);
nor I_38439 (I656204,I656173,I655941);
nor I_38440 (I656221,I656173,I655975);
nand I_38441 (I655824,I655907,I656221);
or I_38442 (I656252,I656173,I656142);
DFFARX1 I_38443  ( .D(I656252), .CLK(I2702), .RSTB(I655856), .Q(I655821) );
not I_38444 (I655827,I656173);
DFFARX1 I_38445  ( .D(I165426), .CLK(I2702), .RSTB(I655856), .Q(I656297) );
not I_38446 (I656314,I656297);
nor I_38447 (I656331,I656314,I655907);
DFFARX1 I_38448  ( .D(I656331), .CLK(I2702), .RSTB(I655856), .Q(I655833) );
nor I_38449 (I655848,I656173,I656314);
nor I_38450 (I655836,I656314,I656077);
not I_38451 (I656390,I656314);
and I_38452 (I656407,I655941,I656390);
nor I_38453 (I655842,I656077,I656407);
nand I_38454 (I655830,I656314,I656204);
not I_38455 (I656485,I2709);
not I_38456 (I656502,I160110);
nor I_38457 (I656519,I160101,I160125);
nand I_38458 (I656536,I656519,I160128);
nor I_38459 (I656553,I656502,I160101);
nand I_38460 (I656570,I656553,I160119);
not I_38461 (I656587,I160101);
not I_38462 (I656604,I656587);
not I_38463 (I656621,I160113);
nor I_38464 (I656638,I656621,I160107);
and I_38465 (I656655,I656638,I160116);
or I_38466 (I656672,I656655,I160104);
DFFARX1 I_38467  ( .D(I656672), .CLK(I2702), .RSTB(I656485), .Q(I656689) );
nand I_38468 (I656706,I656502,I160113);
or I_38469 (I656474,I656706,I656689);
not I_38470 (I656737,I656706);
nor I_38471 (I656754,I656689,I656737);
and I_38472 (I656771,I656587,I656754);
nand I_38473 (I656447,I656706,I656604);
DFFARX1 I_38474  ( .D(I160098), .CLK(I2702), .RSTB(I656485), .Q(I656802) );
or I_38475 (I656468,I656802,I656689);
nor I_38476 (I656833,I656802,I656570);
nor I_38477 (I656850,I656802,I656604);
nand I_38478 (I656453,I656536,I656850);
or I_38479 (I656881,I656802,I656771);
DFFARX1 I_38480  ( .D(I656881), .CLK(I2702), .RSTB(I656485), .Q(I656450) );
not I_38481 (I656456,I656802);
DFFARX1 I_38482  ( .D(I160122), .CLK(I2702), .RSTB(I656485), .Q(I656926) );
not I_38483 (I656943,I656926);
nor I_38484 (I656960,I656943,I656536);
DFFARX1 I_38485  ( .D(I656960), .CLK(I2702), .RSTB(I656485), .Q(I656462) );
nor I_38486 (I656477,I656802,I656943);
nor I_38487 (I656465,I656943,I656706);
not I_38488 (I657019,I656943);
and I_38489 (I657036,I656570,I657019);
nor I_38490 (I656471,I656706,I657036);
nand I_38491 (I656459,I656943,I656833);
not I_38492 (I657114,I2709);
not I_38493 (I657131,I455265);
nor I_38494 (I657148,I455238,I455256);
nand I_38495 (I657165,I657148,I455241);
nor I_38496 (I657182,I657131,I455238);
nand I_38497 (I657199,I657182,I455259);
not I_38498 (I657216,I455238);
not I_38499 (I657233,I657216);
not I_38500 (I657250,I455235);
nor I_38501 (I657267,I657250,I455262);
and I_38502 (I657284,I657267,I455253);
or I_38503 (I657301,I657284,I455244);
DFFARX1 I_38504  ( .D(I657301), .CLK(I2702), .RSTB(I657114), .Q(I657318) );
nand I_38505 (I657335,I657131,I455235);
or I_38506 (I657103,I657335,I657318);
not I_38507 (I657366,I657335);
nor I_38508 (I657383,I657318,I657366);
and I_38509 (I657400,I657216,I657383);
nand I_38510 (I657076,I657335,I657233);
DFFARX1 I_38511  ( .D(I455247), .CLK(I2702), .RSTB(I657114), .Q(I657431) );
or I_38512 (I657097,I657431,I657318);
nor I_38513 (I657462,I657431,I657199);
nor I_38514 (I657479,I657431,I657233);
nand I_38515 (I657082,I657165,I657479);
or I_38516 (I657510,I657431,I657400);
DFFARX1 I_38517  ( .D(I657510), .CLK(I2702), .RSTB(I657114), .Q(I657079) );
not I_38518 (I657085,I657431);
DFFARX1 I_38519  ( .D(I455250), .CLK(I2702), .RSTB(I657114), .Q(I657555) );
not I_38520 (I657572,I657555);
nor I_38521 (I657589,I657572,I657165);
DFFARX1 I_38522  ( .D(I657589), .CLK(I2702), .RSTB(I657114), .Q(I657091) );
nor I_38523 (I657106,I657431,I657572);
nor I_38524 (I657094,I657572,I657335);
not I_38525 (I657648,I657572);
and I_38526 (I657665,I657199,I657648);
nor I_38527 (I657100,I657335,I657665);
nand I_38528 (I657088,I657572,I657462);
not I_38529 (I657743,I2709);
not I_38530 (I657760,I38619);
nor I_38531 (I657777,I38622,I38631);
nand I_38532 (I657794,I657777,I38646);
nor I_38533 (I657811,I657760,I38622);
nand I_38534 (I657828,I657811,I38625);
not I_38535 (I657845,I38622);
not I_38536 (I657862,I657845);
not I_38537 (I657879,I38616);
nor I_38538 (I657896,I657879,I38640);
and I_38539 (I657913,I657896,I38628);
or I_38540 (I657930,I657913,I38634);
DFFARX1 I_38541  ( .D(I657930), .CLK(I2702), .RSTB(I657743), .Q(I657947) );
nand I_38542 (I657964,I657760,I38616);
or I_38543 (I657732,I657964,I657947);
not I_38544 (I657995,I657964);
nor I_38545 (I658012,I657947,I657995);
and I_38546 (I658029,I657845,I658012);
nand I_38547 (I657705,I657964,I657862);
DFFARX1 I_38548  ( .D(I38637), .CLK(I2702), .RSTB(I657743), .Q(I658060) );
or I_38549 (I657726,I658060,I657947);
nor I_38550 (I658091,I658060,I657828);
nor I_38551 (I658108,I658060,I657862);
nand I_38552 (I657711,I657794,I658108);
or I_38553 (I658139,I658060,I658029);
DFFARX1 I_38554  ( .D(I658139), .CLK(I2702), .RSTB(I657743), .Q(I657708) );
not I_38555 (I657714,I658060);
DFFARX1 I_38556  ( .D(I38643), .CLK(I2702), .RSTB(I657743), .Q(I658184) );
not I_38557 (I658201,I658184);
nor I_38558 (I658218,I658201,I657794);
DFFARX1 I_38559  ( .D(I658218), .CLK(I2702), .RSTB(I657743), .Q(I657720) );
nor I_38560 (I657735,I658060,I658201);
nor I_38561 (I657723,I658201,I657964);
not I_38562 (I658277,I658201);
and I_38563 (I658294,I657828,I658277);
nor I_38564 (I657729,I657964,I658294);
nand I_38565 (I657717,I658201,I658091);
not I_38566 (I658372,I2709);
not I_38567 (I658389,I204073);
nor I_38568 (I658406,I204049,I204064);
nand I_38569 (I658423,I658406,I204046);
nor I_38570 (I658440,I658389,I204049);
nand I_38571 (I658457,I658440,I204061);
not I_38572 (I658474,I204049);
not I_38573 (I658491,I658474);
not I_38574 (I658508,I204052);
nor I_38575 (I658525,I658508,I204067);
and I_38576 (I658542,I658525,I204058);
or I_38577 (I658559,I658542,I204043);
DFFARX1 I_38578  ( .D(I658559), .CLK(I2702), .RSTB(I658372), .Q(I658576) );
nand I_38579 (I658593,I658389,I204052);
or I_38580 (I658361,I658593,I658576);
not I_38581 (I658624,I658593);
nor I_38582 (I658641,I658576,I658624);
and I_38583 (I658658,I658474,I658641);
nand I_38584 (I658334,I658593,I658491);
DFFARX1 I_38585  ( .D(I204055), .CLK(I2702), .RSTB(I658372), .Q(I658689) );
or I_38586 (I658355,I658689,I658576);
nor I_38587 (I658720,I658689,I658457);
nor I_38588 (I658737,I658689,I658491);
nand I_38589 (I658340,I658423,I658737);
or I_38590 (I658768,I658689,I658658);
DFFARX1 I_38591  ( .D(I658768), .CLK(I2702), .RSTB(I658372), .Q(I658337) );
not I_38592 (I658343,I658689);
DFFARX1 I_38593  ( .D(I204070), .CLK(I2702), .RSTB(I658372), .Q(I658813) );
not I_38594 (I658830,I658813);
nor I_38595 (I658847,I658830,I658423);
DFFARX1 I_38596  ( .D(I658847), .CLK(I2702), .RSTB(I658372), .Q(I658349) );
nor I_38597 (I658364,I658689,I658830);
nor I_38598 (I658352,I658830,I658593);
not I_38599 (I658906,I658830);
and I_38600 (I658923,I658457,I658906);
nor I_38601 (I658358,I658593,I658923);
nand I_38602 (I658346,I658830,I658720);
not I_38603 (I659001,I2709);
not I_38604 (I659018,I176685);
nor I_38605 (I659035,I176676,I176700);
nand I_38606 (I659052,I659035,I176703);
nor I_38607 (I659069,I659018,I176676);
nand I_38608 (I659086,I659069,I176694);
not I_38609 (I659103,I176676);
not I_38610 (I659120,I659103);
not I_38611 (I659137,I176688);
nor I_38612 (I659154,I659137,I176682);
and I_38613 (I659171,I659154,I176691);
or I_38614 (I659188,I659171,I176679);
DFFARX1 I_38615  ( .D(I659188), .CLK(I2702), .RSTB(I659001), .Q(I659205) );
nand I_38616 (I659222,I659018,I176688);
or I_38617 (I658990,I659222,I659205);
not I_38618 (I659253,I659222);
nor I_38619 (I659270,I659205,I659253);
and I_38620 (I659287,I659103,I659270);
nand I_38621 (I658963,I659222,I659120);
DFFARX1 I_38622  ( .D(I176673), .CLK(I2702), .RSTB(I659001), .Q(I659318) );
or I_38623 (I658984,I659318,I659205);
nor I_38624 (I659349,I659318,I659086);
nor I_38625 (I659366,I659318,I659120);
nand I_38626 (I658969,I659052,I659366);
or I_38627 (I659397,I659318,I659287);
DFFARX1 I_38628  ( .D(I659397), .CLK(I2702), .RSTB(I659001), .Q(I658966) );
not I_38629 (I658972,I659318);
DFFARX1 I_38630  ( .D(I176697), .CLK(I2702), .RSTB(I659001), .Q(I659442) );
not I_38631 (I659459,I659442);
nor I_38632 (I659476,I659459,I659052);
DFFARX1 I_38633  ( .D(I659476), .CLK(I2702), .RSTB(I659001), .Q(I658978) );
nor I_38634 (I658993,I659318,I659459);
nor I_38635 (I658981,I659459,I659222);
not I_38636 (I659535,I659459);
and I_38637 (I659552,I659086,I659535);
nor I_38638 (I658987,I659222,I659552);
nand I_38639 (I658975,I659459,I659349);
not I_38640 (I659630,I2709);
not I_38641 (I659647,I185304);
nor I_38642 (I659664,I185295,I185319);
nand I_38643 (I659681,I659664,I185322);
nor I_38644 (I659698,I659647,I185295);
nand I_38645 (I659715,I659698,I185313);
not I_38646 (I659732,I185295);
not I_38647 (I659749,I659732);
not I_38648 (I659766,I185307);
nor I_38649 (I659783,I659766,I185301);
and I_38650 (I659800,I659783,I185310);
or I_38651 (I659817,I659800,I185298);
DFFARX1 I_38652  ( .D(I659817), .CLK(I2702), .RSTB(I659630), .Q(I659834) );
nand I_38653 (I659851,I659647,I185307);
or I_38654 (I659619,I659851,I659834);
not I_38655 (I659882,I659851);
nor I_38656 (I659899,I659834,I659882);
and I_38657 (I659916,I659732,I659899);
nand I_38658 (I659592,I659851,I659749);
DFFARX1 I_38659  ( .D(I185292), .CLK(I2702), .RSTB(I659630), .Q(I659947) );
or I_38660 (I659613,I659947,I659834);
nor I_38661 (I659978,I659947,I659715);
nor I_38662 (I659995,I659947,I659749);
nand I_38663 (I659598,I659681,I659995);
or I_38664 (I660026,I659947,I659916);
DFFARX1 I_38665  ( .D(I660026), .CLK(I2702), .RSTB(I659630), .Q(I659595) );
not I_38666 (I659601,I659947);
DFFARX1 I_38667  ( .D(I185316), .CLK(I2702), .RSTB(I659630), .Q(I660071) );
not I_38668 (I660088,I660071);
nor I_38669 (I660105,I660088,I659681);
DFFARX1 I_38670  ( .D(I660105), .CLK(I2702), .RSTB(I659630), .Q(I659607) );
nor I_38671 (I659622,I659947,I660088);
nor I_38672 (I659610,I660088,I659851);
not I_38673 (I660164,I660088);
and I_38674 (I660181,I659715,I660164);
nor I_38675 (I659616,I659851,I660181);
nand I_38676 (I659604,I660088,I659978);
not I_38677 (I660259,I2709);
not I_38678 (I660276,I169392);
nor I_38679 (I660293,I169383,I169407);
nand I_38680 (I660310,I660293,I169410);
nor I_38681 (I660327,I660276,I169383);
nand I_38682 (I660344,I660327,I169401);
not I_38683 (I660361,I169383);
not I_38684 (I660378,I660361);
not I_38685 (I660395,I169395);
nor I_38686 (I660412,I660395,I169389);
and I_38687 (I660429,I660412,I169398);
or I_38688 (I660446,I660429,I169386);
DFFARX1 I_38689  ( .D(I660446), .CLK(I2702), .RSTB(I660259), .Q(I660463) );
nand I_38690 (I660480,I660276,I169395);
or I_38691 (I660248,I660480,I660463);
not I_38692 (I660511,I660480);
nor I_38693 (I660528,I660463,I660511);
and I_38694 (I660545,I660361,I660528);
nand I_38695 (I660221,I660480,I660378);
DFFARX1 I_38696  ( .D(I169380), .CLK(I2702), .RSTB(I660259), .Q(I660576) );
or I_38697 (I660242,I660576,I660463);
nor I_38698 (I660607,I660576,I660344);
nor I_38699 (I660624,I660576,I660378);
nand I_38700 (I660227,I660310,I660624);
or I_38701 (I660655,I660576,I660545);
DFFARX1 I_38702  ( .D(I660655), .CLK(I2702), .RSTB(I660259), .Q(I660224) );
not I_38703 (I660230,I660576);
DFFARX1 I_38704  ( .D(I169404), .CLK(I2702), .RSTB(I660259), .Q(I660700) );
not I_38705 (I660717,I660700);
nor I_38706 (I660734,I660717,I660310);
DFFARX1 I_38707  ( .D(I660734), .CLK(I2702), .RSTB(I660259), .Q(I660236) );
nor I_38708 (I660251,I660576,I660717);
nor I_38709 (I660239,I660717,I660480);
not I_38710 (I660793,I660717);
and I_38711 (I660810,I660344,I660793);
nor I_38712 (I660245,I660480,I660810);
nand I_38713 (I660233,I660717,I660607);
not I_38714 (I660888,I2709);
not I_38715 (I660905,I31887);
nor I_38716 (I660922,I31890,I31899);
nand I_38717 (I660939,I660922,I31914);
nor I_38718 (I660956,I660905,I31890);
nand I_38719 (I660973,I660956,I31893);
not I_38720 (I660990,I31890);
not I_38721 (I661007,I660990);
not I_38722 (I661024,I31884);
nor I_38723 (I661041,I661024,I31908);
and I_38724 (I661058,I661041,I31896);
or I_38725 (I661075,I661058,I31902);
DFFARX1 I_38726  ( .D(I661075), .CLK(I2702), .RSTB(I660888), .Q(I661092) );
nand I_38727 (I661109,I660905,I31884);
or I_38728 (I660877,I661109,I661092);
not I_38729 (I661140,I661109);
nor I_38730 (I661157,I661092,I661140);
and I_38731 (I661174,I660990,I661157);
nand I_38732 (I660850,I661109,I661007);
DFFARX1 I_38733  ( .D(I31905), .CLK(I2702), .RSTB(I660888), .Q(I661205) );
or I_38734 (I660871,I661205,I661092);
nor I_38735 (I661236,I661205,I660973);
nor I_38736 (I661253,I661205,I661007);
nand I_38737 (I660856,I660939,I661253);
or I_38738 (I661284,I661205,I661174);
DFFARX1 I_38739  ( .D(I661284), .CLK(I2702), .RSTB(I660888), .Q(I660853) );
not I_38740 (I660859,I661205);
DFFARX1 I_38741  ( .D(I31911), .CLK(I2702), .RSTB(I660888), .Q(I661329) );
not I_38742 (I661346,I661329);
nor I_38743 (I661363,I661346,I660939);
DFFARX1 I_38744  ( .D(I661363), .CLK(I2702), .RSTB(I660888), .Q(I660865) );
nor I_38745 (I660880,I661205,I661346);
nor I_38746 (I660868,I661346,I661109);
not I_38747 (I661422,I661346);
and I_38748 (I661439,I660973,I661422);
nor I_38749 (I660874,I661109,I661439);
nand I_38750 (I660862,I661346,I661236);
not I_38751 (I661517,I2709);
not I_38752 (I661534,I140220);
nor I_38753 (I661551,I140211,I140235);
nand I_38754 (I661568,I661551,I140238);
nor I_38755 (I661585,I661534,I140211);
nand I_38756 (I661602,I661585,I140229);
not I_38757 (I661619,I140211);
not I_38758 (I661636,I661619);
not I_38759 (I661653,I140223);
nor I_38760 (I661670,I661653,I140217);
and I_38761 (I661687,I661670,I140226);
or I_38762 (I661704,I661687,I140214);
DFFARX1 I_38763  ( .D(I661704), .CLK(I2702), .RSTB(I661517), .Q(I661721) );
nand I_38764 (I661738,I661534,I140223);
or I_38765 (I661506,I661738,I661721);
not I_38766 (I661769,I661738);
nor I_38767 (I661786,I661721,I661769);
and I_38768 (I661803,I661619,I661786);
nand I_38769 (I661479,I661738,I661636);
DFFARX1 I_38770  ( .D(I140208), .CLK(I2702), .RSTB(I661517), .Q(I661834) );
or I_38771 (I661500,I661834,I661721);
nor I_38772 (I661865,I661834,I661602);
nor I_38773 (I661882,I661834,I661636);
nand I_38774 (I661485,I661568,I661882);
or I_38775 (I661913,I661834,I661803);
DFFARX1 I_38776  ( .D(I661913), .CLK(I2702), .RSTB(I661517), .Q(I661482) );
not I_38777 (I661488,I661834);
DFFARX1 I_38778  ( .D(I140232), .CLK(I2702), .RSTB(I661517), .Q(I661958) );
not I_38779 (I661975,I661958);
nor I_38780 (I661992,I661975,I661568);
DFFARX1 I_38781  ( .D(I661992), .CLK(I2702), .RSTB(I661517), .Q(I661494) );
nor I_38782 (I661509,I661834,I661975);
nor I_38783 (I661497,I661975,I661738);
not I_38784 (I662051,I661975);
and I_38785 (I662068,I661602,I662051);
nor I_38786 (I661503,I661738,I662068);
nand I_38787 (I661491,I661975,I661865);
not I_38788 (I662146,I2709);
not I_38789 (I662163,I62677);
nor I_38790 (I662180,I62695,I62674);
nand I_38791 (I662197,I662180,I62692);
nor I_38792 (I662214,I662163,I62695);
nand I_38793 (I662231,I662214,I62686);
not I_38794 (I662248,I62695);
not I_38795 (I662265,I662248);
not I_38796 (I662282,I62689);
nor I_38797 (I662299,I662282,I62683);
and I_38798 (I662316,I662299,I62680);
or I_38799 (I662333,I662316,I62671);
DFFARX1 I_38800  ( .D(I662333), .CLK(I2702), .RSTB(I662146), .Q(I662350) );
nand I_38801 (I662367,I662163,I62689);
or I_38802 (I662135,I662367,I662350);
not I_38803 (I662398,I662367);
nor I_38804 (I662415,I662350,I662398);
and I_38805 (I662432,I662248,I662415);
nand I_38806 (I662108,I662367,I662265);
DFFARX1 I_38807  ( .D(I62701), .CLK(I2702), .RSTB(I662146), .Q(I662463) );
or I_38808 (I662129,I662463,I662350);
nor I_38809 (I662494,I662463,I662231);
nor I_38810 (I662511,I662463,I662265);
nand I_38811 (I662114,I662197,I662511);
or I_38812 (I662542,I662463,I662432);
DFFARX1 I_38813  ( .D(I662542), .CLK(I2702), .RSTB(I662146), .Q(I662111) );
not I_38814 (I662117,I662463);
DFFARX1 I_38815  ( .D(I62698), .CLK(I2702), .RSTB(I662146), .Q(I662587) );
not I_38816 (I662604,I662587);
nor I_38817 (I662621,I662604,I662197);
DFFARX1 I_38818  ( .D(I662621), .CLK(I2702), .RSTB(I662146), .Q(I662123) );
nor I_38819 (I662138,I662463,I662604);
nor I_38820 (I662126,I662604,I662367);
not I_38821 (I662680,I662604);
and I_38822 (I662697,I662231,I662680);
nor I_38823 (I662132,I662367,I662697);
nand I_38824 (I662120,I662604,I662494);
not I_38825 (I662775,I2709);
not I_38826 (I662792,I250284);
nor I_38827 (I662809,I250290,I250269);
nand I_38828 (I662826,I662809,I250275);
nor I_38829 (I662843,I662792,I250290);
nand I_38830 (I662860,I662843,I250281);
not I_38831 (I662877,I250290);
not I_38832 (I662894,I662877);
not I_38833 (I662911,I250278);
nor I_38834 (I662928,I662911,I250296);
and I_38835 (I662945,I662928,I250287);
or I_38836 (I662962,I662945,I250266);
DFFARX1 I_38837  ( .D(I662962), .CLK(I2702), .RSTB(I662775), .Q(I662979) );
nand I_38838 (I662996,I662792,I250278);
or I_38839 (I662764,I662996,I662979);
not I_38840 (I663027,I662996);
nor I_38841 (I663044,I662979,I663027);
and I_38842 (I663061,I662877,I663044);
nand I_38843 (I662737,I662996,I662894);
DFFARX1 I_38844  ( .D(I250293), .CLK(I2702), .RSTB(I662775), .Q(I663092) );
or I_38845 (I662758,I663092,I662979);
nor I_38846 (I663123,I663092,I662860);
nor I_38847 (I663140,I663092,I662894);
nand I_38848 (I662743,I662826,I663140);
or I_38849 (I663171,I663092,I663061);
DFFARX1 I_38850  ( .D(I663171), .CLK(I2702), .RSTB(I662775), .Q(I662740) );
not I_38851 (I662746,I663092);
DFFARX1 I_38852  ( .D(I250272), .CLK(I2702), .RSTB(I662775), .Q(I663216) );
not I_38853 (I663233,I663216);
nor I_38854 (I663250,I663233,I662826);
DFFARX1 I_38855  ( .D(I663250), .CLK(I2702), .RSTB(I662775), .Q(I662752) );
nor I_38856 (I662767,I663092,I663233);
nor I_38857 (I662755,I663233,I662996);
not I_38858 (I663309,I663233);
and I_38859 (I663326,I662860,I663309);
nor I_38860 (I662761,I662996,I663326);
nand I_38861 (I662749,I663233,I663123);
not I_38862 (I663404,I2709);
not I_38863 (I663421,I586348);
nor I_38864 (I663438,I586351,I586360);
nand I_38865 (I663455,I663438,I586345);
nor I_38866 (I663472,I663421,I586351);
nand I_38867 (I663489,I663472,I586354);
not I_38868 (I663506,I586351);
not I_38869 (I663523,I663506);
not I_38870 (I663540,I586369);
nor I_38871 (I663557,I663540,I586357);
and I_38872 (I663574,I663557,I586342);
or I_38873 (I663591,I663574,I586339);
DFFARX1 I_38874  ( .D(I663591), .CLK(I2702), .RSTB(I663404), .Q(I663608) );
nand I_38875 (I663625,I663421,I586369);
or I_38876 (I663393,I663625,I663608);
not I_38877 (I663656,I663625);
nor I_38878 (I663673,I663608,I663656);
and I_38879 (I663690,I663506,I663673);
nand I_38880 (I663366,I663625,I663523);
DFFARX1 I_38881  ( .D(I586363), .CLK(I2702), .RSTB(I663404), .Q(I663721) );
or I_38882 (I663387,I663721,I663608);
nor I_38883 (I663752,I663721,I663489);
nor I_38884 (I663769,I663721,I663523);
nand I_38885 (I663372,I663455,I663769);
or I_38886 (I663800,I663721,I663690);
DFFARX1 I_38887  ( .D(I663800), .CLK(I2702), .RSTB(I663404), .Q(I663369) );
not I_38888 (I663375,I663721);
DFFARX1 I_38889  ( .D(I586366), .CLK(I2702), .RSTB(I663404), .Q(I663845) );
not I_38890 (I663862,I663845);
nor I_38891 (I663879,I663862,I663455);
DFFARX1 I_38892  ( .D(I663879), .CLK(I2702), .RSTB(I663404), .Q(I663381) );
nor I_38893 (I663396,I663721,I663862);
nor I_38894 (I663384,I663862,I663625);
not I_38895 (I663938,I663862);
and I_38896 (I663955,I663489,I663938);
nor I_38897 (I663390,I663625,I663955);
nand I_38898 (I663378,I663862,I663752);
not I_38899 (I664033,I2709);
not I_38900 (I664050,I98207);
nor I_38901 (I664067,I98225,I98204);
nand I_38902 (I664084,I664067,I98222);
nor I_38903 (I664101,I664050,I98225);
nand I_38904 (I664118,I664101,I98216);
not I_38905 (I664135,I98225);
not I_38906 (I664152,I664135);
not I_38907 (I664169,I98219);
nor I_38908 (I664186,I664169,I98213);
and I_38909 (I664203,I664186,I98210);
or I_38910 (I664220,I664203,I98201);
DFFARX1 I_38911  ( .D(I664220), .CLK(I2702), .RSTB(I664033), .Q(I664237) );
nand I_38912 (I664254,I664050,I98219);
or I_38913 (I664022,I664254,I664237);
not I_38914 (I664285,I664254);
nor I_38915 (I664302,I664237,I664285);
and I_38916 (I664319,I664135,I664302);
nand I_38917 (I663995,I664254,I664152);
DFFARX1 I_38918  ( .D(I98231), .CLK(I2702), .RSTB(I664033), .Q(I664350) );
or I_38919 (I664016,I664350,I664237);
nor I_38920 (I664381,I664350,I664118);
nor I_38921 (I664398,I664350,I664152);
nand I_38922 (I664001,I664084,I664398);
or I_38923 (I664429,I664350,I664319);
DFFARX1 I_38924  ( .D(I664429), .CLK(I2702), .RSTB(I664033), .Q(I663998) );
not I_38925 (I664004,I664350);
DFFARX1 I_38926  ( .D(I98228), .CLK(I2702), .RSTB(I664033), .Q(I664474) );
not I_38927 (I664491,I664474);
nor I_38928 (I664508,I664491,I664084);
DFFARX1 I_38929  ( .D(I664508), .CLK(I2702), .RSTB(I664033), .Q(I664010) );
nor I_38930 (I664025,I664350,I664491);
nor I_38931 (I664013,I664491,I664254);
not I_38932 (I664567,I664491);
and I_38933 (I664584,I664118,I664567);
nor I_38934 (I664019,I664254,I664584);
nand I_38935 (I664007,I664491,I664381);
not I_38936 (I664662,I2709);
not I_38937 (I664679,I421751);
nor I_38938 (I664696,I421775,I421754);
nand I_38939 (I664713,I664696,I421760);
nor I_38940 (I664730,I664679,I421775);
nand I_38941 (I664747,I664730,I421772);
not I_38942 (I664764,I421775);
not I_38943 (I664781,I664764);
not I_38944 (I664798,I421769);
nor I_38945 (I664815,I664798,I421748);
and I_38946 (I664832,I664815,I421745);
or I_38947 (I664849,I664832,I421757);
DFFARX1 I_38948  ( .D(I664849), .CLK(I2702), .RSTB(I664662), .Q(I664866) );
nand I_38949 (I664883,I664679,I421769);
or I_38950 (I664651,I664883,I664866);
not I_38951 (I664914,I664883);
nor I_38952 (I664931,I664866,I664914);
and I_38953 (I664948,I664764,I664931);
nand I_38954 (I664624,I664883,I664781);
DFFARX1 I_38955  ( .D(I421763), .CLK(I2702), .RSTB(I664662), .Q(I664979) );
or I_38956 (I664645,I664979,I664866);
nor I_38957 (I665010,I664979,I664747);
nor I_38958 (I665027,I664979,I664781);
nand I_38959 (I664630,I664713,I665027);
or I_38960 (I665058,I664979,I664948);
DFFARX1 I_38961  ( .D(I665058), .CLK(I2702), .RSTB(I664662), .Q(I664627) );
not I_38962 (I664633,I664979);
DFFARX1 I_38963  ( .D(I421766), .CLK(I2702), .RSTB(I664662), .Q(I665103) );
not I_38964 (I665120,I665103);
nor I_38965 (I665137,I665120,I664713);
DFFARX1 I_38966  ( .D(I665137), .CLK(I2702), .RSTB(I664662), .Q(I664639) );
nor I_38967 (I664654,I664979,I665120);
nor I_38968 (I664642,I665120,I664883);
not I_38969 (I665196,I665120);
and I_38970 (I665213,I664747,I665196);
nor I_38971 (I664648,I664883,I665213);
nand I_38972 (I664636,I665120,I665010);
not I_38973 (I665291,I2709);
not I_38974 (I665308,I696148);
nor I_38975 (I665325,I696172,I696157);
nand I_38976 (I665342,I665325,I696142);
nor I_38977 (I665359,I665308,I696172);
nand I_38978 (I665376,I665359,I696169);
not I_38979 (I665393,I696172);
not I_38980 (I665410,I665393);
not I_38981 (I665427,I696151);
nor I_38982 (I665444,I665427,I696145);
and I_38983 (I665461,I665444,I696166);
or I_38984 (I665478,I665461,I696154);
DFFARX1 I_38985  ( .D(I665478), .CLK(I2702), .RSTB(I665291), .Q(I665495) );
nand I_38986 (I665512,I665308,I696151);
or I_38987 (I665280,I665512,I665495);
not I_38988 (I665543,I665512);
nor I_38989 (I665560,I665495,I665543);
and I_38990 (I665577,I665393,I665560);
nand I_38991 (I665253,I665512,I665410);
DFFARX1 I_38992  ( .D(I696163), .CLK(I2702), .RSTB(I665291), .Q(I665608) );
or I_38993 (I665274,I665608,I665495);
nor I_38994 (I665639,I665608,I665376);
nor I_38995 (I665656,I665608,I665410);
nand I_38996 (I665259,I665342,I665656);
or I_38997 (I665687,I665608,I665577);
DFFARX1 I_38998  ( .D(I665687), .CLK(I2702), .RSTB(I665291), .Q(I665256) );
not I_38999 (I665262,I665608);
DFFARX1 I_39000  ( .D(I696160), .CLK(I2702), .RSTB(I665291), .Q(I665732) );
not I_39001 (I665749,I665732);
nor I_39002 (I665766,I665749,I665342);
DFFARX1 I_39003  ( .D(I665766), .CLK(I2702), .RSTB(I665291), .Q(I665268) );
nor I_39004 (I665283,I665608,I665749);
nor I_39005 (I665271,I665749,I665512);
not I_39006 (I665825,I665749);
and I_39007 (I665842,I665376,I665825);
nor I_39008 (I665277,I665512,I665842);
nand I_39009 (I665265,I665749,I665639);
not I_39010 (I665920,I2709);
not I_39011 (I665937,I101437);
nor I_39012 (I665954,I101455,I101434);
nand I_39013 (I665971,I665954,I101452);
nor I_39014 (I665988,I665937,I101455);
nand I_39015 (I666005,I665988,I101446);
not I_39016 (I666022,I101455);
not I_39017 (I666039,I666022);
not I_39018 (I666056,I101449);
nor I_39019 (I666073,I666056,I101443);
and I_39020 (I666090,I666073,I101440);
or I_39021 (I666107,I666090,I101431);
DFFARX1 I_39022  ( .D(I666107), .CLK(I2702), .RSTB(I665920), .Q(I666124) );
nand I_39023 (I666141,I665937,I101449);
or I_39024 (I665909,I666141,I666124);
not I_39025 (I666172,I666141);
nor I_39026 (I666189,I666124,I666172);
and I_39027 (I666206,I666022,I666189);
nand I_39028 (I665882,I666141,I666039);
DFFARX1 I_39029  ( .D(I101461), .CLK(I2702), .RSTB(I665920), .Q(I666237) );
or I_39030 (I665903,I666237,I666124);
nor I_39031 (I666268,I666237,I666005);
nor I_39032 (I666285,I666237,I666039);
nand I_39033 (I665888,I665971,I666285);
or I_39034 (I666316,I666237,I666206);
DFFARX1 I_39035  ( .D(I666316), .CLK(I2702), .RSTB(I665920), .Q(I665885) );
not I_39036 (I665891,I666237);
DFFARX1 I_39037  ( .D(I101458), .CLK(I2702), .RSTB(I665920), .Q(I666361) );
not I_39038 (I666378,I666361);
nor I_39039 (I666395,I666378,I665971);
DFFARX1 I_39040  ( .D(I666395), .CLK(I2702), .RSTB(I665920), .Q(I665897) );
nor I_39041 (I665912,I666237,I666378);
nor I_39042 (I665900,I666378,I666141);
not I_39043 (I666454,I666378);
and I_39044 (I666471,I666005,I666454);
nor I_39045 (I665906,I666141,I666471);
nand I_39046 (I665894,I666378,I666268);
not I_39047 (I666549,I2709);
not I_39048 (I666566,I450641);
nor I_39049 (I666583,I450614,I450632);
nand I_39050 (I666600,I666583,I450617);
nor I_39051 (I666617,I666566,I450614);
nand I_39052 (I666634,I666617,I450635);
not I_39053 (I666651,I450614);
not I_39054 (I666668,I666651);
not I_39055 (I666685,I450611);
nor I_39056 (I666702,I666685,I450638);
and I_39057 (I666719,I666702,I450629);
or I_39058 (I666736,I666719,I450620);
DFFARX1 I_39059  ( .D(I666736), .CLK(I2702), .RSTB(I666549), .Q(I666753) );
nand I_39060 (I666770,I666566,I450611);
or I_39061 (I666538,I666770,I666753);
not I_39062 (I666801,I666770);
nor I_39063 (I666818,I666753,I666801);
and I_39064 (I666835,I666651,I666818);
nand I_39065 (I666511,I666770,I666668);
DFFARX1 I_39066  ( .D(I450623), .CLK(I2702), .RSTB(I666549), .Q(I666866) );
or I_39067 (I666532,I666866,I666753);
nor I_39068 (I666897,I666866,I666634);
nor I_39069 (I666914,I666866,I666668);
nand I_39070 (I666517,I666600,I666914);
or I_39071 (I666945,I666866,I666835);
DFFARX1 I_39072  ( .D(I666945), .CLK(I2702), .RSTB(I666549), .Q(I666514) );
not I_39073 (I666520,I666866);
DFFARX1 I_39074  ( .D(I450626), .CLK(I2702), .RSTB(I666549), .Q(I666990) );
not I_39075 (I667007,I666990);
nor I_39076 (I667024,I667007,I666600);
DFFARX1 I_39077  ( .D(I667024), .CLK(I2702), .RSTB(I666549), .Q(I666526) );
nor I_39078 (I666541,I666866,I667007);
nor I_39079 (I666529,I667007,I666770);
not I_39080 (I667083,I667007);
and I_39081 (I667100,I666634,I667083);
nor I_39082 (I666535,I666770,I667100);
nand I_39083 (I666523,I667007,I666897);
not I_39084 (I667178,I2709);
not I_39085 (I667195,I493769);
nor I_39086 (I667212,I493760,I493787);
nand I_39087 (I667229,I667212,I493757);
nor I_39088 (I667246,I667195,I493760);
nand I_39089 (I667263,I667246,I493781);
not I_39090 (I667280,I493760);
not I_39091 (I667297,I667280);
not I_39092 (I667314,I493766);
nor I_39093 (I667331,I667314,I493784);
and I_39094 (I667348,I667331,I493775);
or I_39095 (I667365,I667348,I493772);
DFFARX1 I_39096  ( .D(I667365), .CLK(I2702), .RSTB(I667178), .Q(I667382) );
nand I_39097 (I667399,I667195,I493766);
or I_39098 (I667167,I667399,I667382);
not I_39099 (I667430,I667399);
nor I_39100 (I667447,I667382,I667430);
and I_39101 (I667464,I667280,I667447);
nand I_39102 (I667140,I667399,I667297);
DFFARX1 I_39103  ( .D(I493763), .CLK(I2702), .RSTB(I667178), .Q(I667495) );
or I_39104 (I667161,I667495,I667382);
nor I_39105 (I667526,I667495,I667263);
nor I_39106 (I667543,I667495,I667297);
nand I_39107 (I667146,I667229,I667543);
or I_39108 (I667574,I667495,I667464);
DFFARX1 I_39109  ( .D(I667574), .CLK(I2702), .RSTB(I667178), .Q(I667143) );
not I_39110 (I667149,I667495);
DFFARX1 I_39111  ( .D(I493778), .CLK(I2702), .RSTB(I667178), .Q(I667619) );
not I_39112 (I667636,I667619);
nor I_39113 (I667653,I667636,I667229);
DFFARX1 I_39114  ( .D(I667653), .CLK(I2702), .RSTB(I667178), .Q(I667155) );
nor I_39115 (I667170,I667495,I667636);
nor I_39116 (I667158,I667636,I667399);
not I_39117 (I667712,I667636);
and I_39118 (I667729,I667263,I667712);
nor I_39119 (I667164,I667399,I667729);
nand I_39120 (I667152,I667636,I667526);
not I_39121 (I667807,I2709);
not I_39122 (I667824,I444861);
nor I_39123 (I667841,I444834,I444852);
nand I_39124 (I667858,I667841,I444837);
nor I_39125 (I667875,I667824,I444834);
nand I_39126 (I667892,I667875,I444855);
not I_39127 (I667909,I444834);
not I_39128 (I667926,I667909);
not I_39129 (I667943,I444831);
nor I_39130 (I667960,I667943,I444858);
and I_39131 (I667977,I667960,I444849);
or I_39132 (I667994,I667977,I444840);
DFFARX1 I_39133  ( .D(I667994), .CLK(I2702), .RSTB(I667807), .Q(I668011) );
nand I_39134 (I668028,I667824,I444831);
or I_39135 (I667796,I668028,I668011);
not I_39136 (I668059,I668028);
nor I_39137 (I668076,I668011,I668059);
and I_39138 (I668093,I667909,I668076);
nand I_39139 (I667769,I668028,I667926);
DFFARX1 I_39140  ( .D(I444843), .CLK(I2702), .RSTB(I667807), .Q(I668124) );
or I_39141 (I667790,I668124,I668011);
nor I_39142 (I668155,I668124,I667892);
nor I_39143 (I668172,I668124,I667926);
nand I_39144 (I667775,I667858,I668172);
or I_39145 (I668203,I668124,I668093);
DFFARX1 I_39146  ( .D(I668203), .CLK(I2702), .RSTB(I667807), .Q(I667772) );
not I_39147 (I667778,I668124);
DFFARX1 I_39148  ( .D(I444846), .CLK(I2702), .RSTB(I667807), .Q(I668248) );
not I_39149 (I668265,I668248);
nor I_39150 (I668282,I668265,I667858);
DFFARX1 I_39151  ( .D(I668282), .CLK(I2702), .RSTB(I667807), .Q(I667784) );
nor I_39152 (I667799,I668124,I668265);
nor I_39153 (I667787,I668265,I668028);
not I_39154 (I668341,I668265);
and I_39155 (I668358,I667892,I668341);
nor I_39156 (I667793,I668028,I668358);
nand I_39157 (I667781,I668265,I668155);
not I_39158 (I668436,I2709);
not I_39159 (I668453,I694992);
nor I_39160 (I668470,I695016,I695001);
nand I_39161 (I668487,I668470,I694986);
nor I_39162 (I668504,I668453,I695016);
nand I_39163 (I668521,I668504,I695013);
not I_39164 (I668538,I695016);
not I_39165 (I668555,I668538);
not I_39166 (I668572,I694995);
nor I_39167 (I668589,I668572,I694989);
and I_39168 (I668606,I668589,I695010);
or I_39169 (I668623,I668606,I694998);
DFFARX1 I_39170  ( .D(I668623), .CLK(I2702), .RSTB(I668436), .Q(I668640) );
nand I_39171 (I668657,I668453,I694995);
or I_39172 (I668425,I668657,I668640);
not I_39173 (I668688,I668657);
nor I_39174 (I668705,I668640,I668688);
and I_39175 (I668722,I668538,I668705);
nand I_39176 (I668398,I668657,I668555);
DFFARX1 I_39177  ( .D(I695007), .CLK(I2702), .RSTB(I668436), .Q(I668753) );
or I_39178 (I668419,I668753,I668640);
nor I_39179 (I668784,I668753,I668521);
nor I_39180 (I668801,I668753,I668555);
nand I_39181 (I668404,I668487,I668801);
or I_39182 (I668832,I668753,I668722);
DFFARX1 I_39183  ( .D(I668832), .CLK(I2702), .RSTB(I668436), .Q(I668401) );
not I_39184 (I668407,I668753);
DFFARX1 I_39185  ( .D(I695004), .CLK(I2702), .RSTB(I668436), .Q(I668877) );
not I_39186 (I668894,I668877);
nor I_39187 (I668911,I668894,I668487);
DFFARX1 I_39188  ( .D(I668911), .CLK(I2702), .RSTB(I668436), .Q(I668413) );
nor I_39189 (I668428,I668753,I668894);
nor I_39190 (I668416,I668894,I668657);
not I_39191 (I668970,I668894);
and I_39192 (I668987,I668521,I668970);
nor I_39193 (I668422,I668657,I668987);
nand I_39194 (I668410,I668894,I668784);
not I_39195 (I669065,I2709);
not I_39196 (I669082,I121463);
nor I_39197 (I669099,I121481,I121460);
nand I_39198 (I669116,I669099,I121478);
nor I_39199 (I669133,I669082,I121481);
nand I_39200 (I669150,I669133,I121472);
not I_39201 (I669167,I121481);
not I_39202 (I669184,I669167);
not I_39203 (I669201,I121475);
nor I_39204 (I669218,I669201,I121469);
and I_39205 (I669235,I669218,I121466);
or I_39206 (I669252,I669235,I121457);
DFFARX1 I_39207  ( .D(I669252), .CLK(I2702), .RSTB(I669065), .Q(I669269) );
nand I_39208 (I669286,I669082,I121475);
or I_39209 (I669054,I669286,I669269);
not I_39210 (I669317,I669286);
nor I_39211 (I669334,I669269,I669317);
and I_39212 (I669351,I669167,I669334);
nand I_39213 (I669027,I669286,I669184);
DFFARX1 I_39214  ( .D(I121487), .CLK(I2702), .RSTB(I669065), .Q(I669382) );
or I_39215 (I669048,I669382,I669269);
nor I_39216 (I669413,I669382,I669150);
nor I_39217 (I669430,I669382,I669184);
nand I_39218 (I669033,I669116,I669430);
or I_39219 (I669461,I669382,I669351);
DFFARX1 I_39220  ( .D(I669461), .CLK(I2702), .RSTB(I669065), .Q(I669030) );
not I_39221 (I669036,I669382);
DFFARX1 I_39222  ( .D(I121484), .CLK(I2702), .RSTB(I669065), .Q(I669506) );
not I_39223 (I669523,I669506);
nor I_39224 (I669540,I669523,I669116);
DFFARX1 I_39225  ( .D(I669540), .CLK(I2702), .RSTB(I669065), .Q(I669042) );
nor I_39226 (I669057,I669382,I669523);
nor I_39227 (I669045,I669523,I669286);
not I_39228 (I669599,I669523);
and I_39229 (I669616,I669150,I669599);
nor I_39230 (I669051,I669286,I669616);
nand I_39231 (I669039,I669523,I669413);
not I_39232 (I669694,I2709);
not I_39233 (I669711,I130507);
nor I_39234 (I669728,I130525,I130504);
nand I_39235 (I669745,I669728,I130522);
nor I_39236 (I669762,I669711,I130525);
nand I_39237 (I669779,I669762,I130516);
not I_39238 (I669796,I130525);
not I_39239 (I669813,I669796);
not I_39240 (I669830,I130519);
nor I_39241 (I669847,I669830,I130513);
and I_39242 (I669864,I669847,I130510);
or I_39243 (I669881,I669864,I130501);
DFFARX1 I_39244  ( .D(I669881), .CLK(I2702), .RSTB(I669694), .Q(I669898) );
nand I_39245 (I669915,I669711,I130519);
or I_39246 (I669683,I669915,I669898);
not I_39247 (I669946,I669915);
nor I_39248 (I669963,I669898,I669946);
and I_39249 (I669980,I669796,I669963);
nand I_39250 (I669656,I669915,I669813);
DFFARX1 I_39251  ( .D(I130531), .CLK(I2702), .RSTB(I669694), .Q(I670011) );
or I_39252 (I669677,I670011,I669898);
nor I_39253 (I670042,I670011,I669779);
nor I_39254 (I670059,I670011,I669813);
nand I_39255 (I669662,I669745,I670059);
or I_39256 (I670090,I670011,I669980);
DFFARX1 I_39257  ( .D(I670090), .CLK(I2702), .RSTB(I669694), .Q(I669659) );
not I_39258 (I669665,I670011);
DFFARX1 I_39259  ( .D(I130528), .CLK(I2702), .RSTB(I669694), .Q(I670135) );
not I_39260 (I670152,I670135);
nor I_39261 (I670169,I670152,I669745);
DFFARX1 I_39262  ( .D(I670169), .CLK(I2702), .RSTB(I669694), .Q(I669671) );
nor I_39263 (I669686,I670011,I670152);
nor I_39264 (I669674,I670152,I669915);
not I_39265 (I670228,I670152);
and I_39266 (I670245,I669779,I670228);
nor I_39267 (I669680,I669915,I670245);
nand I_39268 (I669668,I670152,I670042);
not I_39269 (I670323,I2709);
not I_39270 (I670340,I564330);
nor I_39271 (I670357,I564348,I564327);
nand I_39272 (I670374,I670357,I564351);
nor I_39273 (I670391,I670340,I564348);
nand I_39274 (I670408,I670391,I564345);
not I_39275 (I670425,I564348);
not I_39276 (I670442,I670425);
not I_39277 (I670459,I564336);
nor I_39278 (I670476,I670459,I564324);
and I_39279 (I670493,I670476,I564342);
or I_39280 (I670510,I670493,I564354);
DFFARX1 I_39281  ( .D(I670510), .CLK(I2702), .RSTB(I670323), .Q(I670527) );
nand I_39282 (I670544,I670340,I564336);
or I_39283 (I670312,I670544,I670527);
not I_39284 (I670575,I670544);
nor I_39285 (I670592,I670527,I670575);
and I_39286 (I670609,I670425,I670592);
nand I_39287 (I670285,I670544,I670442);
DFFARX1 I_39288  ( .D(I564333), .CLK(I2702), .RSTB(I670323), .Q(I670640) );
or I_39289 (I670306,I670640,I670527);
nor I_39290 (I670671,I670640,I670408);
nor I_39291 (I670688,I670640,I670442);
nand I_39292 (I670291,I670374,I670688);
or I_39293 (I670719,I670640,I670609);
DFFARX1 I_39294  ( .D(I670719), .CLK(I2702), .RSTB(I670323), .Q(I670288) );
not I_39295 (I670294,I670640);
DFFARX1 I_39296  ( .D(I564339), .CLK(I2702), .RSTB(I670323), .Q(I670764) );
not I_39297 (I670781,I670764);
nor I_39298 (I670798,I670781,I670374);
DFFARX1 I_39299  ( .D(I670798), .CLK(I2702), .RSTB(I670323), .Q(I670300) );
nor I_39300 (I670315,I670640,I670781);
nor I_39301 (I670303,I670781,I670544);
not I_39302 (I670857,I670781);
and I_39303 (I670874,I670408,I670857);
nor I_39304 (I670309,I670544,I670874);
nand I_39305 (I670297,I670781,I670671);
not I_39306 (I670952,I2709);
not I_39307 (I670969,I119525);
nor I_39308 (I670986,I119543,I119522);
nand I_39309 (I671003,I670986,I119540);
nor I_39310 (I671020,I670969,I119543);
nand I_39311 (I671037,I671020,I119534);
not I_39312 (I671054,I119543);
not I_39313 (I671071,I671054);
not I_39314 (I671088,I119537);
nor I_39315 (I671105,I671088,I119531);
and I_39316 (I671122,I671105,I119528);
or I_39317 (I671139,I671122,I119519);
DFFARX1 I_39318  ( .D(I671139), .CLK(I2702), .RSTB(I670952), .Q(I671156) );
nand I_39319 (I671173,I670969,I119537);
or I_39320 (I670941,I671173,I671156);
not I_39321 (I671204,I671173);
nor I_39322 (I671221,I671156,I671204);
and I_39323 (I671238,I671054,I671221);
nand I_39324 (I670914,I671173,I671071);
DFFARX1 I_39325  ( .D(I119549), .CLK(I2702), .RSTB(I670952), .Q(I671269) );
or I_39326 (I670935,I671269,I671156);
nor I_39327 (I671300,I671269,I671037);
nor I_39328 (I671317,I671269,I671071);
nand I_39329 (I670920,I671003,I671317);
or I_39330 (I671348,I671269,I671238);
DFFARX1 I_39331  ( .D(I671348), .CLK(I2702), .RSTB(I670952), .Q(I670917) );
not I_39332 (I670923,I671269);
DFFARX1 I_39333  ( .D(I119546), .CLK(I2702), .RSTB(I670952), .Q(I671393) );
not I_39334 (I671410,I671393);
nor I_39335 (I671427,I671410,I671003);
DFFARX1 I_39336  ( .D(I671427), .CLK(I2702), .RSTB(I670952), .Q(I670929) );
nor I_39337 (I670944,I671269,I671410);
nor I_39338 (I670932,I671410,I671173);
not I_39339 (I671486,I671410);
and I_39340 (I671503,I671037,I671486);
nor I_39341 (I670938,I671173,I671503);
nand I_39342 (I670926,I671410,I671300);
not I_39343 (I671581,I2709);
not I_39344 (I671598,I380317);
nor I_39345 (I671615,I380326,I380329);
nand I_39346 (I671632,I671615,I380314);
nor I_39347 (I671649,I671598,I380326);
nand I_39348 (I671666,I671649,I380311);
not I_39349 (I671683,I380326);
not I_39350 (I671700,I671683);
not I_39351 (I671717,I380299);
nor I_39352 (I671734,I671717,I380305);
and I_39353 (I671751,I671734,I380302);
or I_39354 (I671768,I671751,I380323);
DFFARX1 I_39355  ( .D(I671768), .CLK(I2702), .RSTB(I671581), .Q(I671785) );
nand I_39356 (I671802,I671598,I380299);
or I_39357 (I671570,I671802,I671785);
not I_39358 (I671833,I671802);
nor I_39359 (I671850,I671785,I671833);
and I_39360 (I671867,I671683,I671850);
nand I_39361 (I671543,I671802,I671700);
DFFARX1 I_39362  ( .D(I380308), .CLK(I2702), .RSTB(I671581), .Q(I671898) );
or I_39363 (I671564,I671898,I671785);
nor I_39364 (I671929,I671898,I671666);
nor I_39365 (I671946,I671898,I671700);
nand I_39366 (I671549,I671632,I671946);
or I_39367 (I671977,I671898,I671867);
DFFARX1 I_39368  ( .D(I671977), .CLK(I2702), .RSTB(I671581), .Q(I671546) );
not I_39369 (I671552,I671898);
DFFARX1 I_39370  ( .D(I380320), .CLK(I2702), .RSTB(I671581), .Q(I672022) );
not I_39371 (I672039,I672022);
nor I_39372 (I672056,I672039,I671632);
DFFARX1 I_39373  ( .D(I672056), .CLK(I2702), .RSTB(I671581), .Q(I671558) );
nor I_39374 (I671573,I671898,I672039);
nor I_39375 (I671561,I672039,I671802);
not I_39376 (I672115,I672039);
and I_39377 (I672132,I671666,I672115);
nor I_39378 (I671567,I671802,I672132);
nand I_39379 (I671555,I672039,I671929);
not I_39380 (I672210,I2709);
not I_39381 (I672227,I120817);
nor I_39382 (I672244,I120835,I120814);
nand I_39383 (I672261,I672244,I120832);
nor I_39384 (I672278,I672227,I120835);
nand I_39385 (I672295,I672278,I120826);
not I_39386 (I672312,I120835);
not I_39387 (I672329,I672312);
not I_39388 (I672346,I120829);
nor I_39389 (I672363,I672346,I120823);
and I_39390 (I672380,I672363,I120820);
or I_39391 (I672397,I672380,I120811);
DFFARX1 I_39392  ( .D(I672397), .CLK(I2702), .RSTB(I672210), .Q(I672414) );
nand I_39393 (I672431,I672227,I120829);
or I_39394 (I672199,I672431,I672414);
not I_39395 (I672462,I672431);
nor I_39396 (I672479,I672414,I672462);
and I_39397 (I672496,I672312,I672479);
nand I_39398 (I672172,I672431,I672329);
DFFARX1 I_39399  ( .D(I120841), .CLK(I2702), .RSTB(I672210), .Q(I672527) );
or I_39400 (I672193,I672527,I672414);
nor I_39401 (I672558,I672527,I672295);
nor I_39402 (I672575,I672527,I672329);
nand I_39403 (I672178,I672261,I672575);
or I_39404 (I672606,I672527,I672496);
DFFARX1 I_39405  ( .D(I672606), .CLK(I2702), .RSTB(I672210), .Q(I672175) );
not I_39406 (I672181,I672527);
DFFARX1 I_39407  ( .D(I120838), .CLK(I2702), .RSTB(I672210), .Q(I672651) );
not I_39408 (I672668,I672651);
nor I_39409 (I672685,I672668,I672261);
DFFARX1 I_39410  ( .D(I672685), .CLK(I2702), .RSTB(I672210), .Q(I672187) );
nor I_39411 (I672202,I672527,I672668);
nor I_39412 (I672190,I672668,I672431);
not I_39413 (I672744,I672668);
and I_39414 (I672761,I672295,I672744);
nor I_39415 (I672196,I672431,I672761);
nand I_39416 (I672184,I672668,I672558);
not I_39417 (I672839,I2709);
not I_39418 (I672856,I117587);
nor I_39419 (I672873,I117605,I117584);
nand I_39420 (I672890,I672873,I117602);
nor I_39421 (I672907,I672856,I117605);
nand I_39422 (I672924,I672907,I117596);
not I_39423 (I672941,I117605);
not I_39424 (I672958,I672941);
not I_39425 (I672975,I117599);
nor I_39426 (I672992,I672975,I117593);
and I_39427 (I673009,I672992,I117590);
or I_39428 (I673026,I673009,I117581);
DFFARX1 I_39429  ( .D(I673026), .CLK(I2702), .RSTB(I672839), .Q(I673043) );
nand I_39430 (I673060,I672856,I117599);
or I_39431 (I672828,I673060,I673043);
not I_39432 (I673091,I673060);
nor I_39433 (I673108,I673043,I673091);
and I_39434 (I673125,I672941,I673108);
nand I_39435 (I672801,I673060,I672958);
DFFARX1 I_39436  ( .D(I117611), .CLK(I2702), .RSTB(I672839), .Q(I673156) );
or I_39437 (I672822,I673156,I673043);
nor I_39438 (I673187,I673156,I672924);
nor I_39439 (I673204,I673156,I672958);
nand I_39440 (I672807,I672890,I673204);
or I_39441 (I673235,I673156,I673125);
DFFARX1 I_39442  ( .D(I673235), .CLK(I2702), .RSTB(I672839), .Q(I672804) );
not I_39443 (I672810,I673156);
DFFARX1 I_39444  ( .D(I117608), .CLK(I2702), .RSTB(I672839), .Q(I673280) );
not I_39445 (I673297,I673280);
nor I_39446 (I673314,I673297,I672890);
DFFARX1 I_39447  ( .D(I673314), .CLK(I2702), .RSTB(I672839), .Q(I672816) );
nor I_39448 (I672831,I673156,I673297);
nor I_39449 (I672819,I673297,I673060);
not I_39450 (I673373,I673297);
and I_39451 (I673390,I672924,I673373);
nor I_39452 (I672825,I673060,I673390);
nand I_39453 (I672813,I673297,I673187);
not I_39454 (I673468,I2709);
not I_39455 (I673485,I24594);
nor I_39456 (I673502,I24597,I24606);
nand I_39457 (I673519,I673502,I24621);
nor I_39458 (I673536,I673485,I24597);
nand I_39459 (I673553,I673536,I24600);
not I_39460 (I673570,I24597);
not I_39461 (I673587,I673570);
not I_39462 (I673604,I24591);
nor I_39463 (I673621,I673604,I24615);
and I_39464 (I673638,I673621,I24603);
or I_39465 (I673655,I673638,I24609);
DFFARX1 I_39466  ( .D(I673655), .CLK(I2702), .RSTB(I673468), .Q(I673672) );
nand I_39467 (I673689,I673485,I24591);
or I_39468 (I673457,I673689,I673672);
not I_39469 (I673720,I673689);
nor I_39470 (I673737,I673672,I673720);
and I_39471 (I673754,I673570,I673737);
nand I_39472 (I673430,I673689,I673587);
DFFARX1 I_39473  ( .D(I24612), .CLK(I2702), .RSTB(I673468), .Q(I673785) );
or I_39474 (I673451,I673785,I673672);
nor I_39475 (I673816,I673785,I673553);
nor I_39476 (I673833,I673785,I673587);
nand I_39477 (I673436,I673519,I673833);
or I_39478 (I673864,I673785,I673754);
DFFARX1 I_39479  ( .D(I673864), .CLK(I2702), .RSTB(I673468), .Q(I673433) );
not I_39480 (I673439,I673785);
DFFARX1 I_39481  ( .D(I24618), .CLK(I2702), .RSTB(I673468), .Q(I673909) );
not I_39482 (I673926,I673909);
nor I_39483 (I673943,I673926,I673519);
DFFARX1 I_39484  ( .D(I673943), .CLK(I2702), .RSTB(I673468), .Q(I673445) );
nor I_39485 (I673460,I673785,I673926);
nor I_39486 (I673448,I673926,I673689);
not I_39487 (I674002,I673926);
and I_39488 (I674019,I673553,I674002);
nor I_39489 (I673454,I673689,I674019);
nand I_39490 (I673442,I673926,I673816);
not I_39491 (I674097,I2709);
not I_39492 (I674114,I157458);
nor I_39493 (I674131,I157449,I157473);
nand I_39494 (I674148,I674131,I157476);
nor I_39495 (I674165,I674114,I157449);
nand I_39496 (I674182,I674165,I157467);
not I_39497 (I674199,I157449);
not I_39498 (I674216,I674199);
not I_39499 (I674233,I157461);
nor I_39500 (I674250,I674233,I157455);
and I_39501 (I674267,I674250,I157464);
or I_39502 (I674284,I674267,I157452);
DFFARX1 I_39503  ( .D(I674284), .CLK(I2702), .RSTB(I674097), .Q(I674301) );
nand I_39504 (I674318,I674114,I157461);
or I_39505 (I674086,I674318,I674301);
not I_39506 (I674349,I674318);
nor I_39507 (I674366,I674301,I674349);
and I_39508 (I674383,I674199,I674366);
nand I_39509 (I674059,I674318,I674216);
DFFARX1 I_39510  ( .D(I157446), .CLK(I2702), .RSTB(I674097), .Q(I674414) );
or I_39511 (I674080,I674414,I674301);
nor I_39512 (I674445,I674414,I674182);
nor I_39513 (I674462,I674414,I674216);
nand I_39514 (I674065,I674148,I674462);
or I_39515 (I674493,I674414,I674383);
DFFARX1 I_39516  ( .D(I674493), .CLK(I2702), .RSTB(I674097), .Q(I674062) );
not I_39517 (I674068,I674414);
DFFARX1 I_39518  ( .D(I157470), .CLK(I2702), .RSTB(I674097), .Q(I674538) );
not I_39519 (I674555,I674538);
nor I_39520 (I674572,I674555,I674148);
DFFARX1 I_39521  ( .D(I674572), .CLK(I2702), .RSTB(I674097), .Q(I674074) );
nor I_39522 (I674089,I674414,I674555);
nor I_39523 (I674077,I674555,I674318);
not I_39524 (I674631,I674555);
and I_39525 (I674648,I674182,I674631);
nor I_39526 (I674083,I674318,I674648);
nand I_39527 (I674071,I674555,I674445);
not I_39528 (I674726,I2709);
not I_39529 (I674743,I2383);
nor I_39530 (I674760,I1367,I2151);
nand I_39531 (I674777,I674760,I2255);
nor I_39532 (I674794,I674743,I1367);
nand I_39533 (I674811,I674794,I1887);
not I_39534 (I674828,I1367);
not I_39535 (I674845,I674828);
not I_39536 (I674862,I2191);
nor I_39537 (I674879,I674862,I1415);
and I_39538 (I674896,I674879,I2143);
or I_39539 (I674913,I674896,I2559);
DFFARX1 I_39540  ( .D(I674913), .CLK(I2702), .RSTB(I674726), .Q(I674930) );
nand I_39541 (I674947,I674743,I2191);
or I_39542 (I674715,I674947,I674930);
not I_39543 (I674978,I674947);
nor I_39544 (I674995,I674930,I674978);
and I_39545 (I675012,I674828,I674995);
nand I_39546 (I674688,I674947,I674845);
DFFARX1 I_39547  ( .D(I1383), .CLK(I2702), .RSTB(I674726), .Q(I675043) );
or I_39548 (I674709,I675043,I674930);
nor I_39549 (I675074,I675043,I674811);
nor I_39550 (I675091,I675043,I674845);
nand I_39551 (I674694,I674777,I675091);
or I_39552 (I675122,I675043,I675012);
DFFARX1 I_39553  ( .D(I675122), .CLK(I2702), .RSTB(I674726), .Q(I674691) );
not I_39554 (I674697,I675043);
DFFARX1 I_39555  ( .D(I2607), .CLK(I2702), .RSTB(I674726), .Q(I675167) );
not I_39556 (I675184,I675167);
nor I_39557 (I675201,I675184,I674777);
DFFARX1 I_39558  ( .D(I675201), .CLK(I2702), .RSTB(I674726), .Q(I674703) );
nor I_39559 (I674718,I675043,I675184);
nor I_39560 (I674706,I675184,I674947);
not I_39561 (I675260,I675184);
and I_39562 (I675277,I674811,I675260);
nor I_39563 (I674712,I674947,I675277);
nand I_39564 (I674700,I675184,I675074);
not I_39565 (I675355,I2709);
not I_39566 (I675372,I511970);
nor I_39567 (I675389,I511988,I511967);
nand I_39568 (I675406,I675389,I511991);
nor I_39569 (I675423,I675372,I511988);
nand I_39570 (I675440,I675423,I511985);
not I_39571 (I675457,I511988);
not I_39572 (I675474,I675457);
not I_39573 (I675491,I511976);
nor I_39574 (I675508,I675491,I511964);
and I_39575 (I675525,I675508,I511982);
or I_39576 (I675542,I675525,I511994);
DFFARX1 I_39577  ( .D(I675542), .CLK(I2702), .RSTB(I675355), .Q(I675559) );
nand I_39578 (I675576,I675372,I511976);
or I_39579 (I675344,I675576,I675559);
not I_39580 (I675607,I675576);
nor I_39581 (I675624,I675559,I675607);
and I_39582 (I675641,I675457,I675624);
nand I_39583 (I675317,I675576,I675474);
DFFARX1 I_39584  ( .D(I511973), .CLK(I2702), .RSTB(I675355), .Q(I675672) );
or I_39585 (I675338,I675672,I675559);
nor I_39586 (I675703,I675672,I675440);
nor I_39587 (I675720,I675672,I675474);
nand I_39588 (I675323,I675406,I675720);
or I_39589 (I675751,I675672,I675641);
DFFARX1 I_39590  ( .D(I675751), .CLK(I2702), .RSTB(I675355), .Q(I675320) );
not I_39591 (I675326,I675672);
DFFARX1 I_39592  ( .D(I511979), .CLK(I2702), .RSTB(I675355), .Q(I675796) );
not I_39593 (I675813,I675796);
nor I_39594 (I675830,I675813,I675406);
DFFARX1 I_39595  ( .D(I675830), .CLK(I2702), .RSTB(I675355), .Q(I675332) );
nor I_39596 (I675347,I675672,I675813);
nor I_39597 (I675335,I675813,I675576);
not I_39598 (I675889,I675813);
and I_39599 (I675906,I675440,I675889);
nor I_39600 (I675341,I675576,I675906);
nand I_39601 (I675329,I675813,I675703);
not I_39602 (I675984,I2709);
not I_39603 (I676001,I525655);
nor I_39604 (I676018,I525673,I525652);
nand I_39605 (I676035,I676018,I525676);
nor I_39606 (I676052,I676001,I525673);
nand I_39607 (I676069,I676052,I525670);
not I_39608 (I676086,I525673);
not I_39609 (I676103,I676086);
not I_39610 (I676120,I525661);
nor I_39611 (I676137,I676120,I525649);
and I_39612 (I676154,I676137,I525667);
or I_39613 (I676171,I676154,I525679);
DFFARX1 I_39614  ( .D(I676171), .CLK(I2702), .RSTB(I675984), .Q(I676188) );
nand I_39615 (I676205,I676001,I525661);
or I_39616 (I675973,I676205,I676188);
not I_39617 (I676236,I676205);
nor I_39618 (I676253,I676188,I676236);
and I_39619 (I676270,I676086,I676253);
nand I_39620 (I675946,I676205,I676103);
DFFARX1 I_39621  ( .D(I525658), .CLK(I2702), .RSTB(I675984), .Q(I676301) );
or I_39622 (I675967,I676301,I676188);
nor I_39623 (I676332,I676301,I676069);
nor I_39624 (I676349,I676301,I676103);
nand I_39625 (I675952,I676035,I676349);
or I_39626 (I676380,I676301,I676270);
DFFARX1 I_39627  ( .D(I676380), .CLK(I2702), .RSTB(I675984), .Q(I675949) );
not I_39628 (I675955,I676301);
DFFARX1 I_39629  ( .D(I525664), .CLK(I2702), .RSTB(I675984), .Q(I676425) );
not I_39630 (I676442,I676425);
nor I_39631 (I676459,I676442,I676035);
DFFARX1 I_39632  ( .D(I676459), .CLK(I2702), .RSTB(I675984), .Q(I675961) );
nor I_39633 (I675976,I676301,I676442);
nor I_39634 (I675964,I676442,I676205);
not I_39635 (I676518,I676442);
and I_39636 (I676535,I676069,I676518);
nor I_39637 (I675970,I676205,I676535);
nand I_39638 (I675958,I676442,I676332);
not I_39639 (I676613,I2709);
not I_39640 (I676630,I306639);
nor I_39641 (I676647,I306645,I306624);
nand I_39642 (I676664,I676647,I306630);
nor I_39643 (I676681,I676630,I306645);
nand I_39644 (I676698,I676681,I306636);
not I_39645 (I676715,I306645);
not I_39646 (I676732,I676715);
not I_39647 (I676749,I306633);
nor I_39648 (I676766,I676749,I306651);
and I_39649 (I676783,I676766,I306642);
or I_39650 (I676800,I676783,I306621);
DFFARX1 I_39651  ( .D(I676800), .CLK(I2702), .RSTB(I676613), .Q(I676817) );
nand I_39652 (I676834,I676630,I306633);
or I_39653 (I676602,I676834,I676817);
not I_39654 (I676865,I676834);
nor I_39655 (I676882,I676817,I676865);
and I_39656 (I676899,I676715,I676882);
nand I_39657 (I676575,I676834,I676732);
DFFARX1 I_39658  ( .D(I306648), .CLK(I2702), .RSTB(I676613), .Q(I676930) );
or I_39659 (I676596,I676930,I676817);
nor I_39660 (I676961,I676930,I676698);
nor I_39661 (I676978,I676930,I676732);
nand I_39662 (I676581,I676664,I676978);
or I_39663 (I677009,I676930,I676899);
DFFARX1 I_39664  ( .D(I677009), .CLK(I2702), .RSTB(I676613), .Q(I676578) );
not I_39665 (I676584,I676930);
DFFARX1 I_39666  ( .D(I306627), .CLK(I2702), .RSTB(I676613), .Q(I677054) );
not I_39667 (I677071,I677054);
nor I_39668 (I677088,I677071,I676664);
DFFARX1 I_39669  ( .D(I677088), .CLK(I2702), .RSTB(I676613), .Q(I676590) );
nor I_39670 (I676605,I676930,I677071);
nor I_39671 (I676593,I677071,I676834);
not I_39672 (I677147,I677071);
and I_39673 (I677164,I676698,I677147);
nor I_39674 (I676599,I676834,I677164);
nand I_39675 (I676587,I677071,I676961);
not I_39676 (I677242,I2709);
not I_39677 (I677259,I718112);
nor I_39678 (I677276,I718136,I718121);
nand I_39679 (I677293,I677276,I718106);
nor I_39680 (I677310,I677259,I718136);
nand I_39681 (I677327,I677310,I718133);
not I_39682 (I677344,I718136);
not I_39683 (I677361,I677344);
not I_39684 (I677378,I718115);
nor I_39685 (I677395,I677378,I718109);
and I_39686 (I677412,I677395,I718130);
or I_39687 (I677429,I677412,I718118);
DFFARX1 I_39688  ( .D(I677429), .CLK(I2702), .RSTB(I677242), .Q(I677446) );
nand I_39689 (I677463,I677259,I718115);
or I_39690 (I677231,I677463,I677446);
not I_39691 (I677494,I677463);
nor I_39692 (I677511,I677446,I677494);
and I_39693 (I677528,I677344,I677511);
nand I_39694 (I677204,I677463,I677361);
DFFARX1 I_39695  ( .D(I718127), .CLK(I2702), .RSTB(I677242), .Q(I677559) );
or I_39696 (I677225,I677559,I677446);
nor I_39697 (I677590,I677559,I677327);
nor I_39698 (I677607,I677559,I677361);
nand I_39699 (I677210,I677293,I677607);
or I_39700 (I677638,I677559,I677528);
DFFARX1 I_39701  ( .D(I677638), .CLK(I2702), .RSTB(I677242), .Q(I677207) );
not I_39702 (I677213,I677559);
DFFARX1 I_39703  ( .D(I718124), .CLK(I2702), .RSTB(I677242), .Q(I677683) );
not I_39704 (I677700,I677683);
nor I_39705 (I677717,I677700,I677293);
DFFARX1 I_39706  ( .D(I677717), .CLK(I2702), .RSTB(I677242), .Q(I677219) );
nor I_39707 (I677234,I677559,I677700);
nor I_39708 (I677222,I677700,I677463);
not I_39709 (I677776,I677700);
and I_39710 (I677793,I677327,I677776);
nor I_39711 (I677228,I677463,I677793);
nand I_39712 (I677216,I677700,I677590);
not I_39713 (I677871,I2709);
not I_39714 (I677888,I401635);
nor I_39715 (I677905,I401644,I401647);
nand I_39716 (I677922,I677905,I401632);
nor I_39717 (I677939,I677888,I401644);
nand I_39718 (I677956,I677939,I401629);
not I_39719 (I677973,I401644);
not I_39720 (I677990,I677973);
not I_39721 (I678007,I401617);
nor I_39722 (I678024,I678007,I401623);
and I_39723 (I678041,I678024,I401620);
or I_39724 (I678058,I678041,I401641);
DFFARX1 I_39725  ( .D(I678058), .CLK(I2702), .RSTB(I677871), .Q(I678075) );
nand I_39726 (I678092,I677888,I401617);
or I_39727 (I677860,I678092,I678075);
not I_39728 (I678123,I678092);
nor I_39729 (I678140,I678075,I678123);
and I_39730 (I678157,I677973,I678140);
nand I_39731 (I677833,I678092,I677990);
DFFARX1 I_39732  ( .D(I401626), .CLK(I2702), .RSTB(I677871), .Q(I678188) );
or I_39733 (I677854,I678188,I678075);
nor I_39734 (I678219,I678188,I677956);
nor I_39735 (I678236,I678188,I677990);
nand I_39736 (I677839,I677922,I678236);
or I_39737 (I678267,I678188,I678157);
DFFARX1 I_39738  ( .D(I678267), .CLK(I2702), .RSTB(I677871), .Q(I677836) );
not I_39739 (I677842,I678188);
DFFARX1 I_39740  ( .D(I401638), .CLK(I2702), .RSTB(I677871), .Q(I678312) );
not I_39741 (I678329,I678312);
nor I_39742 (I678346,I678329,I677922);
DFFARX1 I_39743  ( .D(I678346), .CLK(I2702), .RSTB(I677871), .Q(I677848) );
nor I_39744 (I677863,I678188,I678329);
nor I_39745 (I677851,I678329,I678092);
not I_39746 (I678405,I678329);
and I_39747 (I678422,I677956,I678405);
nor I_39748 (I677857,I678092,I678422);
nand I_39749 (I677845,I678329,I678219);
not I_39750 (I678500,I2709);
not I_39751 (I678517,I272163);
nor I_39752 (I678534,I272169,I272148);
nand I_39753 (I678551,I678534,I272154);
nor I_39754 (I678568,I678517,I272169);
nand I_39755 (I678585,I678568,I272160);
not I_39756 (I678602,I272169);
not I_39757 (I678619,I678602);
not I_39758 (I678636,I272157);
nor I_39759 (I678653,I678636,I272175);
and I_39760 (I678670,I678653,I272166);
or I_39761 (I678687,I678670,I272145);
DFFARX1 I_39762  ( .D(I678687), .CLK(I2702), .RSTB(I678500), .Q(I678704) );
nand I_39763 (I678721,I678517,I272157);
or I_39764 (I678489,I678721,I678704);
not I_39765 (I678752,I678721);
nor I_39766 (I678769,I678704,I678752);
and I_39767 (I678786,I678602,I678769);
nand I_39768 (I678462,I678721,I678619);
DFFARX1 I_39769  ( .D(I272172), .CLK(I2702), .RSTB(I678500), .Q(I678817) );
or I_39770 (I678483,I678817,I678704);
nor I_39771 (I678848,I678817,I678585);
nor I_39772 (I678865,I678817,I678619);
nand I_39773 (I678468,I678551,I678865);
or I_39774 (I678896,I678817,I678786);
DFFARX1 I_39775  ( .D(I678896), .CLK(I2702), .RSTB(I678500), .Q(I678465) );
not I_39776 (I678471,I678817);
DFFARX1 I_39777  ( .D(I272151), .CLK(I2702), .RSTB(I678500), .Q(I678941) );
not I_39778 (I678958,I678941);
nor I_39779 (I678975,I678958,I678551);
DFFARX1 I_39780  ( .D(I678975), .CLK(I2702), .RSTB(I678500), .Q(I678477) );
nor I_39781 (I678492,I678817,I678958);
nor I_39782 (I678480,I678958,I678721);
not I_39783 (I679034,I678958);
and I_39784 (I679051,I678585,I679034);
nor I_39785 (I678486,I678721,I679051);
nand I_39786 (I678474,I678958,I678848);
not I_39787 (I679129,I2709);
not I_39788 (I679146,I279456);
nor I_39789 (I679163,I279462,I279441);
nand I_39790 (I679180,I679163,I279447);
nor I_39791 (I679197,I679146,I279462);
nand I_39792 (I679214,I679197,I279453);
not I_39793 (I679231,I279462);
not I_39794 (I679248,I679231);
not I_39795 (I679265,I279450);
nor I_39796 (I679282,I679265,I279468);
and I_39797 (I679299,I679282,I279459);
or I_39798 (I679316,I679299,I279438);
DFFARX1 I_39799  ( .D(I679316), .CLK(I2702), .RSTB(I679129), .Q(I679333) );
nand I_39800 (I679350,I679146,I279450);
or I_39801 (I679118,I679350,I679333);
not I_39802 (I679381,I679350);
nor I_39803 (I679398,I679333,I679381);
and I_39804 (I679415,I679231,I679398);
nand I_39805 (I679091,I679350,I679248);
DFFARX1 I_39806  ( .D(I279465), .CLK(I2702), .RSTB(I679129), .Q(I679446) );
or I_39807 (I679112,I679446,I679333);
nor I_39808 (I679477,I679446,I679214);
nor I_39809 (I679494,I679446,I679248);
nand I_39810 (I679097,I679180,I679494);
or I_39811 (I679525,I679446,I679415);
DFFARX1 I_39812  ( .D(I679525), .CLK(I2702), .RSTB(I679129), .Q(I679094) );
not I_39813 (I679100,I679446);
DFFARX1 I_39814  ( .D(I279444), .CLK(I2702), .RSTB(I679129), .Q(I679570) );
not I_39815 (I679587,I679570);
nor I_39816 (I679604,I679587,I679180);
DFFARX1 I_39817  ( .D(I679604), .CLK(I2702), .RSTB(I679129), .Q(I679106) );
nor I_39818 (I679121,I679446,I679587);
nor I_39819 (I679109,I679587,I679350);
not I_39820 (I679663,I679587);
and I_39821 (I679680,I679214,I679663);
nor I_39822 (I679115,I679350,I679680);
nand I_39823 (I679103,I679587,I679477);
not I_39824 (I679758,I2709);
not I_39825 (I679775,I115649);
nor I_39826 (I679792,I115667,I115646);
nand I_39827 (I679809,I679792,I115664);
nor I_39828 (I679826,I679775,I115667);
nand I_39829 (I679843,I679826,I115658);
not I_39830 (I679860,I115667);
not I_39831 (I679877,I679860);
not I_39832 (I679894,I115661);
nor I_39833 (I679911,I679894,I115655);
and I_39834 (I679928,I679911,I115652);
or I_39835 (I679945,I679928,I115643);
DFFARX1 I_39836  ( .D(I679945), .CLK(I2702), .RSTB(I679758), .Q(I679962) );
nand I_39837 (I679979,I679775,I115661);
or I_39838 (I679747,I679979,I679962);
not I_39839 (I680010,I679979);
nor I_39840 (I680027,I679962,I680010);
and I_39841 (I680044,I679860,I680027);
nand I_39842 (I679720,I679979,I679877);
DFFARX1 I_39843  ( .D(I115673), .CLK(I2702), .RSTB(I679758), .Q(I680075) );
or I_39844 (I679741,I680075,I679962);
nor I_39845 (I680106,I680075,I679843);
nor I_39846 (I680123,I680075,I679877);
nand I_39847 (I679726,I679809,I680123);
or I_39848 (I680154,I680075,I680044);
DFFARX1 I_39849  ( .D(I680154), .CLK(I2702), .RSTB(I679758), .Q(I679723) );
not I_39850 (I679729,I680075);
DFFARX1 I_39851  ( .D(I115670), .CLK(I2702), .RSTB(I679758), .Q(I680199) );
not I_39852 (I680216,I680199);
nor I_39853 (I680233,I680216,I679809);
DFFARX1 I_39854  ( .D(I680233), .CLK(I2702), .RSTB(I679758), .Q(I679735) );
nor I_39855 (I679750,I680075,I680216);
nor I_39856 (I679738,I680216,I679979);
not I_39857 (I680292,I680216);
and I_39858 (I680309,I679843,I680292);
nor I_39859 (I679744,I679979,I680309);
nand I_39860 (I679732,I680216,I680106);
not I_39861 (I680387,I2709);
not I_39862 (I680404,I514350);
nor I_39863 (I680421,I514368,I514347);
nand I_39864 (I680438,I680421,I514371);
nor I_39865 (I680455,I680404,I514368);
nand I_39866 (I680472,I680455,I514365);
not I_39867 (I680489,I514368);
not I_39868 (I680506,I680489);
not I_39869 (I680523,I514356);
nor I_39870 (I680540,I680523,I514344);
and I_39871 (I680557,I680540,I514362);
or I_39872 (I680574,I680557,I514374);
DFFARX1 I_39873  ( .D(I680574), .CLK(I2702), .RSTB(I680387), .Q(I680591) );
nand I_39874 (I680608,I680404,I514356);
or I_39875 (I680376,I680608,I680591);
not I_39876 (I680639,I680608);
nor I_39877 (I680656,I680591,I680639);
and I_39878 (I680673,I680489,I680656);
nand I_39879 (I680349,I680608,I680506);
DFFARX1 I_39880  ( .D(I514353), .CLK(I2702), .RSTB(I680387), .Q(I680704) );
or I_39881 (I680370,I680704,I680591);
nor I_39882 (I680735,I680704,I680472);
nor I_39883 (I680752,I680704,I680506);
nand I_39884 (I680355,I680438,I680752);
or I_39885 (I680783,I680704,I680673);
DFFARX1 I_39886  ( .D(I680783), .CLK(I2702), .RSTB(I680387), .Q(I680352) );
not I_39887 (I680358,I680704);
DFFARX1 I_39888  ( .D(I514359), .CLK(I2702), .RSTB(I680387), .Q(I680828) );
not I_39889 (I680845,I680828);
nor I_39890 (I680862,I680845,I680438);
DFFARX1 I_39891  ( .D(I680862), .CLK(I2702), .RSTB(I680387), .Q(I680364) );
nor I_39892 (I680379,I680704,I680845);
nor I_39893 (I680367,I680845,I680608);
not I_39894 (I680921,I680845);
and I_39895 (I680938,I680472,I680921);
nor I_39896 (I680373,I680608,I680938);
nand I_39897 (I680361,I680845,I680735);
not I_39898 (I681016,I2709);
not I_39899 (I681033,I147513);
nor I_39900 (I681050,I147504,I147528);
nand I_39901 (I681067,I681050,I147531);
nor I_39902 (I681084,I681033,I147504);
nand I_39903 (I681101,I681084,I147522);
not I_39904 (I681118,I147504);
not I_39905 (I681135,I681118);
not I_39906 (I681152,I147516);
nor I_39907 (I681169,I681152,I147510);
and I_39908 (I681186,I681169,I147519);
or I_39909 (I681203,I681186,I147507);
DFFARX1 I_39910  ( .D(I681203), .CLK(I2702), .RSTB(I681016), .Q(I681220) );
nand I_39911 (I681237,I681033,I147516);
or I_39912 (I681005,I681237,I681220);
not I_39913 (I681268,I681237);
nor I_39914 (I681285,I681220,I681268);
and I_39915 (I681302,I681118,I681285);
nand I_39916 (I680978,I681237,I681135);
DFFARX1 I_39917  ( .D(I147501), .CLK(I2702), .RSTB(I681016), .Q(I681333) );
or I_39918 (I680999,I681333,I681220);
nor I_39919 (I681364,I681333,I681101);
nor I_39920 (I681381,I681333,I681135);
nand I_39921 (I680984,I681067,I681381);
or I_39922 (I681412,I681333,I681302);
DFFARX1 I_39923  ( .D(I681412), .CLK(I2702), .RSTB(I681016), .Q(I680981) );
not I_39924 (I680987,I681333);
DFFARX1 I_39925  ( .D(I147525), .CLK(I2702), .RSTB(I681016), .Q(I681457) );
not I_39926 (I681474,I681457);
nor I_39927 (I681491,I681474,I681067);
DFFARX1 I_39928  ( .D(I681491), .CLK(I2702), .RSTB(I681016), .Q(I680993) );
nor I_39929 (I681008,I681333,I681474);
nor I_39930 (I680996,I681474,I681237);
not I_39931 (I681550,I681474);
and I_39932 (I681567,I681101,I681550);
nor I_39933 (I681002,I681237,I681567);
nand I_39934 (I680990,I681474,I681364);
not I_39935 (I681645,I2709);
not I_39936 (I681662,I501391);
nor I_39937 (I681679,I501376,I501397);
nand I_39938 (I681696,I681679,I501385);
nor I_39939 (I681713,I681662,I501376);
nand I_39940 (I681730,I681713,I501373);
not I_39941 (I681747,I501376);
not I_39942 (I681764,I681747);
not I_39943 (I681781,I501400);
nor I_39944 (I681798,I681781,I501388);
and I_39945 (I681815,I681798,I501382);
or I_39946 (I681832,I681815,I501379);
DFFARX1 I_39947  ( .D(I681832), .CLK(I2702), .RSTB(I681645), .Q(I681849) );
nand I_39948 (I681866,I681662,I501400);
or I_39949 (I681634,I681866,I681849);
not I_39950 (I681897,I681866);
nor I_39951 (I681914,I681849,I681897);
and I_39952 (I681931,I681747,I681914);
nand I_39953 (I681607,I681866,I681764);
DFFARX1 I_39954  ( .D(I501403), .CLK(I2702), .RSTB(I681645), .Q(I681962) );
or I_39955 (I681628,I681962,I681849);
nor I_39956 (I681993,I681962,I681730);
nor I_39957 (I682010,I681962,I681764);
nand I_39958 (I681613,I681696,I682010);
or I_39959 (I682041,I681962,I681931);
DFFARX1 I_39960  ( .D(I682041), .CLK(I2702), .RSTB(I681645), .Q(I681610) );
not I_39961 (I681616,I681962);
DFFARX1 I_39962  ( .D(I501394), .CLK(I2702), .RSTB(I681645), .Q(I682086) );
not I_39963 (I682103,I682086);
nor I_39964 (I682120,I682103,I681696);
DFFARX1 I_39965  ( .D(I682120), .CLK(I2702), .RSTB(I681645), .Q(I681622) );
nor I_39966 (I681637,I681962,I682103);
nor I_39967 (I681625,I682103,I681866);
not I_39968 (I682179,I682103);
and I_39969 (I682196,I681730,I682179);
nor I_39970 (I681631,I681866,I682196);
nand I_39971 (I681619,I682103,I681993);
not I_39972 (I682274,I2709);
not I_39973 (I682291,I141546);
nor I_39974 (I682308,I141537,I141561);
nand I_39975 (I682325,I682308,I141564);
nor I_39976 (I682342,I682291,I141537);
nand I_39977 (I682359,I682342,I141555);
not I_39978 (I682376,I141537);
not I_39979 (I682393,I682376);
not I_39980 (I682410,I141549);
nor I_39981 (I682427,I682410,I141543);
and I_39982 (I682444,I682427,I141552);
or I_39983 (I682461,I682444,I141540);
DFFARX1 I_39984  ( .D(I682461), .CLK(I2702), .RSTB(I682274), .Q(I682478) );
nand I_39985 (I682495,I682291,I141549);
or I_39986 (I682263,I682495,I682478);
not I_39987 (I682526,I682495);
nor I_39988 (I682543,I682478,I682526);
and I_39989 (I682560,I682376,I682543);
nand I_39990 (I682236,I682495,I682393);
DFFARX1 I_39991  ( .D(I141534), .CLK(I2702), .RSTB(I682274), .Q(I682591) );
or I_39992 (I682257,I682591,I682478);
nor I_39993 (I682622,I682591,I682359);
nor I_39994 (I682639,I682591,I682393);
nand I_39995 (I682242,I682325,I682639);
or I_39996 (I682670,I682591,I682560);
DFFARX1 I_39997  ( .D(I682670), .CLK(I2702), .RSTB(I682274), .Q(I682239) );
not I_39998 (I682245,I682591);
DFFARX1 I_39999  ( .D(I141558), .CLK(I2702), .RSTB(I682274), .Q(I682715) );
not I_40000 (I682732,I682715);
nor I_40001 (I682749,I682732,I682325);
DFFARX1 I_40002  ( .D(I682749), .CLK(I2702), .RSTB(I682274), .Q(I682251) );
nor I_40003 (I682266,I682591,I682732);
nor I_40004 (I682254,I682732,I682495);
not I_40005 (I682808,I682732);
and I_40006 (I682825,I682359,I682808);
nor I_40007 (I682260,I682495,I682825);
nand I_40008 (I682248,I682732,I682622);
not I_40009 (I682903,I2709);
not I_40010 (I682920,I564925);
nor I_40011 (I682937,I564943,I564922);
nand I_40012 (I682954,I682937,I564946);
nor I_40013 (I682971,I682920,I564943);
nand I_40014 (I682988,I682971,I564940);
not I_40015 (I683005,I564943);
not I_40016 (I683022,I683005);
not I_40017 (I683039,I564931);
nor I_40018 (I683056,I683039,I564919);
and I_40019 (I683073,I683056,I564937);
or I_40020 (I683090,I683073,I564949);
DFFARX1 I_40021  ( .D(I683090), .CLK(I2702), .RSTB(I682903), .Q(I683107) );
nand I_40022 (I683124,I682920,I564931);
or I_40023 (I682892,I683124,I683107);
not I_40024 (I683155,I683124);
nor I_40025 (I683172,I683107,I683155);
and I_40026 (I683189,I683005,I683172);
nand I_40027 (I682865,I683124,I683022);
DFFARX1 I_40028  ( .D(I564928), .CLK(I2702), .RSTB(I682903), .Q(I683220) );
or I_40029 (I682886,I683220,I683107);
nor I_40030 (I683251,I683220,I682988);
nor I_40031 (I683268,I683220,I683022);
nand I_40032 (I682871,I682954,I683268);
or I_40033 (I683299,I683220,I683189);
DFFARX1 I_40034  ( .D(I683299), .CLK(I2702), .RSTB(I682903), .Q(I682868) );
not I_40035 (I682874,I683220);
DFFARX1 I_40036  ( .D(I564934), .CLK(I2702), .RSTB(I682903), .Q(I683344) );
not I_40037 (I683361,I683344);
nor I_40038 (I683378,I683361,I682954);
DFFARX1 I_40039  ( .D(I683378), .CLK(I2702), .RSTB(I682903), .Q(I682880) );
nor I_40040 (I682895,I683220,I683361);
nor I_40041 (I682883,I683361,I683124);
not I_40042 (I683437,I683361);
and I_40043 (I683454,I682988,I683437);
nor I_40044 (I682889,I683124,I683454);
nand I_40045 (I682877,I683361,I683251);
not I_40046 (I683532,I2709);
not I_40047 (I683549,I608363);
nor I_40048 (I683566,I608366,I608375);
nand I_40049 (I683583,I683566,I608360);
nor I_40050 (I683600,I683549,I608366);
nand I_40051 (I683617,I683600,I608369);
not I_40052 (I683634,I608366);
not I_40053 (I683651,I683634);
not I_40054 (I683668,I608384);
nor I_40055 (I683685,I683668,I608372);
and I_40056 (I683702,I683685,I608357);
or I_40057 (I683719,I683702,I608354);
DFFARX1 I_40058  ( .D(I683719), .CLK(I2702), .RSTB(I683532), .Q(I683736) );
nand I_40059 (I683753,I683549,I608384);
or I_40060 (I683521,I683753,I683736);
not I_40061 (I683784,I683753);
nor I_40062 (I683801,I683736,I683784);
and I_40063 (I683818,I683634,I683801);
nand I_40064 (I683494,I683753,I683651);
DFFARX1 I_40065  ( .D(I608378), .CLK(I2702), .RSTB(I683532), .Q(I683849) );
or I_40066 (I683515,I683849,I683736);
nor I_40067 (I683880,I683849,I683617);
nor I_40068 (I683897,I683849,I683651);
nand I_40069 (I683500,I683583,I683897);
or I_40070 (I683928,I683849,I683818);
DFFARX1 I_40071  ( .D(I683928), .CLK(I2702), .RSTB(I683532), .Q(I683497) );
not I_40072 (I683503,I683849);
DFFARX1 I_40073  ( .D(I608381), .CLK(I2702), .RSTB(I683532), .Q(I683973) );
not I_40074 (I683990,I683973);
nor I_40075 (I684007,I683990,I683583);
DFFARX1 I_40076  ( .D(I684007), .CLK(I2702), .RSTB(I683532), .Q(I683509) );
nor I_40077 (I683524,I683849,I683990);
nor I_40078 (I683512,I683990,I683753);
not I_40079 (I684066,I683990);
and I_40080 (I684083,I683617,I684066);
nor I_40081 (I683518,I683753,I684083);
nand I_40082 (I683506,I683990,I683880);
not I_40083 (I684161,I2709);
not I_40084 (I684178,I395821);
nor I_40085 (I684195,I395830,I395833);
nand I_40086 (I684212,I684195,I395818);
nor I_40087 (I684229,I684178,I395830);
nand I_40088 (I684246,I684229,I395815);
not I_40089 (I684263,I395830);
not I_40090 (I684280,I684263);
not I_40091 (I684297,I395803);
nor I_40092 (I684314,I684297,I395809);
and I_40093 (I684331,I684314,I395806);
or I_40094 (I684348,I684331,I395827);
DFFARX1 I_40095  ( .D(I684348), .CLK(I2702), .RSTB(I684161), .Q(I684365) );
nand I_40096 (I684382,I684178,I395803);
or I_40097 (I684150,I684382,I684365);
not I_40098 (I684413,I684382);
nor I_40099 (I684430,I684365,I684413);
and I_40100 (I684447,I684263,I684430);
nand I_40101 (I684123,I684382,I684280);
DFFARX1 I_40102  ( .D(I395812), .CLK(I2702), .RSTB(I684161), .Q(I684478) );
or I_40103 (I684144,I684478,I684365);
nor I_40104 (I684509,I684478,I684246);
nor I_40105 (I684526,I684478,I684280);
nand I_40106 (I684129,I684212,I684526);
or I_40107 (I684557,I684478,I684447);
DFFARX1 I_40108  ( .D(I684557), .CLK(I2702), .RSTB(I684161), .Q(I684126) );
not I_40109 (I684132,I684478);
DFFARX1 I_40110  ( .D(I395824), .CLK(I2702), .RSTB(I684161), .Q(I684602) );
not I_40111 (I684619,I684602);
nor I_40112 (I684636,I684619,I684212);
DFFARX1 I_40113  ( .D(I684636), .CLK(I2702), .RSTB(I684161), .Q(I684138) );
nor I_40114 (I684153,I684478,I684619);
nor I_40115 (I684141,I684619,I684382);
not I_40116 (I684695,I684619);
and I_40117 (I684712,I684246,I684695);
nor I_40118 (I684147,I684382,I684712);
nand I_40119 (I684135,I684619,I684509);
not I_40120 (I684790,I2709);
not I_40121 (I684807,I268185);
nor I_40122 (I684824,I268191,I268170);
nand I_40123 (I684841,I684824,I268176);
nor I_40124 (I684858,I684807,I268191);
nand I_40125 (I684875,I684858,I268182);
not I_40126 (I684892,I268191);
not I_40127 (I684909,I684892);
not I_40128 (I684926,I268179);
nor I_40129 (I684943,I684926,I268197);
and I_40130 (I684960,I684943,I268188);
or I_40131 (I684977,I684960,I268167);
DFFARX1 I_40132  ( .D(I684977), .CLK(I2702), .RSTB(I684790), .Q(I684994) );
nand I_40133 (I685011,I684807,I268179);
or I_40134 (I684779,I685011,I684994);
not I_40135 (I685042,I685011);
nor I_40136 (I685059,I684994,I685042);
and I_40137 (I685076,I684892,I685059);
nand I_40138 (I684752,I685011,I684909);
DFFARX1 I_40139  ( .D(I268194), .CLK(I2702), .RSTB(I684790), .Q(I685107) );
or I_40140 (I684773,I685107,I684994);
nor I_40141 (I685138,I685107,I684875);
nor I_40142 (I685155,I685107,I684909);
nand I_40143 (I684758,I684841,I685155);
or I_40144 (I685186,I685107,I685076);
DFFARX1 I_40145  ( .D(I685186), .CLK(I2702), .RSTB(I684790), .Q(I684755) );
not I_40146 (I684761,I685107);
DFFARX1 I_40147  ( .D(I268173), .CLK(I2702), .RSTB(I684790), .Q(I685231) );
not I_40148 (I685248,I685231);
nor I_40149 (I685265,I685248,I684841);
DFFARX1 I_40150  ( .D(I685265), .CLK(I2702), .RSTB(I684790), .Q(I684767) );
nor I_40151 (I684782,I685107,I685248);
nor I_40152 (I684770,I685248,I685011);
not I_40153 (I685324,I685248);
and I_40154 (I685341,I684875,I685324);
nor I_40155 (I684776,I685011,I685341);
nand I_40156 (I684764,I685248,I685138);
not I_40157 (I685419,I2709);
not I_40158 (I685436,I207643);
nor I_40159 (I685453,I207619,I207634);
nand I_40160 (I685470,I685453,I207616);
nor I_40161 (I685487,I685436,I207619);
nand I_40162 (I685504,I685487,I207631);
not I_40163 (I685521,I207619);
not I_40164 (I685538,I685521);
not I_40165 (I685555,I207622);
nor I_40166 (I685572,I685555,I207637);
and I_40167 (I685589,I685572,I207628);
or I_40168 (I685606,I685589,I207613);
DFFARX1 I_40169  ( .D(I685606), .CLK(I2702), .RSTB(I685419), .Q(I685623) );
nand I_40170 (I685640,I685436,I207622);
or I_40171 (I685408,I685640,I685623);
not I_40172 (I685671,I685640);
nor I_40173 (I685688,I685623,I685671);
and I_40174 (I685705,I685521,I685688);
nand I_40175 (I685381,I685640,I685538);
DFFARX1 I_40176  ( .D(I207625), .CLK(I2702), .RSTB(I685419), .Q(I685736) );
or I_40177 (I685402,I685736,I685623);
nor I_40178 (I685767,I685736,I685504);
nor I_40179 (I685784,I685736,I685538);
nand I_40180 (I685387,I685470,I685784);
or I_40181 (I685815,I685736,I685705);
DFFARX1 I_40182  ( .D(I685815), .CLK(I2702), .RSTB(I685419), .Q(I685384) );
not I_40183 (I685390,I685736);
DFFARX1 I_40184  ( .D(I207640), .CLK(I2702), .RSTB(I685419), .Q(I685860) );
not I_40185 (I685877,I685860);
nor I_40186 (I685894,I685877,I685470);
DFFARX1 I_40187  ( .D(I685894), .CLK(I2702), .RSTB(I685419), .Q(I685396) );
nor I_40188 (I685411,I685736,I685877);
nor I_40189 (I685399,I685877,I685640);
not I_40190 (I685953,I685877);
and I_40191 (I685970,I685504,I685953);
nor I_40192 (I685405,I685640,I685970);
nand I_40193 (I685393,I685877,I685767);
not I_40194 (I686048,I2709);
not I_40195 (I686065,I268848);
nor I_40196 (I686082,I268854,I268833);
nand I_40197 (I686099,I686082,I268839);
nor I_40198 (I686116,I686065,I268854);
nand I_40199 (I686133,I686116,I268845);
not I_40200 (I686150,I268854);
not I_40201 (I686167,I686150);
not I_40202 (I686184,I268842);
nor I_40203 (I686201,I686184,I268860);
and I_40204 (I686218,I686201,I268851);
or I_40205 (I686235,I686218,I268830);
DFFARX1 I_40206  ( .D(I686235), .CLK(I2702), .RSTB(I686048), .Q(I686252) );
nand I_40207 (I686269,I686065,I268842);
or I_40208 (I686037,I686269,I686252);
not I_40209 (I686300,I686269);
nor I_40210 (I686317,I686252,I686300);
and I_40211 (I686334,I686150,I686317);
nand I_40212 (I686010,I686269,I686167);
DFFARX1 I_40213  ( .D(I268857), .CLK(I2702), .RSTB(I686048), .Q(I686365) );
or I_40214 (I686031,I686365,I686252);
nor I_40215 (I686396,I686365,I686133);
nor I_40216 (I686413,I686365,I686167);
nand I_40217 (I686016,I686099,I686413);
or I_40218 (I686444,I686365,I686334);
DFFARX1 I_40219  ( .D(I686444), .CLK(I2702), .RSTB(I686048), .Q(I686013) );
not I_40220 (I686019,I686365);
DFFARX1 I_40221  ( .D(I268836), .CLK(I2702), .RSTB(I686048), .Q(I686489) );
not I_40222 (I686506,I686489);
nor I_40223 (I686523,I686506,I686099);
DFFARX1 I_40224  ( .D(I686523), .CLK(I2702), .RSTB(I686048), .Q(I686025) );
nor I_40225 (I686040,I686365,I686506);
nor I_40226 (I686028,I686506,I686269);
not I_40227 (I686582,I686506);
and I_40228 (I686599,I686133,I686582);
nor I_40229 (I686034,I686269,I686599);
nand I_40230 (I686022,I686506,I686396);
not I_40231 (I686677,I2709);
not I_40232 (I686694,I579803);
nor I_40233 (I686711,I579806,I579815);
nand I_40234 (I686728,I686711,I579800);
nor I_40235 (I686745,I686694,I579806);
nand I_40236 (I686762,I686745,I579809);
not I_40237 (I686779,I579806);
not I_40238 (I686796,I686779);
not I_40239 (I686813,I579824);
nor I_40240 (I686830,I686813,I579812);
and I_40241 (I686847,I686830,I579797);
or I_40242 (I686864,I686847,I579794);
DFFARX1 I_40243  ( .D(I686864), .CLK(I2702), .RSTB(I686677), .Q(I686881) );
nand I_40244 (I686898,I686694,I579824);
or I_40245 (I686666,I686898,I686881);
not I_40246 (I686929,I686898);
nor I_40247 (I686946,I686881,I686929);
and I_40248 (I686963,I686779,I686946);
nand I_40249 (I686639,I686898,I686796);
DFFARX1 I_40250  ( .D(I579818), .CLK(I2702), .RSTB(I686677), .Q(I686994) );
or I_40251 (I686660,I686994,I686881);
nor I_40252 (I687025,I686994,I686762);
nor I_40253 (I687042,I686994,I686796);
nand I_40254 (I686645,I686728,I687042);
or I_40255 (I687073,I686994,I686963);
DFFARX1 I_40256  ( .D(I687073), .CLK(I2702), .RSTB(I686677), .Q(I686642) );
not I_40257 (I686648,I686994);
DFFARX1 I_40258  ( .D(I579821), .CLK(I2702), .RSTB(I686677), .Q(I687118) );
not I_40259 (I687135,I687118);
nor I_40260 (I687152,I687135,I686728);
DFFARX1 I_40261  ( .D(I687152), .CLK(I2702), .RSTB(I686677), .Q(I686654) );
nor I_40262 (I686669,I686994,I687135);
nor I_40263 (I686657,I687135,I686898);
not I_40264 (I687211,I687135);
and I_40265 (I687228,I686762,I687211);
nor I_40266 (I686663,I686898,I687228);
nand I_40267 (I686651,I687135,I687025);
not I_40268 (I687306,I2709);
not I_40269 (I687323,I134383);
nor I_40270 (I687340,I134401,I134380);
nand I_40271 (I687357,I687340,I134398);
nor I_40272 (I687374,I687323,I134401);
nand I_40273 (I687391,I687374,I134392);
not I_40274 (I687408,I134401);
not I_40275 (I687425,I687408);
not I_40276 (I687442,I134395);
nor I_40277 (I687459,I687442,I134389);
and I_40278 (I687476,I687459,I134386);
or I_40279 (I687493,I687476,I134377);
DFFARX1 I_40280  ( .D(I687493), .CLK(I2702), .RSTB(I687306), .Q(I687510) );
nand I_40281 (I687527,I687323,I134395);
or I_40282 (I687295,I687527,I687510);
not I_40283 (I687558,I687527);
nor I_40284 (I687575,I687510,I687558);
and I_40285 (I687592,I687408,I687575);
nand I_40286 (I687268,I687527,I687425);
DFFARX1 I_40287  ( .D(I134407), .CLK(I2702), .RSTB(I687306), .Q(I687623) );
or I_40288 (I687289,I687623,I687510);
nor I_40289 (I687654,I687623,I687391);
nor I_40290 (I687671,I687623,I687425);
nand I_40291 (I687274,I687357,I687671);
or I_40292 (I687702,I687623,I687592);
DFFARX1 I_40293  ( .D(I687702), .CLK(I2702), .RSTB(I687306), .Q(I687271) );
not I_40294 (I687277,I687623);
DFFARX1 I_40295  ( .D(I134404), .CLK(I2702), .RSTB(I687306), .Q(I687747) );
not I_40296 (I687764,I687747);
nor I_40297 (I687781,I687764,I687357);
DFFARX1 I_40298  ( .D(I687781), .CLK(I2702), .RSTB(I687306), .Q(I687283) );
nor I_40299 (I687298,I687623,I687764);
nor I_40300 (I687286,I687764,I687527);
not I_40301 (I687840,I687764);
and I_40302 (I687857,I687391,I687840);
nor I_40303 (I687292,I687527,I687857);
nand I_40304 (I687280,I687764,I687654);
not I_40305 (I687935,I2709);
not I_40306 (I687952,I545290);
nor I_40307 (I687969,I545308,I545287);
nand I_40308 (I687986,I687969,I545311);
nor I_40309 (I688003,I687952,I545308);
nand I_40310 (I688020,I688003,I545305);
not I_40311 (I688037,I545308);
not I_40312 (I688054,I688037);
not I_40313 (I688071,I545296);
nor I_40314 (I688088,I688071,I545284);
and I_40315 (I688105,I688088,I545302);
or I_40316 (I688122,I688105,I545314);
DFFARX1 I_40317  ( .D(I688122), .CLK(I2702), .RSTB(I687935), .Q(I688139) );
nand I_40318 (I688156,I687952,I545296);
or I_40319 (I687924,I688156,I688139);
not I_40320 (I688187,I688156);
nor I_40321 (I688204,I688139,I688187);
and I_40322 (I688221,I688037,I688204);
nand I_40323 (I687897,I688156,I688054);
DFFARX1 I_40324  ( .D(I545293), .CLK(I2702), .RSTB(I687935), .Q(I688252) );
or I_40325 (I687918,I688252,I688139);
nor I_40326 (I688283,I688252,I688020);
nor I_40327 (I688300,I688252,I688054);
nand I_40328 (I687903,I687986,I688300);
or I_40329 (I688331,I688252,I688221);
DFFARX1 I_40330  ( .D(I688331), .CLK(I2702), .RSTB(I687935), .Q(I687900) );
not I_40331 (I687906,I688252);
DFFARX1 I_40332  ( .D(I545299), .CLK(I2702), .RSTB(I687935), .Q(I688376) );
not I_40333 (I688393,I688376);
nor I_40334 (I688410,I688393,I687986);
DFFARX1 I_40335  ( .D(I688410), .CLK(I2702), .RSTB(I687935), .Q(I687912) );
nor I_40336 (I687927,I688252,I688393);
nor I_40337 (I687915,I688393,I688156);
not I_40338 (I688469,I688393);
and I_40339 (I688486,I688020,I688469);
nor I_40340 (I687921,I688156,I688486);
nand I_40341 (I687909,I688393,I688283);
not I_40342 (I688564,I2709);
not I_40343 (I688581,I500813);
nor I_40344 (I688598,I500798,I500819);
nand I_40345 (I688615,I688598,I500807);
nor I_40346 (I688632,I688581,I500798);
nand I_40347 (I688649,I688632,I500795);
not I_40348 (I688666,I500798);
not I_40349 (I688683,I688666);
not I_40350 (I688700,I500822);
nor I_40351 (I688717,I688700,I500810);
and I_40352 (I688734,I688717,I500804);
or I_40353 (I688751,I688734,I500801);
DFFARX1 I_40354  ( .D(I688751), .CLK(I2702), .RSTB(I688564), .Q(I688768) );
nand I_40355 (I688785,I688581,I500822);
or I_40356 (I688553,I688785,I688768);
not I_40357 (I688816,I688785);
nor I_40358 (I688833,I688768,I688816);
and I_40359 (I688850,I688666,I688833);
nand I_40360 (I688526,I688785,I688683);
DFFARX1 I_40361  ( .D(I500825), .CLK(I2702), .RSTB(I688564), .Q(I688881) );
or I_40362 (I688547,I688881,I688768);
nor I_40363 (I688912,I688881,I688649);
nor I_40364 (I688929,I688881,I688683);
nand I_40365 (I688532,I688615,I688929);
or I_40366 (I688960,I688881,I688850);
DFFARX1 I_40367  ( .D(I688960), .CLK(I2702), .RSTB(I688564), .Q(I688529) );
not I_40368 (I688535,I688881);
DFFARX1 I_40369  ( .D(I500816), .CLK(I2702), .RSTB(I688564), .Q(I689005) );
not I_40370 (I689022,I689005);
nor I_40371 (I689039,I689022,I688615);
DFFARX1 I_40372  ( .D(I689039), .CLK(I2702), .RSTB(I688564), .Q(I688541) );
nor I_40373 (I688556,I688881,I689022);
nor I_40374 (I688544,I689022,I688785);
not I_40375 (I689098,I689022);
and I_40376 (I689115,I688649,I689098);
nor I_40377 (I688550,I688785,I689115);
nand I_40378 (I688538,I689022,I688912);
not I_40379 (I689193,I2709);
not I_40380 (I689210,I214188);
nor I_40381 (I689227,I214164,I214179);
nand I_40382 (I689244,I689227,I214161);
nor I_40383 (I689261,I689210,I214164);
nand I_40384 (I689278,I689261,I214176);
not I_40385 (I689295,I214164);
not I_40386 (I689312,I689295);
not I_40387 (I689329,I214167);
nor I_40388 (I689346,I689329,I214182);
and I_40389 (I689363,I689346,I214173);
or I_40390 (I689380,I689363,I214158);
DFFARX1 I_40391  ( .D(I689380), .CLK(I2702), .RSTB(I689193), .Q(I689397) );
nand I_40392 (I689414,I689210,I214167);
or I_40393 (I689182,I689414,I689397);
not I_40394 (I689445,I689414);
nor I_40395 (I689462,I689397,I689445);
and I_40396 (I689479,I689295,I689462);
nand I_40397 (I689155,I689414,I689312);
DFFARX1 I_40398  ( .D(I214170), .CLK(I2702), .RSTB(I689193), .Q(I689510) );
or I_40399 (I689176,I689510,I689397);
nor I_40400 (I689541,I689510,I689278);
nor I_40401 (I689558,I689510,I689312);
nand I_40402 (I689161,I689244,I689558);
or I_40403 (I689589,I689510,I689479);
DFFARX1 I_40404  ( .D(I689589), .CLK(I2702), .RSTB(I689193), .Q(I689158) );
not I_40405 (I689164,I689510);
DFFARX1 I_40406  ( .D(I214185), .CLK(I2702), .RSTB(I689193), .Q(I689634) );
not I_40407 (I689651,I689634);
nor I_40408 (I689668,I689651,I689244);
DFFARX1 I_40409  ( .D(I689668), .CLK(I2702), .RSTB(I689193), .Q(I689170) );
nor I_40410 (I689185,I689510,I689651);
nor I_40411 (I689173,I689651,I689414);
not I_40412 (I689727,I689651);
and I_40413 (I689744,I689278,I689727);
nor I_40414 (I689179,I689414,I689744);
nand I_40415 (I689167,I689651,I689541);
not I_40416 (I689822,I2709);
nand I_40417 (I689839,I126646,I126631);
and I_40418 (I689856,I689839,I126625);
DFFARX1 I_40419  ( .D(I689856), .CLK(I2702), .RSTB(I689822), .Q(I689873) );
not I_40420 (I689811,I689873);
DFFARX1 I_40421  ( .D(I689873), .CLK(I2702), .RSTB(I689822), .Q(I689904) );
not I_40422 (I689799,I689904);
nor I_40423 (I689935,I126652,I126631);
not I_40424 (I689952,I689935);
nor I_40425 (I689969,I689873,I689952);
DFFARX1 I_40426  ( .D(I126655), .CLK(I2702), .RSTB(I689822), .Q(I689986) );
not I_40427 (I690003,I689986);
nand I_40428 (I689802,I689986,I689952);
DFFARX1 I_40429  ( .D(I689986), .CLK(I2702), .RSTB(I689822), .Q(I690034) );
and I_40430 (I689787,I689873,I690034);
nand I_40431 (I690065,I126637,I126640);
and I_40432 (I690082,I690065,I126643);
DFFARX1 I_40433  ( .D(I690082), .CLK(I2702), .RSTB(I689822), .Q(I690099) );
nor I_40434 (I690116,I690099,I690003);
and I_40435 (I690133,I689935,I690116);
nor I_40436 (I690150,I690099,I689873);
DFFARX1 I_40437  ( .D(I690099), .CLK(I2702), .RSTB(I689822), .Q(I689793) );
DFFARX1 I_40438  ( .D(I126649), .CLK(I2702), .RSTB(I689822), .Q(I690181) );
and I_40439 (I690198,I690181,I126634);
or I_40440 (I690215,I690198,I690133);
DFFARX1 I_40441  ( .D(I690215), .CLK(I2702), .RSTB(I689822), .Q(I689805) );
nand I_40442 (I689814,I690198,I690150);
DFFARX1 I_40443  ( .D(I690198), .CLK(I2702), .RSTB(I689822), .Q(I689784) );
DFFARX1 I_40444  ( .D(I126628), .CLK(I2702), .RSTB(I689822), .Q(I690274) );
nand I_40445 (I689808,I690274,I689969);
DFFARX1 I_40446  ( .D(I690274), .CLK(I2702), .RSTB(I689822), .Q(I689796) );
nand I_40447 (I690319,I690274,I689935);
and I_40448 (I690336,I689986,I690319);
DFFARX1 I_40449  ( .D(I690336), .CLK(I2702), .RSTB(I689822), .Q(I689790) );
not I_40450 (I690400,I2709);
nand I_40451 (I690417,I535190,I535172);
and I_40452 (I690434,I690417,I535187);
DFFARX1 I_40453  ( .D(I690434), .CLK(I2702), .RSTB(I690400), .Q(I690451) );
not I_40454 (I690389,I690451);
DFFARX1 I_40455  ( .D(I690451), .CLK(I2702), .RSTB(I690400), .Q(I690482) );
not I_40456 (I690377,I690482);
nor I_40457 (I690513,I535178,I535172);
not I_40458 (I690530,I690513);
nor I_40459 (I690547,I690451,I690530);
DFFARX1 I_40460  ( .D(I535193), .CLK(I2702), .RSTB(I690400), .Q(I690564) );
not I_40461 (I690581,I690564);
nand I_40462 (I690380,I690564,I690530);
DFFARX1 I_40463  ( .D(I690564), .CLK(I2702), .RSTB(I690400), .Q(I690612) );
and I_40464 (I690365,I690451,I690612);
nand I_40465 (I690643,I535169,I535175);
and I_40466 (I690660,I690643,I535181);
DFFARX1 I_40467  ( .D(I690660), .CLK(I2702), .RSTB(I690400), .Q(I690677) );
nor I_40468 (I690694,I690677,I690581);
and I_40469 (I690711,I690513,I690694);
nor I_40470 (I690728,I690677,I690451);
DFFARX1 I_40471  ( .D(I690677), .CLK(I2702), .RSTB(I690400), .Q(I690371) );
DFFARX1 I_40472  ( .D(I535196), .CLK(I2702), .RSTB(I690400), .Q(I690759) );
and I_40473 (I690776,I690759,I535184);
or I_40474 (I690793,I690776,I690711);
DFFARX1 I_40475  ( .D(I690793), .CLK(I2702), .RSTB(I690400), .Q(I690383) );
nand I_40476 (I690392,I690776,I690728);
DFFARX1 I_40477  ( .D(I690776), .CLK(I2702), .RSTB(I690400), .Q(I690362) );
DFFARX1 I_40478  ( .D(I535199), .CLK(I2702), .RSTB(I690400), .Q(I690852) );
nand I_40479 (I690386,I690852,I690547);
DFFARX1 I_40480  ( .D(I690852), .CLK(I2702), .RSTB(I690400), .Q(I690374) );
nand I_40481 (I690897,I690852,I690513);
and I_40482 (I690914,I690564,I690897);
DFFARX1 I_40483  ( .D(I690914), .CLK(I2702), .RSTB(I690400), .Q(I690368) );
not I_40484 (I690978,I2709);
nand I_40485 (I690995,I687271,I687289);
and I_40486 (I691012,I690995,I687286);
DFFARX1 I_40487  ( .D(I691012), .CLK(I2702), .RSTB(I690978), .Q(I691029) );
not I_40488 (I690967,I691029);
DFFARX1 I_40489  ( .D(I691029), .CLK(I2702), .RSTB(I690978), .Q(I691060) );
not I_40490 (I690955,I691060);
nor I_40491 (I691091,I687292,I687289);
not I_40492 (I691108,I691091);
nor I_40493 (I691125,I691029,I691108);
DFFARX1 I_40494  ( .D(I687295), .CLK(I2702), .RSTB(I690978), .Q(I691142) );
not I_40495 (I691159,I691142);
nand I_40496 (I690958,I691142,I691108);
DFFARX1 I_40497  ( .D(I691142), .CLK(I2702), .RSTB(I690978), .Q(I691190) );
and I_40498 (I690943,I691029,I691190);
nand I_40499 (I691221,I687280,I687274);
and I_40500 (I691238,I691221,I687277);
DFFARX1 I_40501  ( .D(I691238), .CLK(I2702), .RSTB(I690978), .Q(I691255) );
nor I_40502 (I691272,I691255,I691159);
and I_40503 (I691289,I691091,I691272);
nor I_40504 (I691306,I691255,I691029);
DFFARX1 I_40505  ( .D(I691255), .CLK(I2702), .RSTB(I690978), .Q(I690949) );
DFFARX1 I_40506  ( .D(I687283), .CLK(I2702), .RSTB(I690978), .Q(I691337) );
and I_40507 (I691354,I691337,I687268);
or I_40508 (I691371,I691354,I691289);
DFFARX1 I_40509  ( .D(I691371), .CLK(I2702), .RSTB(I690978), .Q(I690961) );
nand I_40510 (I690970,I691354,I691306);
DFFARX1 I_40511  ( .D(I691354), .CLK(I2702), .RSTB(I690978), .Q(I690940) );
DFFARX1 I_40512  ( .D(I687298), .CLK(I2702), .RSTB(I690978), .Q(I691430) );
nand I_40513 (I690964,I691430,I691125);
DFFARX1 I_40514  ( .D(I691430), .CLK(I2702), .RSTB(I690978), .Q(I690952) );
nand I_40515 (I691475,I691430,I691091);
and I_40516 (I691492,I691142,I691475);
DFFARX1 I_40517  ( .D(I691492), .CLK(I2702), .RSTB(I690978), .Q(I690946) );
not I_40518 (I691556,I2709);
nand I_40519 (I691573,I61400,I61385);
and I_40520 (I691590,I691573,I61379);
DFFARX1 I_40521  ( .D(I691590), .CLK(I2702), .RSTB(I691556), .Q(I691607) );
not I_40522 (I691545,I691607);
DFFARX1 I_40523  ( .D(I691607), .CLK(I2702), .RSTB(I691556), .Q(I691638) );
not I_40524 (I691533,I691638);
nor I_40525 (I691669,I61406,I61385);
not I_40526 (I691686,I691669);
nor I_40527 (I691703,I691607,I691686);
DFFARX1 I_40528  ( .D(I61409), .CLK(I2702), .RSTB(I691556), .Q(I691720) );
not I_40529 (I691737,I691720);
nand I_40530 (I691536,I691720,I691686);
DFFARX1 I_40531  ( .D(I691720), .CLK(I2702), .RSTB(I691556), .Q(I691768) );
and I_40532 (I691521,I691607,I691768);
nand I_40533 (I691799,I61391,I61394);
and I_40534 (I691816,I691799,I61397);
DFFARX1 I_40535  ( .D(I691816), .CLK(I2702), .RSTB(I691556), .Q(I691833) );
nor I_40536 (I691850,I691833,I691737);
and I_40537 (I691867,I691669,I691850);
nor I_40538 (I691884,I691833,I691607);
DFFARX1 I_40539  ( .D(I691833), .CLK(I2702), .RSTB(I691556), .Q(I691527) );
DFFARX1 I_40540  ( .D(I61403), .CLK(I2702), .RSTB(I691556), .Q(I691915) );
and I_40541 (I691932,I691915,I61388);
or I_40542 (I691949,I691932,I691867);
DFFARX1 I_40543  ( .D(I691949), .CLK(I2702), .RSTB(I691556), .Q(I691539) );
nand I_40544 (I691548,I691932,I691884);
DFFARX1 I_40545  ( .D(I691932), .CLK(I2702), .RSTB(I691556), .Q(I691518) );
DFFARX1 I_40546  ( .D(I61382), .CLK(I2702), .RSTB(I691556), .Q(I692008) );
nand I_40547 (I691542,I692008,I691703);
DFFARX1 I_40548  ( .D(I692008), .CLK(I2702), .RSTB(I691556), .Q(I691530) );
nand I_40549 (I692053,I692008,I691669);
and I_40550 (I692070,I691720,I692053);
DFFARX1 I_40551  ( .D(I692070), .CLK(I2702), .RSTB(I691556), .Q(I691524) );
not I_40552 (I692134,I2709);
nand I_40553 (I692151,I540545,I540527);
and I_40554 (I692168,I692151,I540542);
DFFARX1 I_40555  ( .D(I692168), .CLK(I2702), .RSTB(I692134), .Q(I692185) );
not I_40556 (I692123,I692185);
DFFARX1 I_40557  ( .D(I692185), .CLK(I2702), .RSTB(I692134), .Q(I692216) );
not I_40558 (I692111,I692216);
nor I_40559 (I692247,I540533,I540527);
not I_40560 (I692264,I692247);
nor I_40561 (I692281,I692185,I692264);
DFFARX1 I_40562  ( .D(I540548), .CLK(I2702), .RSTB(I692134), .Q(I692298) );
not I_40563 (I692315,I692298);
nand I_40564 (I692114,I692298,I692264);
DFFARX1 I_40565  ( .D(I692298), .CLK(I2702), .RSTB(I692134), .Q(I692346) );
and I_40566 (I692099,I692185,I692346);
nand I_40567 (I692377,I540524,I540530);
and I_40568 (I692394,I692377,I540536);
DFFARX1 I_40569  ( .D(I692394), .CLK(I2702), .RSTB(I692134), .Q(I692411) );
nor I_40570 (I692428,I692411,I692315);
and I_40571 (I692445,I692247,I692428);
nor I_40572 (I692462,I692411,I692185);
DFFARX1 I_40573  ( .D(I692411), .CLK(I2702), .RSTB(I692134), .Q(I692105) );
DFFARX1 I_40574  ( .D(I540551), .CLK(I2702), .RSTB(I692134), .Q(I692493) );
and I_40575 (I692510,I692493,I540539);
or I_40576 (I692527,I692510,I692445);
DFFARX1 I_40577  ( .D(I692527), .CLK(I2702), .RSTB(I692134), .Q(I692117) );
nand I_40578 (I692126,I692510,I692462);
DFFARX1 I_40579  ( .D(I692510), .CLK(I2702), .RSTB(I692134), .Q(I692096) );
DFFARX1 I_40580  ( .D(I540554), .CLK(I2702), .RSTB(I692134), .Q(I692586) );
nand I_40581 (I692120,I692586,I692281);
DFFARX1 I_40582  ( .D(I692586), .CLK(I2702), .RSTB(I692134), .Q(I692108) );
nand I_40583 (I692631,I692586,I692247);
and I_40584 (I692648,I692298,I692631);
DFFARX1 I_40585  ( .D(I692648), .CLK(I2702), .RSTB(I692134), .Q(I692102) );
not I_40586 (I692712,I2709);
nand I_40587 (I692729,I299337,I299334);
and I_40588 (I692746,I692729,I299358);
DFFARX1 I_40589  ( .D(I692746), .CLK(I2702), .RSTB(I692712), .Q(I692763) );
not I_40590 (I692701,I692763);
DFFARX1 I_40591  ( .D(I692763), .CLK(I2702), .RSTB(I692712), .Q(I692794) );
not I_40592 (I692689,I692794);
nor I_40593 (I692825,I299340,I299334);
not I_40594 (I692842,I692825);
nor I_40595 (I692859,I692763,I692842);
DFFARX1 I_40596  ( .D(I299355), .CLK(I2702), .RSTB(I692712), .Q(I692876) );
not I_40597 (I692893,I692876);
nand I_40598 (I692692,I692876,I692842);
DFFARX1 I_40599  ( .D(I692876), .CLK(I2702), .RSTB(I692712), .Q(I692924) );
and I_40600 (I692677,I692763,I692924);
nand I_40601 (I692955,I299343,I299328);
and I_40602 (I692972,I692955,I299346);
DFFARX1 I_40603  ( .D(I692972), .CLK(I2702), .RSTB(I692712), .Q(I692989) );
nor I_40604 (I693006,I692989,I692893);
and I_40605 (I693023,I692825,I693006);
nor I_40606 (I693040,I692989,I692763);
DFFARX1 I_40607  ( .D(I692989), .CLK(I2702), .RSTB(I692712), .Q(I692683) );
DFFARX1 I_40608  ( .D(I299349), .CLK(I2702), .RSTB(I692712), .Q(I693071) );
and I_40609 (I693088,I693071,I299352);
or I_40610 (I693105,I693088,I693023);
DFFARX1 I_40611  ( .D(I693105), .CLK(I2702), .RSTB(I692712), .Q(I692695) );
nand I_40612 (I692704,I693088,I693040);
DFFARX1 I_40613  ( .D(I693088), .CLK(I2702), .RSTB(I692712), .Q(I692674) );
DFFARX1 I_40614  ( .D(I299331), .CLK(I2702), .RSTB(I692712), .Q(I693164) );
nand I_40615 (I692698,I693164,I692859);
DFFARX1 I_40616  ( .D(I693164), .CLK(I2702), .RSTB(I692712), .Q(I692686) );
nand I_40617 (I693209,I693164,I692825);
and I_40618 (I693226,I692876,I693209);
DFFARX1 I_40619  ( .D(I693226), .CLK(I2702), .RSTB(I692712), .Q(I692680) );
not I_40620 (I693290,I2709);
nand I_40621 (I693307,I667772,I667790);
and I_40622 (I693324,I693307,I667787);
DFFARX1 I_40623  ( .D(I693324), .CLK(I2702), .RSTB(I693290), .Q(I693341) );
not I_40624 (I693279,I693341);
DFFARX1 I_40625  ( .D(I693341), .CLK(I2702), .RSTB(I693290), .Q(I693372) );
not I_40626 (I693267,I693372);
nor I_40627 (I693403,I667793,I667790);
not I_40628 (I693420,I693403);
nor I_40629 (I693437,I693341,I693420);
DFFARX1 I_40630  ( .D(I667796), .CLK(I2702), .RSTB(I693290), .Q(I693454) );
not I_40631 (I693471,I693454);
nand I_40632 (I693270,I693454,I693420);
DFFARX1 I_40633  ( .D(I693454), .CLK(I2702), .RSTB(I693290), .Q(I693502) );
and I_40634 (I693255,I693341,I693502);
nand I_40635 (I693533,I667781,I667775);
and I_40636 (I693550,I693533,I667778);
DFFARX1 I_40637  ( .D(I693550), .CLK(I2702), .RSTB(I693290), .Q(I693567) );
nor I_40638 (I693584,I693567,I693471);
and I_40639 (I693601,I693403,I693584);
nor I_40640 (I693618,I693567,I693341);
DFFARX1 I_40641  ( .D(I693567), .CLK(I2702), .RSTB(I693290), .Q(I693261) );
DFFARX1 I_40642  ( .D(I667784), .CLK(I2702), .RSTB(I693290), .Q(I693649) );
and I_40643 (I693666,I693649,I667769);
or I_40644 (I693683,I693666,I693601);
DFFARX1 I_40645  ( .D(I693683), .CLK(I2702), .RSTB(I693290), .Q(I693273) );
nand I_40646 (I693282,I693666,I693618);
DFFARX1 I_40647  ( .D(I693666), .CLK(I2702), .RSTB(I693290), .Q(I693252) );
DFFARX1 I_40648  ( .D(I667799), .CLK(I2702), .RSTB(I693290), .Q(I693742) );
nand I_40649 (I693276,I693742,I693437);
DFFARX1 I_40650  ( .D(I693742), .CLK(I2702), .RSTB(I693290), .Q(I693264) );
nand I_40651 (I693787,I693742,I693403);
and I_40652 (I693804,I693454,I693787);
DFFARX1 I_40653  ( .D(I693804), .CLK(I2702), .RSTB(I693290), .Q(I693258) );
not I_40654 (I693868,I2709);
nand I_40655 (I693885,I522695,I522677);
and I_40656 (I693902,I693885,I522692);
DFFARX1 I_40657  ( .D(I693902), .CLK(I2702), .RSTB(I693868), .Q(I693919) );
not I_40658 (I693857,I693919);
DFFARX1 I_40659  ( .D(I693919), .CLK(I2702), .RSTB(I693868), .Q(I693950) );
not I_40660 (I693845,I693950);
nor I_40661 (I693981,I522683,I522677);
not I_40662 (I693998,I693981);
nor I_40663 (I694015,I693919,I693998);
DFFARX1 I_40664  ( .D(I522698), .CLK(I2702), .RSTB(I693868), .Q(I694032) );
not I_40665 (I694049,I694032);
nand I_40666 (I693848,I694032,I693998);
DFFARX1 I_40667  ( .D(I694032), .CLK(I2702), .RSTB(I693868), .Q(I694080) );
and I_40668 (I693833,I693919,I694080);
nand I_40669 (I694111,I522674,I522680);
and I_40670 (I694128,I694111,I522686);
DFFARX1 I_40671  ( .D(I694128), .CLK(I2702), .RSTB(I693868), .Q(I694145) );
nor I_40672 (I694162,I694145,I694049);
and I_40673 (I694179,I693981,I694162);
nor I_40674 (I694196,I694145,I693919);
DFFARX1 I_40675  ( .D(I694145), .CLK(I2702), .RSTB(I693868), .Q(I693839) );
DFFARX1 I_40676  ( .D(I522701), .CLK(I2702), .RSTB(I693868), .Q(I694227) );
and I_40677 (I694244,I694227,I522689);
or I_40678 (I694261,I694244,I694179);
DFFARX1 I_40679  ( .D(I694261), .CLK(I2702), .RSTB(I693868), .Q(I693851) );
nand I_40680 (I693860,I694244,I694196);
DFFARX1 I_40681  ( .D(I694244), .CLK(I2702), .RSTB(I693868), .Q(I693830) );
DFFARX1 I_40682  ( .D(I522704), .CLK(I2702), .RSTB(I693868), .Q(I694320) );
nand I_40683 (I693854,I694320,I694015);
DFFARX1 I_40684  ( .D(I694320), .CLK(I2702), .RSTB(I693868), .Q(I693842) );
nand I_40685 (I694365,I694320,I693981);
and I_40686 (I694382,I694032,I694365);
DFFARX1 I_40687  ( .D(I694382), .CLK(I2702), .RSTB(I693868), .Q(I693836) );
not I_40688 (I694446,I2709);
nand I_40689 (I694463,I327846,I327843);
and I_40690 (I694480,I694463,I327867);
DFFARX1 I_40691  ( .D(I694480), .CLK(I2702), .RSTB(I694446), .Q(I694497) );
not I_40692 (I694435,I694497);
DFFARX1 I_40693  ( .D(I694497), .CLK(I2702), .RSTB(I694446), .Q(I694528) );
not I_40694 (I694423,I694528);
nor I_40695 (I694559,I327849,I327843);
not I_40696 (I694576,I694559);
nor I_40697 (I694593,I694497,I694576);
DFFARX1 I_40698  ( .D(I327864), .CLK(I2702), .RSTB(I694446), .Q(I694610) );
not I_40699 (I694627,I694610);
nand I_40700 (I694426,I694610,I694576);
DFFARX1 I_40701  ( .D(I694610), .CLK(I2702), .RSTB(I694446), .Q(I694658) );
and I_40702 (I694411,I694497,I694658);
nand I_40703 (I694689,I327852,I327837);
and I_40704 (I694706,I694689,I327855);
DFFARX1 I_40705  ( .D(I694706), .CLK(I2702), .RSTB(I694446), .Q(I694723) );
nor I_40706 (I694740,I694723,I694627);
and I_40707 (I694757,I694559,I694740);
nor I_40708 (I694774,I694723,I694497);
DFFARX1 I_40709  ( .D(I694723), .CLK(I2702), .RSTB(I694446), .Q(I694417) );
DFFARX1 I_40710  ( .D(I327858), .CLK(I2702), .RSTB(I694446), .Q(I694805) );
and I_40711 (I694822,I694805,I327861);
or I_40712 (I694839,I694822,I694757);
DFFARX1 I_40713  ( .D(I694839), .CLK(I2702), .RSTB(I694446), .Q(I694429) );
nand I_40714 (I694438,I694822,I694774);
DFFARX1 I_40715  ( .D(I694822), .CLK(I2702), .RSTB(I694446), .Q(I694408) );
DFFARX1 I_40716  ( .D(I327840), .CLK(I2702), .RSTB(I694446), .Q(I694898) );
nand I_40717 (I694432,I694898,I694593);
DFFARX1 I_40718  ( .D(I694898), .CLK(I2702), .RSTB(I694446), .Q(I694420) );
nand I_40719 (I694943,I694898,I694559);
and I_40720 (I694960,I694610,I694943);
DFFARX1 I_40721  ( .D(I694960), .CLK(I2702), .RSTB(I694446), .Q(I694414) );
not I_40722 (I695024,I2709);
nand I_40723 (I695041,I358999,I359002);
and I_40724 (I695058,I695041,I358981);
DFFARX1 I_40725  ( .D(I695058), .CLK(I2702), .RSTB(I695024), .Q(I695075) );
not I_40726 (I695013,I695075);
DFFARX1 I_40727  ( .D(I695075), .CLK(I2702), .RSTB(I695024), .Q(I695106) );
not I_40728 (I695001,I695106);
nor I_40729 (I695137,I358996,I359002);
not I_40730 (I695154,I695137);
nor I_40731 (I695171,I695075,I695154);
DFFARX1 I_40732  ( .D(I359005), .CLK(I2702), .RSTB(I695024), .Q(I695188) );
not I_40733 (I695205,I695188);
nand I_40734 (I695004,I695188,I695154);
DFFARX1 I_40735  ( .D(I695188), .CLK(I2702), .RSTB(I695024), .Q(I695236) );
and I_40736 (I694989,I695075,I695236);
nand I_40737 (I695267,I358993,I359011);
and I_40738 (I695284,I695267,I358987);
DFFARX1 I_40739  ( .D(I695284), .CLK(I2702), .RSTB(I695024), .Q(I695301) );
nor I_40740 (I695318,I695301,I695205);
and I_40741 (I695335,I695137,I695318);
nor I_40742 (I695352,I695301,I695075);
DFFARX1 I_40743  ( .D(I695301), .CLK(I2702), .RSTB(I695024), .Q(I694995) );
DFFARX1 I_40744  ( .D(I358984), .CLK(I2702), .RSTB(I695024), .Q(I695383) );
and I_40745 (I695400,I695383,I358990);
or I_40746 (I695417,I695400,I695335);
DFFARX1 I_40747  ( .D(I695417), .CLK(I2702), .RSTB(I695024), .Q(I695007) );
nand I_40748 (I695016,I695400,I695352);
DFFARX1 I_40749  ( .D(I695400), .CLK(I2702), .RSTB(I695024), .Q(I694986) );
DFFARX1 I_40750  ( .D(I359008), .CLK(I2702), .RSTB(I695024), .Q(I695476) );
nand I_40751 (I695010,I695476,I695171);
DFFARX1 I_40752  ( .D(I695476), .CLK(I2702), .RSTB(I695024), .Q(I694998) );
nand I_40753 (I695521,I695476,I695137);
and I_40754 (I695538,I695188,I695521);
DFFARX1 I_40755  ( .D(I695538), .CLK(I2702), .RSTB(I695024), .Q(I694992) );
not I_40756 (I695602,I2709);
nand I_40757 (I695619,I458128,I458146);
and I_40758 (I695636,I695619,I458137);
DFFARX1 I_40759  ( .D(I695636), .CLK(I2702), .RSTB(I695602), .Q(I695653) );
not I_40760 (I695591,I695653);
DFFARX1 I_40761  ( .D(I695653), .CLK(I2702), .RSTB(I695602), .Q(I695684) );
not I_40762 (I695579,I695684);
nor I_40763 (I695715,I458134,I458146);
not I_40764 (I695732,I695715);
nor I_40765 (I695749,I695653,I695732);
DFFARX1 I_40766  ( .D(I458125), .CLK(I2702), .RSTB(I695602), .Q(I695766) );
not I_40767 (I695783,I695766);
nand I_40768 (I695582,I695766,I695732);
DFFARX1 I_40769  ( .D(I695766), .CLK(I2702), .RSTB(I695602), .Q(I695814) );
and I_40770 (I695567,I695653,I695814);
nand I_40771 (I695845,I458143,I458155);
and I_40772 (I695862,I695845,I458149);
DFFARX1 I_40773  ( .D(I695862), .CLK(I2702), .RSTB(I695602), .Q(I695879) );
nor I_40774 (I695896,I695879,I695783);
and I_40775 (I695913,I695715,I695896);
nor I_40776 (I695930,I695879,I695653);
DFFARX1 I_40777  ( .D(I695879), .CLK(I2702), .RSTB(I695602), .Q(I695573) );
DFFARX1 I_40778  ( .D(I458131), .CLK(I2702), .RSTB(I695602), .Q(I695961) );
and I_40779 (I695978,I695961,I458140);
or I_40780 (I695995,I695978,I695913);
DFFARX1 I_40781  ( .D(I695995), .CLK(I2702), .RSTB(I695602), .Q(I695585) );
nand I_40782 (I695594,I695978,I695930);
DFFARX1 I_40783  ( .D(I695978), .CLK(I2702), .RSTB(I695602), .Q(I695564) );
DFFARX1 I_40784  ( .D(I458152), .CLK(I2702), .RSTB(I695602), .Q(I696054) );
nand I_40785 (I695588,I696054,I695749);
DFFARX1 I_40786  ( .D(I696054), .CLK(I2702), .RSTB(I695602), .Q(I695576) );
nand I_40787 (I696099,I696054,I695715);
and I_40788 (I696116,I695766,I696099);
DFFARX1 I_40789  ( .D(I696116), .CLK(I2702), .RSTB(I695602), .Q(I695570) );
not I_40790 (I696180,I2709);
nand I_40791 (I696197,I554825,I554807);
and I_40792 (I696214,I696197,I554822);
DFFARX1 I_40793  ( .D(I696214), .CLK(I2702), .RSTB(I696180), .Q(I696231) );
not I_40794 (I696169,I696231);
DFFARX1 I_40795  ( .D(I696231), .CLK(I2702), .RSTB(I696180), .Q(I696262) );
not I_40796 (I696157,I696262);
nor I_40797 (I696293,I554813,I554807);
not I_40798 (I696310,I696293);
nor I_40799 (I696327,I696231,I696310);
DFFARX1 I_40800  ( .D(I554828), .CLK(I2702), .RSTB(I696180), .Q(I696344) );
not I_40801 (I696361,I696344);
nand I_40802 (I696160,I696344,I696310);
DFFARX1 I_40803  ( .D(I696344), .CLK(I2702), .RSTB(I696180), .Q(I696392) );
and I_40804 (I696145,I696231,I696392);
nand I_40805 (I696423,I554804,I554810);
and I_40806 (I696440,I696423,I554816);
DFFARX1 I_40807  ( .D(I696440), .CLK(I2702), .RSTB(I696180), .Q(I696457) );
nor I_40808 (I696474,I696457,I696361);
and I_40809 (I696491,I696293,I696474);
nor I_40810 (I696508,I696457,I696231);
DFFARX1 I_40811  ( .D(I696457), .CLK(I2702), .RSTB(I696180), .Q(I696151) );
DFFARX1 I_40812  ( .D(I554831), .CLK(I2702), .RSTB(I696180), .Q(I696539) );
and I_40813 (I696556,I696539,I554819);
or I_40814 (I696573,I696556,I696491);
DFFARX1 I_40815  ( .D(I696573), .CLK(I2702), .RSTB(I696180), .Q(I696163) );
nand I_40816 (I696172,I696556,I696508);
DFFARX1 I_40817  ( .D(I696556), .CLK(I2702), .RSTB(I696180), .Q(I696142) );
DFFARX1 I_40818  ( .D(I554834), .CLK(I2702), .RSTB(I696180), .Q(I696632) );
nand I_40819 (I696166,I696632,I696327);
DFFARX1 I_40820  ( .D(I696632), .CLK(I2702), .RSTB(I696180), .Q(I696154) );
nand I_40821 (I696677,I696632,I696293);
and I_40822 (I696694,I696344,I696677);
DFFARX1 I_40823  ( .D(I696694), .CLK(I2702), .RSTB(I696180), .Q(I696148) );
not I_40824 (I696758,I2709);
nand I_40825 (I696775,I317901,I317898);
and I_40826 (I696792,I696775,I317922);
DFFARX1 I_40827  ( .D(I696792), .CLK(I2702), .RSTB(I696758), .Q(I696809) );
not I_40828 (I696747,I696809);
DFFARX1 I_40829  ( .D(I696809), .CLK(I2702), .RSTB(I696758), .Q(I696840) );
not I_40830 (I696735,I696840);
nor I_40831 (I696871,I317904,I317898);
not I_40832 (I696888,I696871);
nor I_40833 (I696905,I696809,I696888);
DFFARX1 I_40834  ( .D(I317919), .CLK(I2702), .RSTB(I696758), .Q(I696922) );
not I_40835 (I696939,I696922);
nand I_40836 (I696738,I696922,I696888);
DFFARX1 I_40837  ( .D(I696922), .CLK(I2702), .RSTB(I696758), .Q(I696970) );
and I_40838 (I696723,I696809,I696970);
nand I_40839 (I697001,I317907,I317892);
and I_40840 (I697018,I697001,I317910);
DFFARX1 I_40841  ( .D(I697018), .CLK(I2702), .RSTB(I696758), .Q(I697035) );
nor I_40842 (I697052,I697035,I696939);
and I_40843 (I697069,I696871,I697052);
nor I_40844 (I697086,I697035,I696809);
DFFARX1 I_40845  ( .D(I697035), .CLK(I2702), .RSTB(I696758), .Q(I696729) );
DFFARX1 I_40846  ( .D(I317913), .CLK(I2702), .RSTB(I696758), .Q(I697117) );
and I_40847 (I697134,I697117,I317916);
or I_40848 (I697151,I697134,I697069);
DFFARX1 I_40849  ( .D(I697151), .CLK(I2702), .RSTB(I696758), .Q(I696741) );
nand I_40850 (I696750,I697134,I697086);
DFFARX1 I_40851  ( .D(I697134), .CLK(I2702), .RSTB(I696758), .Q(I696720) );
DFFARX1 I_40852  ( .D(I317895), .CLK(I2702), .RSTB(I696758), .Q(I697210) );
nand I_40853 (I696744,I697210,I696905);
DFFARX1 I_40854  ( .D(I697210), .CLK(I2702), .RSTB(I696758), .Q(I696732) );
nand I_40855 (I697255,I697210,I696871);
and I_40856 (I697272,I696922,I697255);
DFFARX1 I_40857  ( .D(I697272), .CLK(I2702), .RSTB(I696758), .Q(I696726) );
not I_40858 (I697336,I2709);
nand I_40859 (I697353,I404219,I404222);
and I_40860 (I697370,I697353,I404201);
DFFARX1 I_40861  ( .D(I697370), .CLK(I2702), .RSTB(I697336), .Q(I697387) );
not I_40862 (I697325,I697387);
DFFARX1 I_40863  ( .D(I697387), .CLK(I2702), .RSTB(I697336), .Q(I697418) );
not I_40864 (I697313,I697418);
nor I_40865 (I697449,I404216,I404222);
not I_40866 (I697466,I697449);
nor I_40867 (I697483,I697387,I697466);
DFFARX1 I_40868  ( .D(I404225), .CLK(I2702), .RSTB(I697336), .Q(I697500) );
not I_40869 (I697517,I697500);
nand I_40870 (I697316,I697500,I697466);
DFFARX1 I_40871  ( .D(I697500), .CLK(I2702), .RSTB(I697336), .Q(I697548) );
and I_40872 (I697301,I697387,I697548);
nand I_40873 (I697579,I404213,I404231);
and I_40874 (I697596,I697579,I404207);
DFFARX1 I_40875  ( .D(I697596), .CLK(I2702), .RSTB(I697336), .Q(I697613) );
nor I_40876 (I697630,I697613,I697517);
and I_40877 (I697647,I697449,I697630);
nor I_40878 (I697664,I697613,I697387);
DFFARX1 I_40879  ( .D(I697613), .CLK(I2702), .RSTB(I697336), .Q(I697307) );
DFFARX1 I_40880  ( .D(I404204), .CLK(I2702), .RSTB(I697336), .Q(I697695) );
and I_40881 (I697712,I697695,I404210);
or I_40882 (I697729,I697712,I697647);
DFFARX1 I_40883  ( .D(I697729), .CLK(I2702), .RSTB(I697336), .Q(I697319) );
nand I_40884 (I697328,I697712,I697664);
DFFARX1 I_40885  ( .D(I697712), .CLK(I2702), .RSTB(I697336), .Q(I697298) );
DFFARX1 I_40886  ( .D(I404228), .CLK(I2702), .RSTB(I697336), .Q(I697788) );
nand I_40887 (I697322,I697788,I697483);
DFFARX1 I_40888  ( .D(I697788), .CLK(I2702), .RSTB(I697336), .Q(I697310) );
nand I_40889 (I697833,I697788,I697449);
and I_40890 (I697850,I697500,I697833);
DFFARX1 I_40891  ( .D(I697850), .CLK(I2702), .RSTB(I697336), .Q(I697304) );
not I_40892 (I697914,I2709);
nand I_40893 (I697931,I143523,I143553);
and I_40894 (I697948,I697931,I143535);
DFFARX1 I_40895  ( .D(I697948), .CLK(I2702), .RSTB(I697914), .Q(I697965) );
not I_40896 (I697903,I697965);
DFFARX1 I_40897  ( .D(I697965), .CLK(I2702), .RSTB(I697914), .Q(I697996) );
not I_40898 (I697891,I697996);
nor I_40899 (I698027,I143532,I143553);
not I_40900 (I698044,I698027);
nor I_40901 (I698061,I697965,I698044);
DFFARX1 I_40902  ( .D(I143526), .CLK(I2702), .RSTB(I697914), .Q(I698078) );
not I_40903 (I698095,I698078);
nand I_40904 (I697894,I698078,I698044);
DFFARX1 I_40905  ( .D(I698078), .CLK(I2702), .RSTB(I697914), .Q(I698126) );
and I_40906 (I697879,I697965,I698126);
nand I_40907 (I698157,I143529,I143544);
and I_40908 (I698174,I698157,I143541);
DFFARX1 I_40909  ( .D(I698174), .CLK(I2702), .RSTB(I697914), .Q(I698191) );
nor I_40910 (I698208,I698191,I698095);
and I_40911 (I698225,I698027,I698208);
nor I_40912 (I698242,I698191,I697965);
DFFARX1 I_40913  ( .D(I698191), .CLK(I2702), .RSTB(I697914), .Q(I697885) );
DFFARX1 I_40914  ( .D(I143538), .CLK(I2702), .RSTB(I697914), .Q(I698273) );
and I_40915 (I698290,I698273,I143550);
or I_40916 (I698307,I698290,I698225);
DFFARX1 I_40917  ( .D(I698307), .CLK(I2702), .RSTB(I697914), .Q(I697897) );
nand I_40918 (I697906,I698290,I698242);
DFFARX1 I_40919  ( .D(I698290), .CLK(I2702), .RSTB(I697914), .Q(I697876) );
DFFARX1 I_40920  ( .D(I143547), .CLK(I2702), .RSTB(I697914), .Q(I698366) );
nand I_40921 (I697900,I698366,I698061);
DFFARX1 I_40922  ( .D(I698366), .CLK(I2702), .RSTB(I697914), .Q(I697888) );
nand I_40923 (I698411,I698366,I698027);
and I_40924 (I698428,I698078,I698411);
DFFARX1 I_40925  ( .D(I698428), .CLK(I2702), .RSTB(I697914), .Q(I697882) );
not I_40926 (I698492,I2709);
nand I_40927 (I698509,I111142,I111127);
and I_40928 (I698526,I698509,I111121);
DFFARX1 I_40929  ( .D(I698526), .CLK(I2702), .RSTB(I698492), .Q(I698543) );
not I_40930 (I698481,I698543);
DFFARX1 I_40931  ( .D(I698543), .CLK(I2702), .RSTB(I698492), .Q(I698574) );
not I_40932 (I698469,I698574);
nor I_40933 (I698605,I111148,I111127);
not I_40934 (I698622,I698605);
nor I_40935 (I698639,I698543,I698622);
DFFARX1 I_40936  ( .D(I111151), .CLK(I2702), .RSTB(I698492), .Q(I698656) );
not I_40937 (I698673,I698656);
nand I_40938 (I698472,I698656,I698622);
DFFARX1 I_40939  ( .D(I698656), .CLK(I2702), .RSTB(I698492), .Q(I698704) );
and I_40940 (I698457,I698543,I698704);
nand I_40941 (I698735,I111133,I111136);
and I_40942 (I698752,I698735,I111139);
DFFARX1 I_40943  ( .D(I698752), .CLK(I2702), .RSTB(I698492), .Q(I698769) );
nor I_40944 (I698786,I698769,I698673);
and I_40945 (I698803,I698605,I698786);
nor I_40946 (I698820,I698769,I698543);
DFFARX1 I_40947  ( .D(I698769), .CLK(I2702), .RSTB(I698492), .Q(I698463) );
DFFARX1 I_40948  ( .D(I111145), .CLK(I2702), .RSTB(I698492), .Q(I698851) );
and I_40949 (I698868,I698851,I111130);
or I_40950 (I698885,I698868,I698803);
DFFARX1 I_40951  ( .D(I698885), .CLK(I2702), .RSTB(I698492), .Q(I698475) );
nand I_40952 (I698484,I698868,I698820);
DFFARX1 I_40953  ( .D(I698868), .CLK(I2702), .RSTB(I698492), .Q(I698454) );
DFFARX1 I_40954  ( .D(I111124), .CLK(I2702), .RSTB(I698492), .Q(I698944) );
nand I_40955 (I698478,I698944,I698639);
DFFARX1 I_40956  ( .D(I698944), .CLK(I2702), .RSTB(I698492), .Q(I698466) );
nand I_40957 (I698989,I698944,I698605);
and I_40958 (I699006,I698656,I698989);
DFFARX1 I_40959  ( .D(I699006), .CLK(I2702), .RSTB(I698492), .Q(I698460) );
not I_40960 (I699070,I2709);
nand I_40961 (I699087,I589335,I589314);
and I_40962 (I699104,I699087,I589332);
DFFARX1 I_40963  ( .D(I699104), .CLK(I2702), .RSTB(I699070), .Q(I699121) );
not I_40964 (I699059,I699121);
DFFARX1 I_40965  ( .D(I699121), .CLK(I2702), .RSTB(I699070), .Q(I699152) );
not I_40966 (I699047,I699152);
nor I_40967 (I699183,I589344,I589314);
not I_40968 (I699200,I699183);
nor I_40969 (I699217,I699121,I699200);
DFFARX1 I_40970  ( .D(I589320), .CLK(I2702), .RSTB(I699070), .Q(I699234) );
not I_40971 (I699251,I699234);
nand I_40972 (I699050,I699234,I699200);
DFFARX1 I_40973  ( .D(I699234), .CLK(I2702), .RSTB(I699070), .Q(I699282) );
and I_40974 (I699035,I699121,I699282);
nand I_40975 (I699313,I589329,I589317);
and I_40976 (I699330,I699313,I589341);
DFFARX1 I_40977  ( .D(I699330), .CLK(I2702), .RSTB(I699070), .Q(I699347) );
nor I_40978 (I699364,I699347,I699251);
and I_40979 (I699381,I699183,I699364);
nor I_40980 (I699398,I699347,I699121);
DFFARX1 I_40981  ( .D(I699347), .CLK(I2702), .RSTB(I699070), .Q(I699041) );
DFFARX1 I_40982  ( .D(I589326), .CLK(I2702), .RSTB(I699070), .Q(I699429) );
and I_40983 (I699446,I699429,I589338);
or I_40984 (I699463,I699446,I699381);
DFFARX1 I_40985  ( .D(I699463), .CLK(I2702), .RSTB(I699070), .Q(I699053) );
nand I_40986 (I699062,I699446,I699398);
DFFARX1 I_40987  ( .D(I699446), .CLK(I2702), .RSTB(I699070), .Q(I699032) );
DFFARX1 I_40988  ( .D(I589323), .CLK(I2702), .RSTB(I699070), .Q(I699522) );
nand I_40989 (I699056,I699522,I699217);
DFFARX1 I_40990  ( .D(I699522), .CLK(I2702), .RSTB(I699070), .Q(I699044) );
nand I_40991 (I699567,I699522,I699183);
and I_40992 (I699584,I699234,I699567);
DFFARX1 I_40993  ( .D(I699584), .CLK(I2702), .RSTB(I699070), .Q(I699038) );
not I_40994 (I699648,I2709);
nand I_40995 (I699665,I654563,I654581);
and I_40996 (I699682,I699665,I654578);
DFFARX1 I_40997  ( .D(I699682), .CLK(I2702), .RSTB(I699648), .Q(I699699) );
not I_40998 (I699637,I699699);
DFFARX1 I_40999  ( .D(I699699), .CLK(I2702), .RSTB(I699648), .Q(I699730) );
not I_41000 (I699625,I699730);
nor I_41001 (I699761,I654584,I654581);
not I_41002 (I699778,I699761);
nor I_41003 (I699795,I699699,I699778);
DFFARX1 I_41004  ( .D(I654587), .CLK(I2702), .RSTB(I699648), .Q(I699812) );
not I_41005 (I699829,I699812);
nand I_41006 (I699628,I699812,I699778);
DFFARX1 I_41007  ( .D(I699812), .CLK(I2702), .RSTB(I699648), .Q(I699860) );
and I_41008 (I699613,I699699,I699860);
nand I_41009 (I699891,I654572,I654566);
and I_41010 (I699908,I699891,I654569);
DFFARX1 I_41011  ( .D(I699908), .CLK(I2702), .RSTB(I699648), .Q(I699925) );
nor I_41012 (I699942,I699925,I699829);
and I_41013 (I699959,I699761,I699942);
nor I_41014 (I699976,I699925,I699699);
DFFARX1 I_41015  ( .D(I699925), .CLK(I2702), .RSTB(I699648), .Q(I699619) );
DFFARX1 I_41016  ( .D(I654575), .CLK(I2702), .RSTB(I699648), .Q(I700007) );
and I_41017 (I700024,I700007,I654560);
or I_41018 (I700041,I700024,I699959);
DFFARX1 I_41019  ( .D(I700041), .CLK(I2702), .RSTB(I699648), .Q(I699631) );
nand I_41020 (I699640,I700024,I699976);
DFFARX1 I_41021  ( .D(I700024), .CLK(I2702), .RSTB(I699648), .Q(I699610) );
DFFARX1 I_41022  ( .D(I654590), .CLK(I2702), .RSTB(I699648), .Q(I700100) );
nand I_41023 (I699634,I700100,I699795);
DFFARX1 I_41024  ( .D(I700100), .CLK(I2702), .RSTB(I699648), .Q(I699622) );
nand I_41025 (I700145,I700100,I699761);
and I_41026 (I700162,I699812,I700145);
DFFARX1 I_41027  ( .D(I700162), .CLK(I2702), .RSTB(I699648), .Q(I699616) );
not I_41028 (I700226,I2709);
nand I_41029 (I700243,I303978,I303975);
and I_41030 (I700260,I700243,I303999);
DFFARX1 I_41031  ( .D(I700260), .CLK(I2702), .RSTB(I700226), .Q(I700277) );
not I_41032 (I700215,I700277);
DFFARX1 I_41033  ( .D(I700277), .CLK(I2702), .RSTB(I700226), .Q(I700308) );
not I_41034 (I700203,I700308);
nor I_41035 (I700339,I303981,I303975);
not I_41036 (I700356,I700339);
nor I_41037 (I700373,I700277,I700356);
DFFARX1 I_41038  ( .D(I303996), .CLK(I2702), .RSTB(I700226), .Q(I700390) );
not I_41039 (I700407,I700390);
nand I_41040 (I700206,I700390,I700356);
DFFARX1 I_41041  ( .D(I700390), .CLK(I2702), .RSTB(I700226), .Q(I700438) );
and I_41042 (I700191,I700277,I700438);
nand I_41043 (I700469,I303984,I303969);
and I_41044 (I700486,I700469,I303987);
DFFARX1 I_41045  ( .D(I700486), .CLK(I2702), .RSTB(I700226), .Q(I700503) );
nor I_41046 (I700520,I700503,I700407);
and I_41047 (I700537,I700339,I700520);
nor I_41048 (I700554,I700503,I700277);
DFFARX1 I_41049  ( .D(I700503), .CLK(I2702), .RSTB(I700226), .Q(I700197) );
DFFARX1 I_41050  ( .D(I303990), .CLK(I2702), .RSTB(I700226), .Q(I700585) );
and I_41051 (I700602,I700585,I303993);
or I_41052 (I700619,I700602,I700537);
DFFARX1 I_41053  ( .D(I700619), .CLK(I2702), .RSTB(I700226), .Q(I700209) );
nand I_41054 (I700218,I700602,I700554);
DFFARX1 I_41055  ( .D(I700602), .CLK(I2702), .RSTB(I700226), .Q(I700188) );
DFFARX1 I_41056  ( .D(I303972), .CLK(I2702), .RSTB(I700226), .Q(I700678) );
nand I_41057 (I700212,I700678,I700373);
DFFARX1 I_41058  ( .D(I700678), .CLK(I2702), .RSTB(I700226), .Q(I700200) );
nand I_41059 (I700723,I700678,I700339);
and I_41060 (I700740,I700390,I700723);
DFFARX1 I_41061  ( .D(I700740), .CLK(I2702), .RSTB(I700226), .Q(I700194) );
not I_41062 (I700804,I2709);
nand I_41063 (I700821,I148164,I148194);
and I_41064 (I700838,I700821,I148176);
DFFARX1 I_41065  ( .D(I700838), .CLK(I2702), .RSTB(I700804), .Q(I700855) );
not I_41066 (I700793,I700855);
DFFARX1 I_41067  ( .D(I700855), .CLK(I2702), .RSTB(I700804), .Q(I700886) );
not I_41068 (I700781,I700886);
nor I_41069 (I700917,I148173,I148194);
not I_41070 (I700934,I700917);
nor I_41071 (I700951,I700855,I700934);
DFFARX1 I_41072  ( .D(I148167), .CLK(I2702), .RSTB(I700804), .Q(I700968) );
not I_41073 (I700985,I700968);
nand I_41074 (I700784,I700968,I700934);
DFFARX1 I_41075  ( .D(I700968), .CLK(I2702), .RSTB(I700804), .Q(I701016) );
and I_41076 (I700769,I700855,I701016);
nand I_41077 (I701047,I148170,I148185);
and I_41078 (I701064,I701047,I148182);
DFFARX1 I_41079  ( .D(I701064), .CLK(I2702), .RSTB(I700804), .Q(I701081) );
nor I_41080 (I701098,I701081,I700985);
and I_41081 (I701115,I700917,I701098);
nor I_41082 (I701132,I701081,I700855);
DFFARX1 I_41083  ( .D(I701081), .CLK(I2702), .RSTB(I700804), .Q(I700775) );
DFFARX1 I_41084  ( .D(I148179), .CLK(I2702), .RSTB(I700804), .Q(I701163) );
and I_41085 (I701180,I701163,I148191);
or I_41086 (I701197,I701180,I701115);
DFFARX1 I_41087  ( .D(I701197), .CLK(I2702), .RSTB(I700804), .Q(I700787) );
nand I_41088 (I700796,I701180,I701132);
DFFARX1 I_41089  ( .D(I701180), .CLK(I2702), .RSTB(I700804), .Q(I700766) );
DFFARX1 I_41090  ( .D(I148188), .CLK(I2702), .RSTB(I700804), .Q(I701256) );
nand I_41091 (I700790,I701256,I700951);
DFFARX1 I_41092  ( .D(I701256), .CLK(I2702), .RSTB(I700804), .Q(I700778) );
nand I_41093 (I701301,I701256,I700917);
and I_41094 (I701318,I700968,I701301);
DFFARX1 I_41095  ( .D(I701318), .CLK(I2702), .RSTB(I700804), .Q(I700772) );
not I_41096 (I701382,I2709);
nand I_41097 (I701399,I545900,I545882);
and I_41098 (I701416,I701399,I545897);
DFFARX1 I_41099  ( .D(I701416), .CLK(I2702), .RSTB(I701382), .Q(I701433) );
not I_41100 (I701371,I701433);
DFFARX1 I_41101  ( .D(I701433), .CLK(I2702), .RSTB(I701382), .Q(I701464) );
not I_41102 (I701359,I701464);
nor I_41103 (I701495,I545888,I545882);
not I_41104 (I701512,I701495);
nor I_41105 (I701529,I701433,I701512);
DFFARX1 I_41106  ( .D(I545903), .CLK(I2702), .RSTB(I701382), .Q(I701546) );
not I_41107 (I701563,I701546);
nand I_41108 (I701362,I701546,I701512);
DFFARX1 I_41109  ( .D(I701546), .CLK(I2702), .RSTB(I701382), .Q(I701594) );
and I_41110 (I701347,I701433,I701594);
nand I_41111 (I701625,I545879,I545885);
and I_41112 (I701642,I701625,I545891);
DFFARX1 I_41113  ( .D(I701642), .CLK(I2702), .RSTB(I701382), .Q(I701659) );
nor I_41114 (I701676,I701659,I701563);
and I_41115 (I701693,I701495,I701676);
nor I_41116 (I701710,I701659,I701433);
DFFARX1 I_41117  ( .D(I701659), .CLK(I2702), .RSTB(I701382), .Q(I701353) );
DFFARX1 I_41118  ( .D(I545906), .CLK(I2702), .RSTB(I701382), .Q(I701741) );
and I_41119 (I701758,I701741,I545894);
or I_41120 (I701775,I701758,I701693);
DFFARX1 I_41121  ( .D(I701775), .CLK(I2702), .RSTB(I701382), .Q(I701365) );
nand I_41122 (I701374,I701758,I701710);
DFFARX1 I_41123  ( .D(I701758), .CLK(I2702), .RSTB(I701382), .Q(I701344) );
DFFARX1 I_41124  ( .D(I545909), .CLK(I2702), .RSTB(I701382), .Q(I701834) );
nand I_41125 (I701368,I701834,I701529);
DFFARX1 I_41126  ( .D(I701834), .CLK(I2702), .RSTB(I701382), .Q(I701356) );
nand I_41127 (I701879,I701834,I701495);
and I_41128 (I701896,I701546,I701879);
DFFARX1 I_41129  ( .D(I701896), .CLK(I2702), .RSTB(I701382), .Q(I701350) );
not I_41130 (I701960,I2709);
nand I_41131 (I701977,I323868,I323865);
and I_41132 (I701994,I701977,I323889);
DFFARX1 I_41133  ( .D(I701994), .CLK(I2702), .RSTB(I701960), .Q(I702011) );
not I_41134 (I701949,I702011);
DFFARX1 I_41135  ( .D(I702011), .CLK(I2702), .RSTB(I701960), .Q(I702042) );
not I_41136 (I701937,I702042);
nor I_41137 (I702073,I323871,I323865);
not I_41138 (I702090,I702073);
nor I_41139 (I702107,I702011,I702090);
DFFARX1 I_41140  ( .D(I323886), .CLK(I2702), .RSTB(I701960), .Q(I702124) );
not I_41141 (I702141,I702124);
nand I_41142 (I701940,I702124,I702090);
DFFARX1 I_41143  ( .D(I702124), .CLK(I2702), .RSTB(I701960), .Q(I702172) );
and I_41144 (I701925,I702011,I702172);
nand I_41145 (I702203,I323874,I323859);
and I_41146 (I702220,I702203,I323877);
DFFARX1 I_41147  ( .D(I702220), .CLK(I2702), .RSTB(I701960), .Q(I702237) );
nor I_41148 (I702254,I702237,I702141);
and I_41149 (I702271,I702073,I702254);
nor I_41150 (I702288,I702237,I702011);
DFFARX1 I_41151  ( .D(I702237), .CLK(I2702), .RSTB(I701960), .Q(I701931) );
DFFARX1 I_41152  ( .D(I323880), .CLK(I2702), .RSTB(I701960), .Q(I702319) );
and I_41153 (I702336,I702319,I323883);
or I_41154 (I702353,I702336,I702271);
DFFARX1 I_41155  ( .D(I702353), .CLK(I2702), .RSTB(I701960), .Q(I701943) );
nand I_41156 (I701952,I702336,I702288);
DFFARX1 I_41157  ( .D(I702336), .CLK(I2702), .RSTB(I701960), .Q(I701922) );
DFFARX1 I_41158  ( .D(I323862), .CLK(I2702), .RSTB(I701960), .Q(I702412) );
nand I_41159 (I701946,I702412,I702107);
DFFARX1 I_41160  ( .D(I702412), .CLK(I2702), .RSTB(I701960), .Q(I701934) );
nand I_41161 (I702457,I702412,I702073);
and I_41162 (I702474,I702124,I702457);
DFFARX1 I_41163  ( .D(I702474), .CLK(I2702), .RSTB(I701960), .Q(I701928) );
not I_41164 (I702538,I2709);
nand I_41165 (I702555,I48738,I48723);
and I_41166 (I702572,I702555,I48732);
DFFARX1 I_41167  ( .D(I702572), .CLK(I2702), .RSTB(I702538), .Q(I702589) );
not I_41168 (I702527,I702589);
DFFARX1 I_41169  ( .D(I702589), .CLK(I2702), .RSTB(I702538), .Q(I702620) );
not I_41170 (I702515,I702620);
nor I_41171 (I702651,I48744,I48723);
not I_41172 (I702668,I702651);
nor I_41173 (I702685,I702589,I702668);
DFFARX1 I_41174  ( .D(I48735), .CLK(I2702), .RSTB(I702538), .Q(I702702) );
not I_41175 (I702719,I702702);
nand I_41176 (I702518,I702702,I702668);
DFFARX1 I_41177  ( .D(I702702), .CLK(I2702), .RSTB(I702538), .Q(I702750) );
and I_41178 (I702503,I702589,I702750);
nand I_41179 (I702781,I48720,I48714);
and I_41180 (I702798,I702781,I48729);
DFFARX1 I_41181  ( .D(I702798), .CLK(I2702), .RSTB(I702538), .Q(I702815) );
nor I_41182 (I702832,I702815,I702719);
and I_41183 (I702849,I702651,I702832);
nor I_41184 (I702866,I702815,I702589);
DFFARX1 I_41185  ( .D(I702815), .CLK(I2702), .RSTB(I702538), .Q(I702509) );
DFFARX1 I_41186  ( .D(I48717), .CLK(I2702), .RSTB(I702538), .Q(I702897) );
and I_41187 (I702914,I702897,I48741);
or I_41188 (I702931,I702914,I702849);
DFFARX1 I_41189  ( .D(I702931), .CLK(I2702), .RSTB(I702538), .Q(I702521) );
nand I_41190 (I702530,I702914,I702866);
DFFARX1 I_41191  ( .D(I702914), .CLK(I2702), .RSTB(I702538), .Q(I702500) );
DFFARX1 I_41192  ( .D(I48726), .CLK(I2702), .RSTB(I702538), .Q(I702990) );
nand I_41193 (I702524,I702990,I702685);
DFFARX1 I_41194  ( .D(I702990), .CLK(I2702), .RSTB(I702538), .Q(I702512) );
nand I_41195 (I703035,I702990,I702651);
and I_41196 (I703052,I702702,I703035);
DFFARX1 I_41197  ( .D(I703052), .CLK(I2702), .RSTB(I702538), .Q(I702506) );
not I_41198 (I703116,I2709);
nand I_41199 (I703133,I634435,I634453);
and I_41200 (I703150,I703133,I634450);
DFFARX1 I_41201  ( .D(I703150), .CLK(I2702), .RSTB(I703116), .Q(I703167) );
not I_41202 (I703105,I703167);
DFFARX1 I_41203  ( .D(I703167), .CLK(I2702), .RSTB(I703116), .Q(I703198) );
not I_41204 (I703093,I703198);
nor I_41205 (I703229,I634456,I634453);
not I_41206 (I703246,I703229);
nor I_41207 (I703263,I703167,I703246);
DFFARX1 I_41208  ( .D(I634459), .CLK(I2702), .RSTB(I703116), .Q(I703280) );
not I_41209 (I703297,I703280);
nand I_41210 (I703096,I703280,I703246);
DFFARX1 I_41211  ( .D(I703280), .CLK(I2702), .RSTB(I703116), .Q(I703328) );
and I_41212 (I703081,I703167,I703328);
nand I_41213 (I703359,I634444,I634438);
and I_41214 (I703376,I703359,I634441);
DFFARX1 I_41215  ( .D(I703376), .CLK(I2702), .RSTB(I703116), .Q(I703393) );
nor I_41216 (I703410,I703393,I703297);
and I_41217 (I703427,I703229,I703410);
nor I_41218 (I703444,I703393,I703167);
DFFARX1 I_41219  ( .D(I703393), .CLK(I2702), .RSTB(I703116), .Q(I703087) );
DFFARX1 I_41220  ( .D(I634447), .CLK(I2702), .RSTB(I703116), .Q(I703475) );
and I_41221 (I703492,I703475,I634432);
or I_41222 (I703509,I703492,I703427);
DFFARX1 I_41223  ( .D(I703509), .CLK(I2702), .RSTB(I703116), .Q(I703099) );
nand I_41224 (I703108,I703492,I703444);
DFFARX1 I_41225  ( .D(I703492), .CLK(I2702), .RSTB(I703116), .Q(I703078) );
DFFARX1 I_41226  ( .D(I634462), .CLK(I2702), .RSTB(I703116), .Q(I703568) );
nand I_41227 (I703102,I703568,I703263);
DFFARX1 I_41228  ( .D(I703568), .CLK(I2702), .RSTB(I703116), .Q(I703090) );
nand I_41229 (I703613,I703568,I703229);
and I_41230 (I703630,I703280,I703613);
DFFARX1 I_41231  ( .D(I703630), .CLK(I2702), .RSTB(I703116), .Q(I703084) );
not I_41232 (I703694,I2709);
nand I_41233 (I703711,I630032,I630050);
and I_41234 (I703728,I703711,I630047);
DFFARX1 I_41235  ( .D(I703728), .CLK(I2702), .RSTB(I703694), .Q(I703745) );
not I_41236 (I703683,I703745);
DFFARX1 I_41237  ( .D(I703745), .CLK(I2702), .RSTB(I703694), .Q(I703776) );
not I_41238 (I703671,I703776);
nor I_41239 (I703807,I630053,I630050);
not I_41240 (I703824,I703807);
nor I_41241 (I703841,I703745,I703824);
DFFARX1 I_41242  ( .D(I630056), .CLK(I2702), .RSTB(I703694), .Q(I703858) );
not I_41243 (I703875,I703858);
nand I_41244 (I703674,I703858,I703824);
DFFARX1 I_41245  ( .D(I703858), .CLK(I2702), .RSTB(I703694), .Q(I703906) );
and I_41246 (I703659,I703745,I703906);
nand I_41247 (I703937,I630041,I630035);
and I_41248 (I703954,I703937,I630038);
DFFARX1 I_41249  ( .D(I703954), .CLK(I2702), .RSTB(I703694), .Q(I703971) );
nor I_41250 (I703988,I703971,I703875);
and I_41251 (I704005,I703807,I703988);
nor I_41252 (I704022,I703971,I703745);
DFFARX1 I_41253  ( .D(I703971), .CLK(I2702), .RSTB(I703694), .Q(I703665) );
DFFARX1 I_41254  ( .D(I630044), .CLK(I2702), .RSTB(I703694), .Q(I704053) );
and I_41255 (I704070,I704053,I630029);
or I_41256 (I704087,I704070,I704005);
DFFARX1 I_41257  ( .D(I704087), .CLK(I2702), .RSTB(I703694), .Q(I703677) );
nand I_41258 (I703686,I704070,I704022);
DFFARX1 I_41259  ( .D(I704070), .CLK(I2702), .RSTB(I703694), .Q(I703656) );
DFFARX1 I_41260  ( .D(I630059), .CLK(I2702), .RSTB(I703694), .Q(I704146) );
nand I_41261 (I703680,I704146,I703841);
DFFARX1 I_41262  ( .D(I704146), .CLK(I2702), .RSTB(I703694), .Q(I703668) );
nand I_41263 (I704191,I704146,I703807);
and I_41264 (I704208,I703858,I704191);
DFFARX1 I_41265  ( .D(I704208), .CLK(I2702), .RSTB(I703694), .Q(I703662) );
not I_41266 (I704272,I2709);
nand I_41267 (I704289,I558990,I558972);
and I_41268 (I704306,I704289,I558987);
DFFARX1 I_41269  ( .D(I704306), .CLK(I2702), .RSTB(I704272), .Q(I704323) );
not I_41270 (I704261,I704323);
DFFARX1 I_41271  ( .D(I704323), .CLK(I2702), .RSTB(I704272), .Q(I704354) );
not I_41272 (I704249,I704354);
nor I_41273 (I704385,I558978,I558972);
not I_41274 (I704402,I704385);
nor I_41275 (I704419,I704323,I704402);
DFFARX1 I_41276  ( .D(I558993), .CLK(I2702), .RSTB(I704272), .Q(I704436) );
not I_41277 (I704453,I704436);
nand I_41278 (I704252,I704436,I704402);
DFFARX1 I_41279  ( .D(I704436), .CLK(I2702), .RSTB(I704272), .Q(I704484) );
and I_41280 (I704237,I704323,I704484);
nand I_41281 (I704515,I558969,I558975);
and I_41282 (I704532,I704515,I558981);
DFFARX1 I_41283  ( .D(I704532), .CLK(I2702), .RSTB(I704272), .Q(I704549) );
nor I_41284 (I704566,I704549,I704453);
and I_41285 (I704583,I704385,I704566);
nor I_41286 (I704600,I704549,I704323);
DFFARX1 I_41287  ( .D(I704549), .CLK(I2702), .RSTB(I704272), .Q(I704243) );
DFFARX1 I_41288  ( .D(I558996), .CLK(I2702), .RSTB(I704272), .Q(I704631) );
and I_41289 (I704648,I704631,I558984);
or I_41290 (I704665,I704648,I704583);
DFFARX1 I_41291  ( .D(I704665), .CLK(I2702), .RSTB(I704272), .Q(I704255) );
nand I_41292 (I704264,I704648,I704600);
DFFARX1 I_41293  ( .D(I704648), .CLK(I2702), .RSTB(I704272), .Q(I704234) );
DFFARX1 I_41294  ( .D(I558999), .CLK(I2702), .RSTB(I704272), .Q(I704724) );
nand I_41295 (I704258,I704724,I704419);
DFFARX1 I_41296  ( .D(I704724), .CLK(I2702), .RSTB(I704272), .Q(I704246) );
nand I_41297 (I704769,I704724,I704385);
and I_41298 (I704786,I704436,I704769);
DFFARX1 I_41299  ( .D(I704786), .CLK(I2702), .RSTB(I704272), .Q(I704240) );
not I_41300 (I704850,I2709);
nand I_41301 (I704867,I188607,I188637);
and I_41302 (I704884,I704867,I188619);
DFFARX1 I_41303  ( .D(I704884), .CLK(I2702), .RSTB(I704850), .Q(I704901) );
not I_41304 (I704839,I704901);
DFFARX1 I_41305  ( .D(I704901), .CLK(I2702), .RSTB(I704850), .Q(I704932) );
not I_41306 (I704827,I704932);
nor I_41307 (I704963,I188616,I188637);
not I_41308 (I704980,I704963);
nor I_41309 (I704997,I704901,I704980);
DFFARX1 I_41310  ( .D(I188610), .CLK(I2702), .RSTB(I704850), .Q(I705014) );
not I_41311 (I705031,I705014);
nand I_41312 (I704830,I705014,I704980);
DFFARX1 I_41313  ( .D(I705014), .CLK(I2702), .RSTB(I704850), .Q(I705062) );
and I_41314 (I704815,I704901,I705062);
nand I_41315 (I705093,I188613,I188628);
and I_41316 (I705110,I705093,I188625);
DFFARX1 I_41317  ( .D(I705110), .CLK(I2702), .RSTB(I704850), .Q(I705127) );
nor I_41318 (I705144,I705127,I705031);
and I_41319 (I705161,I704963,I705144);
nor I_41320 (I705178,I705127,I704901);
DFFARX1 I_41321  ( .D(I705127), .CLK(I2702), .RSTB(I704850), .Q(I704821) );
DFFARX1 I_41322  ( .D(I188622), .CLK(I2702), .RSTB(I704850), .Q(I705209) );
and I_41323 (I705226,I705209,I188634);
or I_41324 (I705243,I705226,I705161);
DFFARX1 I_41325  ( .D(I705243), .CLK(I2702), .RSTB(I704850), .Q(I704833) );
nand I_41326 (I704842,I705226,I705178);
DFFARX1 I_41327  ( .D(I705226), .CLK(I2702), .RSTB(I704850), .Q(I704812) );
DFFARX1 I_41328  ( .D(I188631), .CLK(I2702), .RSTB(I704850), .Q(I705302) );
nand I_41329 (I704836,I705302,I704997);
DFFARX1 I_41330  ( .D(I705302), .CLK(I2702), .RSTB(I704850), .Q(I704824) );
nand I_41331 (I705347,I705302,I704963);
and I_41332 (I705364,I705014,I705347);
DFFARX1 I_41333  ( .D(I705364), .CLK(I2702), .RSTB(I704850), .Q(I704818) );
not I_41334 (I705428,I2709);
nand I_41335 (I705445,I332487,I332484);
and I_41336 (I705462,I705445,I332508);
DFFARX1 I_41337  ( .D(I705462), .CLK(I2702), .RSTB(I705428), .Q(I705479) );
not I_41338 (I705417,I705479);
DFFARX1 I_41339  ( .D(I705479), .CLK(I2702), .RSTB(I705428), .Q(I705510) );
not I_41340 (I705405,I705510);
nor I_41341 (I705541,I332490,I332484);
not I_41342 (I705558,I705541);
nor I_41343 (I705575,I705479,I705558);
DFFARX1 I_41344  ( .D(I332505), .CLK(I2702), .RSTB(I705428), .Q(I705592) );
not I_41345 (I705609,I705592);
nand I_41346 (I705408,I705592,I705558);
DFFARX1 I_41347  ( .D(I705592), .CLK(I2702), .RSTB(I705428), .Q(I705640) );
and I_41348 (I705393,I705479,I705640);
nand I_41349 (I705671,I332493,I332478);
and I_41350 (I705688,I705671,I332496);
DFFARX1 I_41351  ( .D(I705688), .CLK(I2702), .RSTB(I705428), .Q(I705705) );
nor I_41352 (I705722,I705705,I705609);
and I_41353 (I705739,I705541,I705722);
nor I_41354 (I705756,I705705,I705479);
DFFARX1 I_41355  ( .D(I705705), .CLK(I2702), .RSTB(I705428), .Q(I705399) );
DFFARX1 I_41356  ( .D(I332499), .CLK(I2702), .RSTB(I705428), .Q(I705787) );
and I_41357 (I705804,I705787,I332502);
or I_41358 (I705821,I705804,I705739);
DFFARX1 I_41359  ( .D(I705821), .CLK(I2702), .RSTB(I705428), .Q(I705411) );
nand I_41360 (I705420,I705804,I705756);
DFFARX1 I_41361  ( .D(I705804), .CLK(I2702), .RSTB(I705428), .Q(I705390) );
DFFARX1 I_41362  ( .D(I332481), .CLK(I2702), .RSTB(I705428), .Q(I705880) );
nand I_41363 (I705414,I705880,I705575);
DFFARX1 I_41364  ( .D(I705880), .CLK(I2702), .RSTB(I705428), .Q(I705402) );
nand I_41365 (I705925,I705880,I705541);
and I_41366 (I705942,I705592,I705925);
DFFARX1 I_41367  ( .D(I705942), .CLK(I2702), .RSTB(I705428), .Q(I705396) );
not I_41368 (I706006,I2709);
nand I_41369 (I706023,I665256,I665274);
and I_41370 (I706040,I706023,I665271);
DFFARX1 I_41371  ( .D(I706040), .CLK(I2702), .RSTB(I706006), .Q(I706057) );
not I_41372 (I705995,I706057);
DFFARX1 I_41373  ( .D(I706057), .CLK(I2702), .RSTB(I706006), .Q(I706088) );
not I_41374 (I705983,I706088);
nor I_41375 (I706119,I665277,I665274);
not I_41376 (I706136,I706119);
nor I_41377 (I706153,I706057,I706136);
DFFARX1 I_41378  ( .D(I665280), .CLK(I2702), .RSTB(I706006), .Q(I706170) );
not I_41379 (I706187,I706170);
nand I_41380 (I705986,I706170,I706136);
DFFARX1 I_41381  ( .D(I706170), .CLK(I2702), .RSTB(I706006), .Q(I706218) );
and I_41382 (I705971,I706057,I706218);
nand I_41383 (I706249,I665265,I665259);
and I_41384 (I706266,I706249,I665262);
DFFARX1 I_41385  ( .D(I706266), .CLK(I2702), .RSTB(I706006), .Q(I706283) );
nor I_41386 (I706300,I706283,I706187);
and I_41387 (I706317,I706119,I706300);
nor I_41388 (I706334,I706283,I706057);
DFFARX1 I_41389  ( .D(I706283), .CLK(I2702), .RSTB(I706006), .Q(I705977) );
DFFARX1 I_41390  ( .D(I665268), .CLK(I2702), .RSTB(I706006), .Q(I706365) );
and I_41391 (I706382,I706365,I665253);
or I_41392 (I706399,I706382,I706317);
DFFARX1 I_41393  ( .D(I706399), .CLK(I2702), .RSTB(I706006), .Q(I705989) );
nand I_41394 (I705998,I706382,I706334);
DFFARX1 I_41395  ( .D(I706382), .CLK(I2702), .RSTB(I706006), .Q(I705968) );
DFFARX1 I_41396  ( .D(I665283), .CLK(I2702), .RSTB(I706006), .Q(I706458) );
nand I_41397 (I705992,I706458,I706153);
DFFARX1 I_41398  ( .D(I706458), .CLK(I2702), .RSTB(I706006), .Q(I705980) );
nand I_41399 (I706503,I706458,I706119);
and I_41400 (I706520,I706170,I706503);
DFFARX1 I_41401  ( .D(I706520), .CLK(I2702), .RSTB(I706006), .Q(I705974) );
not I_41402 (I706584,I2709);
nand I_41403 (I706601,I209407,I209404);
and I_41404 (I706618,I706601,I209416);
DFFARX1 I_41405  ( .D(I706618), .CLK(I2702), .RSTB(I706584), .Q(I706635) );
not I_41406 (I706573,I706635);
DFFARX1 I_41407  ( .D(I706635), .CLK(I2702), .RSTB(I706584), .Q(I706666) );
not I_41408 (I706561,I706666);
nor I_41409 (I706697,I209419,I209404);
not I_41410 (I706714,I706697);
nor I_41411 (I706731,I706635,I706714);
DFFARX1 I_41412  ( .D(I209425), .CLK(I2702), .RSTB(I706584), .Q(I706748) );
not I_41413 (I706765,I706748);
nand I_41414 (I706564,I706748,I706714);
DFFARX1 I_41415  ( .D(I706748), .CLK(I2702), .RSTB(I706584), .Q(I706796) );
and I_41416 (I706549,I706635,I706796);
nand I_41417 (I706827,I209398,I209401);
and I_41418 (I706844,I706827,I209410);
DFFARX1 I_41419  ( .D(I706844), .CLK(I2702), .RSTB(I706584), .Q(I706861) );
nor I_41420 (I706878,I706861,I706765);
and I_41421 (I706895,I706697,I706878);
nor I_41422 (I706912,I706861,I706635);
DFFARX1 I_41423  ( .D(I706861), .CLK(I2702), .RSTB(I706584), .Q(I706555) );
DFFARX1 I_41424  ( .D(I209428), .CLK(I2702), .RSTB(I706584), .Q(I706943) );
and I_41425 (I706960,I706943,I209422);
or I_41426 (I706977,I706960,I706895);
DFFARX1 I_41427  ( .D(I706977), .CLK(I2702), .RSTB(I706584), .Q(I706567) );
nand I_41428 (I706576,I706960,I706912);
DFFARX1 I_41429  ( .D(I706960), .CLK(I2702), .RSTB(I706584), .Q(I706546) );
DFFARX1 I_41430  ( .D(I209413), .CLK(I2702), .RSTB(I706584), .Q(I707036) );
nand I_41431 (I706570,I707036,I706731);
DFFARX1 I_41432  ( .D(I707036), .CLK(I2702), .RSTB(I706584), .Q(I706558) );
nand I_41433 (I707081,I707036,I706697);
and I_41434 (I707098,I706748,I707081);
DFFARX1 I_41435  ( .D(I707098), .CLK(I2702), .RSTB(I706584), .Q(I706552) );
not I_41436 (I707162,I2709);
nand I_41437 (I707179,I376441,I376444);
and I_41438 (I707196,I707179,I376423);
DFFARX1 I_41439  ( .D(I707196), .CLK(I2702), .RSTB(I707162), .Q(I707213) );
not I_41440 (I707151,I707213);
DFFARX1 I_41441  ( .D(I707213), .CLK(I2702), .RSTB(I707162), .Q(I707244) );
not I_41442 (I707139,I707244);
nor I_41443 (I707275,I376438,I376444);
not I_41444 (I707292,I707275);
nor I_41445 (I707309,I707213,I707292);
DFFARX1 I_41446  ( .D(I376447), .CLK(I2702), .RSTB(I707162), .Q(I707326) );
not I_41447 (I707343,I707326);
nand I_41448 (I707142,I707326,I707292);
DFFARX1 I_41449  ( .D(I707326), .CLK(I2702), .RSTB(I707162), .Q(I707374) );
and I_41450 (I707127,I707213,I707374);
nand I_41451 (I707405,I376435,I376453);
and I_41452 (I707422,I707405,I376429);
DFFARX1 I_41453  ( .D(I707422), .CLK(I2702), .RSTB(I707162), .Q(I707439) );
nor I_41454 (I707456,I707439,I707343);
and I_41455 (I707473,I707275,I707456);
nor I_41456 (I707490,I707439,I707213);
DFFARX1 I_41457  ( .D(I707439), .CLK(I2702), .RSTB(I707162), .Q(I707133) );
DFFARX1 I_41458  ( .D(I376426), .CLK(I2702), .RSTB(I707162), .Q(I707521) );
and I_41459 (I707538,I707521,I376432);
or I_41460 (I707555,I707538,I707473);
DFFARX1 I_41461  ( .D(I707555), .CLK(I2702), .RSTB(I707162), .Q(I707145) );
nand I_41462 (I707154,I707538,I707490);
DFFARX1 I_41463  ( .D(I707538), .CLK(I2702), .RSTB(I707162), .Q(I707124) );
DFFARX1 I_41464  ( .D(I376450), .CLK(I2702), .RSTB(I707162), .Q(I707614) );
nand I_41465 (I707148,I707614,I707309);
DFFARX1 I_41466  ( .D(I707614), .CLK(I2702), .RSTB(I707162), .Q(I707136) );
nand I_41467 (I707659,I707614,I707275);
and I_41468 (I707676,I707326,I707659);
DFFARX1 I_41469  ( .D(I707676), .CLK(I2702), .RSTB(I707162), .Q(I707130) );
not I_41470 (I707740,I2709);
nand I_41471 (I707757,I476046,I476064);
and I_41472 (I707774,I707757,I476055);
DFFARX1 I_41473  ( .D(I707774), .CLK(I2702), .RSTB(I707740), .Q(I707791) );
not I_41474 (I707729,I707791);
DFFARX1 I_41475  ( .D(I707791), .CLK(I2702), .RSTB(I707740), .Q(I707822) );
not I_41476 (I707717,I707822);
nor I_41477 (I707853,I476052,I476064);
not I_41478 (I707870,I707853);
nor I_41479 (I707887,I707791,I707870);
DFFARX1 I_41480  ( .D(I476043), .CLK(I2702), .RSTB(I707740), .Q(I707904) );
not I_41481 (I707921,I707904);
nand I_41482 (I707720,I707904,I707870);
DFFARX1 I_41483  ( .D(I707904), .CLK(I2702), .RSTB(I707740), .Q(I707952) );
and I_41484 (I707705,I707791,I707952);
nand I_41485 (I707983,I476061,I476073);
and I_41486 (I708000,I707983,I476067);
DFFARX1 I_41487  ( .D(I708000), .CLK(I2702), .RSTB(I707740), .Q(I708017) );
nor I_41488 (I708034,I708017,I707921);
and I_41489 (I708051,I707853,I708034);
nor I_41490 (I708068,I708017,I707791);
DFFARX1 I_41491  ( .D(I708017), .CLK(I2702), .RSTB(I707740), .Q(I707711) );
DFFARX1 I_41492  ( .D(I476049), .CLK(I2702), .RSTB(I707740), .Q(I708099) );
and I_41493 (I708116,I708099,I476058);
or I_41494 (I708133,I708116,I708051);
DFFARX1 I_41495  ( .D(I708133), .CLK(I2702), .RSTB(I707740), .Q(I707723) );
nand I_41496 (I707732,I708116,I708068);
DFFARX1 I_41497  ( .D(I708116), .CLK(I2702), .RSTB(I707740), .Q(I707702) );
DFFARX1 I_41498  ( .D(I476070), .CLK(I2702), .RSTB(I707740), .Q(I708192) );
nand I_41499 (I707726,I708192,I707887);
DFFARX1 I_41500  ( .D(I708192), .CLK(I2702), .RSTB(I707740), .Q(I707714) );
nand I_41501 (I708237,I708192,I707853);
and I_41502 (I708254,I707904,I708237);
DFFARX1 I_41503  ( .D(I708254), .CLK(I2702), .RSTB(I707740), .Q(I707708) );
not I_41504 (I708318,I2709);
nand I_41505 (I708335,I210002,I209999);
and I_41506 (I708352,I708335,I210011);
DFFARX1 I_41507  ( .D(I708352), .CLK(I2702), .RSTB(I708318), .Q(I708369) );
not I_41508 (I708307,I708369);
DFFARX1 I_41509  ( .D(I708369), .CLK(I2702), .RSTB(I708318), .Q(I708400) );
not I_41510 (I708295,I708400);
nor I_41511 (I708431,I210014,I209999);
not I_41512 (I708448,I708431);
nor I_41513 (I708465,I708369,I708448);
DFFARX1 I_41514  ( .D(I210020), .CLK(I2702), .RSTB(I708318), .Q(I708482) );
not I_41515 (I708499,I708482);
nand I_41516 (I708298,I708482,I708448);
DFFARX1 I_41517  ( .D(I708482), .CLK(I2702), .RSTB(I708318), .Q(I708530) );
and I_41518 (I708283,I708369,I708530);
nand I_41519 (I708561,I209993,I209996);
and I_41520 (I708578,I708561,I210005);
DFFARX1 I_41521  ( .D(I708578), .CLK(I2702), .RSTB(I708318), .Q(I708595) );
nor I_41522 (I708612,I708595,I708499);
and I_41523 (I708629,I708431,I708612);
nor I_41524 (I708646,I708595,I708369);
DFFARX1 I_41525  ( .D(I708595), .CLK(I2702), .RSTB(I708318), .Q(I708289) );
DFFARX1 I_41526  ( .D(I210023), .CLK(I2702), .RSTB(I708318), .Q(I708677) );
and I_41527 (I708694,I708677,I210017);
or I_41528 (I708711,I708694,I708629);
DFFARX1 I_41529  ( .D(I708711), .CLK(I2702), .RSTB(I708318), .Q(I708301) );
nand I_41530 (I708310,I708694,I708646);
DFFARX1 I_41531  ( .D(I708694), .CLK(I2702), .RSTB(I708318), .Q(I708280) );
DFFARX1 I_41532  ( .D(I210008), .CLK(I2702), .RSTB(I708318), .Q(I708770) );
nand I_41533 (I708304,I708770,I708465);
DFFARX1 I_41534  ( .D(I708770), .CLK(I2702), .RSTB(I708318), .Q(I708292) );
nand I_41535 (I708815,I708770,I708431);
and I_41536 (I708832,I708482,I708815);
DFFARX1 I_41537  ( .D(I708832), .CLK(I2702), .RSTB(I708318), .Q(I708286) );
not I_41538 (I708896,I2709);
nand I_41539 (I708913,I333805,I333808);
and I_41540 (I708930,I708913,I333787);
DFFARX1 I_41541  ( .D(I708930), .CLK(I2702), .RSTB(I708896), .Q(I708947) );
not I_41542 (I708885,I708947);
DFFARX1 I_41543  ( .D(I708947), .CLK(I2702), .RSTB(I708896), .Q(I708978) );
not I_41544 (I708873,I708978);
nor I_41545 (I709009,I333802,I333808);
not I_41546 (I709026,I709009);
nor I_41547 (I709043,I708947,I709026);
DFFARX1 I_41548  ( .D(I333811), .CLK(I2702), .RSTB(I708896), .Q(I709060) );
not I_41549 (I709077,I709060);
nand I_41550 (I708876,I709060,I709026);
DFFARX1 I_41551  ( .D(I709060), .CLK(I2702), .RSTB(I708896), .Q(I709108) );
and I_41552 (I708861,I708947,I709108);
nand I_41553 (I709139,I333799,I333817);
and I_41554 (I709156,I709139,I333793);
DFFARX1 I_41555  ( .D(I709156), .CLK(I2702), .RSTB(I708896), .Q(I709173) );
nor I_41556 (I709190,I709173,I709077);
and I_41557 (I709207,I709009,I709190);
nor I_41558 (I709224,I709173,I708947);
DFFARX1 I_41559  ( .D(I709173), .CLK(I2702), .RSTB(I708896), .Q(I708867) );
DFFARX1 I_41560  ( .D(I333790), .CLK(I2702), .RSTB(I708896), .Q(I709255) );
and I_41561 (I709272,I709255,I333796);
or I_41562 (I709289,I709272,I709207);
DFFARX1 I_41563  ( .D(I709289), .CLK(I2702), .RSTB(I708896), .Q(I708879) );
nand I_41564 (I708888,I709272,I709224);
DFFARX1 I_41565  ( .D(I709272), .CLK(I2702), .RSTB(I708896), .Q(I708858) );
DFFARX1 I_41566  ( .D(I333814), .CLK(I2702), .RSTB(I708896), .Q(I709348) );
nand I_41567 (I708882,I709348,I709043);
DFFARX1 I_41568  ( .D(I709348), .CLK(I2702), .RSTB(I708896), .Q(I708870) );
nand I_41569 (I709393,I709348,I709009);
and I_41570 (I709410,I709060,I709393);
DFFARX1 I_41571  ( .D(I709410), .CLK(I2702), .RSTB(I708896), .Q(I708864) );
not I_41572 (I709474,I2709);
nand I_41573 (I709491,I20127,I20112);
and I_41574 (I709508,I709491,I20121);
DFFARX1 I_41575  ( .D(I709508), .CLK(I2702), .RSTB(I709474), .Q(I709525) );
not I_41576 (I709463,I709525);
DFFARX1 I_41577  ( .D(I709525), .CLK(I2702), .RSTB(I709474), .Q(I709556) );
not I_41578 (I709451,I709556);
nor I_41579 (I709587,I20133,I20112);
not I_41580 (I709604,I709587);
nor I_41581 (I709621,I709525,I709604);
DFFARX1 I_41582  ( .D(I20124), .CLK(I2702), .RSTB(I709474), .Q(I709638) );
not I_41583 (I709655,I709638);
nand I_41584 (I709454,I709638,I709604);
DFFARX1 I_41585  ( .D(I709638), .CLK(I2702), .RSTB(I709474), .Q(I709686) );
and I_41586 (I709439,I709525,I709686);
nand I_41587 (I709717,I20109,I20103);
and I_41588 (I709734,I709717,I20118);
DFFARX1 I_41589  ( .D(I709734), .CLK(I2702), .RSTB(I709474), .Q(I709751) );
nor I_41590 (I709768,I709751,I709655);
and I_41591 (I709785,I709587,I709768);
nor I_41592 (I709802,I709751,I709525);
DFFARX1 I_41593  ( .D(I709751), .CLK(I2702), .RSTB(I709474), .Q(I709445) );
DFFARX1 I_41594  ( .D(I20106), .CLK(I2702), .RSTB(I709474), .Q(I709833) );
and I_41595 (I709850,I709833,I20130);
or I_41596 (I709867,I709850,I709785);
DFFARX1 I_41597  ( .D(I709867), .CLK(I2702), .RSTB(I709474), .Q(I709457) );
nand I_41598 (I709466,I709850,I709802);
DFFARX1 I_41599  ( .D(I709850), .CLK(I2702), .RSTB(I709474), .Q(I709436) );
DFFARX1 I_41600  ( .D(I20115), .CLK(I2702), .RSTB(I709474), .Q(I709926) );
nand I_41601 (I709460,I709926,I709621);
DFFARX1 I_41602  ( .D(I709926), .CLK(I2702), .RSTB(I709474), .Q(I709448) );
nand I_41603 (I709971,I709926,I709587);
and I_41604 (I709988,I709638,I709971);
DFFARX1 I_41605  ( .D(I709988), .CLK(I2702), .RSTB(I709474), .Q(I709442) );
not I_41606 (I710052,I2709);
nand I_41607 (I710069,I319227,I319224);
and I_41608 (I710086,I710069,I319248);
DFFARX1 I_41609  ( .D(I710086), .CLK(I2702), .RSTB(I710052), .Q(I710103) );
not I_41610 (I710041,I710103);
DFFARX1 I_41611  ( .D(I710103), .CLK(I2702), .RSTB(I710052), .Q(I710134) );
not I_41612 (I710029,I710134);
nor I_41613 (I710165,I319230,I319224);
not I_41614 (I710182,I710165);
nor I_41615 (I710199,I710103,I710182);
DFFARX1 I_41616  ( .D(I319245), .CLK(I2702), .RSTB(I710052), .Q(I710216) );
not I_41617 (I710233,I710216);
nand I_41618 (I710032,I710216,I710182);
DFFARX1 I_41619  ( .D(I710216), .CLK(I2702), .RSTB(I710052), .Q(I710264) );
and I_41620 (I710017,I710103,I710264);
nand I_41621 (I710295,I319233,I319218);
and I_41622 (I710312,I710295,I319236);
DFFARX1 I_41623  ( .D(I710312), .CLK(I2702), .RSTB(I710052), .Q(I710329) );
nor I_41624 (I710346,I710329,I710233);
and I_41625 (I710363,I710165,I710346);
nor I_41626 (I710380,I710329,I710103);
DFFARX1 I_41627  ( .D(I710329), .CLK(I2702), .RSTB(I710052), .Q(I710023) );
DFFARX1 I_41628  ( .D(I319239), .CLK(I2702), .RSTB(I710052), .Q(I710411) );
and I_41629 (I710428,I710411,I319242);
or I_41630 (I710445,I710428,I710363);
DFFARX1 I_41631  ( .D(I710445), .CLK(I2702), .RSTB(I710052), .Q(I710035) );
nand I_41632 (I710044,I710428,I710380);
DFFARX1 I_41633  ( .D(I710428), .CLK(I2702), .RSTB(I710052), .Q(I710014) );
DFFARX1 I_41634  ( .D(I319221), .CLK(I2702), .RSTB(I710052), .Q(I710504) );
nand I_41635 (I710038,I710504,I710199);
DFFARX1 I_41636  ( .D(I710504), .CLK(I2702), .RSTB(I710052), .Q(I710026) );
nand I_41637 (I710549,I710504,I710165);
and I_41638 (I710566,I710216,I710549);
DFFARX1 I_41639  ( .D(I710566), .CLK(I2702), .RSTB(I710052), .Q(I710020) );
not I_41640 (I710630,I2709);
nand I_41641 (I710647,I18444,I18429);
and I_41642 (I710664,I710647,I18438);
DFFARX1 I_41643  ( .D(I710664), .CLK(I2702), .RSTB(I710630), .Q(I710681) );
not I_41644 (I710619,I710681);
DFFARX1 I_41645  ( .D(I710681), .CLK(I2702), .RSTB(I710630), .Q(I710712) );
not I_41646 (I710607,I710712);
nor I_41647 (I710743,I18450,I18429);
not I_41648 (I710760,I710743);
nor I_41649 (I710777,I710681,I710760);
DFFARX1 I_41650  ( .D(I18441), .CLK(I2702), .RSTB(I710630), .Q(I710794) );
not I_41651 (I710811,I710794);
nand I_41652 (I710610,I710794,I710760);
DFFARX1 I_41653  ( .D(I710794), .CLK(I2702), .RSTB(I710630), .Q(I710842) );
and I_41654 (I710595,I710681,I710842);
nand I_41655 (I710873,I18426,I18420);
and I_41656 (I710890,I710873,I18435);
DFFARX1 I_41657  ( .D(I710890), .CLK(I2702), .RSTB(I710630), .Q(I710907) );
nor I_41658 (I710924,I710907,I710811);
and I_41659 (I710941,I710743,I710924);
nor I_41660 (I710958,I710907,I710681);
DFFARX1 I_41661  ( .D(I710907), .CLK(I2702), .RSTB(I710630), .Q(I710601) );
DFFARX1 I_41662  ( .D(I18423), .CLK(I2702), .RSTB(I710630), .Q(I710989) );
and I_41663 (I711006,I710989,I18447);
or I_41664 (I711023,I711006,I710941);
DFFARX1 I_41665  ( .D(I711023), .CLK(I2702), .RSTB(I710630), .Q(I710613) );
nand I_41666 (I710622,I711006,I710958);
DFFARX1 I_41667  ( .D(I711006), .CLK(I2702), .RSTB(I710630), .Q(I710592) );
DFFARX1 I_41668  ( .D(I18432), .CLK(I2702), .RSTB(I710630), .Q(I711082) );
nand I_41669 (I710616,I711082,I710777);
DFFARX1 I_41670  ( .D(I711082), .CLK(I2702), .RSTB(I710630), .Q(I710604) );
nand I_41671 (I711127,I711082,I710743);
and I_41672 (I711144,I710794,I711127);
DFFARX1 I_41673  ( .D(I711144), .CLK(I2702), .RSTB(I710630), .Q(I710598) );
not I_41674 (I711208,I2709);
nand I_41675 (I711225,I31347,I31332);
and I_41676 (I711242,I711225,I31341);
DFFARX1 I_41677  ( .D(I711242), .CLK(I2702), .RSTB(I711208), .Q(I711259) );
not I_41678 (I711197,I711259);
DFFARX1 I_41679  ( .D(I711259), .CLK(I2702), .RSTB(I711208), .Q(I711290) );
not I_41680 (I711185,I711290);
nor I_41681 (I711321,I31353,I31332);
not I_41682 (I711338,I711321);
nor I_41683 (I711355,I711259,I711338);
DFFARX1 I_41684  ( .D(I31344), .CLK(I2702), .RSTB(I711208), .Q(I711372) );
not I_41685 (I711389,I711372);
nand I_41686 (I711188,I711372,I711338);
DFFARX1 I_41687  ( .D(I711372), .CLK(I2702), .RSTB(I711208), .Q(I711420) );
and I_41688 (I711173,I711259,I711420);
nand I_41689 (I711451,I31329,I31323);
and I_41690 (I711468,I711451,I31338);
DFFARX1 I_41691  ( .D(I711468), .CLK(I2702), .RSTB(I711208), .Q(I711485) );
nor I_41692 (I711502,I711485,I711389);
and I_41693 (I711519,I711321,I711502);
nor I_41694 (I711536,I711485,I711259);
DFFARX1 I_41695  ( .D(I711485), .CLK(I2702), .RSTB(I711208), .Q(I711179) );
DFFARX1 I_41696  ( .D(I31326), .CLK(I2702), .RSTB(I711208), .Q(I711567) );
and I_41697 (I711584,I711567,I31350);
or I_41698 (I711601,I711584,I711519);
DFFARX1 I_41699  ( .D(I711601), .CLK(I2702), .RSTB(I711208), .Q(I711191) );
nand I_41700 (I711200,I711584,I711536);
DFFARX1 I_41701  ( .D(I711584), .CLK(I2702), .RSTB(I711208), .Q(I711170) );
DFFARX1 I_41702  ( .D(I31335), .CLK(I2702), .RSTB(I711208), .Q(I711660) );
nand I_41703 (I711194,I711660,I711355);
DFFARX1 I_41704  ( .D(I711660), .CLK(I2702), .RSTB(I711208), .Q(I711182) );
nand I_41705 (I711705,I711660,I711321);
and I_41706 (I711722,I711372,I711705);
DFFARX1 I_41707  ( .D(I711722), .CLK(I2702), .RSTB(I711208), .Q(I711176) );
not I_41708 (I711786,I2709);
nand I_41709 (I711803,I458706,I458724);
and I_41710 (I711820,I711803,I458715);
DFFARX1 I_41711  ( .D(I711820), .CLK(I2702), .RSTB(I711786), .Q(I711837) );
not I_41712 (I711775,I711837);
DFFARX1 I_41713  ( .D(I711837), .CLK(I2702), .RSTB(I711786), .Q(I711868) );
not I_41714 (I711763,I711868);
nor I_41715 (I711899,I458712,I458724);
not I_41716 (I711916,I711899);
nor I_41717 (I711933,I711837,I711916);
DFFARX1 I_41718  ( .D(I458703), .CLK(I2702), .RSTB(I711786), .Q(I711950) );
not I_41719 (I711967,I711950);
nand I_41720 (I711766,I711950,I711916);
DFFARX1 I_41721  ( .D(I711950), .CLK(I2702), .RSTB(I711786), .Q(I711998) );
and I_41722 (I711751,I711837,I711998);
nand I_41723 (I712029,I458721,I458733);
and I_41724 (I712046,I712029,I458727);
DFFARX1 I_41725  ( .D(I712046), .CLK(I2702), .RSTB(I711786), .Q(I712063) );
nor I_41726 (I712080,I712063,I711967);
and I_41727 (I712097,I711899,I712080);
nor I_41728 (I712114,I712063,I711837);
DFFARX1 I_41729  ( .D(I712063), .CLK(I2702), .RSTB(I711786), .Q(I711757) );
DFFARX1 I_41730  ( .D(I458709), .CLK(I2702), .RSTB(I711786), .Q(I712145) );
and I_41731 (I712162,I712145,I458718);
or I_41732 (I712179,I712162,I712097);
DFFARX1 I_41733  ( .D(I712179), .CLK(I2702), .RSTB(I711786), .Q(I711769) );
nand I_41734 (I711778,I712162,I712114);
DFFARX1 I_41735  ( .D(I712162), .CLK(I2702), .RSTB(I711786), .Q(I711748) );
DFFARX1 I_41736  ( .D(I458730), .CLK(I2702), .RSTB(I711786), .Q(I712238) );
nand I_41737 (I711772,I712238,I711933);
DFFARX1 I_41738  ( .D(I712238), .CLK(I2702), .RSTB(I711786), .Q(I711760) );
nand I_41739 (I712283,I712238,I711899);
and I_41740 (I712300,I711950,I712283);
DFFARX1 I_41741  ( .D(I712300), .CLK(I2702), .RSTB(I711786), .Q(I711754) );
not I_41742 (I712364,I2709);
nand I_41743 (I712381,I75612,I75597);
and I_41744 (I712398,I712381,I75591);
DFFARX1 I_41745  ( .D(I712398), .CLK(I2702), .RSTB(I712364), .Q(I712415) );
not I_41746 (I712353,I712415);
DFFARX1 I_41747  ( .D(I712415), .CLK(I2702), .RSTB(I712364), .Q(I712446) );
not I_41748 (I712341,I712446);
nor I_41749 (I712477,I75618,I75597);
not I_41750 (I712494,I712477);
nor I_41751 (I712511,I712415,I712494);
DFFARX1 I_41752  ( .D(I75621), .CLK(I2702), .RSTB(I712364), .Q(I712528) );
not I_41753 (I712545,I712528);
nand I_41754 (I712344,I712528,I712494);
DFFARX1 I_41755  ( .D(I712528), .CLK(I2702), .RSTB(I712364), .Q(I712576) );
and I_41756 (I712329,I712415,I712576);
nand I_41757 (I712607,I75603,I75606);
and I_41758 (I712624,I712607,I75609);
DFFARX1 I_41759  ( .D(I712624), .CLK(I2702), .RSTB(I712364), .Q(I712641) );
nor I_41760 (I712658,I712641,I712545);
and I_41761 (I712675,I712477,I712658);
nor I_41762 (I712692,I712641,I712415);
DFFARX1 I_41763  ( .D(I712641), .CLK(I2702), .RSTB(I712364), .Q(I712335) );
DFFARX1 I_41764  ( .D(I75615), .CLK(I2702), .RSTB(I712364), .Q(I712723) );
and I_41765 (I712740,I712723,I75600);
or I_41766 (I712757,I712740,I712675);
DFFARX1 I_41767  ( .D(I712757), .CLK(I2702), .RSTB(I712364), .Q(I712347) );
nand I_41768 (I712356,I712740,I712692);
DFFARX1 I_41769  ( .D(I712740), .CLK(I2702), .RSTB(I712364), .Q(I712326) );
DFFARX1 I_41770  ( .D(I75594), .CLK(I2702), .RSTB(I712364), .Q(I712816) );
nand I_41771 (I712350,I712816,I712511);
DFFARX1 I_41772  ( .D(I712816), .CLK(I2702), .RSTB(I712364), .Q(I712338) );
nand I_41773 (I712861,I712816,I712477);
and I_41774 (I712878,I712528,I712861);
DFFARX1 I_41775  ( .D(I712878), .CLK(I2702), .RSTB(I712364), .Q(I712332) );
not I_41776 (I712942,I2709);
nand I_41777 (I712959,I252264,I252261);
and I_41778 (I712976,I712959,I252285);
DFFARX1 I_41779  ( .D(I712976), .CLK(I2702), .RSTB(I712942), .Q(I712993) );
not I_41780 (I712931,I712993);
DFFARX1 I_41781  ( .D(I712993), .CLK(I2702), .RSTB(I712942), .Q(I713024) );
not I_41782 (I712919,I713024);
nor I_41783 (I713055,I252267,I252261);
not I_41784 (I713072,I713055);
nor I_41785 (I713089,I712993,I713072);
DFFARX1 I_41786  ( .D(I252282), .CLK(I2702), .RSTB(I712942), .Q(I713106) );
not I_41787 (I713123,I713106);
nand I_41788 (I712922,I713106,I713072);
DFFARX1 I_41789  ( .D(I713106), .CLK(I2702), .RSTB(I712942), .Q(I713154) );
and I_41790 (I712907,I712993,I713154);
nand I_41791 (I713185,I252270,I252255);
and I_41792 (I713202,I713185,I252273);
DFFARX1 I_41793  ( .D(I713202), .CLK(I2702), .RSTB(I712942), .Q(I713219) );
nor I_41794 (I713236,I713219,I713123);
and I_41795 (I713253,I713055,I713236);
nor I_41796 (I713270,I713219,I712993);
DFFARX1 I_41797  ( .D(I713219), .CLK(I2702), .RSTB(I712942), .Q(I712913) );
DFFARX1 I_41798  ( .D(I252276), .CLK(I2702), .RSTB(I712942), .Q(I713301) );
and I_41799 (I713318,I713301,I252279);
or I_41800 (I713335,I713318,I713253);
DFFARX1 I_41801  ( .D(I713335), .CLK(I2702), .RSTB(I712942), .Q(I712925) );
nand I_41802 (I712934,I713318,I713270);
DFFARX1 I_41803  ( .D(I713318), .CLK(I2702), .RSTB(I712942), .Q(I712904) );
DFFARX1 I_41804  ( .D(I252258), .CLK(I2702), .RSTB(I712942), .Q(I713394) );
nand I_41805 (I712928,I713394,I713089);
DFFARX1 I_41806  ( .D(I713394), .CLK(I2702), .RSTB(I712942), .Q(I712916) );
nand I_41807 (I713439,I713394,I713055);
and I_41808 (I713456,I713106,I713439);
DFFARX1 I_41809  ( .D(I713456), .CLK(I2702), .RSTB(I712942), .Q(I712910) );
not I_41810 (I713520,I2709);
nand I_41811 (I713537,I472000,I472018);
and I_41812 (I713554,I713537,I472009);
DFFARX1 I_41813  ( .D(I713554), .CLK(I2702), .RSTB(I713520), .Q(I713571) );
not I_41814 (I713509,I713571);
DFFARX1 I_41815  ( .D(I713571), .CLK(I2702), .RSTB(I713520), .Q(I713602) );
not I_41816 (I713497,I713602);
nor I_41817 (I713633,I472006,I472018);
not I_41818 (I713650,I713633);
nor I_41819 (I713667,I713571,I713650);
DFFARX1 I_41820  ( .D(I471997), .CLK(I2702), .RSTB(I713520), .Q(I713684) );
not I_41821 (I713701,I713684);
nand I_41822 (I713500,I713684,I713650);
DFFARX1 I_41823  ( .D(I713684), .CLK(I2702), .RSTB(I713520), .Q(I713732) );
and I_41824 (I713485,I713571,I713732);
nand I_41825 (I713763,I472015,I472027);
and I_41826 (I713780,I713763,I472021);
DFFARX1 I_41827  ( .D(I713780), .CLK(I2702), .RSTB(I713520), .Q(I713797) );
nor I_41828 (I713814,I713797,I713701);
and I_41829 (I713831,I713633,I713814);
nor I_41830 (I713848,I713797,I713571);
DFFARX1 I_41831  ( .D(I713797), .CLK(I2702), .RSTB(I713520), .Q(I713491) );
DFFARX1 I_41832  ( .D(I472003), .CLK(I2702), .RSTB(I713520), .Q(I713879) );
and I_41833 (I713896,I713879,I472012);
or I_41834 (I713913,I713896,I713831);
DFFARX1 I_41835  ( .D(I713913), .CLK(I2702), .RSTB(I713520), .Q(I713503) );
nand I_41836 (I713512,I713896,I713848);
DFFARX1 I_41837  ( .D(I713896), .CLK(I2702), .RSTB(I713520), .Q(I713482) );
DFFARX1 I_41838  ( .D(I472024), .CLK(I2702), .RSTB(I713520), .Q(I713972) );
nand I_41839 (I713506,I713972,I713667);
DFFARX1 I_41840  ( .D(I713972), .CLK(I2702), .RSTB(I713520), .Q(I713494) );
nand I_41841 (I714017,I713972,I713633);
and I_41842 (I714034,I713684,I714017);
DFFARX1 I_41843  ( .D(I714034), .CLK(I2702), .RSTB(I713520), .Q(I713488) );
not I_41844 (I714098,I2709);
nand I_41845 (I714115,I567915,I567897);
and I_41846 (I714132,I714115,I567912);
DFFARX1 I_41847  ( .D(I714132), .CLK(I2702), .RSTB(I714098), .Q(I714149) );
not I_41848 (I714087,I714149);
DFFARX1 I_41849  ( .D(I714149), .CLK(I2702), .RSTB(I714098), .Q(I714180) );
not I_41850 (I714075,I714180);
nor I_41851 (I714211,I567903,I567897);
not I_41852 (I714228,I714211);
nor I_41853 (I714245,I714149,I714228);
DFFARX1 I_41854  ( .D(I567918), .CLK(I2702), .RSTB(I714098), .Q(I714262) );
not I_41855 (I714279,I714262);
nand I_41856 (I714078,I714262,I714228);
DFFARX1 I_41857  ( .D(I714262), .CLK(I2702), .RSTB(I714098), .Q(I714310) );
and I_41858 (I714063,I714149,I714310);
nand I_41859 (I714341,I567894,I567900);
and I_41860 (I714358,I714341,I567906);
DFFARX1 I_41861  ( .D(I714358), .CLK(I2702), .RSTB(I714098), .Q(I714375) );
nor I_41862 (I714392,I714375,I714279);
and I_41863 (I714409,I714211,I714392);
nor I_41864 (I714426,I714375,I714149);
DFFARX1 I_41865  ( .D(I714375), .CLK(I2702), .RSTB(I714098), .Q(I714069) );
DFFARX1 I_41866  ( .D(I567921), .CLK(I2702), .RSTB(I714098), .Q(I714457) );
and I_41867 (I714474,I714457,I567909);
or I_41868 (I714491,I714474,I714409);
DFFARX1 I_41869  ( .D(I714491), .CLK(I2702), .RSTB(I714098), .Q(I714081) );
nand I_41870 (I714090,I714474,I714426);
DFFARX1 I_41871  ( .D(I714474), .CLK(I2702), .RSTB(I714098), .Q(I714060) );
DFFARX1 I_41872  ( .D(I567924), .CLK(I2702), .RSTB(I714098), .Q(I714550) );
nand I_41873 (I714084,I714550,I714245);
DFFARX1 I_41874  ( .D(I714550), .CLK(I2702), .RSTB(I714098), .Q(I714072) );
nand I_41875 (I714595,I714550,I714211);
and I_41876 (I714612,I714262,I714595);
DFFARX1 I_41877  ( .D(I714612), .CLK(I2702), .RSTB(I714098), .Q(I714066) );
not I_41878 (I714676,I2709);
nand I_41879 (I714693,I311934,I311931);
and I_41880 (I714710,I714693,I311955);
DFFARX1 I_41881  ( .D(I714710), .CLK(I2702), .RSTB(I714676), .Q(I714727) );
not I_41882 (I714665,I714727);
DFFARX1 I_41883  ( .D(I714727), .CLK(I2702), .RSTB(I714676), .Q(I714758) );
not I_41884 (I714653,I714758);
nor I_41885 (I714789,I311937,I311931);
not I_41886 (I714806,I714789);
nor I_41887 (I714823,I714727,I714806);
DFFARX1 I_41888  ( .D(I311952), .CLK(I2702), .RSTB(I714676), .Q(I714840) );
not I_41889 (I714857,I714840);
nand I_41890 (I714656,I714840,I714806);
DFFARX1 I_41891  ( .D(I714840), .CLK(I2702), .RSTB(I714676), .Q(I714888) );
and I_41892 (I714641,I714727,I714888);
nand I_41893 (I714919,I311940,I311925);
and I_41894 (I714936,I714919,I311943);
DFFARX1 I_41895  ( .D(I714936), .CLK(I2702), .RSTB(I714676), .Q(I714953) );
nor I_41896 (I714970,I714953,I714857);
and I_41897 (I714987,I714789,I714970);
nor I_41898 (I715004,I714953,I714727);
DFFARX1 I_41899  ( .D(I714953), .CLK(I2702), .RSTB(I714676), .Q(I714647) );
DFFARX1 I_41900  ( .D(I311946), .CLK(I2702), .RSTB(I714676), .Q(I715035) );
and I_41901 (I715052,I715035,I311949);
or I_41902 (I715069,I715052,I714987);
DFFARX1 I_41903  ( .D(I715069), .CLK(I2702), .RSTB(I714676), .Q(I714659) );
nand I_41904 (I714668,I715052,I715004);
DFFARX1 I_41905  ( .D(I715052), .CLK(I2702), .RSTB(I714676), .Q(I714638) );
DFFARX1 I_41906  ( .D(I311928), .CLK(I2702), .RSTB(I714676), .Q(I715128) );
nand I_41907 (I714662,I715128,I714823);
DFFARX1 I_41908  ( .D(I715128), .CLK(I2702), .RSTB(I714676), .Q(I714650) );
nand I_41909 (I715173,I715128,I714789);
and I_41910 (I715190,I714840,I715173);
DFFARX1 I_41911  ( .D(I715190), .CLK(I2702), .RSTB(I714676), .Q(I714644) );
not I_41912 (I715254,I2709);
nand I_41913 (I715271,I181977,I182007);
and I_41914 (I715288,I715271,I181989);
DFFARX1 I_41915  ( .D(I715288), .CLK(I2702), .RSTB(I715254), .Q(I715305) );
not I_41916 (I715243,I715305);
DFFARX1 I_41917  ( .D(I715305), .CLK(I2702), .RSTB(I715254), .Q(I715336) );
not I_41918 (I715231,I715336);
nor I_41919 (I715367,I181986,I182007);
not I_41920 (I715384,I715367);
nor I_41921 (I715401,I715305,I715384);
DFFARX1 I_41922  ( .D(I181980), .CLK(I2702), .RSTB(I715254), .Q(I715418) );
not I_41923 (I715435,I715418);
nand I_41924 (I715234,I715418,I715384);
DFFARX1 I_41925  ( .D(I715418), .CLK(I2702), .RSTB(I715254), .Q(I715466) );
and I_41926 (I715219,I715305,I715466);
nand I_41927 (I715497,I181983,I181998);
and I_41928 (I715514,I715497,I181995);
DFFARX1 I_41929  ( .D(I715514), .CLK(I2702), .RSTB(I715254), .Q(I715531) );
nor I_41930 (I715548,I715531,I715435);
and I_41931 (I715565,I715367,I715548);
nor I_41932 (I715582,I715531,I715305);
DFFARX1 I_41933  ( .D(I715531), .CLK(I2702), .RSTB(I715254), .Q(I715225) );
DFFARX1 I_41934  ( .D(I181992), .CLK(I2702), .RSTB(I715254), .Q(I715613) );
and I_41935 (I715630,I715613,I182004);
or I_41936 (I715647,I715630,I715565);
DFFARX1 I_41937  ( .D(I715647), .CLK(I2702), .RSTB(I715254), .Q(I715237) );
nand I_41938 (I715246,I715630,I715582);
DFFARX1 I_41939  ( .D(I715630), .CLK(I2702), .RSTB(I715254), .Q(I715216) );
DFFARX1 I_41940  ( .D(I182001), .CLK(I2702), .RSTB(I715254), .Q(I715706) );
nand I_41941 (I715240,I715706,I715401);
DFFARX1 I_41942  ( .D(I715706), .CLK(I2702), .RSTB(I715254), .Q(I715228) );
nand I_41943 (I715751,I715706,I715367);
and I_41944 (I715768,I715418,I715751);
DFFARX1 I_41945  ( .D(I715768), .CLK(I2702), .RSTB(I715254), .Q(I715222) );
not I_41946 (I715832,I2709);
nand I_41947 (I715849,I8346,I8331);
and I_41948 (I715866,I715849,I8340);
DFFARX1 I_41949  ( .D(I715866), .CLK(I2702), .RSTB(I715832), .Q(I715883) );
not I_41950 (I715821,I715883);
DFFARX1 I_41951  ( .D(I715883), .CLK(I2702), .RSTB(I715832), .Q(I715914) );
not I_41952 (I715809,I715914);
nor I_41953 (I715945,I8352,I8331);
not I_41954 (I715962,I715945);
nor I_41955 (I715979,I715883,I715962);
DFFARX1 I_41956  ( .D(I8343), .CLK(I2702), .RSTB(I715832), .Q(I715996) );
not I_41957 (I716013,I715996);
nand I_41958 (I715812,I715996,I715962);
DFFARX1 I_41959  ( .D(I715996), .CLK(I2702), .RSTB(I715832), .Q(I716044) );
and I_41960 (I715797,I715883,I716044);
nand I_41961 (I716075,I8328,I8322);
and I_41962 (I716092,I716075,I8337);
DFFARX1 I_41963  ( .D(I716092), .CLK(I2702), .RSTB(I715832), .Q(I716109) );
nor I_41964 (I716126,I716109,I716013);
and I_41965 (I716143,I715945,I716126);
nor I_41966 (I716160,I716109,I715883);
DFFARX1 I_41967  ( .D(I716109), .CLK(I2702), .RSTB(I715832), .Q(I715803) );
DFFARX1 I_41968  ( .D(I8325), .CLK(I2702), .RSTB(I715832), .Q(I716191) );
and I_41969 (I716208,I716191,I8349);
or I_41970 (I716225,I716208,I716143);
DFFARX1 I_41971  ( .D(I716225), .CLK(I2702), .RSTB(I715832), .Q(I715815) );
nand I_41972 (I715824,I716208,I716160);
DFFARX1 I_41973  ( .D(I716208), .CLK(I2702), .RSTB(I715832), .Q(I715794) );
DFFARX1 I_41974  ( .D(I8334), .CLK(I2702), .RSTB(I715832), .Q(I716284) );
nand I_41975 (I715818,I716284,I715979);
DFFARX1 I_41976  ( .D(I716284), .CLK(I2702), .RSTB(I715832), .Q(I715806) );
nand I_41977 (I716329,I716284,I715945);
and I_41978 (I716346,I715996,I716329);
DFFARX1 I_41979  ( .D(I716346), .CLK(I2702), .RSTB(I715832), .Q(I715800) );
not I_41980 (I716410,I2709);
nand I_41981 (I716427,I234403,I234391);
and I_41982 (I716444,I716427,I234415);
DFFARX1 I_41983  ( .D(I716444), .CLK(I2702), .RSTB(I716410), .Q(I716461) );
not I_41984 (I716399,I716461);
DFFARX1 I_41985  ( .D(I716461), .CLK(I2702), .RSTB(I716410), .Q(I716492) );
not I_41986 (I716387,I716492);
nor I_41987 (I716523,I234409,I234391);
not I_41988 (I716540,I716523);
nor I_41989 (I716557,I716461,I716540);
DFFARX1 I_41990  ( .D(I234388), .CLK(I2702), .RSTB(I716410), .Q(I716574) );
not I_41991 (I716591,I716574);
nand I_41992 (I716390,I716574,I716540);
DFFARX1 I_41993  ( .D(I716574), .CLK(I2702), .RSTB(I716410), .Q(I716622) );
and I_41994 (I716375,I716461,I716622);
nand I_41995 (I716653,I234418,I234400);
and I_41996 (I716670,I716653,I234406);
DFFARX1 I_41997  ( .D(I716670), .CLK(I2702), .RSTB(I716410), .Q(I716687) );
nor I_41998 (I716704,I716687,I716591);
and I_41999 (I716721,I716523,I716704);
nor I_42000 (I716738,I716687,I716461);
DFFARX1 I_42001  ( .D(I716687), .CLK(I2702), .RSTB(I716410), .Q(I716381) );
DFFARX1 I_42002  ( .D(I234394), .CLK(I2702), .RSTB(I716410), .Q(I716769) );
and I_42003 (I716786,I716769,I234412);
or I_42004 (I716803,I716786,I716721);
DFFARX1 I_42005  ( .D(I716803), .CLK(I2702), .RSTB(I716410), .Q(I716393) );
nand I_42006 (I716402,I716786,I716738);
DFFARX1 I_42007  ( .D(I716786), .CLK(I2702), .RSTB(I716410), .Q(I716372) );
DFFARX1 I_42008  ( .D(I234397), .CLK(I2702), .RSTB(I716410), .Q(I716862) );
nand I_42009 (I716396,I716862,I716557);
DFFARX1 I_42010  ( .D(I716862), .CLK(I2702), .RSTB(I716410), .Q(I716384) );
nand I_42011 (I716907,I716862,I716523);
and I_42012 (I716924,I716574,I716907);
DFFARX1 I_42013  ( .D(I716924), .CLK(I2702), .RSTB(I716410), .Q(I716378) );
not I_42014 (I716988,I2709);
nand I_42015 (I717005,I344141,I344144);
and I_42016 (I717022,I717005,I344123);
DFFARX1 I_42017  ( .D(I717022), .CLK(I2702), .RSTB(I716988), .Q(I717039) );
not I_42018 (I716977,I717039);
DFFARX1 I_42019  ( .D(I717039), .CLK(I2702), .RSTB(I716988), .Q(I717070) );
not I_42020 (I716965,I717070);
nor I_42021 (I717101,I344138,I344144);
not I_42022 (I717118,I717101);
nor I_42023 (I717135,I717039,I717118);
DFFARX1 I_42024  ( .D(I344147), .CLK(I2702), .RSTB(I716988), .Q(I717152) );
not I_42025 (I717169,I717152);
nand I_42026 (I716968,I717152,I717118);
DFFARX1 I_42027  ( .D(I717152), .CLK(I2702), .RSTB(I716988), .Q(I717200) );
and I_42028 (I716953,I717039,I717200);
nand I_42029 (I717231,I344135,I344153);
and I_42030 (I717248,I717231,I344129);
DFFARX1 I_42031  ( .D(I717248), .CLK(I2702), .RSTB(I716988), .Q(I717265) );
nor I_42032 (I717282,I717265,I717169);
and I_42033 (I717299,I717101,I717282);
nor I_42034 (I717316,I717265,I717039);
DFFARX1 I_42035  ( .D(I717265), .CLK(I2702), .RSTB(I716988), .Q(I716959) );
DFFARX1 I_42036  ( .D(I344126), .CLK(I2702), .RSTB(I716988), .Q(I717347) );
and I_42037 (I717364,I717347,I344132);
or I_42038 (I717381,I717364,I717299);
DFFARX1 I_42039  ( .D(I717381), .CLK(I2702), .RSTB(I716988), .Q(I716971) );
nand I_42040 (I716980,I717364,I717316);
DFFARX1 I_42041  ( .D(I717364), .CLK(I2702), .RSTB(I716988), .Q(I716950) );
DFFARX1 I_42042  ( .D(I344150), .CLK(I2702), .RSTB(I716988), .Q(I717440) );
nand I_42043 (I716974,I717440,I717135);
DFFARX1 I_42044  ( .D(I717440), .CLK(I2702), .RSTB(I716988), .Q(I716962) );
nand I_42045 (I717485,I717440,I717101);
and I_42046 (I717502,I717152,I717485);
DFFARX1 I_42047  ( .D(I717502), .CLK(I2702), .RSTB(I716988), .Q(I716956) );
not I_42048 (I717566,I2709);
nand I_42049 (I717583,I387423,I387426);
and I_42050 (I717600,I717583,I387405);
DFFARX1 I_42051  ( .D(I717600), .CLK(I2702), .RSTB(I717566), .Q(I717617) );
not I_42052 (I717555,I717617);
DFFARX1 I_42053  ( .D(I717617), .CLK(I2702), .RSTB(I717566), .Q(I717648) );
not I_42054 (I717543,I717648);
nor I_42055 (I717679,I387420,I387426);
not I_42056 (I717696,I717679);
nor I_42057 (I717713,I717617,I717696);
DFFARX1 I_42058  ( .D(I387429), .CLK(I2702), .RSTB(I717566), .Q(I717730) );
not I_42059 (I717747,I717730);
nand I_42060 (I717546,I717730,I717696);
DFFARX1 I_42061  ( .D(I717730), .CLK(I2702), .RSTB(I717566), .Q(I717778) );
and I_42062 (I717531,I717617,I717778);
nand I_42063 (I717809,I387417,I387435);
and I_42064 (I717826,I717809,I387411);
DFFARX1 I_42065  ( .D(I717826), .CLK(I2702), .RSTB(I717566), .Q(I717843) );
nor I_42066 (I717860,I717843,I717747);
and I_42067 (I717877,I717679,I717860);
nor I_42068 (I717894,I717843,I717617);
DFFARX1 I_42069  ( .D(I717843), .CLK(I2702), .RSTB(I717566), .Q(I717537) );
DFFARX1 I_42070  ( .D(I387408), .CLK(I2702), .RSTB(I717566), .Q(I717925) );
and I_42071 (I717942,I717925,I387414);
or I_42072 (I717959,I717942,I717877);
DFFARX1 I_42073  ( .D(I717959), .CLK(I2702), .RSTB(I717566), .Q(I717549) );
nand I_42074 (I717558,I717942,I717894);
DFFARX1 I_42075  ( .D(I717942), .CLK(I2702), .RSTB(I717566), .Q(I717528) );
DFFARX1 I_42076  ( .D(I387432), .CLK(I2702), .RSTB(I717566), .Q(I718018) );
nand I_42077 (I717552,I718018,I717713);
DFFARX1 I_42078  ( .D(I718018), .CLK(I2702), .RSTB(I717566), .Q(I717540) );
nand I_42079 (I718063,I718018,I717679);
and I_42080 (I718080,I717730,I718063);
DFFARX1 I_42081  ( .D(I718080), .CLK(I2702), .RSTB(I717566), .Q(I717534) );
not I_42082 (I718144,I2709);
nand I_42083 (I718161,I65276,I65261);
and I_42084 (I718178,I718161,I65255);
DFFARX1 I_42085  ( .D(I718178), .CLK(I2702), .RSTB(I718144), .Q(I718195) );
not I_42086 (I718133,I718195);
DFFARX1 I_42087  ( .D(I718195), .CLK(I2702), .RSTB(I718144), .Q(I718226) );
not I_42088 (I718121,I718226);
nor I_42089 (I718257,I65282,I65261);
not I_42090 (I718274,I718257);
nor I_42091 (I718291,I718195,I718274);
DFFARX1 I_42092  ( .D(I65285), .CLK(I2702), .RSTB(I718144), .Q(I718308) );
not I_42093 (I718325,I718308);
nand I_42094 (I718124,I718308,I718274);
DFFARX1 I_42095  ( .D(I718308), .CLK(I2702), .RSTB(I718144), .Q(I718356) );
and I_42096 (I718109,I718195,I718356);
nand I_42097 (I718387,I65267,I65270);
and I_42098 (I718404,I718387,I65273);
DFFARX1 I_42099  ( .D(I718404), .CLK(I2702), .RSTB(I718144), .Q(I718421) );
nor I_42100 (I718438,I718421,I718325);
and I_42101 (I718455,I718257,I718438);
nor I_42102 (I718472,I718421,I718195);
DFFARX1 I_42103  ( .D(I718421), .CLK(I2702), .RSTB(I718144), .Q(I718115) );
DFFARX1 I_42104  ( .D(I65279), .CLK(I2702), .RSTB(I718144), .Q(I718503) );
and I_42105 (I718520,I718503,I65264);
or I_42106 (I718537,I718520,I718455);
DFFARX1 I_42107  ( .D(I718537), .CLK(I2702), .RSTB(I718144), .Q(I718127) );
nand I_42108 (I718136,I718520,I718472);
DFFARX1 I_42109  ( .D(I718520), .CLK(I2702), .RSTB(I718144), .Q(I718106) );
DFFARX1 I_42110  ( .D(I65258), .CLK(I2702), .RSTB(I718144), .Q(I718596) );
nand I_42111 (I718130,I718596,I718291);
DFFARX1 I_42112  ( .D(I718596), .CLK(I2702), .RSTB(I718144), .Q(I718118) );
nand I_42113 (I718641,I718596,I718257);
and I_42114 (I718658,I718308,I718641);
DFFARX1 I_42115  ( .D(I718658), .CLK(I2702), .RSTB(I718144), .Q(I718112) );
not I_42116 (I718722,I2709);
nand I_42117 (I718739,I192585,I192615);
and I_42118 (I718756,I718739,I192597);
DFFARX1 I_42119  ( .D(I718756), .CLK(I2702), .RSTB(I718722), .Q(I718773) );
not I_42120 (I718711,I718773);
DFFARX1 I_42121  ( .D(I718773), .CLK(I2702), .RSTB(I718722), .Q(I718804) );
not I_42122 (I718699,I718804);
nor I_42123 (I718835,I192594,I192615);
not I_42124 (I718852,I718835);
nor I_42125 (I718869,I718773,I718852);
DFFARX1 I_42126  ( .D(I192588), .CLK(I2702), .RSTB(I718722), .Q(I718886) );
not I_42127 (I718903,I718886);
nand I_42128 (I718702,I718886,I718852);
DFFARX1 I_42129  ( .D(I718886), .CLK(I2702), .RSTB(I718722), .Q(I718934) );
and I_42130 (I718687,I718773,I718934);
nand I_42131 (I718965,I192591,I192606);
and I_42132 (I718982,I718965,I192603);
DFFARX1 I_42133  ( .D(I718982), .CLK(I2702), .RSTB(I718722), .Q(I718999) );
nor I_42134 (I719016,I718999,I718903);
and I_42135 (I719033,I718835,I719016);
nor I_42136 (I719050,I718999,I718773);
DFFARX1 I_42137  ( .D(I718999), .CLK(I2702), .RSTB(I718722), .Q(I718693) );
DFFARX1 I_42138  ( .D(I192600), .CLK(I2702), .RSTB(I718722), .Q(I719081) );
and I_42139 (I719098,I719081,I192612);
or I_42140 (I719115,I719098,I719033);
DFFARX1 I_42141  ( .D(I719115), .CLK(I2702), .RSTB(I718722), .Q(I718705) );
nand I_42142 (I718714,I719098,I719050);
DFFARX1 I_42143  ( .D(I719098), .CLK(I2702), .RSTB(I718722), .Q(I718684) );
DFFARX1 I_42144  ( .D(I192609), .CLK(I2702), .RSTB(I718722), .Q(I719174) );
nand I_42145 (I718708,I719174,I718869);
DFFARX1 I_42146  ( .D(I719174), .CLK(I2702), .RSTB(I718722), .Q(I718696) );
nand I_42147 (I719219,I719174,I718835);
and I_42148 (I719236,I718886,I719219);
DFFARX1 I_42149  ( .D(I719236), .CLK(I2702), .RSTB(I718722), .Q(I718690) );
not I_42150 (I719300,I2709);
nand I_42151 (I719317,I1919,I2423);
and I_42152 (I719334,I719317,I2655);
DFFARX1 I_42153  ( .D(I719334), .CLK(I2702), .RSTB(I719300), .Q(I719351) );
not I_42154 (I719289,I719351);
DFFARX1 I_42155  ( .D(I719351), .CLK(I2702), .RSTB(I719300), .Q(I719382) );
not I_42156 (I719277,I719382);
nor I_42157 (I719413,I2095,I2423);
not I_42158 (I719430,I719413);
nor I_42159 (I719447,I719351,I719430);
DFFARX1 I_42160  ( .D(I2311), .CLK(I2702), .RSTB(I719300), .Q(I719464) );
not I_42161 (I719481,I719464);
nand I_42162 (I719280,I719464,I719430);
DFFARX1 I_42163  ( .D(I719464), .CLK(I2702), .RSTB(I719300), .Q(I719512) );
and I_42164 (I719265,I719351,I719512);
nand I_42165 (I719543,I2063,I2439);
and I_42166 (I719560,I719543,I1519);
DFFARX1 I_42167  ( .D(I719560), .CLK(I2702), .RSTB(I719300), .Q(I719577) );
nor I_42168 (I719594,I719577,I719481);
and I_42169 (I719611,I719413,I719594);
nor I_42170 (I719628,I719577,I719351);
DFFARX1 I_42171  ( .D(I719577), .CLK(I2702), .RSTB(I719300), .Q(I719271) );
DFFARX1 I_42172  ( .D(I1671), .CLK(I2702), .RSTB(I719300), .Q(I719659) );
and I_42173 (I719676,I719659,I1335);
or I_42174 (I719693,I719676,I719611);
DFFARX1 I_42175  ( .D(I719693), .CLK(I2702), .RSTB(I719300), .Q(I719283) );
nand I_42176 (I719292,I719676,I719628);
DFFARX1 I_42177  ( .D(I719676), .CLK(I2702), .RSTB(I719300), .Q(I719262) );
DFFARX1 I_42178  ( .D(I2335), .CLK(I2702), .RSTB(I719300), .Q(I719752) );
nand I_42179 (I719286,I719752,I719447);
DFFARX1 I_42180  ( .D(I719752), .CLK(I2702), .RSTB(I719300), .Q(I719274) );
nand I_42181 (I719797,I719752,I719413);
and I_42182 (I719814,I719464,I719797);
DFFARX1 I_42183  ( .D(I719814), .CLK(I2702), .RSTB(I719300), .Q(I719268) );
not I_42184 (I719878,I2709);
nand I_42185 (I719895,I658966,I658984);
and I_42186 (I719912,I719895,I658981);
DFFARX1 I_42187  ( .D(I719912), .CLK(I2702), .RSTB(I719878), .Q(I719929) );
not I_42188 (I719867,I719929);
DFFARX1 I_42189  ( .D(I719929), .CLK(I2702), .RSTB(I719878), .Q(I719960) );
not I_42190 (I719855,I719960);
nor I_42191 (I719991,I658987,I658984);
not I_42192 (I720008,I719991);
nor I_42193 (I720025,I719929,I720008);
DFFARX1 I_42194  ( .D(I658990), .CLK(I2702), .RSTB(I719878), .Q(I720042) );
not I_42195 (I720059,I720042);
nand I_42196 (I719858,I720042,I720008);
DFFARX1 I_42197  ( .D(I720042), .CLK(I2702), .RSTB(I719878), .Q(I720090) );
and I_42198 (I719843,I719929,I720090);
nand I_42199 (I720121,I658975,I658969);
and I_42200 (I720138,I720121,I658972);
DFFARX1 I_42201  ( .D(I720138), .CLK(I2702), .RSTB(I719878), .Q(I720155) );
nor I_42202 (I720172,I720155,I720059);
and I_42203 (I720189,I719991,I720172);
nor I_42204 (I720206,I720155,I719929);
DFFARX1 I_42205  ( .D(I720155), .CLK(I2702), .RSTB(I719878), .Q(I719849) );
DFFARX1 I_42206  ( .D(I658978), .CLK(I2702), .RSTB(I719878), .Q(I720237) );
and I_42207 (I720254,I720237,I658963);
or I_42208 (I720271,I720254,I720189);
DFFARX1 I_42209  ( .D(I720271), .CLK(I2702), .RSTB(I719878), .Q(I719861) );
nand I_42210 (I719870,I720254,I720206);
DFFARX1 I_42211  ( .D(I720254), .CLK(I2702), .RSTB(I719878), .Q(I719840) );
DFFARX1 I_42212  ( .D(I658993), .CLK(I2702), .RSTB(I719878), .Q(I720330) );
nand I_42213 (I719864,I720330,I720025);
DFFARX1 I_42214  ( .D(I720330), .CLK(I2702), .RSTB(I719878), .Q(I719852) );
nand I_42215 (I720375,I720330,I719991);
and I_42216 (I720392,I720042,I720375);
DFFARX1 I_42217  ( .D(I720392), .CLK(I2702), .RSTB(I719878), .Q(I719846) );
not I_42218 (I720456,I2709);
nand I_42219 (I720473,I655192,I655210);
and I_42220 (I720490,I720473,I655207);
DFFARX1 I_42221  ( .D(I720490), .CLK(I2702), .RSTB(I720456), .Q(I720507) );
not I_42222 (I720445,I720507);
DFFARX1 I_42223  ( .D(I720507), .CLK(I2702), .RSTB(I720456), .Q(I720538) );
not I_42224 (I720433,I720538);
nor I_42225 (I720569,I655213,I655210);
not I_42226 (I720586,I720569);
nor I_42227 (I720603,I720507,I720586);
DFFARX1 I_42228  ( .D(I655216), .CLK(I2702), .RSTB(I720456), .Q(I720620) );
not I_42229 (I720637,I720620);
nand I_42230 (I720436,I720620,I720586);
DFFARX1 I_42231  ( .D(I720620), .CLK(I2702), .RSTB(I720456), .Q(I720668) );
and I_42232 (I720421,I720507,I720668);
nand I_42233 (I720699,I655201,I655195);
and I_42234 (I720716,I720699,I655198);
DFFARX1 I_42235  ( .D(I720716), .CLK(I2702), .RSTB(I720456), .Q(I720733) );
nor I_42236 (I720750,I720733,I720637);
and I_42237 (I720767,I720569,I720750);
nor I_42238 (I720784,I720733,I720507);
DFFARX1 I_42239  ( .D(I720733), .CLK(I2702), .RSTB(I720456), .Q(I720427) );
DFFARX1 I_42240  ( .D(I655204), .CLK(I2702), .RSTB(I720456), .Q(I720815) );
and I_42241 (I720832,I720815,I655189);
or I_42242 (I720849,I720832,I720767);
DFFARX1 I_42243  ( .D(I720849), .CLK(I2702), .RSTB(I720456), .Q(I720439) );
nand I_42244 (I720448,I720832,I720784);
DFFARX1 I_42245  ( .D(I720832), .CLK(I2702), .RSTB(I720456), .Q(I720418) );
DFFARX1 I_42246  ( .D(I655219), .CLK(I2702), .RSTB(I720456), .Q(I720908) );
nand I_42247 (I720442,I720908,I720603);
DFFARX1 I_42248  ( .D(I720908), .CLK(I2702), .RSTB(I720456), .Q(I720430) );
nand I_42249 (I720953,I720908,I720569);
and I_42250 (I720970,I720620,I720953);
DFFARX1 I_42251  ( .D(I720970), .CLK(I2702), .RSTB(I720456), .Q(I720424) );
not I_42252 (I721034,I2709);
nand I_42253 (I721051,I146175,I146205);
and I_42254 (I721068,I721051,I146187);
DFFARX1 I_42255  ( .D(I721068), .CLK(I2702), .RSTB(I721034), .Q(I721085) );
not I_42256 (I721023,I721085);
DFFARX1 I_42257  ( .D(I721085), .CLK(I2702), .RSTB(I721034), .Q(I721116) );
not I_42258 (I721011,I721116);
nor I_42259 (I721147,I146184,I146205);
not I_42260 (I721164,I721147);
nor I_42261 (I721181,I721085,I721164);
DFFARX1 I_42262  ( .D(I146178), .CLK(I2702), .RSTB(I721034), .Q(I721198) );
not I_42263 (I721215,I721198);
nand I_42264 (I721014,I721198,I721164);
DFFARX1 I_42265  ( .D(I721198), .CLK(I2702), .RSTB(I721034), .Q(I721246) );
and I_42266 (I720999,I721085,I721246);
nand I_42267 (I721277,I146181,I146196);
and I_42268 (I721294,I721277,I146193);
DFFARX1 I_42269  ( .D(I721294), .CLK(I2702), .RSTB(I721034), .Q(I721311) );
nor I_42270 (I721328,I721311,I721215);
and I_42271 (I721345,I721147,I721328);
nor I_42272 (I721362,I721311,I721085);
DFFARX1 I_42273  ( .D(I721311), .CLK(I2702), .RSTB(I721034), .Q(I721005) );
DFFARX1 I_42274  ( .D(I146190), .CLK(I2702), .RSTB(I721034), .Q(I721393) );
and I_42275 (I721410,I721393,I146202);
or I_42276 (I721427,I721410,I721345);
DFFARX1 I_42277  ( .D(I721427), .CLK(I2702), .RSTB(I721034), .Q(I721017) );
nand I_42278 (I721026,I721410,I721362);
DFFARX1 I_42279  ( .D(I721410), .CLK(I2702), .RSTB(I721034), .Q(I720996) );
DFFARX1 I_42280  ( .D(I146199), .CLK(I2702), .RSTB(I721034), .Q(I721486) );
nand I_42281 (I721020,I721486,I721181);
DFFARX1 I_42282  ( .D(I721486), .CLK(I2702), .RSTB(I721034), .Q(I721008) );
nand I_42283 (I721531,I721486,I721147);
and I_42284 (I721548,I721198,I721531);
DFFARX1 I_42285  ( .D(I721548), .CLK(I2702), .RSTB(I721034), .Q(I721002) );
not I_42286 (I721612,I2709);
nand I_42287 (I721629,I60108,I60093);
and I_42288 (I721646,I721629,I60087);
DFFARX1 I_42289  ( .D(I721646), .CLK(I2702), .RSTB(I721612), .Q(I721663) );
not I_42290 (I721601,I721663);
DFFARX1 I_42291  ( .D(I721663), .CLK(I2702), .RSTB(I721612), .Q(I721694) );
not I_42292 (I721589,I721694);
nor I_42293 (I721725,I60114,I60093);
not I_42294 (I721742,I721725);
nor I_42295 (I721759,I721663,I721742);
DFFARX1 I_42296  ( .D(I60117), .CLK(I2702), .RSTB(I721612), .Q(I721776) );
not I_42297 (I721793,I721776);
nand I_42298 (I721592,I721776,I721742);
DFFARX1 I_42299  ( .D(I721776), .CLK(I2702), .RSTB(I721612), .Q(I721824) );
and I_42300 (I721577,I721663,I721824);
nand I_42301 (I721855,I60099,I60102);
and I_42302 (I721872,I721855,I60105);
DFFARX1 I_42303  ( .D(I721872), .CLK(I2702), .RSTB(I721612), .Q(I721889) );
nor I_42304 (I721906,I721889,I721793);
and I_42305 (I721923,I721725,I721906);
nor I_42306 (I721940,I721889,I721663);
DFFARX1 I_42307  ( .D(I721889), .CLK(I2702), .RSTB(I721612), .Q(I721583) );
DFFARX1 I_42308  ( .D(I60111), .CLK(I2702), .RSTB(I721612), .Q(I721971) );
and I_42309 (I721988,I721971,I60096);
or I_42310 (I722005,I721988,I721923);
DFFARX1 I_42311  ( .D(I722005), .CLK(I2702), .RSTB(I721612), .Q(I721595) );
nand I_42312 (I721604,I721988,I721940);
DFFARX1 I_42313  ( .D(I721988), .CLK(I2702), .RSTB(I721612), .Q(I721574) );
DFFARX1 I_42314  ( .D(I60090), .CLK(I2702), .RSTB(I721612), .Q(I722064) );
nand I_42315 (I721598,I722064,I721759);
DFFARX1 I_42316  ( .D(I722064), .CLK(I2702), .RSTB(I721612), .Q(I721586) );
nand I_42317 (I722109,I722064,I721725);
and I_42318 (I722126,I721776,I722109);
DFFARX1 I_42319  ( .D(I722126), .CLK(I2702), .RSTB(I721612), .Q(I721580) );
not I_42320 (I722190,I2709);
nand I_42321 (I722207,I89824,I89809);
and I_42322 (I722224,I722207,I89803);
DFFARX1 I_42323  ( .D(I722224), .CLK(I2702), .RSTB(I722190), .Q(I722241) );
not I_42324 (I722179,I722241);
DFFARX1 I_42325  ( .D(I722241), .CLK(I2702), .RSTB(I722190), .Q(I722272) );
not I_42326 (I722167,I722272);
nor I_42327 (I722303,I89830,I89809);
not I_42328 (I722320,I722303);
nor I_42329 (I722337,I722241,I722320);
DFFARX1 I_42330  ( .D(I89833), .CLK(I2702), .RSTB(I722190), .Q(I722354) );
not I_42331 (I722371,I722354);
nand I_42332 (I722170,I722354,I722320);
DFFARX1 I_42333  ( .D(I722354), .CLK(I2702), .RSTB(I722190), .Q(I722402) );
and I_42334 (I722155,I722241,I722402);
nand I_42335 (I722433,I89815,I89818);
and I_42336 (I722450,I722433,I89821);
DFFARX1 I_42337  ( .D(I722450), .CLK(I2702), .RSTB(I722190), .Q(I722467) );
nor I_42338 (I722484,I722467,I722371);
and I_42339 (I722501,I722303,I722484);
nor I_42340 (I722518,I722467,I722241);
DFFARX1 I_42341  ( .D(I722467), .CLK(I2702), .RSTB(I722190), .Q(I722161) );
DFFARX1 I_42342  ( .D(I89827), .CLK(I2702), .RSTB(I722190), .Q(I722549) );
and I_42343 (I722566,I722549,I89812);
or I_42344 (I722583,I722566,I722501);
DFFARX1 I_42345  ( .D(I722583), .CLK(I2702), .RSTB(I722190), .Q(I722173) );
nand I_42346 (I722182,I722566,I722518);
DFFARX1 I_42347  ( .D(I722566), .CLK(I2702), .RSTB(I722190), .Q(I722152) );
DFFARX1 I_42348  ( .D(I89806), .CLK(I2702), .RSTB(I722190), .Q(I722642) );
nand I_42349 (I722176,I722642,I722337);
DFFARX1 I_42350  ( .D(I722642), .CLK(I2702), .RSTB(I722190), .Q(I722164) );
nand I_42351 (I722687,I722642,I722303);
and I_42352 (I722704,I722354,I722687);
DFFARX1 I_42353  ( .D(I722704), .CLK(I2702), .RSTB(I722190), .Q(I722158) );
not I_42354 (I722768,I2709);
nand I_42355 (I722785,I381609,I381612);
and I_42356 (I722802,I722785,I381591);
DFFARX1 I_42357  ( .D(I722802), .CLK(I2702), .RSTB(I722768), .Q(I722819) );
not I_42358 (I722757,I722819);
DFFARX1 I_42359  ( .D(I722819), .CLK(I2702), .RSTB(I722768), .Q(I722850) );
not I_42360 (I722745,I722850);
nor I_42361 (I722881,I381606,I381612);
not I_42362 (I722898,I722881);
nor I_42363 (I722915,I722819,I722898);
DFFARX1 I_42364  ( .D(I381615), .CLK(I2702), .RSTB(I722768), .Q(I722932) );
not I_42365 (I722949,I722932);
nand I_42366 (I722748,I722932,I722898);
DFFARX1 I_42367  ( .D(I722932), .CLK(I2702), .RSTB(I722768), .Q(I722980) );
and I_42368 (I722733,I722819,I722980);
nand I_42369 (I723011,I381603,I381621);
and I_42370 (I723028,I723011,I381597);
DFFARX1 I_42371  ( .D(I723028), .CLK(I2702), .RSTB(I722768), .Q(I723045) );
nor I_42372 (I723062,I723045,I722949);
and I_42373 (I723079,I722881,I723062);
nor I_42374 (I723096,I723045,I722819);
DFFARX1 I_42375  ( .D(I723045), .CLK(I2702), .RSTB(I722768), .Q(I722739) );
DFFARX1 I_42376  ( .D(I381594), .CLK(I2702), .RSTB(I722768), .Q(I723127) );
and I_42377 (I723144,I723127,I381600);
or I_42378 (I723161,I723144,I723079);
DFFARX1 I_42379  ( .D(I723161), .CLK(I2702), .RSTB(I722768), .Q(I722751) );
nand I_42380 (I722760,I723144,I723096);
DFFARX1 I_42381  ( .D(I723144), .CLK(I2702), .RSTB(I722768), .Q(I722730) );
DFFARX1 I_42382  ( .D(I381618), .CLK(I2702), .RSTB(I722768), .Q(I723220) );
nand I_42383 (I722754,I723220,I722915);
DFFARX1 I_42384  ( .D(I723220), .CLK(I2702), .RSTB(I722768), .Q(I722742) );
nand I_42385 (I723265,I723220,I722881);
and I_42386 (I723282,I722932,I723265);
DFFARX1 I_42387  ( .D(I723282), .CLK(I2702), .RSTB(I722768), .Q(I722736) );
not I_42388 (I723346,I2709);
nand I_42389 (I723363,I16761,I16746);
and I_42390 (I723380,I723363,I16755);
DFFARX1 I_42391  ( .D(I723380), .CLK(I2702), .RSTB(I723346), .Q(I723397) );
not I_42392 (I723335,I723397);
DFFARX1 I_42393  ( .D(I723397), .CLK(I2702), .RSTB(I723346), .Q(I723428) );
not I_42394 (I723323,I723428);
nor I_42395 (I723459,I16767,I16746);
not I_42396 (I723476,I723459);
nor I_42397 (I723493,I723397,I723476);
DFFARX1 I_42398  ( .D(I16758), .CLK(I2702), .RSTB(I723346), .Q(I723510) );
not I_42399 (I723527,I723510);
nand I_42400 (I723326,I723510,I723476);
DFFARX1 I_42401  ( .D(I723510), .CLK(I2702), .RSTB(I723346), .Q(I723558) );
and I_42402 (I723311,I723397,I723558);
nand I_42403 (I723589,I16743,I16737);
and I_42404 (I723606,I723589,I16752);
DFFARX1 I_42405  ( .D(I723606), .CLK(I2702), .RSTB(I723346), .Q(I723623) );
nor I_42406 (I723640,I723623,I723527);
and I_42407 (I723657,I723459,I723640);
nor I_42408 (I723674,I723623,I723397);
DFFARX1 I_42409  ( .D(I723623), .CLK(I2702), .RSTB(I723346), .Q(I723317) );
DFFARX1 I_42410  ( .D(I16740), .CLK(I2702), .RSTB(I723346), .Q(I723705) );
and I_42411 (I723722,I723705,I16764);
or I_42412 (I723739,I723722,I723657);
DFFARX1 I_42413  ( .D(I723739), .CLK(I2702), .RSTB(I723346), .Q(I723329) );
nand I_42414 (I723338,I723722,I723674);
DFFARX1 I_42415  ( .D(I723722), .CLK(I2702), .RSTB(I723346), .Q(I723308) );
DFFARX1 I_42416  ( .D(I16749), .CLK(I2702), .RSTB(I723346), .Q(I723798) );
nand I_42417 (I723332,I723798,I723493);
DFFARX1 I_42418  ( .D(I723798), .CLK(I2702), .RSTB(I723346), .Q(I723320) );
nand I_42419 (I723843,I723798,I723459);
and I_42420 (I723860,I723510,I723843);
DFFARX1 I_42421  ( .D(I723860), .CLK(I2702), .RSTB(I723346), .Q(I723314) );
not I_42422 (I723924,I2709);
nand I_42423 (I723941,I499082,I499088);
and I_42424 (I723958,I723941,I499067);
DFFARX1 I_42425  ( .D(I723958), .CLK(I2702), .RSTB(I723924), .Q(I723975) );
not I_42426 (I723913,I723975);
DFFARX1 I_42427  ( .D(I723975), .CLK(I2702), .RSTB(I723924), .Q(I724006) );
not I_42428 (I723901,I724006);
nor I_42429 (I724037,I499070,I499088);
not I_42430 (I724054,I724037);
nor I_42431 (I724071,I723975,I724054);
DFFARX1 I_42432  ( .D(I499064), .CLK(I2702), .RSTB(I723924), .Q(I724088) );
not I_42433 (I724105,I724088);
nand I_42434 (I723904,I724088,I724054);
DFFARX1 I_42435  ( .D(I724088), .CLK(I2702), .RSTB(I723924), .Q(I724136) );
and I_42436 (I723889,I723975,I724136);
nand I_42437 (I724167,I499061,I499076);
and I_42438 (I724184,I724167,I499085);
DFFARX1 I_42439  ( .D(I724184), .CLK(I2702), .RSTB(I723924), .Q(I724201) );
nor I_42440 (I724218,I724201,I724105);
and I_42441 (I724235,I724037,I724218);
nor I_42442 (I724252,I724201,I723975);
DFFARX1 I_42443  ( .D(I724201), .CLK(I2702), .RSTB(I723924), .Q(I723895) );
DFFARX1 I_42444  ( .D(I499091), .CLK(I2702), .RSTB(I723924), .Q(I724283) );
and I_42445 (I724300,I724283,I499073);
or I_42446 (I724317,I724300,I724235);
DFFARX1 I_42447  ( .D(I724317), .CLK(I2702), .RSTB(I723924), .Q(I723907) );
nand I_42448 (I723916,I724300,I724252);
DFFARX1 I_42449  ( .D(I724300), .CLK(I2702), .RSTB(I723924), .Q(I723886) );
DFFARX1 I_42450  ( .D(I499079), .CLK(I2702), .RSTB(I723924), .Q(I724376) );
nand I_42451 (I723910,I724376,I724071);
DFFARX1 I_42452  ( .D(I724376), .CLK(I2702), .RSTB(I723924), .Q(I723898) );
nand I_42453 (I724421,I724376,I724037);
and I_42454 (I724438,I724088,I724421);
DFFARX1 I_42455  ( .D(I724438), .CLK(I2702), .RSTB(I723924), .Q(I723892) );
not I_42456 (I724502,I2709);
nand I_42457 (I724519,I33030,I33015);
and I_42458 (I724536,I724519,I33024);
DFFARX1 I_42459  ( .D(I724536), .CLK(I2702), .RSTB(I724502), .Q(I724553) );
not I_42460 (I724491,I724553);
DFFARX1 I_42461  ( .D(I724553), .CLK(I2702), .RSTB(I724502), .Q(I724584) );
not I_42462 (I724479,I724584);
nor I_42463 (I724615,I33036,I33015);
not I_42464 (I724632,I724615);
nor I_42465 (I724649,I724553,I724632);
DFFARX1 I_42466  ( .D(I33027), .CLK(I2702), .RSTB(I724502), .Q(I724666) );
not I_42467 (I724683,I724666);
nand I_42468 (I724482,I724666,I724632);
DFFARX1 I_42469  ( .D(I724666), .CLK(I2702), .RSTB(I724502), .Q(I724714) );
and I_42470 (I724467,I724553,I724714);
nand I_42471 (I724745,I33012,I33006);
and I_42472 (I724762,I724745,I33021);
DFFARX1 I_42473  ( .D(I724762), .CLK(I2702), .RSTB(I724502), .Q(I724779) );
nor I_42474 (I724796,I724779,I724683);
and I_42475 (I724813,I724615,I724796);
nor I_42476 (I724830,I724779,I724553);
DFFARX1 I_42477  ( .D(I724779), .CLK(I2702), .RSTB(I724502), .Q(I724473) );
DFFARX1 I_42478  ( .D(I33009), .CLK(I2702), .RSTB(I724502), .Q(I724861) );
and I_42479 (I724878,I724861,I33033);
or I_42480 (I724895,I724878,I724813);
DFFARX1 I_42481  ( .D(I724895), .CLK(I2702), .RSTB(I724502), .Q(I724485) );
nand I_42482 (I724494,I724878,I724830);
DFFARX1 I_42483  ( .D(I724878), .CLK(I2702), .RSTB(I724502), .Q(I724464) );
DFFARX1 I_42484  ( .D(I33018), .CLK(I2702), .RSTB(I724502), .Q(I724954) );
nand I_42485 (I724488,I724954,I724649);
DFFARX1 I_42486  ( .D(I724954), .CLK(I2702), .RSTB(I724502), .Q(I724476) );
nand I_42487 (I724999,I724954,I724615);
and I_42488 (I725016,I724666,I724999);
DFFARX1 I_42489  ( .D(I725016), .CLK(I2702), .RSTB(I724502), .Q(I724470) );
not I_42490 (I725080,I2709);
nand I_42491 (I725097,I41445,I41430);
and I_42492 (I725114,I725097,I41439);
DFFARX1 I_42493  ( .D(I725114), .CLK(I2702), .RSTB(I725080), .Q(I725131) );
not I_42494 (I725069,I725131);
DFFARX1 I_42495  ( .D(I725131), .CLK(I2702), .RSTB(I725080), .Q(I725162) );
not I_42496 (I725057,I725162);
nor I_42497 (I725193,I41451,I41430);
not I_42498 (I725210,I725193);
nor I_42499 (I725227,I725131,I725210);
DFFARX1 I_42500  ( .D(I41442), .CLK(I2702), .RSTB(I725080), .Q(I725244) );
not I_42501 (I725261,I725244);
nand I_42502 (I725060,I725244,I725210);
DFFARX1 I_42503  ( .D(I725244), .CLK(I2702), .RSTB(I725080), .Q(I725292) );
and I_42504 (I725045,I725131,I725292);
nand I_42505 (I725323,I41427,I41421);
and I_42506 (I725340,I725323,I41436);
DFFARX1 I_42507  ( .D(I725340), .CLK(I2702), .RSTB(I725080), .Q(I725357) );
nor I_42508 (I725374,I725357,I725261);
and I_42509 (I725391,I725193,I725374);
nor I_42510 (I725408,I725357,I725131);
DFFARX1 I_42511  ( .D(I725357), .CLK(I2702), .RSTB(I725080), .Q(I725051) );
DFFARX1 I_42512  ( .D(I41424), .CLK(I2702), .RSTB(I725080), .Q(I725439) );
and I_42513 (I725456,I725439,I41448);
or I_42514 (I725473,I725456,I725391);
DFFARX1 I_42515  ( .D(I725473), .CLK(I2702), .RSTB(I725080), .Q(I725063) );
nand I_42516 (I725072,I725456,I725408);
DFFARX1 I_42517  ( .D(I725456), .CLK(I2702), .RSTB(I725080), .Q(I725042) );
DFFARX1 I_42518  ( .D(I41433), .CLK(I2702), .RSTB(I725080), .Q(I725532) );
nand I_42519 (I725066,I725532,I725227);
DFFARX1 I_42520  ( .D(I725532), .CLK(I2702), .RSTB(I725080), .Q(I725054) );
nand I_42521 (I725577,I725532,I725193);
and I_42522 (I725594,I725244,I725577);
DFFARX1 I_42523  ( .D(I725594), .CLK(I2702), .RSTB(I725080), .Q(I725048) );
not I_42524 (I725658,I2709);
nand I_42525 (I725675,I641354,I641372);
and I_42526 (I725692,I725675,I641369);
DFFARX1 I_42527  ( .D(I725692), .CLK(I2702), .RSTB(I725658), .Q(I725709) );
not I_42528 (I725647,I725709);
DFFARX1 I_42529  ( .D(I725709), .CLK(I2702), .RSTB(I725658), .Q(I725740) );
not I_42530 (I725635,I725740);
nor I_42531 (I725771,I641375,I641372);
not I_42532 (I725788,I725771);
nor I_42533 (I725805,I725709,I725788);
DFFARX1 I_42534  ( .D(I641378), .CLK(I2702), .RSTB(I725658), .Q(I725822) );
not I_42535 (I725839,I725822);
nand I_42536 (I725638,I725822,I725788);
DFFARX1 I_42537  ( .D(I725822), .CLK(I2702), .RSTB(I725658), .Q(I725870) );
and I_42538 (I725623,I725709,I725870);
nand I_42539 (I725901,I641363,I641357);
and I_42540 (I725918,I725901,I641360);
DFFARX1 I_42541  ( .D(I725918), .CLK(I2702), .RSTB(I725658), .Q(I725935) );
nor I_42542 (I725952,I725935,I725839);
and I_42543 (I725969,I725771,I725952);
nor I_42544 (I725986,I725935,I725709);
DFFARX1 I_42545  ( .D(I725935), .CLK(I2702), .RSTB(I725658), .Q(I725629) );
DFFARX1 I_42546  ( .D(I641366), .CLK(I2702), .RSTB(I725658), .Q(I726017) );
and I_42547 (I726034,I726017,I641351);
or I_42548 (I726051,I726034,I725969);
DFFARX1 I_42549  ( .D(I726051), .CLK(I2702), .RSTB(I725658), .Q(I725641) );
nand I_42550 (I725650,I726034,I725986);
DFFARX1 I_42551  ( .D(I726034), .CLK(I2702), .RSTB(I725658), .Q(I725620) );
DFFARX1 I_42552  ( .D(I641381), .CLK(I2702), .RSTB(I725658), .Q(I726110) );
nand I_42553 (I725644,I726110,I725805);
DFFARX1 I_42554  ( .D(I726110), .CLK(I2702), .RSTB(I725658), .Q(I725632) );
nand I_42555 (I726155,I726110,I725771);
and I_42556 (I726172,I725822,I726155);
DFFARX1 I_42557  ( .D(I726172), .CLK(I2702), .RSTB(I725658), .Q(I725626) );
not I_42558 (I726236,I2709);
nand I_42559 (I726253,I325857,I325854);
and I_42560 (I726270,I726253,I325878);
DFFARX1 I_42561  ( .D(I726270), .CLK(I2702), .RSTB(I726236), .Q(I726287) );
not I_42562 (I726225,I726287);
DFFARX1 I_42563  ( .D(I726287), .CLK(I2702), .RSTB(I726236), .Q(I726318) );
not I_42564 (I726213,I726318);
nor I_42565 (I726349,I325860,I325854);
not I_42566 (I726366,I726349);
nor I_42567 (I726383,I726287,I726366);
DFFARX1 I_42568  ( .D(I325875), .CLK(I2702), .RSTB(I726236), .Q(I726400) );
not I_42569 (I726417,I726400);
nand I_42570 (I726216,I726400,I726366);
DFFARX1 I_42571  ( .D(I726400), .CLK(I2702), .RSTB(I726236), .Q(I726448) );
and I_42572 (I726201,I726287,I726448);
nand I_42573 (I726479,I325863,I325848);
and I_42574 (I726496,I726479,I325866);
DFFARX1 I_42575  ( .D(I726496), .CLK(I2702), .RSTB(I726236), .Q(I726513) );
nor I_42576 (I726530,I726513,I726417);
and I_42577 (I726547,I726349,I726530);
nor I_42578 (I726564,I726513,I726287);
DFFARX1 I_42579  ( .D(I726513), .CLK(I2702), .RSTB(I726236), .Q(I726207) );
DFFARX1 I_42580  ( .D(I325869), .CLK(I2702), .RSTB(I726236), .Q(I726595) );
and I_42581 (I726612,I726595,I325872);
or I_42582 (I726629,I726612,I726547);
DFFARX1 I_42583  ( .D(I726629), .CLK(I2702), .RSTB(I726236), .Q(I726219) );
nand I_42584 (I726228,I726612,I726564);
DFFARX1 I_42585  ( .D(I726612), .CLK(I2702), .RSTB(I726236), .Q(I726198) );
DFFARX1 I_42586  ( .D(I325851), .CLK(I2702), .RSTB(I726236), .Q(I726688) );
nand I_42587 (I726222,I726688,I726383);
DFFARX1 I_42588  ( .D(I726688), .CLK(I2702), .RSTB(I726236), .Q(I726210) );
nand I_42589 (I726733,I726688,I726349);
and I_42590 (I726750,I726400,I726733);
DFFARX1 I_42591  ( .D(I726750), .CLK(I2702), .RSTB(I726236), .Q(I726204) );
not I_42592 (I726814,I2709);
nand I_42593 (I726831,I673433,I673451);
and I_42594 (I726848,I726831,I673448);
DFFARX1 I_42595  ( .D(I726848), .CLK(I2702), .RSTB(I726814), .Q(I726865) );
not I_42596 (I726803,I726865);
DFFARX1 I_42597  ( .D(I726865), .CLK(I2702), .RSTB(I726814), .Q(I726896) );
not I_42598 (I726791,I726896);
nor I_42599 (I726927,I673454,I673451);
not I_42600 (I726944,I726927);
nor I_42601 (I726961,I726865,I726944);
DFFARX1 I_42602  ( .D(I673457), .CLK(I2702), .RSTB(I726814), .Q(I726978) );
not I_42603 (I726995,I726978);
nand I_42604 (I726794,I726978,I726944);
DFFARX1 I_42605  ( .D(I726978), .CLK(I2702), .RSTB(I726814), .Q(I727026) );
and I_42606 (I726779,I726865,I727026);
nand I_42607 (I727057,I673442,I673436);
and I_42608 (I727074,I727057,I673439);
DFFARX1 I_42609  ( .D(I727074), .CLK(I2702), .RSTB(I726814), .Q(I727091) );
nor I_42610 (I727108,I727091,I726995);
and I_42611 (I727125,I726927,I727108);
nor I_42612 (I727142,I727091,I726865);
DFFARX1 I_42613  ( .D(I727091), .CLK(I2702), .RSTB(I726814), .Q(I726785) );
DFFARX1 I_42614  ( .D(I673445), .CLK(I2702), .RSTB(I726814), .Q(I727173) );
and I_42615 (I727190,I727173,I673430);
or I_42616 (I727207,I727190,I727125);
DFFARX1 I_42617  ( .D(I727207), .CLK(I2702), .RSTB(I726814), .Q(I726797) );
nand I_42618 (I726806,I727190,I727142);
DFFARX1 I_42619  ( .D(I727190), .CLK(I2702), .RSTB(I726814), .Q(I726776) );
DFFARX1 I_42620  ( .D(I673460), .CLK(I2702), .RSTB(I726814), .Q(I727266) );
nand I_42621 (I726800,I727266,I726961);
DFFARX1 I_42622  ( .D(I727266), .CLK(I2702), .RSTB(I726814), .Q(I726788) );
nand I_42623 (I727311,I727266,I726927);
and I_42624 (I727328,I726978,I727311);
DFFARX1 I_42625  ( .D(I727328), .CLK(I2702), .RSTB(I726814), .Q(I726782) );
not I_42626 (I727392,I2709);
nand I_42627 (I727409,I267513,I267510);
and I_42628 (I727426,I727409,I267534);
DFFARX1 I_42629  ( .D(I727426), .CLK(I2702), .RSTB(I727392), .Q(I727443) );
not I_42630 (I727381,I727443);
DFFARX1 I_42631  ( .D(I727443), .CLK(I2702), .RSTB(I727392), .Q(I727474) );
not I_42632 (I727369,I727474);
nor I_42633 (I727505,I267516,I267510);
not I_42634 (I727522,I727505);
nor I_42635 (I727539,I727443,I727522);
DFFARX1 I_42636  ( .D(I267531), .CLK(I2702), .RSTB(I727392), .Q(I727556) );
not I_42637 (I727573,I727556);
nand I_42638 (I727372,I727556,I727522);
DFFARX1 I_42639  ( .D(I727556), .CLK(I2702), .RSTB(I727392), .Q(I727604) );
and I_42640 (I727357,I727443,I727604);
nand I_42641 (I727635,I267519,I267504);
and I_42642 (I727652,I727635,I267522);
DFFARX1 I_42643  ( .D(I727652), .CLK(I2702), .RSTB(I727392), .Q(I727669) );
nor I_42644 (I727686,I727669,I727573);
and I_42645 (I727703,I727505,I727686);
nor I_42646 (I727720,I727669,I727443);
DFFARX1 I_42647  ( .D(I727669), .CLK(I2702), .RSTB(I727392), .Q(I727363) );
DFFARX1 I_42648  ( .D(I267525), .CLK(I2702), .RSTB(I727392), .Q(I727751) );
and I_42649 (I727768,I727751,I267528);
or I_42650 (I727785,I727768,I727703);
DFFARX1 I_42651  ( .D(I727785), .CLK(I2702), .RSTB(I727392), .Q(I727375) );
nand I_42652 (I727384,I727768,I727720);
DFFARX1 I_42653  ( .D(I727768), .CLK(I2702), .RSTB(I727392), .Q(I727354) );
DFFARX1 I_42654  ( .D(I267507), .CLK(I2702), .RSTB(I727392), .Q(I727844) );
nand I_42655 (I727378,I727844,I727539);
DFFARX1 I_42656  ( .D(I727844), .CLK(I2702), .RSTB(I727392), .Q(I727366) );
nand I_42657 (I727889,I727844,I727505);
and I_42658 (I727906,I727556,I727889);
DFFARX1 I_42659  ( .D(I727906), .CLK(I2702), .RSTB(I727392), .Q(I727360) );
endmodule


