module test_I9459(I9672,I1477,I1470,I8315,I9459);
input I9672,I1477,I1470,I8315;
output I9459;
wire I8187,I8216,I8753,I9720,I9754,I9771,I9737,I8178,I8205,I9621,I9689,I8736,I9491;
DFFARX1 I_0(I8315,I1470,I8216,,,I8187,);
not I_1(I8216,I1477);
not I_2(I8753,I8736);
not I_3(I9720,I9689);
DFFARX1 I_4(I8187,I1470,I9491,,,I9754,);
and I_5(I9771,I9754,I8178);
nor I_6(I9737,I9621,I9720);
nand I_7(I9459,I9771,I9737);
DFFARX1 I_8(I8753,I1470,I8216,,,I8178,);
not I_9(I8205,I8315);
DFFARX1 I_10(I8205,I1470,I9491,,,I9621,);
DFFARX1 I_11(I9672,I1470,I9491,,,I9689,);
DFFARX1 I_12(I1470,I8216,,,I8736,);
not I_13(I9491,I1477);
endmodule


