module test_final(IN_1_0_l_6,IN_2_0_l_6,IN_3_0_l_6,IN_4_0_l_6,IN_1_1_l_6,IN_2_1_l_6,IN_3_1_l_6,IN_1_10_l_6,IN_2_10_l_6,IN_3_10_l_6,IN_4_10_l_6,blif_clk_net_8_r_1,blif_reset_net_8_r_1,N6147_3_r_1,N1372_4_r_1,N1508_4_r_1,n_42_8_r_1,G199_8_r_1,N6147_9_r_1,N6134_9_r_1,N1372_10_r_1,N1508_10_r_1);
input IN_1_0_l_6,IN_2_0_l_6,IN_3_0_l_6,IN_4_0_l_6,IN_1_1_l_6,IN_2_1_l_6,IN_3_1_l_6,IN_1_10_l_6,IN_2_10_l_6,IN_3_10_l_6,IN_4_10_l_6,blif_clk_net_8_r_1,blif_reset_net_8_r_1;
output N6147_3_r_1,N1372_4_r_1,N1508_4_r_1,n_42_8_r_1,G199_8_r_1,N6147_9_r_1,N6134_9_r_1,N1372_10_r_1,N1508_10_r_1;
wire N1371_0_r_6,N1508_0_r_6,N6147_3_r_6,n_429_or_0_5_r_6,G78_5_r_6,n_576_5_r_6,n_102_5_r_6,n_547_5_r_6,N1372_10_r_6,N1508_10_r_6,n_431_5_r_6,n24_6,n25_6,n26_6,n27_6,n28_6,n29_6,n30_6,n31_6,n32_6,n33_6,n34_6,n35_6,n36_6,n37_6,n38_6,n39_6,n40_6,n41_6,n42_6,I_BUFF_1_9_r_1,N3_8_l_1,n7_1,n38_1,n22_1,N3_8_r_1,n23_1,n24_1,n25_1,n26_1,n27_1,n28_1,n29_1,n30_1,n31_1,n32_1,n33_1,n34_1,n35_1,n36_1,n37_1;
nor I_0(N1371_0_r_6,n26_6,n38_6);
not I_1(N1508_0_r_6,n38_6);
nor I_2(N6147_3_r_6,n30_6,n35_6);
nand I_3(n_429_or_0_5_r_6,n30_6,n32_6);
DFFARX1 I_4(n_431_5_r_6,blif_clk_net_8_r_1,n7_1,G78_5_r_6,);
nand I_5(n_576_5_r_6,n24_6,n25_6);
not I_6(n_102_5_r_6,n26_6);
or I_7(n_547_5_r_6,n_429_or_0_5_r_6,n26_6);
not I_8(N1372_10_r_6,n37_6);
nor I_9(N1508_10_r_6,n36_6,n37_6);
nand I_10(n_431_5_r_6,n_102_5_r_6,n28_6);
nor I_11(n24_6,n33_6,n34_6);
nor I_12(n25_6,n26_6,n27_6);
nor I_13(n26_6,IN_2_0_l_6,n40_6);
nand I_14(n27_6,IN_1_1_l_6,IN_2_1_l_6);
nand I_15(n28_6,n29_6,n30_6);
nor I_16(n29_6,IN_3_1_l_6,n31_6);
not I_17(n30_6,n27_6);
nor I_18(n31_6,n39_6,n40_6);
nor I_19(n32_6,IN_3_1_l_6,n24_6);
not I_20(n33_6,IN_1_10_l_6);
not I_21(n34_6,IN_2_10_l_6);
or I_22(n35_6,n26_6,n31_6);
and I_23(n36_6,IN_3_1_l_6,n38_6);
nand I_24(n37_6,n30_6,n31_6);
nand I_25(n38_6,IN_2_10_l_6,n41_6);
nor I_26(n39_6,IN_3_0_l_6,IN_4_0_l_6);
not I_27(n40_6,IN_1_0_l_6);
nor I_28(n41_6,n33_6,n42_6);
nor I_29(n42_6,IN_3_10_l_6,IN_4_10_l_6);
nor I_30(N6147_3_r_1,n26_1,n27_1);
not I_31(N1372_4_r_1,n34_1);
nor I_32(N1508_4_r_1,n30_1,n34_1);
nor I_33(n_42_8_r_1,n23_1,n24_1);
DFFARX1 I_34(N3_8_r_1,blif_clk_net_8_r_1,n7_1,G199_8_r_1,);
nor I_35(N6147_9_r_1,n22_1,n25_1);
nor I_36(N6134_9_r_1,n29_1,n30_1);
not I_37(I_BUFF_1_9_r_1,n32_1);
not I_38(N1372_10_r_1,n36_1);
nor I_39(N1508_10_r_1,n35_1,n36_1);
and I_40(N3_8_l_1,n33_1,N1508_10_r_6);
not I_41(n7_1,blif_reset_net_8_r_1);
DFFARX1 I_42(N3_8_l_1,blif_clk_net_8_r_1,n7_1,n38_1,);
not I_43(n22_1,n38_1);
nor I_44(N3_8_r_1,n31_1,n32_1);
nor I_45(n23_1,n28_1,N1371_0_r_6);
nor I_46(n24_1,n_576_5_r_6,N1372_10_r_6);
nor I_47(n25_1,n23_1,n26_1);
not I_48(n26_1,n30_1);
nand I_49(n27_1,n22_1,n28_1);
nand I_50(n28_1,N1508_0_r_6,N6147_3_r_6);
not I_51(n29_1,n28_1);
nand I_52(n30_1,N1371_0_r_6,N1508_0_r_6);
and I_53(n31_1,n38_1,n24_1);
nand I_54(n32_1,n26_1,n37_1);
nand I_55(n33_1,N1372_10_r_6,N6147_3_r_6);
nand I_56(n34_1,n24_1,n29_1);
nor I_57(n35_1,n38_1,n24_1);
nand I_58(n36_1,I_BUFF_1_9_r_1,n23_1);
or I_59(n37_1,G78_5_r_6,n_547_5_r_6);
endmodule


