module test_final(IN_1_0_l_8,IN_2_0_l_8,IN_4_0_l_8,IN_1_1_l_8,IN_2_1_l_8,IN_3_1_l_8,IN_6_1_l_8,IN_1_5_l_8,IN_2_5_l_8,IN_3_5_l_8,IN_6_5_l_8,blif_clk_net_3_r_13,blif_reset_net_3_r_13,n_429_or_0_3_r_13,G78_3_r_13,n_576_3_r_13,n_102_3_r_13,n_547_3_r_13,G42_4_r_13,n_572_4_r_13,n_573_4_r_13,n_549_4_r_13,n_569_4_r_13,n_452_4_r_13);
input IN_1_0_l_8,IN_2_0_l_8,IN_4_0_l_8,IN_1_1_l_8,IN_2_1_l_8,IN_3_1_l_8,IN_6_1_l_8,IN_1_5_l_8,IN_2_5_l_8,IN_3_5_l_8,IN_6_5_l_8,blif_clk_net_3_r_13,blif_reset_net_3_r_13;
output n_429_or_0_3_r_13,G78_3_r_13,n_576_3_r_13,n_102_3_r_13,n_547_3_r_13,G42_4_r_13,n_572_4_r_13,n_573_4_r_13,n_549_4_r_13,n_569_4_r_13,n_452_4_r_13;
wire ACVQN2_0_r_8,n_266_and_0_0_r_8,ACVQN1_2_r_8,P6_2_r_8,n_429_or_0_3_r_8,G78_3_r_8,n_576_3_r_8,n_102_3_r_8,n_547_3_r_8,n_42_5_r_8,G199_5_r_8,ACVQN2_0_l_8,n_266_and_0_0_l_8,ACVQN1_0_l_8,N1_1_l_8,G199_1_l_8,G214_1_l_8,n3_1_l_8,n_42_5_l_8,N3_5_l_8,G199_5_l_8,n3_5_l_8,ACVQN1_0_r_8,P6_internal_2_r_8,n12_3_r_8,n_431_3_r_8,n11_3_r_8,n13_3_r_8,n14_3_r_8,n15_3_r_8,n16_3_r_8,N3_5_r_8,n3_5_r_8,n2_3_r_13,ACVQN1_2_l_13,P6_2_l_13,P6_internal_2_l_13,n_429_or_0_3_l_13,n12_3_l_13,n_431_3_l_13,G78_3_l_13,n_576_3_l_13,n11_3_l_13,n_102_3_l_13,n_547_3_l_13,n13_3_l_13,n14_3_l_13,n15_3_l_13,n16_3_l_13,n12_3_r_13,n_431_3_r_13,n11_3_r_13,n13_3_r_13,n14_3_r_13,n15_3_r_13,n16_3_r_13,n4_4_r_13,n_87_4_r_13,n7_4_r_13;
DFFARX1 I_0(n_266_and_0_0_l_8,blif_clk_net_3_r_13,n2_3_r_13,ACVQN2_0_r_8,);
and I_1(n_266_and_0_0_r_8,G199_5_l_8,ACVQN1_0_r_8);
DFFARX1 I_2(G199_5_l_8,blif_clk_net_3_r_13,n2_3_r_13,ACVQN1_2_r_8,);
not I_3(P6_2_r_8,P6_internal_2_r_8);
nand I_4(n_429_or_0_3_r_8,G199_5_l_8,n12_3_r_8);
DFFARX1 I_5(n_431_3_r_8,blif_clk_net_3_r_13,n2_3_r_13,G78_3_r_8,);
nand I_6(n_576_3_r_8,n_42_5_l_8,n11_3_r_8);
not I_7(n_102_3_r_8,n_266_and_0_0_l_8);
nand I_8(n_547_3_r_8,ACVQN2_0_l_8,n13_3_r_8);
nor I_9(n_42_5_r_8,ACVQN2_0_l_8,n_266_and_0_0_l_8);
DFFARX1 I_10(N3_5_r_8,blif_clk_net_3_r_13,n2_3_r_13,G199_5_r_8,);
DFFARX1 I_11(IN_1_0_l_8,blif_clk_net_3_r_13,n2_3_r_13,ACVQN2_0_l_8,);
and I_12(n_266_and_0_0_l_8,IN_4_0_l_8,ACVQN1_0_l_8);
DFFARX1 I_13(IN_2_0_l_8,blif_clk_net_3_r_13,n2_3_r_13,ACVQN1_0_l_8,);
and I_14(N1_1_l_8,IN_6_1_l_8,n3_1_l_8);
DFFARX1 I_15(N1_1_l_8,blif_clk_net_3_r_13,n2_3_r_13,G199_1_l_8,);
DFFARX1 I_16(IN_3_1_l_8,blif_clk_net_3_r_13,n2_3_r_13,G214_1_l_8,);
nand I_17(n3_1_l_8,IN_1_1_l_8,IN_2_1_l_8);
nor I_18(n_42_5_l_8,IN_1_5_l_8,IN_3_5_l_8);
and I_19(N3_5_l_8,IN_6_5_l_8,n3_5_l_8);
DFFARX1 I_20(N3_5_l_8,blif_clk_net_3_r_13,n2_3_r_13,G199_5_l_8,);
nand I_21(n3_5_l_8,IN_2_5_l_8,IN_3_5_l_8);
DFFARX1 I_22(G214_1_l_8,blif_clk_net_3_r_13,n2_3_r_13,ACVQN1_0_r_8,);
DFFARX1 I_23(G214_1_l_8,blif_clk_net_3_r_13,n2_3_r_13,P6_internal_2_r_8,);
not I_24(n12_3_r_8,G199_1_l_8);
or I_25(n_431_3_r_8,n_42_5_l_8,n14_3_r_8);
nor I_26(n11_3_r_8,n_266_and_0_0_l_8,n12_3_r_8);
nor I_27(n13_3_r_8,n_266_and_0_0_l_8,G199_1_l_8);
and I_28(n14_3_r_8,ACVQN2_0_l_8,n15_3_r_8);
nor I_29(n15_3_r_8,G199_1_l_8,n16_3_r_8);
not I_30(n16_3_r_8,G199_5_l_8);
and I_31(N3_5_r_8,n_42_5_l_8,n3_5_r_8);
nand I_32(n3_5_r_8,ACVQN2_0_l_8,G214_1_l_8);
nand I_33(n_429_or_0_3_r_13,n_429_or_0_3_l_13,n12_3_r_13);
DFFARX1 I_34(n_431_3_r_13,blif_clk_net_3_r_13,n2_3_r_13,G78_3_r_13,);
nand I_35(n_576_3_r_13,n_547_3_l_13,n11_3_r_13);
not I_36(n_102_3_r_13,ACVQN1_2_l_13);
nand I_37(n_547_3_r_13,P6_2_l_13,n13_3_r_13);
DFFARX1 I_38(n4_4_r_13,blif_clk_net_3_r_13,n2_3_r_13,G42_4_r_13,);
nor I_39(n_572_4_r_13,P6_2_l_13,n_429_or_0_3_l_13);
or I_40(n_573_4_r_13,ACVQN1_2_l_13,G78_3_l_13);
nor I_41(n_549_4_r_13,n_429_or_0_3_l_13,n7_4_r_13);
or I_42(n_569_4_r_13,n_429_or_0_3_l_13,G78_3_l_13);
nor I_43(n_452_4_r_13,ACVQN1_2_l_13,P6_2_l_13);
not I_44(n2_3_r_13,blif_reset_net_3_r_13);
DFFARX1 I_45(n_429_or_0_3_r_8,blif_clk_net_3_r_13,n2_3_r_13,ACVQN1_2_l_13,);
not I_46(P6_2_l_13,P6_internal_2_l_13);
DFFARX1 I_47(G78_3_r_8,blif_clk_net_3_r_13,n2_3_r_13,P6_internal_2_l_13,);
nand I_48(n_429_or_0_3_l_13,n12_3_l_13,ACVQN2_0_r_8);
not I_49(n12_3_l_13,G199_5_r_8);
or I_50(n_431_3_l_13,n14_3_l_13,P6_2_r_8);
DFFARX1 I_51(n_431_3_l_13,blif_clk_net_3_r_13,n2_3_r_13,G78_3_l_13,);
nand I_52(n_576_3_l_13,n11_3_l_13,n_547_3_r_8);
nor I_53(n11_3_l_13,n12_3_l_13,n_266_and_0_0_r_8);
not I_54(n_102_3_l_13,n_266_and_0_0_r_8);
nand I_55(n_547_3_l_13,n13_3_l_13,ACVQN1_2_r_8);
nor I_56(n13_3_l_13,n_266_and_0_0_r_8,n_102_3_r_8);
and I_57(n14_3_l_13,n15_3_l_13,n_576_3_r_8);
nor I_58(n15_3_l_13,n16_3_l_13,n_42_5_r_8);
not I_59(n16_3_l_13,ACVQN2_0_r_8);
not I_60(n12_3_r_13,n_102_3_l_13);
or I_61(n_431_3_r_13,ACVQN1_2_l_13,n14_3_r_13);
nor I_62(n11_3_r_13,ACVQN1_2_l_13,n12_3_r_13);
nor I_63(n13_3_r_13,ACVQN1_2_l_13,n_576_3_l_13);
and I_64(n14_3_r_13,n_102_3_l_13,n15_3_r_13);
nor I_65(n15_3_r_13,G78_3_l_13,n16_3_r_13);
not I_66(n16_3_r_13,n_429_or_0_3_l_13);
nor I_67(n4_4_r_13,P6_2_l_13,n_547_3_l_13);
not I_68(n_87_4_r_13,P6_2_l_13);
and I_69(n7_4_r_13,n_576_3_l_13,n_87_4_r_13);
endmodule


