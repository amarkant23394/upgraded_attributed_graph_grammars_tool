module test_I8623(I4629,I1477,I6011,I1470,I5785,I4824,I8623);
input I4629,I1477,I6011,I1470,I5785,I4824;
output I8623;
wire I8216,I5751,I6110,I5743,I6028,I6127,I6079,I4533,I5802,I4509;
not I_0(I8216,I1477);
not I_1(I5751,I1477);
DFFARX1 I_2(I4509,I1470,I5751,,,I6110,);
DFFARX1 I_3(I5743,I1470,I8216,,,I8623,);
nand I_4(I5743,I6127,I6079);
DFFARX1 I_5(I6011,I1470,I5751,,,I6028,);
and I_6(I6127,I6110,I4533);
nor I_7(I6079,I6028,I5802);
or I_8(I4533,I4824,I4629);
DFFARX1 I_9(I5785,I1470,I5751,,,I5802,);
DFFARX1 I_10(I1470,,,I4509,);
endmodule


