module test_final(G18_1_l_3,G15_1_l_3,IN_1_1_l_3,IN_4_1_l_3,IN_5_1_l_3,IN_7_1_l_3,IN_9_1_l_3,IN_10_1_l_3,IN_1_3_l_3,IN_2_3_l_3,IN_4_3_l_3,blif_clk_net_1_r_7,blif_reset_net_1_r_7,G42_1_r_7,n_572_1_r_7,n_573_1_r_7,n_549_1_r_7,n_569_1_r_7,G199_4_r_7,G214_4_r_7,ACVQN1_5_r_7,P6_5_r_7);
input G18_1_l_3,G15_1_l_3,IN_1_1_l_3,IN_4_1_l_3,IN_5_1_l_3,IN_7_1_l_3,IN_9_1_l_3,IN_10_1_l_3,IN_1_3_l_3,IN_2_3_l_3,IN_4_3_l_3,blif_clk_net_1_r_7,blif_reset_net_1_r_7;
output G42_1_r_7,n_572_1_r_7,n_573_1_r_7,n_549_1_r_7,n_569_1_r_7,G199_4_r_7,G214_4_r_7,ACVQN1_5_r_7,P6_5_r_7;
wire G42_1_r_3,n_572_1_r_3,n_573_1_r_3,n_549_1_r_3,n_569_1_r_3,n_452_1_r_3,n_42_2_r_3,G199_2_r_3,ACVQN2_3_r_3,n_266_and_0_3_r_3,n4_1_l_3,G42_1_l_3,n22_3,n40_3,n25_internal_3,n25_3,n4_1_r_3,N3_2_r_3,n_572_1_l_3,ACVQN1_3_r_3,n26_3,n27_3,n28_3,n29_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3,n_431_0_l_7,n8_7,n43_7,n27_7,ACVQN1_5_l_7,n44_7,n4_1_r_7,N1_4_r_7,n26_7,n5_7,P6_5_r_internal_7,n28_7,n29_7,n30_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7;
DFFARX1 I_0(n4_1_r_3,blif_clk_net_1_r_7,n8_7,G42_1_r_3,);
nor I_1(n_572_1_r_3,G42_1_l_3,n28_3);
nand I_2(n_573_1_r_3,n26_3,n27_3);
nor I_3(n_549_1_r_3,n40_3,n32_3);
nand I_4(n_569_1_r_3,n27_3,n31_3);
and I_5(n_452_1_r_3,G18_1_l_3,n26_3);
nor I_6(n_42_2_r_3,n_572_1_l_3,n34_3);
DFFARX1 I_7(N3_2_r_3,blif_clk_net_1_r_7,n8_7,G199_2_r_3,);
DFFARX1 I_8(n_572_1_l_3,blif_clk_net_1_r_7,n8_7,ACVQN2_3_r_3,);
nor I_9(n_266_and_0_3_r_3,n25_3,n35_3);
nor I_10(n4_1_l_3,G18_1_l_3,IN_1_1_l_3);
DFFARX1 I_11(n4_1_l_3,blif_clk_net_1_r_7,n8_7,G42_1_l_3,);
not I_12(n22_3,G42_1_l_3);
DFFARX1 I_13(IN_1_3_l_3,blif_clk_net_1_r_7,n8_7,n40_3,);
DFFARX1 I_14(IN_2_3_l_3,blif_clk_net_1_r_7,n8_7,n25_internal_3,);
not I_15(n25_3,n25_internal_3);
nor I_16(n4_1_r_3,n40_3,n36_3);
nor I_17(N3_2_r_3,n26_3,n37_3);
nor I_18(n_572_1_l_3,G15_1_l_3,IN_7_1_l_3);
DFFARX1 I_19(G42_1_l_3,blif_clk_net_1_r_7,n8_7,ACVQN1_3_r_3,);
nor I_20(n26_3,IN_5_1_l_3,IN_9_1_l_3);
not I_21(n27_3,IN_10_1_l_3);
nor I_22(n28_3,IN_10_1_l_3,n29_3);
nor I_23(n29_3,G15_1_l_3,n30_3);
not I_24(n30_3,IN_4_1_l_3);
nor I_25(n31_3,IN_9_1_l_3,n40_3);
nor I_26(n32_3,n25_3,n33_3);
nand I_27(n33_3,IN_4_3_l_3,n22_3);
or I_28(n34_3,IN_9_1_l_3,IN_10_1_l_3);
nand I_29(n35_3,IN_4_3_l_3,ACVQN1_3_r_3);
nor I_30(n36_3,G18_1_l_3,IN_5_1_l_3);
nor I_31(n37_3,n38_3,n39_3);
not I_32(n38_3,n_572_1_l_3);
nand I_33(n39_3,n27_3,n30_3);
DFFARX1 I_34(n4_1_r_7,blif_clk_net_1_r_7,n8_7,G42_1_r_7,);
nor I_35(n_572_1_r_7,n30_7,n31_7);
nand I_36(n_573_1_r_7,n28_7,n_569_1_r_3);
nor I_37(n_549_1_r_7,ACVQN1_5_l_7,n35_7);
nand I_38(n_569_1_r_7,n32_7,n33_7);
DFFARX1 I_39(N1_4_r_7,blif_clk_net_1_r_7,n8_7,G199_4_r_7,);
DFFARX1 I_40(n26_7,blif_clk_net_1_r_7,n8_7,G214_4_r_7,);
DFFARX1 I_41(n5_7,blif_clk_net_1_r_7,n8_7,ACVQN1_5_r_7,);
not I_42(P6_5_r_7,P6_5_r_internal_7);
or I_43(n_431_0_l_7,n36_7,n_549_1_r_3);
not I_44(n8_7,blif_reset_net_1_r_7);
DFFARX1 I_45(n_431_0_l_7,blif_clk_net_1_r_7,n8_7,n43_7,);
not I_46(n27_7,n43_7);
DFFARX1 I_47(n_42_2_r_3,blif_clk_net_1_r_7,n8_7,ACVQN1_5_l_7,);
DFFARX1 I_48(n_573_1_r_3,blif_clk_net_1_r_7,n8_7,n44_7,);
nor I_49(n4_1_r_7,n30_7,n38_7);
nor I_50(N1_4_r_7,n27_7,n40_7);
nand I_51(n26_7,n39_7,n_266_and_0_3_r_3);
not I_52(n5_7,G199_2_r_3);
DFFARX1 I_53(ACVQN1_5_l_7,blif_clk_net_1_r_7,n8_7,P6_5_r_internal_7,);
nor I_54(n28_7,n26_7,n29_7);
not I_55(n29_7,n_572_1_r_3);
not I_56(n30_7,n_452_1_r_3);
nand I_57(n31_7,n27_7,n29_7);
nor I_58(n32_7,ACVQN1_5_l_7,n34_7);
nor I_59(n33_7,n29_7,G199_2_r_3);
not I_60(n34_7,n_569_1_r_3);
nor I_61(n35_7,n43_7,n44_7);
and I_62(n36_7,n37_7,ACVQN2_3_r_3);
nor I_63(n37_7,n30_7,G42_1_r_3);
nand I_64(n38_7,n29_7,G199_2_r_3);
nor I_65(n39_7,G199_2_r_3,G42_1_r_3);
nor I_66(n40_7,n44_7,n41_7);
nor I_67(n41_7,n34_7,n42_7);
nand I_68(n42_7,n5_7,n_572_1_r_3);
endmodule


