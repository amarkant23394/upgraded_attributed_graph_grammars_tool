module test_I16240(I1477,I16240);
input I1477;
output I16240;
wire ;
not I_0(I16240,I1477);
endmodule


