module test_I2149(I1231,I1477,I1470,I1239,I1375,I1287,I2149);
input I1231,I1477,I1470,I1239,I1375,I1287;
output I2149;
wire I2181,I2294,I2678,I2345,I2633,I2695;
not I_0(I2181,I1477);
nor I_1(I2294,I1287,I1231);
DFFARX1 I_2(I2695,I1470,I2181,,,I2149,);
nand I_3(I2678,I2633,I2294);
DFFARX1 I_4(I1375,I1470,I2181,,,I2345,);
DFFARX1 I_5(I1239,I1470,I2181,,,I2633,);
and I_6(I2695,I2345,I2678);
endmodule


