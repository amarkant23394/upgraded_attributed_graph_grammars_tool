module test_I2583(I1301,I2583);
input I1301;
output I2583;
wire ;
not I_0(I2583,I1301);
endmodule


