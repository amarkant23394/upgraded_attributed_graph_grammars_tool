module test_I6144(I2167,I1477,I6011,I2173,I1470,I6144);
input I2167,I1477,I6011,I2173,I1470;
output I6144;
wire I4629,I6045,I6110,I6028,I4544,I4869,I4595,I5932,I6062,I2143,I4536,I5751,I4533,I5013,I5915,I4807,I5864,I4515,I6127,I4824,I4509;
nor I_0(I4629,I2167,I2173);
nor I_1(I6045,I6028,I5932);
DFFARX1 I_2(I4509,I1470,I5751,,,I6110,);
DFFARX1 I_3(I6011,I1470,I5751,,,I6028,);
not I_4(I4544,I1477);
DFFARX1 I_5(I1470,I4544,,,I4869,);
DFFARX1 I_6(I1470,I4544,,,I4595,);
not I_7(I5932,I5915);
or I_8(I6144,I6127,I6062);
and I_9(I6062,I5864,I6045);
DFFARX1 I_10(I1470,,,I2143,);
nor I_11(I4536,I4869,I4595);
not I_12(I5751,I1477);
or I_13(I4533,I4824,I4629);
or I_14(I5013,I4824);
DFFARX1 I_15(I1470,I5751,,,I5915,);
DFFARX1 I_16(I1470,I4544,,,I4807,);
nor I_17(I5864,I4536,I4515);
not I_18(I4515,I4629);
and I_19(I6127,I6110,I4533);
and I_20(I4824,I4807,I2143);
DFFARX1 I_21(I5013,I1470,I4544,,,I4509,);
endmodule


