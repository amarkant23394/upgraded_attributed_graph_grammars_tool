module test_I11593(I8824,I11508,I1477,I1470,I11593);
input I8824,I11508,I1477,I1470;
output I11593;
wire I11542,I11525,I8833,I9179,I11559,I11310;
or I_0(I11542,I11525,I8833);
DFFARX1 I_1(I11559,I1470,I11310,,,I11593,);
and I_2(I11525,I11508,I8824);
not I_3(I8833,I9179);
DFFARX1 I_4(I1470,,,I9179,);
DFFARX1 I_5(I11542,I1470,I11310,,,I11559,);
not I_6(I11310,I1477);
endmodule


