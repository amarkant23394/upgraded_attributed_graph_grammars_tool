module test_I15276(I10961,I1477,I13102,I1470,I15276);
input I10961,I1477,I13102,I1470;
output I15276;
wire I10647,I12930,I12596,I10639,I12848,I12718,I13119,I12964,I12619,I12913,I14982,I12599,I12882,I10615,I11201,I10609;
not I_0(I10647,I1477);
and I_1(I12930,I12913,I10609);
DFFARX1 I_2(I13119,I1470,I12619,,,I12596,);
DFFARX1 I_3(I11201,I1470,I10647,,,I10639,);
nand I_4(I15276,I14982,I12599);
DFFARX1 I_5(I1470,I12619,,,I12848,);
nor I_6(I12718,I10615,I10639);
or I_7(I13119,I12718,I13102);
nor I_8(I12964,I12930,I12882);
not I_9(I12619,I1477);
DFFARX1 I_10(I1470,I12619,,,I12913,);
not I_11(I14982,I12596);
nand I_12(I12599,I12718,I12964);
not I_13(I12882,I12848);
DFFARX1 I_14(I10961,I1470,I10647,,,I10615,);
and I_15(I11201,I10961);
DFFARX1 I_16(I1470,I10647,,,I10609,);
endmodule


