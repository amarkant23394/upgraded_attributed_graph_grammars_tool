module test_I1492(I1207,I1492);
input I1207;
output I1492;
wire ;
not I_0(I1492,I1207);
endmodule


