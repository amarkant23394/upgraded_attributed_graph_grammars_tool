module test_I12587(I11167,I1477,I11057,I1470,I12587);
input I11167,I1477,I11057,I1470;
output I12587;
wire I12619,I12670,I10612,I10627,I10639,I12653,I12636;
not I_0(I12619,I1477);
DFFARX1 I_1(I12653,I1470,I12619,,,I12670,);
DFFARX1 I_2(I1470,,,I10612,);
nand I_3(I10627,I11167,I11057);
DFFARX1 I_4(I1470,,,I10639,);
and I_5(I12653,I12636,I10627);
DFFARX1 I_6(I12670,I1470,I12619,,,I12587,);
nand I_7(I12636,I10612,I10639);
endmodule


