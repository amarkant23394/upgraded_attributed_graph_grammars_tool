module test_final(IN_1_0_l_15,IN_2_0_l_15,IN_3_0_l_15,IN_4_0_l_15,IN_1_1_l_15,IN_2_1_l_15,IN_3_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_3_3_l_15,IN_1_6_l_15,IN_2_6_l_15,IN_3_6_l_15,IN_4_6_l_15,IN_5_6_l_15,blif_clk_net_5_r_9,blif_reset_net_5_r_9,N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,G78_5_r_9,n_576_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9);
input IN_1_0_l_15,IN_2_0_l_15,IN_3_0_l_15,IN_4_0_l_15,IN_1_1_l_15,IN_2_1_l_15,IN_3_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_3_3_l_15,IN_1_6_l_15,IN_2_6_l_15,IN_3_6_l_15,IN_4_6_l_15,IN_5_6_l_15,blif_clk_net_5_r_9,blif_reset_net_5_r_9;
output N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,G78_5_r_9,n_576_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9;
wire N1371_0_r_15,N1508_0_r_15,N1372_1_r_15,N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_102_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15,n_431_5_r_15,n31_15,n32_15,n33_15,n34_15,n35_15,n36_15,n37_15,n38_15,n39_15,n40_15,n41_15,n42_15,n43_15,n44_15,n45_15,n46_15,n47_15,n48_15,n49_15,n50_15,n51_15,n52_15,n53_15,n54_15,n55_15,n_429_or_0_5_r_9,n_102_5_r_9,I_BUFF_1_9_r_9,n4_7_l_9,n10_9,n62_9,N3_8_l_9,n63_9,n38_9,n_431_5_r_9,N3_8_r_9,n39_9,n40_9,n41_9,n42_9,n43_9,n44_9,n45_9,n46_9,n47_9,n48_9,n49_9,n50_9,n51_9,n52_9,n53_9,n54_9,n55_9,n56_9,n57_9,n58_9,n59_9,n60_9,n61_9;
and I_0(N1371_0_r_15,N1508_0_r_15,n_102_5_r_15);
nor I_1(N1508_0_r_15,IN_2_0_l_15,n55_15);
nor I_2(N1372_1_r_15,n_102_5_r_15,n46_15);
nor I_3(N1508_1_r_15,N1508_0_r_15,n45_15);
not I_4(N1372_4_r_15,n39_15);
nor I_5(N1508_4_r_15,n39_15,n43_15);
nand I_6(n_429_or_0_5_r_15,n36_15,n38_15);
DFFARX1 I_7(n_431_5_r_15,blif_clk_net_5_r_9,n10_9,G78_5_r_15,);
nand I_8(n_576_5_r_15,n31_15,n32_15);
not I_9(n_102_5_r_15,n33_15);
nand I_10(n_547_5_r_15,N1371_0_r_15,n35_15);
nor I_11(N1507_6_r_15,n42_15,n46_15);
nand I_12(N1508_6_r_15,n39_15,n40_15);
nand I_13(n_431_5_r_15,n36_15,n37_15);
nor I_14(n31_15,n33_15,n34_15);
nor I_15(n32_15,IN_1_3_l_15,n44_15);
nor I_16(n33_15,n54_15,n55_15);
nand I_17(n34_15,IN_2_6_l_15,n49_15);
nand I_18(n35_15,IN_1_1_l_15,IN_2_1_l_15);
not I_19(n36_15,n32_15);
nand I_20(n37_15,n34_15,n38_15);
not I_21(n38_15,n46_15);
nand I_22(n39_15,n38_15,n41_15);
nand I_23(n40_15,n41_15,n42_15);
and I_24(n41_15,IN_5_6_l_15,n51_15);
and I_25(n42_15,IN_2_1_l_15,n47_15);
and I_26(n43_15,n34_15,n36_15);
or I_27(n44_15,IN_2_3_l_15,IN_3_3_l_15);
not I_28(n45_15,N1372_1_r_15);
nand I_29(n46_15,IN_2_1_l_15,n53_15);
nor I_30(n47_15,n34_15,n48_15);
not I_31(n48_15,IN_1_1_l_15);
and I_32(n49_15,IN_1_6_l_15,n50_15);
nand I_33(n50_15,n51_15,n52_15);
nand I_34(n51_15,IN_3_6_l_15,IN_4_6_l_15);
not I_35(n52_15,IN_5_6_l_15);
nor I_36(n53_15,IN_3_1_l_15,n48_15);
nor I_37(n54_15,IN_3_0_l_15,IN_4_0_l_15);
not I_38(n55_15,IN_1_0_l_15);
nor I_39(N6147_2_r_9,n62_9,n46_9);
not I_40(N1372_4_r_9,n59_9);
nor I_41(N1508_4_r_9,n58_9,n59_9);
nand I_42(n_429_or_0_5_r_9,n_431_5_r_9,n42_9);
DFFARX1 I_43(n_431_5_r_9,blif_clk_net_5_r_9,n10_9,G78_5_r_9,);
nand I_44(n_576_5_r_9,n39_9,n40_9);
not I_45(n_102_5_r_9,I_BUFF_1_9_r_9);
nand I_46(n_547_5_r_9,n43_9,N1372_4_r_15);
and I_47(n_42_8_r_9,n44_9,N1508_1_r_15);
DFFARX1 I_48(N3_8_r_9,blif_clk_net_5_r_9,n10_9,G199_8_r_9,);
nor I_49(N6147_9_r_9,n41_9,n45_9);
nor I_50(N6134_9_r_9,n45_9,n51_9);
nor I_51(I_BUFF_1_9_r_9,n41_9,N1372_4_r_15);
nor I_52(n4_7_l_9,N1508_1_r_15,G78_5_r_15);
not I_53(n10_9,blif_reset_net_5_r_9);
DFFARX1 I_54(n4_7_l_9,blif_clk_net_5_r_9,n10_9,n62_9,);
and I_55(N3_8_l_9,n57_9,n_547_5_r_15);
DFFARX1 I_56(N3_8_l_9,blif_clk_net_5_r_9,n10_9,n63_9,);
not I_57(n38_9,n63_9);
nor I_58(n_431_5_r_9,N1508_4_r_15,n_429_or_0_5_r_15);
nor I_59(N3_8_r_9,n_102_5_r_9,n53_9);
nor I_60(n39_9,I_BUFF_1_9_r_9,n42_9);
not I_61(n40_9,n41_9);
nand I_62(n41_9,n_429_or_0_5_r_15,N1508_1_r_15);
nor I_63(n42_9,G78_5_r_15,N1507_6_r_15);
nor I_64(n43_9,n63_9,n41_9);
nor I_65(n44_9,G78_5_r_15,N1372_4_r_15);
and I_66(n45_9,n52_9,N1508_4_r_15);
nor I_67(n46_9,n47_9,n48_9);
nor I_68(n47_9,n49_9,n50_9);
not I_69(n48_9,n_429_or_0_5_r_9);
not I_70(n49_9,n42_9);
or I_71(n50_9,n63_9,n51_9);
nor I_72(n51_9,n_576_5_r_15,N1508_6_r_15);
nor I_73(n52_9,n49_9,n_429_or_0_5_r_15);
nor I_74(n53_9,n54_9,n55_9);
nor I_75(n54_9,n56_9,n_429_or_0_5_r_15);
or I_76(n55_9,n44_9,N1507_6_r_15);
not I_77(n56_9,N1508_4_r_15);
nand I_78(n57_9,N1508_6_r_15,n_576_5_r_15);
nor I_79(n58_9,n62_9,n60_9);
nand I_80(n59_9,n51_9,n61_9);
nor I_81(n60_9,n38_9,n44_9);
nor I_82(n61_9,N1508_1_r_15,N1372_4_r_15);
endmodule


