module test_final(IN_1_0_l,IN_2_0_l,IN_4_0_l,G18_4_l,G15_4_l,IN_1_4_l,IN_4_4_l,IN_5_4_l,IN_7_4_l,IN_9_4_l,IN_10_4_l,blif_clk_net_1_r,blif_reset_net_1_r,G199_1_r,G214_1_r,ACVQN1_2_r,P6_2_r,n_429_or_0_3_r,G78_3_r,n_576_3_r,n_102_3_r,n_547_3_r,n_42_5_r,G199_5_r);
input IN_1_0_l,IN_2_0_l,IN_4_0_l,G18_4_l,G15_4_l,IN_1_4_l,IN_4_4_l,IN_5_4_l,IN_7_4_l,IN_9_4_l,IN_10_4_l,blif_clk_net_1_r,blif_reset_net_1_r;
output G199_1_r,G214_1_r,ACVQN1_2_r,P6_2_r,n_429_or_0_3_r,G78_3_r,n_576_3_r,n_102_3_r,n_547_3_r,n_42_5_r,G199_5_r;
wire ACVQN2_0_l,n_266_and_0_0_l,ACVQN1_0_l,G42_4_l,n_87_4_l,n_572_4_l,n_573_4_l,n_549_4_l,n_569_4_l,n_452_4_l,n4_4_l,n7_4_l,N1_1_r,n1_1_r,n3_1_r,P6_internal_2_r,n_431_3_r,n11_3_r,n12_3_r,n13_3_r,n14_3_r,n15_3_r,n16_3_r,N3_5_r,n3_5_r;
DFFARX1 I_0 ( .D(IN_1_0_l), .CLK(blif_clk_net_1_r), .RSTB(n1_1_r), .Q(ACVQN2_0_l) );
and I_1(n_266_and_0_0_l,IN_4_0_l,ACVQN1_0_l);
DFFARX1 I_2 ( .D(IN_2_0_l), .CLK(blif_clk_net_1_r), .RSTB(n1_1_r), .Q(ACVQN1_0_l) );
DFFARX1 I_3 ( .D(n4_4_l), .CLK(blif_clk_net_1_r), .RSTB(n1_1_r), .Q(G42_4_l) );
not I_4(n_87_4_l,G15_4_l);
nor I_5(n_572_4_l,G15_4_l,IN_7_4_l);
or I_6(n_573_4_l,IN_5_4_l,IN_9_4_l);
nor I_7(n_549_4_l,IN_10_4_l,n7_4_l);
or I_8(n_569_4_l,IN_9_4_l,IN_10_4_l);
nor I_9(n_452_4_l,G18_4_l,IN_5_4_l);
nor I_10(n4_4_l,G18_4_l,IN_1_4_l);
and I_11(n7_4_l,IN_4_4_l,n_87_4_l);
DFFARX1 I_12 ( .D(N1_1_r), .CLK(blif_clk_net_1_r), .RSTB(n1_1_r), .Q(G199_1_r) );
DFFARX1 I_13 ( .D(G42_4_l), .CLK(blif_clk_net_1_r), .RSTB(n1_1_r), .Q(G214_1_r) );
and I_14(N1_1_r,n3_1_r,n_266_and_0_0_l);
not I_15(n1_1_r,blif_reset_net_1_r);
nand I_16(n3_1_r,n_569_4_l,n_572_4_l);
DFFARX1 I_17 ( .D(n_572_4_l), .CLK(blif_clk_net_1_r), .RSTB(n1_1_r), .Q(ACVQN1_2_r) );
not I_18(P6_2_r,P6_internal_2_r);
DFFARX1 I_19 ( .D(n_266_and_0_0_l), .CLK(blif_clk_net_1_r), .RSTB(n1_1_r), .Q(P6_internal_2_r) );
nand I_20(n_429_or_0_3_r,n12_3_r,n_572_4_l);
DFFARX1 I_21 ( .D(n_431_3_r), .CLK(blif_clk_net_1_r), .RSTB(n1_1_r), .Q(G78_3_r) );
nand I_22(n_576_3_r,n11_3_r,n_573_4_l);
not I_23(n_102_3_r,n_266_and_0_0_l);
nand I_24(n_547_3_r,n13_3_r,n_549_4_l);
or I_25(n_431_3_r,n14_3_r,n_549_4_l);
nor I_26(n11_3_r,n12_3_r,ACVQN2_0_l);
not I_27(n12_3_r,G42_4_l);
nor I_28(n13_3_r,ACVQN2_0_l,n_266_and_0_0_l);
and I_29(n14_3_r,n15_3_r,n_452_4_l);
nor I_30(n15_3_r,n16_3_r,G42_4_l);
not I_31(n16_3_r,n_572_4_l);
nor I_32(n_42_5_r,n_452_4_l,n_569_4_l);
DFFARX1 I_33 ( .D(N3_5_r), .CLK(blif_clk_net_1_r), .RSTB(n1_1_r), .Q(G199_5_r) );
and I_34(N3_5_r,n3_5_r,ACVQN2_0_l);
nand I_35(n3_5_r,n_573_4_l,n_452_4_l);
endmodule


