module test_I17645(I15713,I1477,I15628,I13749,I1470,I16069,I17645);
input I15713,I1477,I15628,I13749,I1470,I16069;
output I17645;
wire I17594,I15582,I14083,I15591,I17628,I15730,I15832,I15576,I13746,I15611,I15573,I15928,I17611;
not I_0(I17594,I15576);
not I_1(I15582,I15928);
DFFARX1 I_2(I1470,,,I14083,);
nor I_3(I15591,I16069,I15832);
and I_4(I17628,I17611,I15573);
not I_5(I15730,I15713);
nand I_6(I15832,I15628,I13749);
DFFARX1 I_7(I1470,I15611,,,I15576,);
not I_8(I13746,I14083);
or I_9(I17645,I17628,I15582);
not I_10(I15611,I1477);
nand I_11(I15573,I15832,I15730);
DFFARX1 I_12(I13746,I1470,I15611,,,I15928,);
nor I_13(I17611,I17594,I15591);
endmodule


