module test_I11959(I1477,I10507,I10202,I10120,I10032,I10349,I1470,I11959);
input I1477,I10507,I10202,I10120,I10032,I10349,I1470;
output I11959;
wire I12058,I12024,I10287,I12380,I10029,I10219,I12041,I10041,I10052,I10026,I12349,I12007,I10044,I10020,I10397,I11990,I11973;
nand I_0(I12058,I12041,I10026);
nand I_1(I12024,I12007,I10044);
and I_2(I10287,I10219);
nor I_3(I12380,I12349,I12024);
DFFARX1 I_4(I1470,I10052,,,I10029,);
DFFARX1 I_5(I10202,I1470,I10052,,,I10219,);
nor I_6(I12041,I11990,I10020);
nor I_7(I10041,I10349,I10120);
not I_8(I10052,I1477);
nand I_9(I10026,I10219,I10397);
DFFARX1 I_10(I10041,I1470,I11973,,,I12349,);
nor I_11(I12007,I10020,I10029);
DFFARX1 I_12(I10507,I1470,I10052,,,I10044,);
DFFARX1 I_13(I10287,I1470,I10052,,,I10020,);
not I_14(I10397,I10349);
not I_15(I11990,I10032);
not I_16(I11973,I1477);
nand I_17(I11959,I12058,I12380);
endmodule


