module test_I1322(I1231,I1263,I1207,I1294,I1359,I1301,I1322);
input I1231,I1263,I1207,I1294,I1359,I1301;
output I1322;
wire I1704,I1622,I1376,I1342,I1427,I1393,I1639,I1687;
nor I_0(I1704,I1393,I1687);
DFFARX1 I_1(I1294,I1342,,,I1622,);
nand I_2(I1322,I1427,I1704);
and I_3(I1376,I1359,I1231);
not I_4(I1342,I1301);
DFFARX1 I_5(I1263,I1294,I1342,,,I1427,);
DFFARX1 I_6(I1376,I1294,I1342,,,I1393,);
and I_7(I1639,I1622,I1207);
not I_8(I1687,I1639);
endmodule


