module test_I8964(I7122,I5085,I1477,I6975,I1470,I5097,I8964);
input I7122,I5085,I1477,I6975,I1470,I5097;
output I8964;
wire I6893,I7156,I7286,I6992,I5067,I6907,I7269,I7139;
nand I_0(I6893,I7156,I7286);
DFFARX1 I_1(I7139,I1470,I6907,,,I7156,);
nor I_2(I7286,I7269,I6992);
nand I_3(I6992,I6975,I5097);
DFFARX1 I_4(I1470,,,I5067,);
not I_5(I6907,I1477);
DFFARX1 I_6(I5067,I1470,I6907,,,I7269,);
or I_7(I7139,I7122,I5085);
not I_8(I8964,I6893);
endmodule


