module test_I12058(I1477,I10185,I7550,I1470,I12058);
input I1477,I10185,I7550,I1470;
output I12058;
wire I10154,I10202,I10032,I10219,I12041,I10052,I10026,I10349,I10414,I7541,I10332,I10020,I10397,I11990,I10137,I10287;
nand I_0(I10154,I10137);
nand I_1(I12058,I12041,I10026);
and I_2(I10202,I10185,I7541);
nand I_3(I10032,I10137,I10414);
DFFARX1 I_4(I10202,I1470,I10052,,,I10219,);
nor I_5(I12041,I11990,I10020);
not I_6(I10052,I1477);
nand I_7(I10026,I10219,I10397);
and I_8(I10349,I10332,I7550);
nor I_9(I10414,I10397);
DFFARX1 I_10(I1470,,,I7541,);
DFFARX1 I_11(I1470,I10052,,,I10332,);
DFFARX1 I_12(I10287,I1470,I10052,,,I10020,);
not I_13(I10397,I10349);
not I_14(I11990,I10032);
DFFARX1 I_15(I1470,I10052,,,I10137,);
and I_16(I10287,I10219,I10154);
endmodule


