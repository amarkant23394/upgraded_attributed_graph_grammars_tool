module test_I1507(I1423,I1215,I1455,I1507);
input I1423,I1215,I1455;
output I1507;
wire I1603,I1637,I1586,I1535;
nand I_0(I1603,I1586,I1423);
nor I_1(I1507,I1603,I1637);
not I_2(I1637,I1215);
nor I_3(I1586,I1535,I1215);
not I_4(I1535,I1455);
endmodule


