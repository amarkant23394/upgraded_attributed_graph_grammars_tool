module test_I2234(I1687,I1263,I1475,I1294,I1279,I1301,I2234);
input I1687,I1263,I1475,I1294,I1279,I1301;
output I2234;
wire I1704,I1322,I1342,I1427,I1509,I1304,I1954,I1393,I1492;
nor I_0(I1704,I1393,I1687);
nand I_1(I1322,I1427,I1704);
not I_2(I1342,I1301);
nand I_3(I2234,I1954,I1304);
DFFARX1 I_4(I1263,I1294,I1342,,,I1427,);
DFFARX1 I_5(I1492,I1294,I1342,,,I1509,);
DFFARX1 I_6(I1509,I1294,I1342,,,I1304,);
not I_7(I1954,I1322);
DFFARX1 I_8(I1294,I1342,,,I1393,);
and I_9(I1492,I1475,I1279);
endmodule


