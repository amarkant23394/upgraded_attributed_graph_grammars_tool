module test_I17126(I1477,I15064,I15276,I1470,I17126);
input I1477,I15064,I15276,I1470;
output I17126;
wire I14933,I15293,I17092,I16818,I14954,I15310,I14965,I17109;
DFFARX1 I_0(I15310,I1470,I14965,,,I14933,);
DFFARX1 I_1(I17109,I1470,I16818,,,I17126,);
nand I_2(I15293,I15276);
DFFARX1 I_3(I14954,I1470,I16818,,,I17092,);
not I_4(I16818,I1477);
not I_5(I14954,I15064);
and I_6(I15310,I15276,I15293);
not I_7(I14965,I1477);
and I_8(I17109,I17092,I14933);
endmodule


