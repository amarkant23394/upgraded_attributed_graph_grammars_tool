module test_final(G18_1_l_13,G15_1_l_13,IN_1_1_l_13,IN_4_1_l_13,IN_5_1_l_13,IN_7_1_l_13,IN_9_1_l_13,IN_10_1_l_13,IN_1_3_l_13,IN_2_3_l_13,IN_4_3_l_13,blif_clk_net_1_r_1,blif_reset_net_1_r_1,G42_1_r_1,n_572_1_r_1,n_573_1_r_1,n_549_1_r_1,n_452_1_r_1,ACVQN2_3_r_1,n_266_and_0_3_r_1,G199_4_r_1,G214_4_r_1);
input G18_1_l_13,G15_1_l_13,IN_1_1_l_13,IN_4_1_l_13,IN_5_1_l_13,IN_7_1_l_13,IN_9_1_l_13,IN_10_1_l_13,IN_1_3_l_13,IN_2_3_l_13,IN_4_3_l_13,blif_clk_net_1_r_1,blif_reset_net_1_r_1;
output G42_1_r_1,n_572_1_r_1,n_573_1_r_1,n_549_1_r_1,n_452_1_r_1,ACVQN2_3_r_1,n_266_and_0_3_r_1,G199_4_r_1,G214_4_r_1;
wire G42_1_r_13,n_572_1_r_13,n_573_1_r_13,n_549_1_r_13,n_569_1_r_13,n_452_1_r_13,ACVQN2_3_r_13,n_266_and_0_3_r_13,ACVQN1_5_r_13,P6_5_r_13,n4_1_l_13,n17_internal_13,n17_13,n28_13,ACVQN1_3_l_13,n4_1_r_13,n_266_and_0_3_l_13,n_573_1_l_13,n14_internal_13,n14_13,n_549_1_l_13,n_569_1_l_13,P6_5_r_internal_13,n18_13,n19_13,n20_13,n21_13,n22_13,n23_13,n24_13,n25_13,n26_13,n27_13,N3_2_l_1,n5_1,n26_1,n17_1,n16_internal_1,n16_1,ACVQN1_3_l_1,N1_4_l_1,G199_4_l_1,G214_4_l_1,n4_1_r_1,n14_internal_1,n14_1,N1_4_r_1,n18_1,n19_1,n20_1,n21_1,n22_1,n23_1,n24_1,n25_1;
DFFARX1 I_0(n4_1_r_13,blif_clk_net_1_r_1,n5_1,G42_1_r_13,);
nor I_1(n_572_1_r_13,n28_13,n_569_1_l_13);
nand I_2(n_573_1_r_13,n18_13,n19_13);
nand I_3(n_549_1_r_13,n_569_1_r_13,n22_13);
nand I_4(n_569_1_r_13,n17_13,n18_13);
nor I_5(n_452_1_r_13,n_573_1_l_13,n25_13);
DFFARX1 I_6(n_266_and_0_3_l_13,blif_clk_net_1_r_1,n5_1,ACVQN2_3_r_13,);
nor I_7(n_266_and_0_3_r_13,n17_13,n14_13);
DFFARX1 I_8(n_549_1_l_13,blif_clk_net_1_r_1,n5_1,ACVQN1_5_r_13,);
not I_9(P6_5_r_13,P6_5_r_internal_13);
nor I_10(n4_1_l_13,G18_1_l_13,IN_1_1_l_13);
DFFARX1 I_11(n4_1_l_13,blif_clk_net_1_r_1,n5_1,n17_internal_13,);
not I_12(n17_13,n17_internal_13);
DFFARX1 I_13(IN_1_3_l_13,blif_clk_net_1_r_1,n5_1,n28_13,);
DFFARX1 I_14(IN_2_3_l_13,blif_clk_net_1_r_1,n5_1,ACVQN1_3_l_13,);
nor I_15(n4_1_r_13,n_573_1_l_13,n_549_1_l_13);
and I_16(n_266_and_0_3_l_13,IN_4_3_l_13,ACVQN1_3_l_13);
nand I_17(n_573_1_l_13,n20_13,n24_13);
DFFARX1 I_18(n_573_1_l_13,blif_clk_net_1_r_1,n5_1,n14_internal_13,);
not I_19(n14_13,n14_internal_13);
and I_20(n_549_1_l_13,n21_13,n26_13);
nand I_21(n_569_1_l_13,n20_13,n21_13);
DFFARX1 I_22(n_569_1_l_13,blif_clk_net_1_r_1,n5_1,P6_5_r_internal_13,);
nand I_23(n18_13,n23_13,n24_13);
or I_24(n19_13,G15_1_l_13,IN_7_1_l_13);
not I_25(n20_13,IN_9_1_l_13);
not I_26(n21_13,IN_10_1_l_13);
nand I_27(n22_13,n17_13,n28_13);
not I_28(n23_13,G18_1_l_13);
not I_29(n24_13,IN_5_1_l_13);
nor I_30(n25_13,G15_1_l_13,IN_7_1_l_13);
nand I_31(n26_13,IN_4_1_l_13,n27_13);
not I_32(n27_13,G15_1_l_13);
DFFARX1 I_33(n4_1_r_1,blif_clk_net_1_r_1,n5_1,G42_1_r_1,);
nor I_34(n_572_1_r_1,n26_1,n19_1);
nand I_35(n_573_1_r_1,n16_1,n18_1);
nor I_36(n_549_1_r_1,n20_1,n21_1);
nor I_37(n_452_1_r_1,G214_4_l_1,n20_1);
DFFARX1 I_38(G199_4_l_1,blif_clk_net_1_r_1,n5_1,ACVQN2_3_r_1,);
nor I_39(n_266_and_0_3_r_1,n16_1,n14_1);
DFFARX1 I_40(N1_4_r_1,blif_clk_net_1_r_1,n5_1,G199_4_r_1,);
DFFARX1 I_41(G199_4_l_1,blif_clk_net_1_r_1,n5_1,G214_4_r_1,);
and I_42(N3_2_l_1,n23_1,ACVQN1_5_r_13);
not I_43(n5_1,blif_reset_net_1_r_1);
DFFARX1 I_44(N3_2_l_1,blif_clk_net_1_r_1,n5_1,n26_1,);
not I_45(n17_1,n26_1);
DFFARX1 I_46(ACVQN2_3_r_13,blif_clk_net_1_r_1,n5_1,n16_internal_1,);
not I_47(n16_1,n16_internal_1);
DFFARX1 I_48(n_573_1_r_13,blif_clk_net_1_r_1,n5_1,ACVQN1_3_l_1,);
and I_49(N1_4_l_1,n25_1,G42_1_r_13);
DFFARX1 I_50(N1_4_l_1,blif_clk_net_1_r_1,n5_1,G199_4_l_1,);
DFFARX1 I_51(P6_5_r_13,blif_clk_net_1_r_1,n5_1,G214_4_l_1,);
nor I_52(n4_1_r_1,n26_1,G214_4_l_1);
DFFARX1 I_53(G214_4_l_1,blif_clk_net_1_r_1,n5_1,n14_internal_1,);
not I_54(n14_1,n14_internal_1);
nor I_55(N1_4_r_1,n17_1,n24_1);
nand I_56(n18_1,ACVQN1_3_l_1,n_266_and_0_3_r_13);
nor I_57(n19_1,G42_1_r_13,n_572_1_r_13);
not I_58(n20_1,n18_1);
nor I_59(n21_1,n26_1,n22_1);
not I_60(n22_1,n19_1);
nand I_61(n23_1,n_549_1_r_13,n_572_1_r_13);
nor I_62(n24_1,n18_1,n22_1);
nand I_63(n25_1,n_572_1_r_13,n_452_1_r_13);
endmodule


