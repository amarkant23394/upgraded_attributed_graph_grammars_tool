module test_final(G18_1_l_13,G15_1_l_13,IN_1_1_l_13,IN_4_1_l_13,IN_5_1_l_13,IN_7_1_l_13,IN_9_1_l_13,IN_10_1_l_13,IN_1_3_l_13,IN_2_3_l_13,IN_4_3_l_13,blif_clk_net_1_r_12,blif_reset_net_1_r_12,G42_1_r_12,n_572_1_r_12,n_573_1_r_12,n_549_1_r_12,n_42_2_r_12,G199_2_r_12,ACVQN1_5_r_12,P6_5_r_12);
input G18_1_l_13,G15_1_l_13,IN_1_1_l_13,IN_4_1_l_13,IN_5_1_l_13,IN_7_1_l_13,IN_9_1_l_13,IN_10_1_l_13,IN_1_3_l_13,IN_2_3_l_13,IN_4_3_l_13,blif_clk_net_1_r_12,blif_reset_net_1_r_12;
output G42_1_r_12,n_572_1_r_12,n_573_1_r_12,n_549_1_r_12,n_42_2_r_12,G199_2_r_12,ACVQN1_5_r_12,P6_5_r_12;
wire G42_1_r_13,n_572_1_r_13,n_573_1_r_13,n_549_1_r_13,n_569_1_r_13,n_452_1_r_13,ACVQN2_3_r_13,n_266_and_0_3_r_13,ACVQN1_5_r_13,P6_5_r_13,n4_1_l_13,n17_internal_13,n17_13,n28_13,ACVQN1_3_l_13,n4_1_r_13,n_266_and_0_3_l_13,n_573_1_l_13,n14_internal_13,n14_13,n_549_1_l_13,n_569_1_l_13,P6_5_r_internal_13,n18_13,n19_13,n20_13,n21_13,n22_13,n23_13,n24_13,n25_13,n26_13,n27_13,n_431_0_l_12,n8_12,n41_12,ACVQN1_5_l_12,n22_12,n42_12,n4_1_r_12,N3_2_r_12,n3_12,P6_5_r_internal_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12;
DFFARX1 I_0(n4_1_r_13,blif_clk_net_1_r_12,n8_12,G42_1_r_13,);
nor I_1(n_572_1_r_13,n28_13,n_569_1_l_13);
nand I_2(n_573_1_r_13,n18_13,n19_13);
nand I_3(n_549_1_r_13,n_569_1_r_13,n22_13);
nand I_4(n_569_1_r_13,n17_13,n18_13);
nor I_5(n_452_1_r_13,n_573_1_l_13,n25_13);
DFFARX1 I_6(n_266_and_0_3_l_13,blif_clk_net_1_r_12,n8_12,ACVQN2_3_r_13,);
nor I_7(n_266_and_0_3_r_13,n17_13,n14_13);
DFFARX1 I_8(n_549_1_l_13,blif_clk_net_1_r_12,n8_12,ACVQN1_5_r_13,);
not I_9(P6_5_r_13,P6_5_r_internal_13);
nor I_10(n4_1_l_13,G18_1_l_13,IN_1_1_l_13);
DFFARX1 I_11(n4_1_l_13,blif_clk_net_1_r_12,n8_12,n17_internal_13,);
not I_12(n17_13,n17_internal_13);
DFFARX1 I_13(IN_1_3_l_13,blif_clk_net_1_r_12,n8_12,n28_13,);
DFFARX1 I_14(IN_2_3_l_13,blif_clk_net_1_r_12,n8_12,ACVQN1_3_l_13,);
nor I_15(n4_1_r_13,n_573_1_l_13,n_549_1_l_13);
and I_16(n_266_and_0_3_l_13,IN_4_3_l_13,ACVQN1_3_l_13);
nand I_17(n_573_1_l_13,n20_13,n24_13);
DFFARX1 I_18(n_573_1_l_13,blif_clk_net_1_r_12,n8_12,n14_internal_13,);
not I_19(n14_13,n14_internal_13);
and I_20(n_549_1_l_13,n21_13,n26_13);
nand I_21(n_569_1_l_13,n20_13,n21_13);
DFFARX1 I_22(n_569_1_l_13,blif_clk_net_1_r_12,n8_12,P6_5_r_internal_13,);
nand I_23(n18_13,n23_13,n24_13);
or I_24(n19_13,G15_1_l_13,IN_7_1_l_13);
not I_25(n20_13,IN_9_1_l_13);
not I_26(n21_13,IN_10_1_l_13);
nand I_27(n22_13,n17_13,n28_13);
not I_28(n23_13,G18_1_l_13);
not I_29(n24_13,IN_5_1_l_13);
nor I_30(n25_13,G15_1_l_13,IN_7_1_l_13);
nand I_31(n26_13,IN_4_1_l_13,n27_13);
not I_32(n27_13,G15_1_l_13);
DFFARX1 I_33(n4_1_r_12,blif_clk_net_1_r_12,n8_12,G42_1_r_12,);
nor I_34(n_572_1_r_12,n29_12,n30_12);
nand I_35(n_573_1_r_12,n26_12,n27_12);
nor I_36(n_549_1_r_12,n33_12,n34_12);
and I_37(n_42_2_r_12,n42_12,n39_12);
DFFARX1 I_38(N3_2_r_12,blif_clk_net_1_r_12,n8_12,G199_2_r_12,);
DFFARX1 I_39(n3_12,blif_clk_net_1_r_12,n8_12,ACVQN1_5_r_12,);
not I_40(P6_5_r_12,P6_5_r_internal_12);
or I_41(n_431_0_l_12,n36_12,n_572_1_r_13);
not I_42(n8_12,blif_reset_net_1_r_12);
DFFARX1 I_43(n_431_0_l_12,blif_clk_net_1_r_12,n8_12,n41_12,);
DFFARX1 I_44(n_266_and_0_3_r_13,blif_clk_net_1_r_12,n8_12,ACVQN1_5_l_12,);
not I_45(n22_12,ACVQN1_5_l_12);
DFFARX1 I_46(n_549_1_r_13,blif_clk_net_1_r_12,n8_12,n42_12,);
nor I_47(n4_1_r_12,n41_12,n31_12);
nor I_48(N3_2_r_12,n22_12,n40_12);
not I_49(n3_12,n39_12);
DFFARX1 I_50(ACVQN1_5_l_12,blif_clk_net_1_r_12,n8_12,P6_5_r_internal_12,);
and I_51(n26_12,P6_5_r_13,n_572_1_r_13);
nor I_52(n27_12,n28_12,n29_12);
not I_53(n28_12,n_573_1_r_13);
nand I_54(n29_12,n31_12,n32_12);
nand I_55(n30_12,n42_12,n_573_1_r_13);
not I_56(n31_12,G42_1_r_13);
not I_57(n32_12,n_452_1_r_13);
nand I_58(n33_12,n31_12,n35_12);
nand I_59(n34_12,P6_5_r_13,n_572_1_r_13);
nand I_60(n35_12,n41_12,n42_12);
and I_61(n36_12,n37_12,ACVQN2_3_r_13);
nor I_62(n37_12,n38_12,ACVQN1_5_r_13);
not I_63(n38_12,G42_1_r_13);
nor I_64(n39_12,n38_12,P6_5_r_13);
nor I_65(n40_12,n39_12,G42_1_r_13);
endmodule


