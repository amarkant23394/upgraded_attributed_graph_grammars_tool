module test_I3504(I1750,I1477,I1470,I1535,I1207,I3504);
input I1750,I1477,I1470,I1535,I1207;
output I3504;
wire I1518,I1486,I1801,I1489,I1832,I3487,I1767;
not I_0(I1518,I1477);
DFFARX1 I_1(I1832,I1470,I1518,,,I1486,);
DFFARX1 I_2(I1767,I1470,I1518,,,I1801,);
and I_3(I3504,I3487,I1489);
not I_4(I1489,I1801);
nand I_5(I1832,I1535,I1207);
not I_6(I3487,I1486);
DFFARX1 I_7(I1750,I1470,I1518,,,I1767,);
endmodule


