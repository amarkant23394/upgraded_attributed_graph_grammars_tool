module test_I7850(I7765,I1477,I6843,I1470,I7850);
input I7765,I1477,I6843,I1470;
output I7850;
wire I6297,I7799,I7816,I7570,I7714,I6329,I7731,I7782,I6312,I6411,I6306;
DFFARX1 I_0(I6843,I1470,I6329,,,I6297,);
or I_1(I7799,I7782,I6306);
DFFARX1 I_2(I7799,I1470,I7570,,,I7816,);
not I_3(I7570,I1477);
not I_4(I7714,I6297);
nor I_5(I7850,I7816,I7731);
not I_6(I6329,I1477);
not I_7(I7731,I7714);
and I_8(I7782,I7765,I6312);
DFFARX1 I_9(I1470,I6329,,,I6312,);
DFFARX1 I_10(I1470,I6329,,,I6411,);
not I_11(I6306,I6411);
endmodule


