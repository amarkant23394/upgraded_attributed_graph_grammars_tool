module test_I4521(I1477,I1470,I2695,I4521);
input I1477,I1470,I2695;
output I4521;
wire I4917,I2181,I4544,I4869,I2149,I4674,I2155,I2633;
nor I_0(I4917,I4869,I4674);
not I_1(I2181,I1477);
not I_2(I4544,I1477);
DFFARX1 I_3(I4917,I1470,I4544,,,I4521,);
DFFARX1 I_4(I2149,I1470,I4544,,,I4869,);
DFFARX1 I_5(I2695,I1470,I2181,,,I2149,);
DFFARX1 I_6(I2155,I1470,I4544,,,I4674,);
DFFARX1 I_7(I2633,I1470,I2181,,,I2155,);
DFFARX1 I_8(I1470,I2181,,,I2633,);
endmodule


