module test_final(G1_0_l_12,G2_0_l_12,IN_2_0_l_12,IN_4_0_l_12,IN_5_0_l_12,IN_7_0_l_12,IN_8_0_l_12,IN_10_0_l_12,IN_11_0_l_12,IN_1_5_l_12,IN_2_5_l_12,blif_clk_net_1_r_4,blif_reset_net_1_r_4,G42_1_r_4,n_572_1_r_4,n_573_1_r_4,n_549_1_r_4,n_569_1_r_4,ACVQN2_3_r_4,n_266_and_0_3_r_4,ACVQN1_5_r_4,P6_5_r_4);
input G1_0_l_12,G2_0_l_12,IN_2_0_l_12,IN_4_0_l_12,IN_5_0_l_12,IN_7_0_l_12,IN_8_0_l_12,IN_10_0_l_12,IN_11_0_l_12,IN_1_5_l_12,IN_2_5_l_12,blif_clk_net_1_r_4,blif_reset_net_1_r_4;
output G42_1_r_4,n_572_1_r_4,n_573_1_r_4,n_549_1_r_4,n_569_1_r_4,ACVQN2_3_r_4,n_266_and_0_3_r_4,ACVQN1_5_r_4,P6_5_r_4;
wire G42_1_r_12,n_572_1_r_12,n_573_1_r_12,n_549_1_r_12,n_42_2_r_12,G199_2_r_12,ACVQN1_5_r_12,P6_5_r_12,n_431_0_l_12,n41_12,ACVQN1_5_l_12,n22_12,n42_12,n4_1_r_12,N3_2_r_12,n3_12,P6_5_r_internal_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12,n_431_0_l_4,n6_4,G78_0_l_4,ACVQN1_5_l_4,n16_4,n17_internal_4,n17_4,n4_1_r_4,n19_4,n15_internal_4,n15_4,P6_5_r_internal_4,n20_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4;
DFFARX1 I_0(n4_1_r_12,blif_clk_net_1_r_4,n6_4,G42_1_r_12,);
nor I_1(n_572_1_r_12,n29_12,n30_12);
nand I_2(n_573_1_r_12,n26_12,n27_12);
nor I_3(n_549_1_r_12,n33_12,n34_12);
and I_4(n_42_2_r_12,n42_12,n39_12);
DFFARX1 I_5(N3_2_r_12,blif_clk_net_1_r_4,n6_4,G199_2_r_12,);
DFFARX1 I_6(n3_12,blif_clk_net_1_r_4,n6_4,ACVQN1_5_r_12,);
not I_7(P6_5_r_12,P6_5_r_internal_12);
or I_8(n_431_0_l_12,IN_8_0_l_12,n36_12);
DFFARX1 I_9(n_431_0_l_12,blif_clk_net_1_r_4,n6_4,n41_12,);
DFFARX1 I_10(IN_2_5_l_12,blif_clk_net_1_r_4,n6_4,ACVQN1_5_l_12,);
not I_11(n22_12,ACVQN1_5_l_12);
DFFARX1 I_12(IN_1_5_l_12,blif_clk_net_1_r_4,n6_4,n42_12,);
nor I_13(n4_1_r_12,n41_12,n31_12);
nor I_14(N3_2_r_12,n22_12,n40_12);
not I_15(n3_12,n39_12);
DFFARX1 I_16(ACVQN1_5_l_12,blif_clk_net_1_r_4,n6_4,P6_5_r_internal_12,);
and I_17(n26_12,IN_5_0_l_12,IN_7_0_l_12);
nor I_18(n27_12,n28_12,n29_12);
not I_19(n28_12,IN_11_0_l_12);
nand I_20(n29_12,n31_12,n32_12);
nand I_21(n30_12,IN_11_0_l_12,n42_12);
not I_22(n31_12,G2_0_l_12);
not I_23(n32_12,IN_10_0_l_12);
nand I_24(n33_12,n31_12,n35_12);
nand I_25(n34_12,IN_5_0_l_12,IN_7_0_l_12);
nand I_26(n35_12,n41_12,n42_12);
and I_27(n36_12,IN_2_0_l_12,n37_12);
nor I_28(n37_12,IN_4_0_l_12,n38_12);
not I_29(n38_12,G1_0_l_12);
nor I_30(n39_12,IN_5_0_l_12,n38_12);
nor I_31(n40_12,G2_0_l_12,n39_12);
DFFARX1 I_32(n4_1_r_4,blif_clk_net_1_r_4,n6_4,G42_1_r_4,);
nor I_33(n_572_1_r_4,G78_0_l_4,n17_4);
nand I_34(n_573_1_r_4,n16_4,P6_5_r_12);
nor I_35(n_549_1_r_4,n22_4,n23_4);
nand I_36(n_569_1_r_4,n20_4,n21_4);
DFFARX1 I_37(n19_4,blif_clk_net_1_r_4,n6_4,ACVQN2_3_r_4,);
nor I_38(n_266_and_0_3_r_4,n15_4,n29_4);
DFFARX1 I_39(n19_4,blif_clk_net_1_r_4,n6_4,ACVQN1_5_r_4,);
not I_40(P6_5_r_4,P6_5_r_internal_4);
or I_41(n_431_0_l_4,n26_4,ACVQN1_5_r_12);
not I_42(n6_4,blif_reset_net_1_r_4);
DFFARX1 I_43(n_431_0_l_4,blif_clk_net_1_r_4,n6_4,G78_0_l_4,);
DFFARX1 I_44(n_572_1_r_12,blif_clk_net_1_r_4,n6_4,ACVQN1_5_l_4,);
not I_45(n16_4,ACVQN1_5_l_4);
DFFARX1 I_46(n_549_1_r_12,blif_clk_net_1_r_4,n6_4,n17_internal_4,);
not I_47(n17_4,n17_internal_4);
nor I_48(n4_1_r_4,n30_4,n31_4);
nand I_49(n19_4,n33_4,G42_1_r_12);
DFFARX1 I_50(G78_0_l_4,blif_clk_net_1_r_4,n6_4,n15_internal_4,);
not I_51(n15_4,n15_internal_4);
DFFARX1 I_52(ACVQN1_5_l_4,blif_clk_net_1_r_4,n6_4,P6_5_r_internal_4,);
and I_53(n20_4,n16_4,n_42_2_r_12);
nor I_54(n21_4,P6_5_r_12,n_572_1_r_12);
nand I_55(n22_4,G78_0_l_4,n25_4);
nand I_56(n23_4,n24_4,n_42_2_r_12);
not I_57(n24_4,P6_5_r_12);
not I_58(n25_4,n_572_1_r_12);
and I_59(n26_4,n27_4,G199_2_r_12);
nor I_60(n27_4,n28_4,n_573_1_r_12);
not I_61(n28_4,G42_1_r_12);
not I_62(n29_4,n30_4);
nand I_63(n30_4,n32_4,G42_1_r_12);
nand I_64(n31_4,n25_4,n_42_2_r_12);
nor I_65(n32_4,n33_4,P6_5_r_12);
not I_66(n33_4,n_573_1_r_12);
endmodule


