module test_final(IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_6_2_l_6,IN_1_3_l_6,IN_2_3_l_6,IN_4_3_l_6,IN_1_4_l_6,IN_2_4_l_6,IN_3_4_l_6,IN_6_4_l_6,blif_clk_net_1_r_16,blif_reset_net_1_r_16,G42_1_r_16,n_572_1_r_16,n_573_1_r_16,n_549_1_r_16,n_569_1_r_16,n_452_1_r_16,G199_4_r_16,G214_4_r_16,ACVQN1_5_r_16,P6_5_r_16);
input IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_6_2_l_6,IN_1_3_l_6,IN_2_3_l_6,IN_4_3_l_6,IN_1_4_l_6,IN_2_4_l_6,IN_3_4_l_6,IN_6_4_l_6,blif_clk_net_1_r_16,blif_reset_net_1_r_16;
output G42_1_r_16,n_572_1_r_16,n_573_1_r_16,n_549_1_r_16,n_569_1_r_16,n_452_1_r_16,G199_4_r_16,G214_4_r_16,ACVQN1_5_r_16,P6_5_r_16;
wire G42_1_r_6,n_572_1_r_6,n_573_1_r_6,n_549_1_r_6,n_569_1_r_6,n_452_1_r_6,G199_4_r_6,G214_4_r_6,ACVQN1_5_r_6,P6_5_r_6,N3_2_l_6,n27_6,n17_6,n28_6,n26_6,N1_4_l_6,n29_6,n18_6,G214_4_l_6,n12_6,n4_1_r_6,N1_4_r_6,n_42_2_l_6,P6_5_r_internal_6,n19_6,n20_6,n21_6,n22_6,n23_6,n24_6,n25_6,n4_1_l_16,n7_16,n29_16,n16_internal_16,n16_16,ACVQN1_3_l_16,n4_1_r_16,N1_4_r_16,n6_16,n_573_1_l_16,n_452_1_l_16,P6_5_r_internal_16,n18_16,n19_16,n20_16,n21_16,n22_16,n23_16,n24_16,n25_16,n26_16,n27_16,n28_16;
DFFARX1 I_0(n4_1_r_6,blif_clk_net_1_r_16,n7_16,G42_1_r_6,);
nor I_1(n_572_1_r_6,n27_6,n28_6);
nand I_2(n_573_1_r_6,n18_6,n19_6);
nor I_3(n_549_1_r_6,n_42_2_l_6,n21_6);
nand I_4(n_569_1_r_6,n19_6,n20_6);
nor I_5(n_452_1_r_6,n28_6,n29_6);
DFFARX1 I_6(N1_4_r_6,blif_clk_net_1_r_16,n7_16,G199_4_r_6,);
DFFARX1 I_7(n_42_2_l_6,blif_clk_net_1_r_16,n7_16,G214_4_r_6,);
DFFARX1 I_8(n_42_2_l_6,blif_clk_net_1_r_16,n7_16,ACVQN1_5_r_6,);
not I_9(P6_5_r_6,P6_5_r_internal_6);
and I_10(N3_2_l_6,IN_6_2_l_6,n23_6);
DFFARX1 I_11(N3_2_l_6,blif_clk_net_1_r_16,n7_16,n27_6,);
not I_12(n17_6,n27_6);
DFFARX1 I_13(IN_1_3_l_6,blif_clk_net_1_r_16,n7_16,n28_6,);
DFFARX1 I_14(IN_2_3_l_6,blif_clk_net_1_r_16,n7_16,n26_6,);
and I_15(N1_4_l_6,IN_6_4_l_6,n25_6);
DFFARX1 I_16(N1_4_l_6,blif_clk_net_1_r_16,n7_16,n29_6,);
not I_17(n18_6,n29_6);
DFFARX1 I_18(IN_3_4_l_6,blif_clk_net_1_r_16,n7_16,G214_4_l_6,);
not I_19(n12_6,G214_4_l_6);
nor I_20(n4_1_r_6,n28_6,n22_6);
nor I_21(N1_4_r_6,n12_6,n24_6);
nor I_22(n_42_2_l_6,IN_1_2_l_6,IN_3_2_l_6);
DFFARX1 I_23(G214_4_l_6,blif_clk_net_1_r_16,n7_16,P6_5_r_internal_6,);
nand I_24(n19_6,IN_4_3_l_6,n26_6);
not I_25(n20_6,n_42_2_l_6);
nor I_26(n21_6,n17_6,n28_6);
and I_27(n22_6,IN_4_3_l_6,n26_6);
nand I_28(n23_6,IN_2_2_l_6,IN_3_2_l_6);
nor I_29(n24_6,n17_6,n18_6);
nand I_30(n25_6,IN_1_4_l_6,IN_2_4_l_6);
DFFARX1 I_31(n4_1_r_16,blif_clk_net_1_r_16,n7_16,G42_1_r_16,);
nor I_32(n_572_1_r_16,n20_16,n21_16);
nand I_33(n_573_1_r_16,n18_16,n19_16);
nor I_34(n_549_1_r_16,n23_16,n24_16);
nand I_35(n_569_1_r_16,n18_16,n22_16);
nor I_36(n_452_1_r_16,n29_16,n6_16);
DFFARX1 I_37(N1_4_r_16,blif_clk_net_1_r_16,n7_16,G199_4_r_16,);
DFFARX1 I_38(n6_16,blif_clk_net_1_r_16,n7_16,G214_4_r_16,);
DFFARX1 I_39(n_573_1_l_16,blif_clk_net_1_r_16,n7_16,ACVQN1_5_r_16,);
not I_40(P6_5_r_16,P6_5_r_internal_16);
nor I_41(n4_1_l_16,G199_4_r_6,ACVQN1_5_r_6);
not I_42(n7_16,blif_reset_net_1_r_16);
DFFARX1 I_43(n4_1_l_16,blif_clk_net_1_r_16,n7_16,n29_16,);
DFFARX1 I_44(G42_1_r_6,blif_clk_net_1_r_16,n7_16,n16_internal_16,);
not I_45(n16_16,n16_internal_16);
DFFARX1 I_46(G214_4_r_6,blif_clk_net_1_r_16,n7_16,ACVQN1_3_l_16,);
nor I_47(n4_1_r_16,n29_16,n21_16);
nor I_48(N1_4_r_16,n27_16,n28_16);
not I_49(n6_16,n19_16);
or I_50(n_573_1_l_16,n_573_1_r_6,n_549_1_r_6);
nor I_51(n_452_1_l_16,n_549_1_r_6,G199_4_r_6);
DFFARX1 I_52(n_452_1_l_16,blif_clk_net_1_r_16,n7_16,P6_5_r_internal_16,);
not I_53(n18_16,n20_16);
nor I_54(n19_16,n_573_1_r_6,G42_1_r_6);
nor I_55(n20_16,n_569_1_r_6,P6_5_r_6);
nor I_56(n21_16,n25_16,G42_1_r_6);
nand I_57(n22_16,ACVQN1_3_l_16,n_572_1_r_6);
not I_58(n23_16,n22_16);
nor I_59(n24_16,n16_16,n20_16);
nor I_60(n25_16,n26_16,P6_5_r_6);
not I_61(n26_16,n_452_1_r_6);
and I_62(n27_16,n29_16,n_573_1_r_6);
not I_63(n28_16,n_452_1_l_16);
endmodule


