module test_final(IN_1_2_l_13,IN_2_2_l_13,G1_3_l_13,G2_3_l_13,IN_2_3_l_13,IN_4_3_l_13,IN_5_3_l_13,IN_7_3_l_13,IN_8_3_l_13,IN_10_3_l_13,IN_11_3_l_13,blif_clk_net_3_r_10,blif_reset_net_3_r_10,n_429_or_0_3_r_10,G78_3_r_10,n_576_3_r_10,n_102_3_r_10,n_547_3_r_10,G42_4_r_10,n_572_4_r_10,n_573_4_r_10,n_549_4_r_10,n_569_4_r_10,n_452_4_r_10);
input IN_1_2_l_13,IN_2_2_l_13,G1_3_l_13,G2_3_l_13,IN_2_3_l_13,IN_4_3_l_13,IN_5_3_l_13,IN_7_3_l_13,IN_8_3_l_13,IN_10_3_l_13,IN_11_3_l_13,blif_clk_net_3_r_10,blif_reset_net_3_r_10;
output n_429_or_0_3_r_10,G78_3_r_10,n_576_3_r_10,n_102_3_r_10,n_547_3_r_10,G42_4_r_10,n_572_4_r_10,n_573_4_r_10,n_549_4_r_10,n_569_4_r_10,n_452_4_r_10;
wire n_429_or_0_3_r_13,G78_3_r_13,n_576_3_r_13,n_102_3_r_13,n_547_3_r_13,G42_4_r_13,n_572_4_r_13,n_573_4_r_13,n_549_4_r_13,n_569_4_r_13,n_452_4_r_13,ACVQN1_2_l_13,P6_2_l_13,P6_internal_2_l_13,n_429_or_0_3_l_13,n12_3_l_13,n_431_3_l_13,G78_3_l_13,n_576_3_l_13,n11_3_l_13,n_102_3_l_13,n_547_3_l_13,n13_3_l_13,n14_3_l_13,n15_3_l_13,n16_3_l_13,n12_3_r_13,n_431_3_r_13,n11_3_r_13,n13_3_r_13,n14_3_r_13,n15_3_r_13,n16_3_r_13,n4_4_r_13,n_87_4_r_13,n7_4_r_13,n2_3_r_10,ACVQN2_0_l_10,n_266_and_0_0_l_10,ACVQN1_0_l_10,n4_4_l_10,G42_4_l_10,n_87_4_l_10,n_572_4_l_10,n_573_4_l_10,n_549_4_l_10,n7_4_l_10,n_569_4_l_10,n_452_4_l_10,n12_3_r_10,n_431_3_r_10,n11_3_r_10,n13_3_r_10,n14_3_r_10,n15_3_r_10,n16_3_r_10,n4_4_r_10,n_87_4_r_10,n7_4_r_10;
nand I_0(n_429_or_0_3_r_13,n_429_or_0_3_l_13,n12_3_r_13);
DFFARX1 I_1(n_431_3_r_13,blif_clk_net_3_r_10,n2_3_r_10,G78_3_r_13,);
nand I_2(n_576_3_r_13,n_547_3_l_13,n11_3_r_13);
not I_3(n_102_3_r_13,ACVQN1_2_l_13);
nand I_4(n_547_3_r_13,P6_2_l_13,n13_3_r_13);
DFFARX1 I_5(n4_4_r_13,blif_clk_net_3_r_10,n2_3_r_10,G42_4_r_13,);
nor I_6(n_572_4_r_13,P6_2_l_13,n_429_or_0_3_l_13);
or I_7(n_573_4_r_13,ACVQN1_2_l_13,G78_3_l_13);
nor I_8(n_549_4_r_13,n_429_or_0_3_l_13,n7_4_r_13);
or I_9(n_569_4_r_13,n_429_or_0_3_l_13,G78_3_l_13);
nor I_10(n_452_4_r_13,ACVQN1_2_l_13,P6_2_l_13);
DFFARX1 I_11(IN_2_2_l_13,blif_clk_net_3_r_10,n2_3_r_10,ACVQN1_2_l_13,);
not I_12(P6_2_l_13,P6_internal_2_l_13);
DFFARX1 I_13(IN_1_2_l_13,blif_clk_net_3_r_10,n2_3_r_10,P6_internal_2_l_13,);
nand I_14(n_429_or_0_3_l_13,G1_3_l_13,n12_3_l_13);
not I_15(n12_3_l_13,IN_5_3_l_13);
or I_16(n_431_3_l_13,IN_8_3_l_13,n14_3_l_13);
DFFARX1 I_17(n_431_3_l_13,blif_clk_net_3_r_10,n2_3_r_10,G78_3_l_13,);
nand I_18(n_576_3_l_13,IN_7_3_l_13,n11_3_l_13);
nor I_19(n11_3_l_13,G2_3_l_13,n12_3_l_13);
not I_20(n_102_3_l_13,G2_3_l_13);
nand I_21(n_547_3_l_13,IN_11_3_l_13,n13_3_l_13);
nor I_22(n13_3_l_13,G2_3_l_13,IN_10_3_l_13);
and I_23(n14_3_l_13,IN_2_3_l_13,n15_3_l_13);
nor I_24(n15_3_l_13,IN_4_3_l_13,n16_3_l_13);
not I_25(n16_3_l_13,G1_3_l_13);
not I_26(n12_3_r_13,n_102_3_l_13);
or I_27(n_431_3_r_13,ACVQN1_2_l_13,n14_3_r_13);
nor I_28(n11_3_r_13,ACVQN1_2_l_13,n12_3_r_13);
nor I_29(n13_3_r_13,ACVQN1_2_l_13,n_576_3_l_13);
and I_30(n14_3_r_13,n_102_3_l_13,n15_3_r_13);
nor I_31(n15_3_r_13,G78_3_l_13,n16_3_r_13);
not I_32(n16_3_r_13,n_429_or_0_3_l_13);
nor I_33(n4_4_r_13,P6_2_l_13,n_547_3_l_13);
not I_34(n_87_4_r_13,P6_2_l_13);
and I_35(n7_4_r_13,n_576_3_l_13,n_87_4_r_13);
nand I_36(n_429_or_0_3_r_10,n_266_and_0_0_l_10,n12_3_r_10);
DFFARX1 I_37(n_431_3_r_10,blif_clk_net_3_r_10,n2_3_r_10,G78_3_r_10,);
nand I_38(n_576_3_r_10,ACVQN2_0_l_10,n11_3_r_10);
not I_39(n_102_3_r_10,G42_4_l_10);
nand I_40(n_547_3_r_10,n_569_4_l_10,n13_3_r_10);
DFFARX1 I_41(n4_4_r_10,blif_clk_net_3_r_10,n2_3_r_10,G42_4_r_10,);
nor I_42(n_572_4_r_10,ACVQN2_0_l_10,n_573_4_l_10);
or I_43(n_573_4_r_10,n_569_4_l_10,n_452_4_l_10);
nor I_44(n_549_4_r_10,n_572_4_l_10,n7_4_r_10);
or I_45(n_569_4_r_10,n_572_4_l_10,n_569_4_l_10);
nor I_46(n_452_4_r_10,n_266_and_0_0_l_10,n_452_4_l_10);
not I_47(n2_3_r_10,blif_reset_net_3_r_10);
DFFARX1 I_48(n_102_3_r_13,blif_clk_net_3_r_10,n2_3_r_10,ACVQN2_0_l_10,);
and I_49(n_266_and_0_0_l_10,ACVQN1_0_l_10,n_573_4_r_13);
DFFARX1 I_50(n_547_3_r_13,blif_clk_net_3_r_10,n2_3_r_10,ACVQN1_0_l_10,);
nor I_51(n4_4_l_10,n_429_or_0_3_r_13,G42_4_r_13);
DFFARX1 I_52(n4_4_l_10,blif_clk_net_3_r_10,n2_3_r_10,G42_4_l_10,);
not I_53(n_87_4_l_10,n_572_4_r_13);
nor I_54(n_572_4_l_10,n_572_4_r_13,n_569_4_r_13);
or I_55(n_573_4_l_10,G78_3_r_13,n_549_4_r_13);
nor I_56(n_549_4_l_10,n7_4_l_10,n_576_3_r_13);
and I_57(n7_4_l_10,n_87_4_l_10,n_452_4_r_13);
or I_58(n_569_4_l_10,G78_3_r_13,n_576_3_r_13);
nor I_59(n_452_4_l_10,G42_4_r_13,n_549_4_r_13);
not I_60(n12_3_r_10,n_549_4_l_10);
or I_61(n_431_3_r_10,n_572_4_l_10,n14_3_r_10);
nor I_62(n11_3_r_10,G42_4_l_10,n12_3_r_10);
nor I_63(n13_3_r_10,G42_4_l_10,n_549_4_l_10);
and I_64(n14_3_r_10,ACVQN2_0_l_10,n15_3_r_10);
nor I_65(n15_3_r_10,n_573_4_l_10,n16_3_r_10);
not I_66(n16_3_r_10,n_266_and_0_0_l_10);
nor I_67(n4_4_r_10,n_266_and_0_0_l_10,G42_4_l_10);
not I_68(n_87_4_r_10,ACVQN2_0_l_10);
and I_69(n7_4_r_10,n_452_4_l_10,n_87_4_r_10);
endmodule


