module test_final(IN_1_0_l_11,IN_2_0_l_11,IN_4_0_l_11,IN_1_1_l_11,IN_2_1_l_11,IN_3_1_l_11,IN_6_1_l_11,IN_1_5_l_11,IN_2_5_l_11,IN_3_5_l_11,IN_6_5_l_11,blif_clk_net_3_r_10,blif_reset_net_3_r_10,n_429_or_0_3_r_10,G78_3_r_10,n_576_3_r_10,n_102_3_r_10,n_547_3_r_10,G42_4_r_10,n_572_4_r_10,n_573_4_r_10,n_549_4_r_10,n_569_4_r_10,n_452_4_r_10);
input IN_1_0_l_11,IN_2_0_l_11,IN_4_0_l_11,IN_1_1_l_11,IN_2_1_l_11,IN_3_1_l_11,IN_6_1_l_11,IN_1_5_l_11,IN_2_5_l_11,IN_3_5_l_11,IN_6_5_l_11,blif_clk_net_3_r_10,blif_reset_net_3_r_10;
output n_429_or_0_3_r_10,G78_3_r_10,n_576_3_r_10,n_102_3_r_10,n_547_3_r_10,G42_4_r_10,n_572_4_r_10,n_573_4_r_10,n_549_4_r_10,n_569_4_r_10,n_452_4_r_10;
wire G199_1_r_11,G214_1_r_11,ACVQN1_2_r_11,P6_2_r_11,n_429_or_0_3_r_11,G78_3_r_11,n_576_3_r_11,n_102_3_r_11,n_547_3_r_11,n_42_5_r_11,G199_5_r_11,ACVQN2_0_l_11,n_266_and_0_0_l_11,ACVQN1_0_l_11,N1_1_l_11,G199_1_l_11,G214_1_l_11,n3_1_l_11,n_42_5_l_11,N3_5_l_11,G199_5_l_11,n3_5_l_11,N1_1_r_11,n3_1_r_11,P6_internal_2_r_11,n12_3_r_11,n_431_3_r_11,n11_3_r_11,n13_3_r_11,n14_3_r_11,n15_3_r_11,n16_3_r_11,N3_5_r_11,n3_5_r_11,n2_3_r_10,ACVQN2_0_l_10,n_266_and_0_0_l_10,ACVQN1_0_l_10,n4_4_l_10,G42_4_l_10,n_87_4_l_10,n_572_4_l_10,n_573_4_l_10,n_549_4_l_10,n7_4_l_10,n_569_4_l_10,n_452_4_l_10,n12_3_r_10,n_431_3_r_10,n11_3_r_10,n13_3_r_10,n14_3_r_10,n15_3_r_10,n16_3_r_10,n4_4_r_10,n_87_4_r_10,n7_4_r_10;
DFFARX1 I_0(N1_1_r_11,blif_clk_net_3_r_10,n2_3_r_10,G199_1_r_11,);
DFFARX1 I_1(ACVQN2_0_l_11,blif_clk_net_3_r_10,n2_3_r_10,G214_1_r_11,);
DFFARX1 I_2(G214_1_l_11,blif_clk_net_3_r_10,n2_3_r_10,ACVQN1_2_r_11,);
not I_3(P6_2_r_11,P6_internal_2_r_11);
nand I_4(n_429_or_0_3_r_11,ACVQN2_0_l_11,n12_3_r_11);
DFFARX1 I_5(n_431_3_r_11,blif_clk_net_3_r_10,n2_3_r_10,G78_3_r_11,);
nand I_6(n_576_3_r_11,G199_1_l_11,n11_3_r_11);
not I_7(n_102_3_r_11,n_42_5_l_11);
nand I_8(n_547_3_r_11,G214_1_l_11,n13_3_r_11);
nor I_9(n_42_5_r_11,G199_1_l_11,G199_5_l_11);
DFFARX1 I_10(N3_5_r_11,blif_clk_net_3_r_10,n2_3_r_10,G199_5_r_11,);
DFFARX1 I_11(IN_1_0_l_11,blif_clk_net_3_r_10,n2_3_r_10,ACVQN2_0_l_11,);
and I_12(n_266_and_0_0_l_11,IN_4_0_l_11,ACVQN1_0_l_11);
DFFARX1 I_13(IN_2_0_l_11,blif_clk_net_3_r_10,n2_3_r_10,ACVQN1_0_l_11,);
and I_14(N1_1_l_11,IN_6_1_l_11,n3_1_l_11);
DFFARX1 I_15(N1_1_l_11,blif_clk_net_3_r_10,n2_3_r_10,G199_1_l_11,);
DFFARX1 I_16(IN_3_1_l_11,blif_clk_net_3_r_10,n2_3_r_10,G214_1_l_11,);
nand I_17(n3_1_l_11,IN_1_1_l_11,IN_2_1_l_11);
nor I_18(n_42_5_l_11,IN_1_5_l_11,IN_3_5_l_11);
and I_19(N3_5_l_11,IN_6_5_l_11,n3_5_l_11);
DFFARX1 I_20(N3_5_l_11,blif_clk_net_3_r_10,n2_3_r_10,G199_5_l_11,);
nand I_21(n3_5_l_11,IN_2_5_l_11,IN_3_5_l_11);
and I_22(N1_1_r_11,G199_5_l_11,n3_1_r_11);
nand I_23(n3_1_r_11,n_266_and_0_0_l_11,G199_1_l_11);
DFFARX1 I_24(n_266_and_0_0_l_11,blif_clk_net_3_r_10,n2_3_r_10,P6_internal_2_r_11,);
not I_25(n12_3_r_11,G214_1_l_11);
or I_26(n_431_3_r_11,n_266_and_0_0_l_11,n14_3_r_11);
nor I_27(n11_3_r_11,n_42_5_l_11,n12_3_r_11);
nor I_28(n13_3_r_11,n_42_5_l_11,G199_5_l_11);
and I_29(n14_3_r_11,ACVQN2_0_l_11,n15_3_r_11);
nor I_30(n15_3_r_11,n_42_5_l_11,n16_3_r_11);
not I_31(n16_3_r_11,ACVQN2_0_l_11);
and I_32(N3_5_r_11,G199_1_l_11,n3_5_r_11);
nand I_33(n3_5_r_11,ACVQN2_0_l_11,G199_5_l_11);
nand I_34(n_429_or_0_3_r_10,n_266_and_0_0_l_10,n12_3_r_10);
DFFARX1 I_35(n_431_3_r_10,blif_clk_net_3_r_10,n2_3_r_10,G78_3_r_10,);
nand I_36(n_576_3_r_10,ACVQN2_0_l_10,n11_3_r_10);
not I_37(n_102_3_r_10,G42_4_l_10);
nand I_38(n_547_3_r_10,n_569_4_l_10,n13_3_r_10);
DFFARX1 I_39(n4_4_r_10,blif_clk_net_3_r_10,n2_3_r_10,G42_4_r_10,);
nor I_40(n_572_4_r_10,ACVQN2_0_l_10,n_573_4_l_10);
or I_41(n_573_4_r_10,n_569_4_l_10,n_452_4_l_10);
nor I_42(n_549_4_r_10,n_572_4_l_10,n7_4_r_10);
or I_43(n_569_4_r_10,n_572_4_l_10,n_569_4_l_10);
nor I_44(n_452_4_r_10,n_266_and_0_0_l_10,n_452_4_l_10);
not I_45(n2_3_r_10,blif_reset_net_3_r_10);
DFFARX1 I_46(n_429_or_0_3_r_11,blif_clk_net_3_r_10,n2_3_r_10,ACVQN2_0_l_10,);
and I_47(n_266_and_0_0_l_10,ACVQN1_0_l_10,n_547_3_r_11);
DFFARX1 I_48(n_42_5_r_11,blif_clk_net_3_r_10,n2_3_r_10,ACVQN1_0_l_10,);
nor I_49(n4_4_l_10,G199_1_r_11,ACVQN1_2_r_11);
DFFARX1 I_50(n4_4_l_10,blif_clk_net_3_r_10,n2_3_r_10,G42_4_l_10,);
not I_51(n_87_4_l_10,G199_5_r_11);
nor I_52(n_572_4_l_10,n_576_3_r_11,G199_5_r_11);
or I_53(n_573_4_l_10,P6_2_r_11,n_102_3_r_11);
nor I_54(n_549_4_l_10,n7_4_l_10,G78_3_r_11);
and I_55(n7_4_l_10,n_87_4_l_10,G214_1_r_11);
or I_56(n_569_4_l_10,G78_3_r_11,n_102_3_r_11);
nor I_57(n_452_4_l_10,ACVQN1_2_r_11,P6_2_r_11);
not I_58(n12_3_r_10,n_549_4_l_10);
or I_59(n_431_3_r_10,n_572_4_l_10,n14_3_r_10);
nor I_60(n11_3_r_10,G42_4_l_10,n12_3_r_10);
nor I_61(n13_3_r_10,G42_4_l_10,n_549_4_l_10);
and I_62(n14_3_r_10,ACVQN2_0_l_10,n15_3_r_10);
nor I_63(n15_3_r_10,n_573_4_l_10,n16_3_r_10);
not I_64(n16_3_r_10,n_266_and_0_0_l_10);
nor I_65(n4_4_r_10,n_266_and_0_0_l_10,G42_4_l_10);
not I_66(n_87_4_r_10,ACVQN2_0_l_10);
and I_67(n7_4_r_10,n_452_4_l_10,n_87_4_r_10);
endmodule


