module test_I8360(I5864,I1477,I4527,I1470,I8360);
input I5864,I1477,I4527,I1470;
output I8360;
wire I6265,I6248,I5751,I6203,I5915,I5719;
and I_0(I6265,I5915,I6248);
nand I_1(I6248,I6203,I5864);
not I_2(I8360,I5719);
not I_3(I5751,I1477);
DFFARX1 I_4(I1470,I5751,,,I6203,);
DFFARX1 I_5(I4527,I1470,I5751,,,I5915,);
DFFARX1 I_6(I6265,I1470,I5751,,,I5719,);
endmodule


