module test_final(IN_1_1_l_7,IN_2_1_l_7,IN_3_1_l_7,G18_7_l_7,G15_7_l_7,IN_1_7_l_7,IN_4_7_l_7,IN_5_7_l_7,IN_7_7_l_7,IN_9_7_l_7,IN_10_7_l_7,IN_1_8_l_7,IN_2_8_l_7,IN_3_8_l_7,IN_6_8_l_7,blif_clk_net_8_r_6,blif_reset_net_8_r_6,N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,N1372_10_r_6,N1508_10_r_6);
input IN_1_1_l_7,IN_2_1_l_7,IN_3_1_l_7,G18_7_l_7,G15_7_l_7,IN_1_7_l_7,IN_4_7_l_7,IN_5_7_l_7,IN_7_7_l_7,IN_9_7_l_7,IN_10_7_l_7,IN_1_8_l_7,IN_2_8_l_7,IN_3_8_l_7,IN_6_8_l_7,blif_clk_net_8_r_6,blif_reset_net_8_r_6;
output N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,N1372_10_r_6,N1508_10_r_6;
wire N1371_0_r_7,N1508_0_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_102_5_r_7,n_547_5_r_7,G42_7_r_7,n_572_7_r_7,n_573_7_r_7,n_549_7_r_7,n_569_7_r_7,n_452_7_r_7,n4_7_l_7,n53_7,n30_7,N3_8_l_7,n54_7,n_431_5_r_7,n4_7_r_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7,n43_7,n44_7,n45_7,n46_7,n47_7,n48_7,n49_7,n50_7,n51_7,n52_7,I_BUFF_1_9_r_6,N3_8_r_6,n9_6,n30_6,n31_6,n32_6,n33_6,n34_6,n35_6,n36_6,n37_6,n38_6,n39_6,n40_6,n41_6,n42_6,n43_6,n44_6,n45_6,n46_6,n47_6,n48_6,n49_6,n50_6,n51_6,n52_6,n53_6,n54_6;
nor I_0(N1371_0_r_7,n53_7,n52_7);
nor I_1(N1508_0_r_7,n51_7,n52_7);
nand I_2(n_429_or_0_5_r_7,n43_7,n48_7);
DFFARX1 I_3(n_431_5_r_7,blif_clk_net_8_r_6,n9_6,G78_5_r_7,);
nand I_4(n_576_5_r_7,n31_7,n32_7);
nor I_5(n_102_5_r_7,IN_5_7_l_7,IN_9_7_l_7);
nand I_6(n_547_5_r_7,n31_7,n38_7);
DFFARX1 I_7(n4_7_r_7,blif_clk_net_8_r_6,n9_6,G42_7_r_7,);
nor I_8(n_572_7_r_7,n54_7,n33_7);
nand I_9(n_573_7_r_7,n_102_5_r_7,n_452_7_r_7);
nor I_10(n_549_7_r_7,n53_7,n36_7);
nand I_11(n_569_7_r_7,n_102_5_r_7,n30_7);
nand I_12(n_452_7_r_7,IN_1_1_l_7,IN_2_1_l_7);
nor I_13(n4_7_l_7,G18_7_l_7,IN_1_7_l_7);
DFFARX1 I_14(n4_7_l_7,blif_clk_net_8_r_6,n9_6,n53_7,);
not I_15(n30_7,n53_7);
and I_16(N3_8_l_7,IN_6_8_l_7,n50_7);
DFFARX1 I_17(N3_8_l_7,blif_clk_net_8_r_6,n9_6,n54_7,);
nand I_18(n_431_5_r_7,n40_7,n41_7);
nor I_19(n4_7_r_7,n54_7,n49_7);
and I_20(n31_7,n_102_5_r_7,n39_7);
not I_21(n32_7,G18_7_l_7);
nor I_22(n33_7,IN_10_7_l_7,n34_7);
and I_23(n34_7,IN_4_7_l_7,n35_7);
not I_24(n35_7,G15_7_l_7);
nor I_25(n36_7,G18_7_l_7,n37_7);
or I_26(n37_7,IN_5_7_l_7,n54_7);
or I_27(n38_7,IN_1_8_l_7,IN_3_8_l_7);
nor I_28(n39_7,IN_3_1_l_7,n_452_7_r_7);
nand I_29(n40_7,n46_7,n47_7);
nand I_30(n41_7,n42_7,n43_7);
nor I_31(n42_7,n44_7,n45_7);
nor I_32(n43_7,IN_1_8_l_7,IN_3_8_l_7);
nor I_33(n44_7,G15_7_l_7,IN_7_7_l_7);
nor I_34(n45_7,IN_9_7_l_7,IN_10_7_l_7);
nand I_35(n46_7,IN_4_7_l_7,n35_7);
not I_36(n47_7,IN_10_7_l_7);
or I_37(n48_7,IN_3_1_l_7,n_452_7_r_7);
not I_38(n49_7,n_452_7_r_7);
nand I_39(n50_7,IN_2_8_l_7,IN_3_8_l_7);
and I_40(n51_7,n_452_7_r_7,n45_7);
not I_41(n52_7,n44_7);
nor I_42(N1371_0_r_6,n30_6,n33_6);
nor I_43(N1508_0_r_6,n33_6,n44_6);
not I_44(N1372_1_r_6,n41_6);
nor I_45(N1508_1_r_6,n40_6,n41_6);
nor I_46(N1507_6_r_6,n39_6,n45_6);
nor I_47(N1508_6_r_6,n37_6,n38_6);
nor I_48(n_42_8_r_6,n30_6,n31_6);
DFFARX1 I_49(N3_8_r_6,blif_clk_net_8_r_6,n9_6,G199_8_r_6,);
nor I_50(N6147_9_r_6,n32_6,n33_6);
nor I_51(N6134_9_r_6,I_BUFF_1_9_r_6,n35_6);
not I_52(I_BUFF_1_9_r_6,n37_6);
not I_53(N1372_10_r_6,n43_6);
nor I_54(N1508_10_r_6,n42_6,n43_6);
nor I_55(N3_8_r_6,n36_6,N1371_0_r_7);
not I_56(n9_6,blif_reset_net_8_r_6);
nor I_57(n30_6,n53_6,n_569_7_r_7);
not I_58(n31_6,n36_6);
nor I_59(n32_6,I_BUFF_1_9_r_6,n34_6);
not I_60(n33_6,N1371_0_r_7);
not I_61(n34_6,n35_6);
nand I_62(n35_6,n49_6,N1371_0_r_7);
nand I_63(n36_6,n51_6,n_549_7_r_7);
nand I_64(n37_6,n54_6,N1508_0_r_7);
or I_65(n38_6,n35_6,n39_6);
nor I_66(n39_6,n40_6,n45_6);
and I_67(n40_6,n46_6,n47_6);
nand I_68(n41_6,n30_6,n31_6);
nor I_69(n42_6,n34_6,n40_6);
nand I_70(n43_6,n30_6,N1371_0_r_7);
nor I_71(n44_6,n31_6,n40_6);
nor I_72(n45_6,n35_6,n36_6);
nor I_73(n46_6,n_572_7_r_7,n_429_or_0_5_r_7);
or I_74(n47_6,n48_6,G42_7_r_7);
nor I_75(n48_6,G78_5_r_7,N1508_0_r_7);
and I_76(n49_6,n50_6,n_429_or_0_5_r_7);
nand I_77(n50_6,n51_6,n52_6);
nand I_78(n51_6,n_547_5_r_7,G78_5_r_7);
not I_79(n52_6,n_549_7_r_7);
nor I_80(n53_6,n_576_5_r_7,n_573_7_r_7);
or I_81(n54_6,n_576_5_r_7,n_573_7_r_7);
endmodule


