module test_final(IN_1_1_l,IN_2_1_l,IN_3_1_l,IN_1_3_l,IN_2_3_l,IN_3_3_l,IN_1_6_l,IN_2_6_l,IN_3_6_l,IN_4_6_l,IN_5_6_l,IN_1_8_l,IN_2_8_l,IN_3_8_l,IN_6_8_l,blif_clk_net_7_r,blif_reset_net_7_r,N6147_2_r,N6147_3_r,N1507_6_r,N1508_6_r,G42_7_r,n_572_7_r,n_573_7_r,n_549_7_r,n_569_7_r,n_452_7_r,N6147_9_r,N6134_9_r,I_BUFF_1_9_r);
input IN_1_1_l,IN_2_1_l,IN_3_1_l,IN_1_3_l,IN_2_3_l,IN_3_3_l,IN_1_6_l,IN_2_6_l,IN_3_6_l,IN_4_6_l,IN_5_6_l,IN_1_8_l,IN_2_8_l,IN_3_8_l,IN_6_8_l,blif_clk_net_7_r,blif_reset_net_7_r;
output N6147_2_r,N6147_3_r,N1507_6_r,N1508_6_r,G42_7_r,n_572_7_r,n_573_7_r,n_549_7_r,n_569_7_r,n_452_7_r,N6147_9_r,N6134_9_r,I_BUFF_1_9_r;
wire N1372_1_l,N1508_1_l,n4_1_l,N6147_3_l,n3_3_l,N6138_3_l,N1507_6_l,N1508_6_l,n6_6_l,n7_6_l,n8_6_l,n9_6_l,n_42_8_l,G199_8_l,N3_8_l,n3_8_l,n5_2_r,n6_2_r,N6138_2_r,n7_2_r,n3_3_r,N6138_3_r,n6_6_r,n7_6_r,n8_6_r,n9_6_r,n_87_7_r,n4_7_r,n2_7_r,n7_7_r,N6150_9_r,n3_9_r;
not I_0(N1372_1_l,n4_1_l);
nor I_1(N1508_1_l,IN_3_1_l,n4_1_l);
nand I_2(n4_1_l,IN_1_1_l,IN_2_1_l);
nor I_3(N6147_3_l,IN_3_3_l,n3_3_l);
not I_4(n3_3_l,N6138_3_l);
nor I_5(N6138_3_l,IN_1_3_l,IN_2_3_l);
nor I_6(N1507_6_l,n8_6_l,n9_6_l);
and I_7(N1508_6_l,IN_2_6_l,n6_6_l);
nor I_8(n6_6_l,n7_6_l,n8_6_l);
not I_9(n7_6_l,IN_1_6_l);
nor I_10(n8_6_l,IN_5_6_l,n9_6_l);
and I_11(n9_6_l,IN_3_6_l,IN_4_6_l);
nor I_12(n_42_8_l,IN_1_8_l,IN_3_8_l);
DFFARX1 I_13(N3_8_l,blif_clk_net_7_r,n2_7_r,G199_8_l,);
and I_14(N3_8_l,IN_6_8_l,n3_8_l);
nand I_15(n3_8_l,IN_2_8_l,IN_3_8_l);
nor I_16(N6147_2_r,n5_2_r,n6_2_r);
nor I_17(n5_2_r,n7_2_r,N1372_1_l);
not I_18(n6_2_r,N6138_2_r);
nor I_19(N6138_2_r,N1507_6_l,N1508_6_l);
nor I_20(n7_2_r,N1508_6_l,G199_8_l);
nor I_21(N6147_3_r,n3_3_r,N1508_6_l);
not I_22(n3_3_r,N6138_3_r);
nor I_23(N6138_3_r,N6147_3_l,N1508_1_l);
nor I_24(N1507_6_r,n8_6_r,n9_6_r);
and I_25(N1508_6_r,n6_6_r,N1507_6_l);
nor I_26(n6_6_r,n7_6_r,n8_6_r);
not I_27(n7_6_r,N1508_1_l);
nor I_28(n8_6_r,n9_6_r,G199_8_l);
and I_29(n9_6_r,N1508_1_l,N6147_3_l);
DFFARX1 I_30(n4_7_r,blif_clk_net_7_r,n2_7_r,G42_7_r,);
not I_31(n_87_7_r,N1372_1_l);
nor I_32(n_572_7_r,N1508_6_l,N1372_1_l);
or I_33(n_573_7_r,n_42_8_l,N1507_6_l);
nor I_34(n_549_7_r,n7_7_r,G199_8_l);
or I_35(n_569_7_r,n_42_8_l,G199_8_l);
nor I_36(n_452_7_r,N1508_1_l,N1507_6_l);
nor I_37(n4_7_r,N1508_1_l,n_42_8_l);
not I_38(n2_7_r,blif_reset_net_7_r);
and I_39(n7_7_r,n_87_7_r,N1372_1_l);
not I_40(N6150_9_r,N1372_1_l);
nor I_41(N6147_9_r,N6150_9_r,n3_9_r);
nor I_42(N6134_9_r,n3_9_r,N6147_3_l);
nor I_43(n3_9_r,n_42_8_l,N6147_3_l);
buf I_44(I_BUFF_1_9_r,N1507_6_l);
endmodule


