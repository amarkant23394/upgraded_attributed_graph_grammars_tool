module test_I1489(I1733,I1477,I1279,I1470,I1489);
input I1733,I1477,I1279,I1470;
output I1489;
wire I1518,I1750,I1801,I1767;
not I_0(I1518,I1477);
or I_1(I1750,I1733,I1279);
DFFARX1 I_2(I1767,I1470,I1518,,,I1801,);
not I_3(I1489,I1801);
DFFARX1 I_4(I1750,I1470,I1518,,,I1767,);
endmodule


