module test_I12913(I9462,I10715,I9465,I10862,I1477,I1470,I12913);
input I9462,I10715,I9465,I10862,I1477,I1470;
output I12913;
wire I12619,I10879,I10647,I10633,I9468,I10896,I11009,I10732,I11026;
not I_0(I12619,I1477);
or I_1(I10879,I10862,I9462);
not I_2(I10647,I1477);
DFFARX1 I_3(I10633,I1470,I12619,,,I12913,);
nand I_4(I10633,I10896,I11026);
DFFARX1 I_5(I1470,,,I9468,);
DFFARX1 I_6(I10879,I1470,I10647,,,I10896,);
DFFARX1 I_7(I9468,I1470,I10647,,,I11009,);
nand I_8(I10732,I10715,I9465);
nor I_9(I11026,I11009,I10732);
endmodule


