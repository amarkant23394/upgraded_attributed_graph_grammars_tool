module Benchmark_testing1000(I76,I84,I92,I100,I108,I116,I124,I132,I140,I148,I156,I164,I172,I180,I188,I196,I204,I212,I220,I228,I236,I244,I251,I258,I11292,I11373,I11391,I11427,I11445,I11517,I11634,I11652,I11724,I22785,I22902,I22992,I23019,I23082,I23109,I23127,I23145,I23172);
input I76,I84,I92,I100,I108,I116,I124,I132,I140,I148,I156,I164,I172,I180,I188,I196,I204,I212,I220,I228,I236,I244,I251,I258;
output I11292,I11373,I11391,I11427,I11445,I11517,I11634,I11652,I11724,I22785,I22902,I22992,I23019,I23082,I23109,I23127,I23145,I23172;
wire I76,I84,I92,I100,I108,I116,I124,I132,I140,I148,I156,I164,I172,I180,I188,I196,I204,I212,I220,I228,I236,I244,I251,I258,I267,I294,I303,I321,I339,I366,I384,I402,I411,I429,I456,I465,I483,I510,I519,I537,I555,I573,I600,I609,I627,I645,I663,I681,I699,I726,I735,I762,I771,I789,I807,I825,I852,I861,I879,I897,I924,I933,I960,I969,I987,I1005,I1023,I1041,I1068,I1077,I1095,I1113,I1131,I1158,I1167,I1185,I1212,I1221,I1248,I1257,I1275,I1293,I1311,I1338,I1347,I1365,I1383,I1401,I1428,I1437,I1464,I1482,I1491,I1509,I1536,I1545,I1563,I1581,I1599,I1617,I1635,I1653,I1671,I1698,I1707,I1725,I1743,I1761,I1779,I1797,I1815,I1842,I1860,I1869,I1887,I1905,I1923,I1950,I1959,I1977,I1995,I2022,I2031,I2049,I2067,I2094,I2112,I2121,I2139,I2166,I2175,I2193,I2211,I2229,I2247,I2265,I2283,I2310,I2319,I2337,I2355,I2382,I2391,I2409,I2427,I2454,I2463,I2490,I2499,I2517,I2535,I2553,I2571,I2598,I2607,I2625,I2643,I2661,I2679,I2697,I2724,I2733,I2760,I2778,I2787,I2805,I2823,I2841,I2868,I2877,I2895,I2913,I2940,I2949,I2967,I2985,I3003,I3021,I3048,I3066,I3075,I3093,I3111,I3129,I3156,I3165,I3183,I3201,I3219,I3237,I3255,I3273,I3291,I3309,I3336,I3354,I3363,I3381,I3408,I3417,I3435,I3453,I3471,I3489,I3507,I3525,I3543,I3570,I3579,I3597,I3615,I3633,I3651,I3669,I3687,I3714,I3732,I3741,I3759,I3777,I3795,I3822,I3831,I3849,I3867,I3894,I3903,I3921,I3939,I3966,I3975,I3993,I4020,I4029,I4047,I4074,I4083,I4101,I4128,I4137,I4155,I4173,I4200,I4218,I4227,I4245,I4263,I4281,I4299,I4326,I4335,I4362,I4380,I4389,I4407,I4425,I4443,I4461,I4488,I4497,I4524,I4542,I4551,I4569,I4596,I4605,I4623,I4641,I4659,I4677,I4695,I4713,I4740,I4749,I4767,I4785,I4812,I4821,I4839,I4857,I4884,I4893,I4920,I4929,I4947,I4965,I4983,I5001,I5028,I5037,I5055,I5073,I5091,I5109,I5127,I5154,I5163,I5181,I5199,I5226,I5244,I5253,I5271,I5298,I5307,I5325,I5343,I5370,I5388,I5397,I5415,I5442,I5460,I5469,I5487,I5505,I5523,I5541,I5559,I5577,I5604,I5613,I5631,I5649,I5667,I5685,I5712,I5730,I5739,I5757,I5784,I5793,I5811,I5829,I5847,I5865,I5883,I5901,I5928,I5937,I5955,I5973,I6000,I6009,I6027,I6045,I6072,I6081,I6108,I6117,I6135,I6153,I6171,I6189,I6216,I6225,I6243,I6261,I6279,I6297,I6315,I6342,I6360,I6369,I6387,I6414,I6423,I6441,I6459,I6477,I6495,I6513,I6531,I6549,I6567,I6585,I6603,I6621,I6639,I6657,I6684,I6693,I6720,I6729,I6747,I6765,I6783,I6810,I6819,I6846,I6855,I6873,I6891,I6909,I6936,I6954,I6963,I6981,I6999,I7017,I7035,I7053,I7080,I7089,I7107,I7134,I7143,I7161,I7179,I7206,I7215,I7233,I7260,I7269,I7287,I7305,I7323,I7341,I7359,I7377,I7395,I7422,I7431,I7449,I7467,I7485,I7503,I7521,I7539,I7557,I7575,I7593,I7620,I7629,I7647,I7674,I7683,I7701,I7728,I7737,I7755,I7782,I7791,I7809,I7827,I7854,I7872,I7881,I7899,I7917,I7935,I7953,I7980,I7989,I8016,I8034,I8043,I8061,I8079,I8097,I8115,I8142,I8151,I8178,I8196,I8205,I8223,I8250,I8259,I8277,I8295,I8313,I8331,I8349,I8367,I8394,I8403,I8421,I8439,I8466,I8475,I8493,I8511,I8538,I8547,I8574,I8583,I8601,I8619,I8637,I8655,I8682,I8691,I8709,I8727,I8745,I8763,I8781,I8808,I8817,I8835,I8853,I8880,I8889,I8916,I8925,I8943,I8961,I8979,I8997,I9024,I9033,I9051,I9069,I9087,I9114,I9123,I9141,I9168,I9177,I9204,I9213,I9231,I9249,I9267,I9294,I9303,I9321,I9339,I9357,I9384,I9393,I9420,I9429,I9447,I9474,I9483,I9501,I9528,I9537,I9555,I9582,I9591,I9609,I9627,I9654,I9672,I9681,I9699,I9717,I9735,I9753,I9780,I9789,I9816,I9834,I9843,I9861,I9879,I9897,I9915,I9942,I9951,I9978,I9987,I10005,I10023,I10050,I10059,I10086,I10095,I10113,I10131,I10149,I10167,I10194,I10203,I10221,I10239,I10257,I10284,I10293,I10311,I10338,I10347,I10374,I10383,I10401,I10419,I10437,I10464,I10473,I10491,I10509,I10527,I10554,I10563,I10590,I10599,I10617,I10635,I10662,I10680,I10689,I10707,I10734,I10743,I10761,I10779,I10806,I10824,I10833,I10851,I10878,I10896,I10905,I10923,I10941,I10959,I10977,I10995,I11013,I11040,I11049,I11067,I11085,I11103,I11121,I11148,I11157,I11184,I11193,I11211,I11229,I11247,I11265,I11301,I11319,I11337,I11355,I11409,I11463,I11481,I11499,I11535,I11553,I11571,I11598,I11607,I11661,I11679,I11697,I11733,I11760,I11769,I11787,I11814,I11823,I11841,I11859,I11877,I11895,I11922,I11931,I11949,I11967,I11985,I12003,I12021,I12039,I12066,I12075,I12093,I12111,I12129,I12147,I12165,I12192,I12201,I12228,I12237,I12264,I12282,I12291,I12309,I12327,I12345,I12372,I12381,I12408,I12426,I12435,I12453,I12471,I12489,I12516,I12525,I12543,I12561,I12588,I12597,I12615,I12633,I12651,I12669,I12696,I12714,I12723,I12741,I12759,I12777,I12804,I12813,I12831,I12849,I12867,I12885,I12903,I12921,I12939,I12957,I12984,I12993,I13011,I13029,I13056,I13065,I13092,I13101,I13119,I13137,I13155,I13173,I13200,I13209,I13227,I13245,I13263,I13290,I13299,I13317,I13344,I13353,I13380,I13389,I13407,I13425,I13443,I13470,I13479,I13497,I13515,I13533,I13560,I13569,I13596,I13605,I13623,I13650,I13659,I13677,I13704,I13713,I13731,I13758,I13767,I13785,I13803,I13830,I13848,I13857,I13875,I13893,I13911,I13929,I13956,I13965,I13992,I14010,I14019,I14037,I14055,I14073,I14091,I14118,I14127,I14154,I14172,I14181,I14199,I14226,I14235,I14253,I14271,I14289,I14307,I14325,I14343,I14370,I14379,I14397,I14415,I14442,I14451,I14469,I14487,I14514,I14523,I14550,I14559,I14577,I14595,I14613,I14631,I14658,I14667,I14685,I14703,I14721,I14739,I14757,I14784,I14802,I14811,I14829,I14847,I14865,I14892,I14901,I14928,I14937,I14955,I14973,I15000,I15009,I15036,I15045,I15063,I15081,I15108,I15117,I15135,I15153,I15171,I15198,I15207,I15225,I15243,I15261,I15279,I15306,I15324,I15333,I15360,I15378,I15387,I15405,I15432,I15441,I15459,I15477,I15495,I15513,I15531,I15549,I15576,I15585,I15603,I15621,I15648,I15657,I15675,I15693,I15720,I15729,I15756,I15765,I15783,I15801,I15819,I15837,I15864,I15873,I15891,I15909,I15927,I15945,I15963,I15990,I15999,I16017,I16035,I16062,I16071,I16098,I16107,I16125,I16143,I16161,I16179,I16206,I16215,I16233,I16251,I16269,I16296,I16305,I16323,I16350,I16359,I16386,I16395,I16413,I16431,I16449,I16476,I16485,I16503,I16521,I16539,I16566,I16575,I16602,I16620,I16629,I16656,I16665,I16683,I16701,I16719,I16737,I16755,I16773,I16800,I16809,I16827,I16845,I16863,I16890,I16899,I16917,I16935,I16953,I16971,I16998,I17007,I17025,I17043,I17070,I17079,I17097,I17115,I17133,I17160,I17169,I17187,I17205,I17232,I17241,I17268,I17286,I17295,I17313,I17331,I17349,I17376,I17385,I17403,I17421,I17448,I17457,I17475,I17493,I17511,I17529,I17556,I17574,I17583,I17601,I17619,I17637,I17664,I17673,I17691,I17709,I17727,I17745,I17763,I17781,I17799,I17817,I17844,I17853,I17871,I17889,I17916,I17925,I17952,I17961,I17979,I17997,I18015,I18033,I18060,I18069,I18087,I18105,I18123,I18150,I18159,I18177,I18204,I18213,I18240,I18249,I18267,I18285,I18303,I18330,I18339,I18357,I18375,I18393,I18420,I18429,I18456,I18465,I18483,I18510,I18519,I18537,I18564,I18573,I18591,I18618,I18627,I18645,I18663,I18690,I18708,I18717,I18735,I18753,I18771,I18789,I18816,I18825,I18852,I18870,I18879,I18897,I18915,I18933,I18951,I18978,I18987,I19014,I19032,I19041,I19059,I19077,I19095,I19122,I19131,I19158,I19167,I19185,I19203,I19230,I19239,I19266,I19275,I19293,I19311,I19338,I19347,I19365,I19383,I19401,I19428,I19437,I19455,I19473,I19491,I19509,I19536,I19554,I19563,I19590,I19599,I19617,I19644,I19653,I19671,I19698,I19707,I19725,I19752,I19761,I19779,I19797,I19824,I19842,I19851,I19869,I19887,I19905,I19923,I19950,I19959,I19986,I20004,I20013,I20031,I20049,I20067,I20085,I20112,I20121,I20148,I20157,I20184,I20202,I20211,I20229,I20247,I20265,I20283,I20301,I20319,I20337,I20355,I20373,I20391,I20409,I20436,I20445,I20463,I20481,I20508,I20517,I20535,I20553,I20580,I20589,I20607,I20625,I20652,I20661,I20679,I20697,I20724,I20733,I20751,I20769,I20796,I20814,I20832,I20841,I20859,I20886,I20895,I20913,I20940,I20949,I20967,I20985,I21003,I21030,I21039,I21057,I21075,I21093,I21111,I21129,I21156,I21165,I21192,I21201,I21219,I21237,I21255,I21282,I21300,I21309,I21327,I21345,I21363,I21381,I21399,I21426,I21435,I21453,I21480,I21489,I21507,I21525,I21552,I21561,I21579,I21606,I21615,I21633,I21651,I21669,I21687,I21705,I21723,I21741,I21768,I21777,I21795,I21813,I21831,I21849,I21867,I21885,I21903,I21921,I21939,I21966,I21984,I21993,I22011,I22038,I22047,I22065,I22083,I22101,I22119,I22137,I22155,I22182,I22191,I22209,I22227,I22254,I22263,I22281,I22299,I22326,I22335,I22362,I22371,I22389,I22407,I22425,I22443,I22470,I22479,I22497,I22515,I22533,I22551,I22569,I22596,I22605,I22623,I22641,I22668,I22677,I22704,I22713,I22731,I22749,I22767,I22812,I22821,I22839,I22857,I22875,I22911,I22929,I22956,I22965,I23001,I23037,I23055,I23091;
not I_0 (I267,I258);
DFFARX1 I_1 (I100,I251,I267,I294,);
not I_2 (I303,I294);
nand I_3 (I321,I140,I148);
and I_4 (I339,I321,I164);
DFFARX1 I_5 (I339,I251,I267,I366,);
DFFARX1 I_6 (I366,I251,I267,I384,);
DFFARX1 I_7 (I204,I251,I267,I402,);
nand I_8 (I411,I402,I196);
not I_9 (I429,I411);
DFFARX1 I_10 (I429,I251,I267,I456,);
not I_11 (I465,I456);
nor I_12 (I483,I303,I465);
DFFARX1 I_13 (I228,I251,I267,I510,);
nor I_14 (I519,I510,I366);
nor I_15 (I537,I510,I429);
nand I_16 (I555,I188,I116);
and I_17 (I573,I555,I156);
DFFARX1 I_18 (I573,I251,I267,I600,);
not I_19 (I609,I600);
nand I_20 (I627,I609,I510);
nand I_21 (I645,I609,I411);
nor I_22 (I663,I132,I116);
and I_23 (I681,I510,I663);
nor I_24 (I699,I609,I681);
DFFARX1 I_25 (I699,I251,I267,I726,);
nor I_26 (I735,I294,I663);
DFFARX1 I_27 (I735,I251,I267,I762,);
nor I_28 (I771,I600,I663);
not I_29 (I789,I771);
nand I_30 (I807,I789,I627);
not I_31 (I825,I258);
DFFARX1 I_32 (I726,I251,I825,I852,);
not I_33 (I861,I852);
nand I_34 (I879,I537,I483);
and I_35 (I897,I879,I384);
DFFARX1 I_36 (I897,I251,I825,I924,);
not I_37 (I933,I807);
DFFARX1 I_38 (I645,I251,I825,I960,);
not I_39 (I969,I960);
nor I_40 (I987,I969,I861);
and I_41 (I1005,I987,I807);
nor I_42 (I1023,I969,I933);
nor I_43 (I1041,I924,I1023);
DFFARX1 I_44 (I762,I251,I825,I1068,);
nor I_45 (I1077,I1068,I924);
not I_46 (I1095,I1077);
not I_47 (I1113,I1068);
nor I_48 (I1131,I1113,I1005);
DFFARX1 I_49 (I1131,I251,I825,I1158,);
nand I_50 (I1167,I762,I537);
and I_51 (I1185,I1167,I645);
DFFARX1 I_52 (I1185,I251,I825,I1212,);
nor I_53 (I1221,I1212,I1068);
DFFARX1 I_54 (I1221,I251,I825,I1248,);
nand I_55 (I1257,I1212,I1113);
nand I_56 (I1275,I1095,I1257);
not I_57 (I1293,I1212);
nor I_58 (I1311,I1293,I1005);
DFFARX1 I_59 (I1311,I251,I825,I1338,);
nor I_60 (I1347,I519,I537);
or I_61 (I1365,I1068,I1347);
nor I_62 (I1383,I1212,I1347);
or I_63 (I1401,I924,I1347);
DFFARX1 I_64 (I1347,I251,I825,I1428,);
not I_65 (I1437,I258);
DFFARX1 I_66 (I1365,I251,I1437,I1464,);
DFFARX1 I_67 (I1464,I251,I1437,I1482,);
not I_68 (I1491,I1482);
not I_69 (I1509,I1464);
DFFARX1 I_70 (I1275,I251,I1437,I1536,);
not I_71 (I1545,I1536);
and I_72 (I1563,I1509,I1041);
not I_73 (I1581,I1248);
nand I_74 (I1599,I1581,I1041);
not I_75 (I1617,I1383);
nor I_76 (I1635,I1617,I1428);
nand I_77 (I1653,I1635,I1338);
nor I_78 (I1671,I1653,I1599);
DFFARX1 I_79 (I1671,I251,I1437,I1698,);
not I_80 (I1707,I1653);
not I_81 (I1725,I1428);
nand I_82 (I1743,I1725,I1041);
nor I_83 (I1761,I1428,I1248);
nand I_84 (I1779,I1563,I1761);
nand I_85 (I1797,I1509,I1428);
nand I_86 (I1815,I1617,I1248);
DFFARX1 I_87 (I1815,I251,I1437,I1842,);
DFFARX1 I_88 (I1815,I251,I1437,I1860,);
not I_89 (I1869,I1248);
nor I_90 (I1887,I1869,I1401);
and I_91 (I1905,I1887,I1158);
or I_92 (I1923,I1905,I1383);
DFFARX1 I_93 (I1923,I251,I1437,I1950,);
nand I_94 (I1959,I1950,I1581);
nor I_95 (I1977,I1959,I1743);
nor I_96 (I1995,I1950,I1545);
DFFARX1 I_97 (I1950,I251,I1437,I2022,);
not I_98 (I2031,I2022);
nor I_99 (I2049,I2031,I1707);
not I_100 (I2067,I258);
DFFARX1 I_101 (I1698,I251,I2067,I2094,);
DFFARX1 I_102 (I1995,I251,I2067,I2112,);
not I_103 (I2121,I2112);
nor I_104 (I2139,I2094,I2121);
DFFARX1 I_105 (I2121,I251,I2067,I2166,);
nor I_106 (I2175,I1977,I1995);
and I_107 (I2193,I2175,I1797);
nor I_108 (I2211,I2193,I1977);
not I_109 (I2229,I1977);
and I_110 (I2247,I2229,I1698);
nand I_111 (I2265,I2247,I2049);
nor I_112 (I2283,I2229,I2265);
DFFARX1 I_113 (I2283,I251,I2067,I2310,);
not I_114 (I2319,I2265);
nand I_115 (I2337,I2121,I2319);
nand I_116 (I2355,I2193,I2319);
DFFARX1 I_117 (I2229,I251,I2067,I2382,);
not I_118 (I2391,I1779);
nor I_119 (I2409,I2391,I1698);
nor I_120 (I2427,I2409,I2211);
DFFARX1 I_121 (I2427,I251,I2067,I2454,);
not I_122 (I2463,I2409);
DFFARX1 I_123 (I2463,I251,I2067,I2490,);
not I_124 (I2499,I2490);
nor I_125 (I2517,I2499,I2409);
nor I_126 (I2535,I2391,I1842);
and I_127 (I2553,I2535,I1860);
or I_128 (I2571,I2553,I1491);
DFFARX1 I_129 (I2571,I251,I2067,I2598,);
not I_130 (I2607,I2598);
nand I_131 (I2625,I2607,I2319);
not I_132 (I2643,I2625);
nand I_133 (I2661,I2625,I2337);
nand I_134 (I2679,I2607,I2193);
not I_135 (I2697,I258);
DFFARX1 I_136 (I2382,I251,I2697,I2724,);
and I_137 (I2733,I2724,I2661);
DFFARX1 I_138 (I2733,I251,I2697,I2760,);
DFFARX1 I_139 (I2310,I251,I2697,I2778,);
not I_140 (I2787,I2643);
not I_141 (I2805,I2139);
nand I_142 (I2823,I2805,I2787);
nor I_143 (I2841,I2778,I2823);
DFFARX1 I_144 (I2823,I251,I2697,I2868,);
not I_145 (I2877,I2868);
not I_146 (I2895,I2355);
nand I_147 (I2913,I2805,I2895);
DFFARX1 I_148 (I2913,I251,I2697,I2940,);
not I_149 (I2949,I2940);
not I_150 (I2967,I2517);
nand I_151 (I2985,I2967,I2310);
and I_152 (I3003,I2787,I2985);
nor I_153 (I3021,I2913,I3003);
DFFARX1 I_154 (I3021,I251,I2697,I3048,);
DFFARX1 I_155 (I3003,I251,I2697,I3066,);
nor I_156 (I3075,I2517,I2454);
nor I_157 (I3093,I2913,I3075);
or I_158 (I3111,I2517,I2454);
nor I_159 (I3129,I2166,I2679);
DFFARX1 I_160 (I3129,I251,I2697,I3156,);
not I_161 (I3165,I3156);
nor I_162 (I3183,I3165,I2949);
nand I_163 (I3201,I3165,I2778);
not I_164 (I3219,I2166);
nand I_165 (I3237,I3219,I2895);
nand I_166 (I3255,I3165,I3237);
nand I_167 (I3273,I3255,I3201);
nand I_168 (I3291,I3237,I3111);
not I_169 (I3309,I258);
DFFARX1 I_170 (I3048,I251,I3309,I3336,);
DFFARX1 I_171 (I3336,I251,I3309,I3354,);
not I_172 (I3363,I3354);
not I_173 (I3381,I3336);
DFFARX1 I_174 (I3048,I251,I3309,I3408,);
not I_175 (I3417,I3408);
and I_176 (I3435,I3381,I2841);
not I_177 (I3453,I2760);
nand I_178 (I3471,I3453,I2841);
not I_179 (I3489,I3066);
nor I_180 (I3507,I3489,I3093);
nand I_181 (I3525,I3507,I3183);
nor I_182 (I3543,I3525,I3471);
DFFARX1 I_183 (I3543,I251,I3309,I3570,);
not I_184 (I3579,I3525);
not I_185 (I3597,I3093);
nand I_186 (I3615,I3597,I2841);
nor I_187 (I3633,I3093,I2760);
nand I_188 (I3651,I3435,I3633);
nand I_189 (I3669,I3381,I3093);
nand I_190 (I3687,I3489,I3273);
DFFARX1 I_191 (I3687,I251,I3309,I3714,);
DFFARX1 I_192 (I3687,I251,I3309,I3732,);
not I_193 (I3741,I3273);
nor I_194 (I3759,I3741,I3291);
and I_195 (I3777,I3759,I2877);
or I_196 (I3795,I3777,I2841);
DFFARX1 I_197 (I3795,I251,I3309,I3822,);
nand I_198 (I3831,I3822,I3453);
nor I_199 (I3849,I3831,I3615);
nor I_200 (I3867,I3822,I3417);
DFFARX1 I_201 (I3822,I251,I3309,I3894,);
not I_202 (I3903,I3894);
nor I_203 (I3921,I3903,I3579);
not I_204 (I3939,I258);
DFFARX1 I_205 (I3570,I251,I3939,I3966,);
nand I_206 (I3975,I3570,I3669);
and I_207 (I3993,I3975,I3363);
DFFARX1 I_208 (I3993,I251,I3939,I4020,);
nor I_209 (I4029,I4020,I3966);
not I_210 (I4047,I4020);
DFFARX1 I_211 (I3651,I251,I3939,I4074,);
nand I_212 (I4083,I4074,I3849);
not I_213 (I4101,I4083);
DFFARX1 I_214 (I4101,I251,I3939,I4128,);
not I_215 (I4137,I4128);
nor I_216 (I4155,I3966,I4083);
nor I_217 (I4173,I4020,I4155);
DFFARX1 I_218 (I3921,I251,I3939,I4200,);
DFFARX1 I_219 (I4200,I251,I3939,I4218,);
not I_220 (I4227,I4218);
not I_221 (I4245,I4200);
nand I_222 (I4263,I4245,I4047);
nand I_223 (I4281,I3867,I3867);
and I_224 (I4299,I4281,I3714);
DFFARX1 I_225 (I4299,I251,I3939,I4326,);
nor I_226 (I4335,I4326,I3966);
DFFARX1 I_227 (I4335,I251,I3939,I4362,);
DFFARX1 I_228 (I4326,I251,I3939,I4380,);
nor I_229 (I4389,I3732,I3867);
not I_230 (I4407,I4389);
nor I_231 (I4425,I4227,I4407);
nand I_232 (I4443,I4245,I4407);
nor I_233 (I4461,I3966,I4389);
DFFARX1 I_234 (I4389,I251,I3939,I4488,);
not I_235 (I4497,I258);
DFFARX1 I_236 (I4425,I251,I4497,I4524,);
DFFARX1 I_237 (I4461,I251,I4497,I4542,);
not I_238 (I4551,I4542);
nor I_239 (I4569,I4524,I4551);
DFFARX1 I_240 (I4551,I251,I4497,I4596,);
nor I_241 (I4605,I4029,I4488);
and I_242 (I4623,I4605,I4380);
nor I_243 (I4641,I4623,I4029);
not I_244 (I4659,I4029);
and I_245 (I4677,I4659,I4362);
nand I_246 (I4695,I4677,I4263);
nor I_247 (I4713,I4659,I4695);
DFFARX1 I_248 (I4713,I251,I4497,I4740,);
not I_249 (I4749,I4695);
nand I_250 (I4767,I4551,I4749);
nand I_251 (I4785,I4623,I4749);
DFFARX1 I_252 (I4659,I251,I4497,I4812,);
not I_253 (I4821,I4137);
nor I_254 (I4839,I4821,I4362);
nor I_255 (I4857,I4839,I4641);
DFFARX1 I_256 (I4857,I251,I4497,I4884,);
not I_257 (I4893,I4839);
DFFARX1 I_258 (I4893,I251,I4497,I4920,);
not I_259 (I4929,I4920);
nor I_260 (I4947,I4929,I4839);
nor I_261 (I4965,I4821,I4173);
and I_262 (I4983,I4965,I4443);
or I_263 (I5001,I4983,I4362);
DFFARX1 I_264 (I5001,I251,I4497,I5028,);
not I_265 (I5037,I5028);
nand I_266 (I5055,I5037,I4749);
not I_267 (I5073,I5055);
nand I_268 (I5091,I5055,I4767);
nand I_269 (I5109,I5037,I4623);
not I_270 (I5127,I258);
DFFARX1 I_271 (I4785,I251,I5127,I5154,);
not I_272 (I5163,I5154);
nand I_273 (I5181,I5109,I4812);
and I_274 (I5199,I5181,I4569);
DFFARX1 I_275 (I5199,I251,I5127,I5226,);
DFFARX1 I_276 (I4884,I251,I5127,I5244,);
and I_277 (I5253,I5244,I4947);
nor I_278 (I5271,I5226,I5253);
DFFARX1 I_279 (I5271,I251,I5127,I5298,);
nand I_280 (I5307,I5244,I4947);
nand I_281 (I5325,I5163,I5307);
not I_282 (I5343,I5325);
DFFARX1 I_283 (I5091,I251,I5127,I5370,);
DFFARX1 I_284 (I5370,I251,I5127,I5388,);
nand I_285 (I5397,I4596,I5073);
and I_286 (I5415,I5397,I4740);
DFFARX1 I_287 (I5415,I251,I5127,I5442,);
DFFARX1 I_288 (I5442,I251,I5127,I5460,);
not I_289 (I5469,I5460);
not I_290 (I5487,I5442);
nand I_291 (I5505,I5487,I5307);
nor I_292 (I5523,I4740,I5073);
not I_293 (I5541,I5523);
nor I_294 (I5559,I5487,I5541);
nor I_295 (I5577,I5163,I5559);
DFFARX1 I_296 (I5577,I251,I5127,I5604,);
nor I_297 (I5613,I5226,I5541);
nor I_298 (I5631,I5442,I5613);
nor I_299 (I5649,I5370,I5523);
nor I_300 (I5667,I5226,I5523);
not I_301 (I5685,I258);
DFFARX1 I_302 (I5388,I251,I5685,I5712,);
DFFARX1 I_303 (I5505,I251,I5685,I5730,);
not I_304 (I5739,I5730);
nor I_305 (I5757,I5712,I5739);
DFFARX1 I_306 (I5739,I251,I5685,I5784,);
nor I_307 (I5793,I5298,I5469);
and I_308 (I5811,I5793,I5667);
nor I_309 (I5829,I5811,I5298);
not I_310 (I5847,I5298);
and I_311 (I5865,I5847,I5631);
nand I_312 (I5883,I5865,I5604);
nor I_313 (I5901,I5847,I5883);
DFFARX1 I_314 (I5901,I251,I5685,I5928,);
not I_315 (I5937,I5883);
nand I_316 (I5955,I5739,I5937);
nand I_317 (I5973,I5811,I5937);
DFFARX1 I_318 (I5847,I251,I5685,I6000,);
not I_319 (I6009,I5298);
nor I_320 (I6027,I6009,I5631);
nor I_321 (I6045,I6027,I5829);
DFFARX1 I_322 (I6045,I251,I5685,I6072,);
not I_323 (I6081,I6027);
DFFARX1 I_324 (I6081,I251,I5685,I6108,);
not I_325 (I6117,I6108);
nor I_326 (I6135,I6117,I6027);
nor I_327 (I6153,I6009,I5667);
and I_328 (I6171,I6153,I5343);
or I_329 (I6189,I6171,I5649);
DFFARX1 I_330 (I6189,I251,I5685,I6216,);
not I_331 (I6225,I6216);
nand I_332 (I6243,I6225,I5937);
not I_333 (I6261,I6243);
nand I_334 (I6279,I6243,I5955);
nand I_335 (I6297,I6225,I5811);
not I_336 (I6315,I258);
DFFARX1 I_337 (I6261,I251,I6315,I6342,);
DFFARX1 I_338 (I6342,I251,I6315,I6360,);
not I_339 (I6369,I6360);
not I_340 (I6387,I6342);
DFFARX1 I_341 (I6279,I251,I6315,I6414,);
nand I_342 (I6423,I6414,I5928);
not I_343 (I6441,I5928);
not I_344 (I6459,I6000);
nand I_345 (I6477,I5973,I6135);
and I_346 (I6495,I5973,I6135);
not I_347 (I6513,I6297);
nand I_348 (I6531,I6513,I6459);
nor I_349 (I6549,I6531,I6423);
nor I_350 (I6567,I6441,I6531);
nand I_351 (I6585,I6495,I6567);
not I_352 (I6603,I6072);
nor I_353 (I6621,I6603,I5973);
nor I_354 (I6639,I6621,I6297);
nor I_355 (I6657,I6387,I6639);
DFFARX1 I_356 (I6657,I251,I6315,I6684,);
not I_357 (I6693,I6621);
DFFARX1 I_358 (I6693,I251,I6315,I6720,);
and I_359 (I6729,I6414,I6621);
nor I_360 (I6747,I6603,I5784);
and I_361 (I6765,I6747,I5928);
or I_362 (I6783,I6765,I5757);
DFFARX1 I_363 (I6783,I251,I6315,I6810,);
nor I_364 (I6819,I6810,I6513);
DFFARX1 I_365 (I6819,I251,I6315,I6846,);
nand I_366 (I6855,I6810,I6414);
nand I_367 (I6873,I6513,I6855);
nor I_368 (I6891,I6873,I6477);
not I_369 (I6909,I258);
DFFARX1 I_370 (I6846,I251,I6909,I6936,);
DFFARX1 I_371 (I6549,I251,I6909,I6954,);
not I_372 (I6963,I6954);
not I_373 (I6981,I6846);
nor I_374 (I6999,I6981,I6729);
not I_375 (I7017,I6369);
nor I_376 (I7035,I6999,I6891);
nor I_377 (I7053,I6954,I7035);
DFFARX1 I_378 (I7053,I251,I6909,I7080,);
nor I_379 (I7089,I6891,I6729);
nand I_380 (I7107,I7089,I6846);
DFFARX1 I_381 (I7107,I251,I6909,I7134,);
nor I_382 (I7143,I7017,I6891);
nand I_383 (I7161,I7143,I6684);
nor I_384 (I7179,I6936,I7161);
DFFARX1 I_385 (I7179,I251,I6909,I7206,);
not I_386 (I7215,I7161);
nand I_387 (I7233,I6954,I7215);
DFFARX1 I_388 (I7161,I251,I6909,I7260,);
not I_389 (I7269,I7260);
not I_390 (I7287,I6891);
not I_391 (I7305,I6585);
nor I_392 (I7323,I7305,I6369);
nor I_393 (I7341,I7269,I7323);
nor I_394 (I7359,I7305,I6720);
and I_395 (I7377,I7359,I6585);
or I_396 (I7395,I7377,I6549);
DFFARX1 I_397 (I7395,I251,I6909,I7422,);
nor I_398 (I7431,I7422,I6936);
not I_399 (I7449,I7422);
and I_400 (I7467,I7449,I6936);
nor I_401 (I7485,I6963,I7467);
nand I_402 (I7503,I7449,I7017);
nor I_403 (I7521,I7305,I7503);
nand I_404 (I7539,I7449,I7215);
nand I_405 (I7557,I7017,I6585);
nor I_406 (I7575,I7287,I7557);
not I_407 (I7593,I258);
DFFARX1 I_408 (I7521,I251,I7593,I7620,);
nand I_409 (I7629,I7206,I7575);
and I_410 (I7647,I7629,I7485);
DFFARX1 I_411 (I7647,I251,I7593,I7674,);
nor I_412 (I7683,I7674,I7620);
not I_413 (I7701,I7674);
DFFARX1 I_414 (I7134,I251,I7593,I7728,);
nand I_415 (I7737,I7728,I7539);
not I_416 (I7755,I7737);
DFFARX1 I_417 (I7755,I251,I7593,I7782,);
not I_418 (I7791,I7782);
nor I_419 (I7809,I7620,I7737);
nor I_420 (I7827,I7674,I7809);
DFFARX1 I_421 (I7233,I251,I7593,I7854,);
DFFARX1 I_422 (I7854,I251,I7593,I7872,);
not I_423 (I7881,I7872);
not I_424 (I7899,I7854);
nand I_425 (I7917,I7899,I7701);
nand I_426 (I7935,I7206,I7341);
and I_427 (I7953,I7935,I7431);
DFFARX1 I_428 (I7953,I251,I7593,I7980,);
nor I_429 (I7989,I7980,I7620);
DFFARX1 I_430 (I7989,I251,I7593,I8016,);
DFFARX1 I_431 (I7980,I251,I7593,I8034,);
nor I_432 (I8043,I7080,I7341);
not I_433 (I8061,I8043);
nor I_434 (I8079,I7881,I8061);
nand I_435 (I8097,I7899,I8061);
nor I_436 (I8115,I7620,I8043);
DFFARX1 I_437 (I8043,I251,I7593,I8142,);
not I_438 (I8151,I258);
DFFARX1 I_439 (I8079,I251,I8151,I8178,);
DFFARX1 I_440 (I8115,I251,I8151,I8196,);
not I_441 (I8205,I8196);
nor I_442 (I8223,I8178,I8205);
DFFARX1 I_443 (I8205,I251,I8151,I8250,);
nor I_444 (I8259,I7683,I8142);
and I_445 (I8277,I8259,I8034);
nor I_446 (I8295,I8277,I7683);
not I_447 (I8313,I7683);
and I_448 (I8331,I8313,I8016);
nand I_449 (I8349,I8331,I7917);
nor I_450 (I8367,I8313,I8349);
DFFARX1 I_451 (I8367,I251,I8151,I8394,);
not I_452 (I8403,I8349);
nand I_453 (I8421,I8205,I8403);
nand I_454 (I8439,I8277,I8403);
DFFARX1 I_455 (I8313,I251,I8151,I8466,);
not I_456 (I8475,I7791);
nor I_457 (I8493,I8475,I8016);
nor I_458 (I8511,I8493,I8295);
DFFARX1 I_459 (I8511,I251,I8151,I8538,);
not I_460 (I8547,I8493);
DFFARX1 I_461 (I8547,I251,I8151,I8574,);
not I_462 (I8583,I8574);
nor I_463 (I8601,I8583,I8493);
nor I_464 (I8619,I8475,I7827);
and I_465 (I8637,I8619,I8097);
or I_466 (I8655,I8637,I8016);
DFFARX1 I_467 (I8655,I251,I8151,I8682,);
not I_468 (I8691,I8682);
nand I_469 (I8709,I8691,I8403);
not I_470 (I8727,I8709);
nand I_471 (I8745,I8709,I8421);
nand I_472 (I8763,I8691,I8277);
not I_473 (I8781,I258);
DFFARX1 I_474 (I8466,I251,I8781,I8808,);
not I_475 (I8817,I8808);
nand I_476 (I8835,I8439,I8394);
and I_477 (I8853,I8835,I8727);
DFFARX1 I_478 (I8853,I251,I8781,I8880,);
not I_479 (I8889,I8394);
DFFARX1 I_480 (I8250,I251,I8781,I8916,);
not I_481 (I8925,I8916);
nor I_482 (I8943,I8925,I8817);
and I_483 (I8961,I8943,I8394);
nor I_484 (I8979,I8925,I8889);
nor I_485 (I8997,I8880,I8979);
DFFARX1 I_486 (I8763,I251,I8781,I9024,);
nor I_487 (I9033,I9024,I8880);
not I_488 (I9051,I9033);
not I_489 (I9069,I9024);
nor I_490 (I9087,I9069,I8961);
DFFARX1 I_491 (I9087,I251,I8781,I9114,);
nand I_492 (I9123,I8223,I8745);
and I_493 (I9141,I9123,I8538);
DFFARX1 I_494 (I9141,I251,I8781,I9168,);
nor I_495 (I9177,I9168,I9024);
DFFARX1 I_496 (I9177,I251,I8781,I9204,);
nand I_497 (I9213,I9168,I9069);
nand I_498 (I9231,I9051,I9213);
not I_499 (I9249,I9168);
nor I_500 (I9267,I9249,I8961);
DFFARX1 I_501 (I9267,I251,I8781,I9294,);
nor I_502 (I9303,I8601,I8745);
or I_503 (I9321,I9024,I9303);
nor I_504 (I9339,I9168,I9303);
or I_505 (I9357,I8880,I9303);
DFFARX1 I_506 (I9303,I251,I8781,I9384,);
not I_507 (I9393,I258);
DFFARX1 I_508 (I9321,I251,I9393,I9420,);
nand I_509 (I9429,I9339,I9114);
and I_510 (I9447,I9429,I9384);
DFFARX1 I_511 (I9447,I251,I9393,I9474,);
nor I_512 (I9483,I9474,I9420);
not I_513 (I9501,I9474);
DFFARX1 I_514 (I9231,I251,I9393,I9528,);
nand I_515 (I9537,I9528,I9339);
not I_516 (I9555,I9537);
DFFARX1 I_517 (I9555,I251,I9393,I9582,);
not I_518 (I9591,I9582);
nor I_519 (I9609,I9420,I9537);
nor I_520 (I9627,I9474,I9609);
DFFARX1 I_521 (I9357,I251,I9393,I9654,);
DFFARX1 I_522 (I9654,I251,I9393,I9672,);
not I_523 (I9681,I9672);
not I_524 (I9699,I9654);
nand I_525 (I9717,I9699,I9501);
nand I_526 (I9735,I9204,I8997);
and I_527 (I9753,I9735,I9204);
DFFARX1 I_528 (I9753,I251,I9393,I9780,);
nor I_529 (I9789,I9780,I9420);
DFFARX1 I_530 (I9789,I251,I9393,I9816,);
DFFARX1 I_531 (I9780,I251,I9393,I9834,);
nor I_532 (I9843,I9294,I8997);
not I_533 (I9861,I9843);
nor I_534 (I9879,I9681,I9861);
nand I_535 (I9897,I9699,I9861);
nor I_536 (I9915,I9420,I9843);
DFFARX1 I_537 (I9843,I251,I9393,I9942,);
not I_538 (I9951,I258);
DFFARX1 I_539 (I9942,I251,I9951,I9978,);
not I_540 (I9987,I9978);
nand I_541 (I10005,I9591,I9483);
and I_542 (I10023,I10005,I9816);
DFFARX1 I_543 (I10023,I251,I9951,I10050,);
not I_544 (I10059,I9897);
DFFARX1 I_545 (I9816,I251,I9951,I10086,);
not I_546 (I10095,I10086);
nor I_547 (I10113,I10095,I9987);
and I_548 (I10131,I10113,I9897);
nor I_549 (I10149,I10095,I10059);
nor I_550 (I10167,I10050,I10149);
DFFARX1 I_551 (I9627,I251,I9951,I10194,);
nor I_552 (I10203,I10194,I10050);
not I_553 (I10221,I10203);
not I_554 (I10239,I10194);
nor I_555 (I10257,I10239,I10131);
DFFARX1 I_556 (I10257,I251,I9951,I10284,);
nand I_557 (I10293,I9717,I9879);
and I_558 (I10311,I10293,I9834);
DFFARX1 I_559 (I10311,I251,I9951,I10338,);
nor I_560 (I10347,I10338,I10194);
DFFARX1 I_561 (I10347,I251,I9951,I10374,);
nand I_562 (I10383,I10338,I10239);
nand I_563 (I10401,I10221,I10383);
not I_564 (I10419,I10338);
nor I_565 (I10437,I10419,I10131);
DFFARX1 I_566 (I10437,I251,I9951,I10464,);
nor I_567 (I10473,I9915,I9879);
or I_568 (I10491,I10194,I10473);
nor I_569 (I10509,I10338,I10473);
or I_570 (I10527,I10050,I10473);
DFFARX1 I_571 (I10473,I251,I9951,I10554,);
not I_572 (I10563,I258);
DFFARX1 I_573 (I10491,I251,I10563,I10590,);
not I_574 (I10599,I10590);
nand I_575 (I10617,I10509,I10464);
and I_576 (I10635,I10617,I10374);
DFFARX1 I_577 (I10635,I251,I10563,I10662,);
DFFARX1 I_578 (I10509,I251,I10563,I10680,);
and I_579 (I10689,I10680,I10527);
nor I_580 (I10707,I10662,I10689);
DFFARX1 I_581 (I10707,I251,I10563,I10734,);
nand I_582 (I10743,I10680,I10527);
nand I_583 (I10761,I10599,I10743);
not I_584 (I10779,I10761);
DFFARX1 I_585 (I10374,I251,I10563,I10806,);
DFFARX1 I_586 (I10806,I251,I10563,I10824,);
nand I_587 (I10833,I10284,I10401);
and I_588 (I10851,I10833,I10554);
DFFARX1 I_589 (I10851,I251,I10563,I10878,);
DFFARX1 I_590 (I10878,I251,I10563,I10896,);
not I_591 (I10905,I10896);
not I_592 (I10923,I10878);
nand I_593 (I10941,I10923,I10743);
nor I_594 (I10959,I10167,I10401);
not I_595 (I10977,I10959);
nor I_596 (I10995,I10923,I10977);
nor I_597 (I11013,I10599,I10995);
DFFARX1 I_598 (I11013,I251,I10563,I11040,);
nor I_599 (I11049,I10662,I10977);
nor I_600 (I11067,I10878,I11049);
nor I_601 (I11085,I10806,I10959);
nor I_602 (I11103,I10662,I10959);
not I_603 (I11121,I258);
DFFARX1 I_604 (I10905,I251,I11121,I11148,);
not I_605 (I11157,I11148);
DFFARX1 I_606 (I11103,I251,I11121,I11184,);
not I_607 (I11193,I10734);
nand I_608 (I11211,I11193,I11085);
not I_609 (I11229,I11211);
nor I_610 (I11247,I11229,I11103);
nor I_611 (I11265,I11157,I11247);
DFFARX1 I_612 (I11265,I251,I11121,I11292,);
not I_613 (I11301,I11103);
nand I_614 (I11319,I11301,I11229);
and I_615 (I11337,I11301,I11067);
nand I_616 (I11355,I11337,I10824);
nor I_617 (I11373,I11355,I11301);
and I_618 (I11391,I11184,I11355);
not I_619 (I11409,I11355);
nand I_620 (I11427,I11184,I11409);
nor I_621 (I11445,I11148,I11355);
not I_622 (I11463,I10779);
nor I_623 (I11481,I11463,I11067);
nand I_624 (I11499,I11481,I11301);
nor I_625 (I11517,I11211,I11499);
nor I_626 (I11535,I11463,I10734);
and I_627 (I11553,I11535,I10941);
or I_628 (I11571,I11553,I11040);
DFFARX1 I_629 (I11571,I251,I11121,I11598,);
nor I_630 (I11607,I11598,I11319);
DFFARX1 I_631 (I11607,I251,I11121,I11634,);
DFFARX1 I_632 (I11598,I251,I11121,I11652,);
not I_633 (I11661,I11598);
nor I_634 (I11679,I11661,I11184);
nor I_635 (I11697,I11481,I11679);
DFFARX1 I_636 (I11697,I251,I11121,I11724,);
not I_637 (I11733,I258);
DFFARX1 I_638 (I244,I251,I11733,I11760,);
nand I_639 (I11769,I11760,I76);
not I_640 (I11787,I11769);
DFFARX1 I_641 (I236,I251,I11733,I11814,);
not I_642 (I11823,I11814);
not I_643 (I11841,I220);
or I_644 (I11859,I180,I220);
nor I_645 (I11877,I180,I220);
or I_646 (I11895,I172,I180);
DFFARX1 I_647 (I11895,I251,I11733,I11922,);
not I_648 (I11931,I212);
nand I_649 (I11949,I11931,I108);
nand I_650 (I11967,I11841,I11949);
and I_651 (I11985,I11823,I11967);
nor I_652 (I12003,I212,I92);
and I_653 (I12021,I11823,I12003);
nor I_654 (I12039,I11787,I12021);
DFFARX1 I_655 (I12003,I251,I11733,I12066,);
not I_656 (I12075,I12066);
nor I_657 (I12093,I11823,I12075);
or I_658 (I12111,I11895,I84);
nor I_659 (I12129,I84,I172);
nand I_660 (I12147,I11967,I12129);
nand I_661 (I12165,I12111,I12147);
DFFARX1 I_662 (I12165,I251,I11733,I12192,);
nor I_663 (I12201,I12129,I11859);
DFFARX1 I_664 (I12201,I251,I11733,I12228,);
nor I_665 (I12237,I84,I124);
DFFARX1 I_666 (I12237,I251,I11733,I12264,);
DFFARX1 I_667 (I12264,I251,I11733,I12282,);
not I_668 (I12291,I12264);
nand I_669 (I12309,I12291,I11769);
nand I_670 (I12327,I12291,I11877);
not I_671 (I12345,I258);
DFFARX1 I_672 (I11922,I251,I12345,I12372,);
and I_673 (I12381,I12372,I12327);
DFFARX1 I_674 (I12381,I251,I12345,I12408,);
DFFARX1 I_675 (I12282,I251,I12345,I12426,);
not I_676 (I12435,I12228);
not I_677 (I12453,I12309);
nand I_678 (I12471,I12453,I12435);
nor I_679 (I12489,I12426,I12471);
DFFARX1 I_680 (I12471,I251,I12345,I12516,);
not I_681 (I12525,I12516);
not I_682 (I12543,I11985);
nand I_683 (I12561,I12453,I12543);
DFFARX1 I_684 (I12561,I251,I12345,I12588,);
not I_685 (I12597,I12588);
not I_686 (I12615,I12228);
nand I_687 (I12633,I12615,I11985);
and I_688 (I12651,I12435,I12633);
nor I_689 (I12669,I12561,I12651);
DFFARX1 I_690 (I12669,I251,I12345,I12696,);
DFFARX1 I_691 (I12651,I251,I12345,I12714,);
nor I_692 (I12723,I12228,I12192);
nor I_693 (I12741,I12561,I12723);
or I_694 (I12759,I12228,I12192);
nor I_695 (I12777,I12039,I12093);
DFFARX1 I_696 (I12777,I251,I12345,I12804,);
not I_697 (I12813,I12804);
nor I_698 (I12831,I12813,I12597);
nand I_699 (I12849,I12813,I12426);
not I_700 (I12867,I12039);
nand I_701 (I12885,I12867,I12543);
nand I_702 (I12903,I12813,I12885);
nand I_703 (I12921,I12903,I12849);
nand I_704 (I12939,I12885,I12759);
not I_705 (I12957,I258);
DFFARX1 I_706 (I12831,I251,I12957,I12984,);
not I_707 (I12993,I12984);
nand I_708 (I13011,I12696,I12741);
and I_709 (I13029,I13011,I12408);
DFFARX1 I_710 (I13029,I251,I12957,I13056,);
not I_711 (I13065,I12921);
DFFARX1 I_712 (I12939,I251,I12957,I13092,);
not I_713 (I13101,I13092);
nor I_714 (I13119,I13101,I12993);
and I_715 (I13137,I13119,I12921);
nor I_716 (I13155,I13101,I13065);
nor I_717 (I13173,I13056,I13155);
DFFARX1 I_718 (I12525,I251,I12957,I13200,);
nor I_719 (I13209,I13200,I13056);
not I_720 (I13227,I13209);
not I_721 (I13245,I13200);
nor I_722 (I13263,I13245,I13137);
DFFARX1 I_723 (I13263,I251,I12957,I13290,);
nand I_724 (I13299,I12489,I12489);
and I_725 (I13317,I13299,I12696);
DFFARX1 I_726 (I13317,I251,I12957,I13344,);
nor I_727 (I13353,I13344,I13200);
DFFARX1 I_728 (I13353,I251,I12957,I13380,);
nand I_729 (I13389,I13344,I13245);
nand I_730 (I13407,I13227,I13389);
not I_731 (I13425,I13344);
nor I_732 (I13443,I13425,I13137);
DFFARX1 I_733 (I13443,I251,I12957,I13470,);
nor I_734 (I13479,I12714,I12489);
or I_735 (I13497,I13200,I13479);
nor I_736 (I13515,I13344,I13479);
or I_737 (I13533,I13056,I13479);
DFFARX1 I_738 (I13479,I251,I12957,I13560,);
not I_739 (I13569,I258);
DFFARX1 I_740 (I13497,I251,I13569,I13596,);
nand I_741 (I13605,I13515,I13290);
and I_742 (I13623,I13605,I13560);
DFFARX1 I_743 (I13623,I251,I13569,I13650,);
nor I_744 (I13659,I13650,I13596);
not I_745 (I13677,I13650);
DFFARX1 I_746 (I13407,I251,I13569,I13704,);
nand I_747 (I13713,I13704,I13515);
not I_748 (I13731,I13713);
DFFARX1 I_749 (I13731,I251,I13569,I13758,);
not I_750 (I13767,I13758);
nor I_751 (I13785,I13596,I13713);
nor I_752 (I13803,I13650,I13785);
DFFARX1 I_753 (I13533,I251,I13569,I13830,);
DFFARX1 I_754 (I13830,I251,I13569,I13848,);
not I_755 (I13857,I13848);
not I_756 (I13875,I13830);
nand I_757 (I13893,I13875,I13677);
nand I_758 (I13911,I13380,I13173);
and I_759 (I13929,I13911,I13380);
DFFARX1 I_760 (I13929,I251,I13569,I13956,);
nor I_761 (I13965,I13956,I13596);
DFFARX1 I_762 (I13965,I251,I13569,I13992,);
DFFARX1 I_763 (I13956,I251,I13569,I14010,);
nor I_764 (I14019,I13470,I13173);
not I_765 (I14037,I14019);
nor I_766 (I14055,I13857,I14037);
nand I_767 (I14073,I13875,I14037);
nor I_768 (I14091,I13596,I14019);
DFFARX1 I_769 (I14019,I251,I13569,I14118,);
not I_770 (I14127,I258);
DFFARX1 I_771 (I14055,I251,I14127,I14154,);
DFFARX1 I_772 (I14091,I251,I14127,I14172,);
not I_773 (I14181,I14172);
nor I_774 (I14199,I14154,I14181);
DFFARX1 I_775 (I14181,I251,I14127,I14226,);
nor I_776 (I14235,I13659,I14118);
and I_777 (I14253,I14235,I14010);
nor I_778 (I14271,I14253,I13659);
not I_779 (I14289,I13659);
and I_780 (I14307,I14289,I13992);
nand I_781 (I14325,I14307,I13893);
nor I_782 (I14343,I14289,I14325);
DFFARX1 I_783 (I14343,I251,I14127,I14370,);
not I_784 (I14379,I14325);
nand I_785 (I14397,I14181,I14379);
nand I_786 (I14415,I14253,I14379);
DFFARX1 I_787 (I14289,I251,I14127,I14442,);
not I_788 (I14451,I13767);
nor I_789 (I14469,I14451,I13992);
nor I_790 (I14487,I14469,I14271);
DFFARX1 I_791 (I14487,I251,I14127,I14514,);
not I_792 (I14523,I14469);
DFFARX1 I_793 (I14523,I251,I14127,I14550,);
not I_794 (I14559,I14550);
nor I_795 (I14577,I14559,I14469);
nor I_796 (I14595,I14451,I13803);
and I_797 (I14613,I14595,I14073);
or I_798 (I14631,I14613,I13992);
DFFARX1 I_799 (I14631,I251,I14127,I14658,);
not I_800 (I14667,I14658);
nand I_801 (I14685,I14667,I14379);
not I_802 (I14703,I14685);
nand I_803 (I14721,I14685,I14397);
nand I_804 (I14739,I14667,I14253);
not I_805 (I14757,I258);
DFFARX1 I_806 (I14442,I251,I14757,I14784,);
DFFARX1 I_807 (I14784,I251,I14757,I14802,);
not I_808 (I14811,I14802);
not I_809 (I14829,I14784);
nand I_810 (I14847,I14199,I14514);
and I_811 (I14865,I14847,I14577);
DFFARX1 I_812 (I14865,I251,I14757,I14892,);
not I_813 (I14901,I14892);
DFFARX1 I_814 (I14370,I251,I14757,I14928,);
and I_815 (I14937,I14928,I14415);
nand I_816 (I14955,I14928,I14415);
nand I_817 (I14973,I14901,I14955);
DFFARX1 I_818 (I14703,I251,I14757,I15000,);
nor I_819 (I15009,I15000,I14937);
DFFARX1 I_820 (I15009,I251,I14757,I15036,);
nor I_821 (I15045,I15000,I14892);
nand I_822 (I15063,I14226,I14739);
and I_823 (I15081,I15063,I14721);
DFFARX1 I_824 (I15081,I251,I14757,I15108,);
nor I_825 (I15117,I15108,I15000);
not I_826 (I15135,I15108);
nor I_827 (I15153,I15135,I14901);
nor I_828 (I15171,I14829,I15153);
DFFARX1 I_829 (I15171,I251,I14757,I15198,);
nor I_830 (I15207,I15135,I15000);
nor I_831 (I15225,I14370,I14739);
nor I_832 (I15243,I15225,I15207);
not I_833 (I15261,I15225);
nand I_834 (I15279,I14955,I15261);
DFFARX1 I_835 (I15225,I251,I14757,I15306,);
DFFARX1 I_836 (I15225,I251,I14757,I15324,);
not I_837 (I15333,I258);
DFFARX1 I_838 (I15036,I251,I15333,I15360,);
DFFARX1 I_839 (I14973,I251,I15333,I15378,);
not I_840 (I15387,I15378);
nor I_841 (I15405,I15360,I15387);
DFFARX1 I_842 (I15387,I251,I15333,I15432,);
nor I_843 (I15441,I15045,I15036);
and I_844 (I15459,I15441,I14811);
nor I_845 (I15477,I15459,I15045);
not I_846 (I15495,I15045);
and I_847 (I15513,I15495,I15117);
nand I_848 (I15531,I15513,I15306);
nor I_849 (I15549,I15495,I15531);
DFFARX1 I_850 (I15549,I251,I15333,I15576,);
not I_851 (I15585,I15531);
nand I_852 (I15603,I15387,I15585);
nand I_853 (I15621,I15459,I15585);
DFFARX1 I_854 (I15495,I251,I15333,I15648,);
not I_855 (I15657,I15279);
nor I_856 (I15675,I15657,I15117);
nor I_857 (I15693,I15675,I15477);
DFFARX1 I_858 (I15693,I251,I15333,I15720,);
not I_859 (I15729,I15675);
DFFARX1 I_860 (I15729,I251,I15333,I15756,);
not I_861 (I15765,I15756);
nor I_862 (I15783,I15765,I15675);
nor I_863 (I15801,I15657,I15243);
and I_864 (I15819,I15801,I15324);
or I_865 (I15837,I15819,I15198);
DFFARX1 I_866 (I15837,I251,I15333,I15864,);
not I_867 (I15873,I15864);
nand I_868 (I15891,I15873,I15585);
not I_869 (I15909,I15891);
nand I_870 (I15927,I15891,I15603);
nand I_871 (I15945,I15873,I15459);
not I_872 (I15963,I258);
DFFARX1 I_873 (I15648,I251,I15963,I15990,);
not I_874 (I15999,I15990);
nand I_875 (I16017,I15621,I15576);
and I_876 (I16035,I16017,I15909);
DFFARX1 I_877 (I16035,I251,I15963,I16062,);
not I_878 (I16071,I15576);
DFFARX1 I_879 (I15432,I251,I15963,I16098,);
not I_880 (I16107,I16098);
nor I_881 (I16125,I16107,I15999);
and I_882 (I16143,I16125,I15576);
nor I_883 (I16161,I16107,I16071);
nor I_884 (I16179,I16062,I16161);
DFFARX1 I_885 (I15945,I251,I15963,I16206,);
nor I_886 (I16215,I16206,I16062);
not I_887 (I16233,I16215);
not I_888 (I16251,I16206);
nor I_889 (I16269,I16251,I16143);
DFFARX1 I_890 (I16269,I251,I15963,I16296,);
nand I_891 (I16305,I15405,I15927);
and I_892 (I16323,I16305,I15720);
DFFARX1 I_893 (I16323,I251,I15963,I16350,);
nor I_894 (I16359,I16350,I16206);
DFFARX1 I_895 (I16359,I251,I15963,I16386,);
nand I_896 (I16395,I16350,I16251);
nand I_897 (I16413,I16233,I16395);
not I_898 (I16431,I16350);
nor I_899 (I16449,I16431,I16143);
DFFARX1 I_900 (I16449,I251,I15963,I16476,);
nor I_901 (I16485,I15783,I15927);
or I_902 (I16503,I16206,I16485);
nor I_903 (I16521,I16350,I16485);
or I_904 (I16539,I16062,I16485);
DFFARX1 I_905 (I16485,I251,I15963,I16566,);
not I_906 (I16575,I258);
DFFARX1 I_907 (I16413,I251,I16575,I16602,);
DFFARX1 I_908 (I16602,I251,I16575,I16620,);
not I_909 (I16629,I16620);
DFFARX1 I_910 (I16521,I251,I16575,I16656,);
not I_911 (I16665,I16386);
nor I_912 (I16683,I16602,I16665);
not I_913 (I16701,I16503);
not I_914 (I16719,I16179);
nand I_915 (I16737,I16719,I16503);
nor I_916 (I16755,I16665,I16737);
nor I_917 (I16773,I16656,I16755);
DFFARX1 I_918 (I16719,I251,I16575,I16800,);
nor I_919 (I16809,I16179,I16566);
nand I_920 (I16827,I16809,I16296);
nor I_921 (I16845,I16827,I16701);
nand I_922 (I16863,I16845,I16386);
DFFARX1 I_923 (I16827,I251,I16575,I16890,);
nand I_924 (I16899,I16701,I16179);
nor I_925 (I16917,I16701,I16179);
nand I_926 (I16935,I16683,I16917);
not I_927 (I16953,I16539);
nor I_928 (I16971,I16953,I16899);
DFFARX1 I_929 (I16971,I251,I16575,I16998,);
nor I_930 (I17007,I16953,I16476);
and I_931 (I17025,I17007,I16386);
or I_932 (I17043,I17025,I16521);
DFFARX1 I_933 (I17043,I251,I16575,I17070,);
nor I_934 (I17079,I17070,I16656);
nor I_935 (I17097,I16602,I17079);
not I_936 (I17115,I17070);
nor I_937 (I17133,I17115,I16773);
DFFARX1 I_938 (I17133,I251,I16575,I17160,);
nand I_939 (I17169,I17115,I16701);
nor I_940 (I17187,I16953,I17169);
not I_941 (I17205,I258);
DFFARX1 I_942 (I17187,I251,I17205,I17232,);
and I_943 (I17241,I17232,I16890);
DFFARX1 I_944 (I17241,I251,I17205,I17268,);
DFFARX1 I_945 (I17097,I251,I17205,I17286,);
not I_946 (I17295,I17187);
not I_947 (I17313,I16800);
nand I_948 (I17331,I17313,I17295);
nor I_949 (I17349,I17286,I17331);
DFFARX1 I_950 (I17331,I251,I17205,I17376,);
not I_951 (I17385,I17376);
not I_952 (I17403,I16935);
nand I_953 (I17421,I17313,I17403);
DFFARX1 I_954 (I17421,I251,I17205,I17448,);
not I_955 (I17457,I17448);
not I_956 (I17475,I16629);
nand I_957 (I17493,I17475,I16998);
and I_958 (I17511,I17295,I17493);
nor I_959 (I17529,I17421,I17511);
DFFARX1 I_960 (I17529,I251,I17205,I17556,);
DFFARX1 I_961 (I17511,I251,I17205,I17574,);
nor I_962 (I17583,I16629,I16998);
nor I_963 (I17601,I17421,I17583);
or I_964 (I17619,I16629,I16998);
nor I_965 (I17637,I16863,I17160);
DFFARX1 I_966 (I17637,I251,I17205,I17664,);
not I_967 (I17673,I17664);
nor I_968 (I17691,I17673,I17457);
nand I_969 (I17709,I17673,I17286);
not I_970 (I17727,I16863);
nand I_971 (I17745,I17727,I17403);
nand I_972 (I17763,I17673,I17745);
nand I_973 (I17781,I17763,I17709);
nand I_974 (I17799,I17745,I17619);
not I_975 (I17817,I258);
DFFARX1 I_976 (I17691,I251,I17817,I17844,);
not I_977 (I17853,I17844);
nand I_978 (I17871,I17556,I17601);
and I_979 (I17889,I17871,I17268);
DFFARX1 I_980 (I17889,I251,I17817,I17916,);
not I_981 (I17925,I17781);
DFFARX1 I_982 (I17799,I251,I17817,I17952,);
not I_983 (I17961,I17952);
nor I_984 (I17979,I17961,I17853);
and I_985 (I17997,I17979,I17781);
nor I_986 (I18015,I17961,I17925);
nor I_987 (I18033,I17916,I18015);
DFFARX1 I_988 (I17385,I251,I17817,I18060,);
nor I_989 (I18069,I18060,I17916);
not I_990 (I18087,I18069);
not I_991 (I18105,I18060);
nor I_992 (I18123,I18105,I17997);
DFFARX1 I_993 (I18123,I251,I17817,I18150,);
nand I_994 (I18159,I17349,I17349);
and I_995 (I18177,I18159,I17556);
DFFARX1 I_996 (I18177,I251,I17817,I18204,);
nor I_997 (I18213,I18204,I18060);
DFFARX1 I_998 (I18213,I251,I17817,I18240,);
nand I_999 (I18249,I18204,I18105);
nand I_1000 (I18267,I18087,I18249);
not I_1001 (I18285,I18204);
nor I_1002 (I18303,I18285,I17997);
DFFARX1 I_1003 (I18303,I251,I17817,I18330,);
nor I_1004 (I18339,I17574,I17349);
or I_1005 (I18357,I18060,I18339);
nor I_1006 (I18375,I18204,I18339);
or I_1007 (I18393,I17916,I18339);
DFFARX1 I_1008 (I18339,I251,I17817,I18420,);
not I_1009 (I18429,I258);
DFFARX1 I_1010 (I18357,I251,I18429,I18456,);
nand I_1011 (I18465,I18375,I18150);
and I_1012 (I18483,I18465,I18420);
DFFARX1 I_1013 (I18483,I251,I18429,I18510,);
nor I_1014 (I18519,I18510,I18456);
not I_1015 (I18537,I18510);
DFFARX1 I_1016 (I18267,I251,I18429,I18564,);
nand I_1017 (I18573,I18564,I18375);
not I_1018 (I18591,I18573);
DFFARX1 I_1019 (I18591,I251,I18429,I18618,);
not I_1020 (I18627,I18618);
nor I_1021 (I18645,I18456,I18573);
nor I_1022 (I18663,I18510,I18645);
DFFARX1 I_1023 (I18393,I251,I18429,I18690,);
DFFARX1 I_1024 (I18690,I251,I18429,I18708,);
not I_1025 (I18717,I18708);
not I_1026 (I18735,I18690);
nand I_1027 (I18753,I18735,I18537);
nand I_1028 (I18771,I18240,I18033);
and I_1029 (I18789,I18771,I18240);
DFFARX1 I_1030 (I18789,I251,I18429,I18816,);
nor I_1031 (I18825,I18816,I18456);
DFFARX1 I_1032 (I18825,I251,I18429,I18852,);
DFFARX1 I_1033 (I18816,I251,I18429,I18870,);
nor I_1034 (I18879,I18330,I18033);
not I_1035 (I18897,I18879);
nor I_1036 (I18915,I18717,I18897);
nand I_1037 (I18933,I18735,I18897);
nor I_1038 (I18951,I18456,I18879);
DFFARX1 I_1039 (I18879,I251,I18429,I18978,);
not I_1040 (I18987,I258);
DFFARX1 I_1041 (I18915,I251,I18987,I19014,);
DFFARX1 I_1042 (I19014,I251,I18987,I19032,);
not I_1043 (I19041,I19032);
not I_1044 (I19059,I19014);
nand I_1045 (I19077,I18852,I18978);
and I_1046 (I19095,I19077,I18627);
DFFARX1 I_1047 (I19095,I251,I18987,I19122,);
not I_1048 (I19131,I19122);
DFFARX1 I_1049 (I18663,I251,I18987,I19158,);
and I_1050 (I19167,I19158,I18951);
nand I_1051 (I19185,I19158,I18951);
nand I_1052 (I19203,I19131,I19185);
DFFARX1 I_1053 (I18519,I251,I18987,I19230,);
nor I_1054 (I19239,I19230,I19167);
DFFARX1 I_1055 (I19239,I251,I18987,I19266,);
nor I_1056 (I19275,I19230,I19122);
nand I_1057 (I19293,I18753,I18852);
and I_1058 (I19311,I19293,I18933);
DFFARX1 I_1059 (I19311,I251,I18987,I19338,);
nor I_1060 (I19347,I19338,I19230);
not I_1061 (I19365,I19338);
nor I_1062 (I19383,I19365,I19131);
nor I_1063 (I19401,I19059,I19383);
DFFARX1 I_1064 (I19401,I251,I18987,I19428,);
nor I_1065 (I19437,I19365,I19230);
nor I_1066 (I19455,I18870,I18852);
nor I_1067 (I19473,I19455,I19437);
not I_1068 (I19491,I19455);
nand I_1069 (I19509,I19185,I19491);
DFFARX1 I_1070 (I19455,I251,I18987,I19536,);
DFFARX1 I_1071 (I19455,I251,I18987,I19554,);
not I_1072 (I19563,I258);
DFFARX1 I_1073 (I19509,I251,I19563,I19590,);
nand I_1074 (I19599,I19536,I19347);
and I_1075 (I19617,I19599,I19041);
DFFARX1 I_1076 (I19617,I251,I19563,I19644,);
nor I_1077 (I19653,I19644,I19590);
not I_1078 (I19671,I19644);
DFFARX1 I_1079 (I19428,I251,I19563,I19698,);
nand I_1080 (I19707,I19698,I19266);
not I_1081 (I19725,I19707);
DFFARX1 I_1082 (I19725,I251,I19563,I19752,);
not I_1083 (I19761,I19752);
nor I_1084 (I19779,I19590,I19707);
nor I_1085 (I19797,I19644,I19779);
DFFARX1 I_1086 (I19275,I251,I19563,I19824,);
DFFARX1 I_1087 (I19824,I251,I19563,I19842,);
not I_1088 (I19851,I19842);
not I_1089 (I19869,I19824);
nand I_1090 (I19887,I19869,I19671);
nand I_1091 (I19905,I19266,I19203);
and I_1092 (I19923,I19905,I19473);
DFFARX1 I_1093 (I19923,I251,I19563,I19950,);
nor I_1094 (I19959,I19950,I19590);
DFFARX1 I_1095 (I19959,I251,I19563,I19986,);
DFFARX1 I_1096 (I19950,I251,I19563,I20004,);
nor I_1097 (I20013,I19554,I19203);
not I_1098 (I20031,I20013);
nor I_1099 (I20049,I19851,I20031);
nand I_1100 (I20067,I19869,I20031);
nor I_1101 (I20085,I19590,I20013);
DFFARX1 I_1102 (I20013,I251,I19563,I20112,);
not I_1103 (I20121,I258);
DFFARX1 I_1104 (I19887,I251,I20121,I20148,);
nand I_1105 (I20157,I20148,I20085);
DFFARX1 I_1106 (I19797,I251,I20121,I20184,);
DFFARX1 I_1107 (I20184,I251,I20121,I20202,);
not I_1108 (I20211,I20202);
not I_1109 (I20229,I20004);
nor I_1110 (I20247,I20004,I19653);
not I_1111 (I20265,I19761);
nand I_1112 (I20283,I20229,I20265);
nor I_1113 (I20301,I19761,I20004);
and I_1114 (I20319,I20301,I20157);
not I_1115 (I20337,I20067);
nand I_1116 (I20355,I20337,I20112);
nor I_1117 (I20373,I20067,I19986);
not I_1118 (I20391,I20373);
nand I_1119 (I20409,I20247,I20391);
DFFARX1 I_1120 (I20373,I251,I20121,I20436,);
nor I_1121 (I20445,I20049,I19761);
nor I_1122 (I20463,I20445,I19653);
and I_1123 (I20481,I20463,I20355);
DFFARX1 I_1124 (I20481,I251,I20121,I20508,);
nor I_1125 (I20517,I20445,I20283);
or I_1126 (I20535,I20373,I20445);
nor I_1127 (I20553,I20049,I19986);
DFFARX1 I_1128 (I20553,I251,I20121,I20580,);
not I_1129 (I20589,I20580);
nand I_1130 (I20607,I20589,I20229);
nor I_1131 (I20625,I20607,I19653);
DFFARX1 I_1132 (I20625,I251,I20121,I20652,);
nor I_1133 (I20661,I20589,I20283);
nor I_1134 (I20679,I20445,I20661);
not I_1135 (I20697,I258);
DFFARX1 I_1136 (I20535,I251,I20697,I20724,);
not I_1137 (I20733,I20724);
nand I_1138 (I20751,I20508,I20652);
and I_1139 (I20769,I20751,I20679);
DFFARX1 I_1140 (I20769,I251,I20697,I20796,);
DFFARX1 I_1141 (I20796,I251,I20697,I20814,);
DFFARX1 I_1142 (I20517,I251,I20697,I20832,);
nand I_1143 (I20841,I20832,I20319);
not I_1144 (I20859,I20841);
DFFARX1 I_1145 (I20859,I251,I20697,I20886,);
not I_1146 (I20895,I20886);
nor I_1147 (I20913,I20733,I20895);
DFFARX1 I_1148 (I20436,I251,I20697,I20940,);
nor I_1149 (I20949,I20940,I20796);
nor I_1150 (I20967,I20940,I20859);
nand I_1151 (I20985,I20652,I20409);
and I_1152 (I21003,I20985,I20211);
DFFARX1 I_1153 (I21003,I251,I20697,I21030,);
not I_1154 (I21039,I21030);
nand I_1155 (I21057,I21039,I20940);
nand I_1156 (I21075,I21039,I20841);
nor I_1157 (I21093,I20319,I20409);
and I_1158 (I21111,I20940,I21093);
nor I_1159 (I21129,I21039,I21111);
DFFARX1 I_1160 (I21129,I251,I20697,I21156,);
nor I_1161 (I21165,I20724,I21093);
DFFARX1 I_1162 (I21165,I251,I20697,I21192,);
nor I_1163 (I21201,I21030,I21093);
not I_1164 (I21219,I21201);
nand I_1165 (I21237,I21219,I21057);
not I_1166 (I21255,I258);
DFFARX1 I_1167 (I21075,I251,I21255,I21282,);
DFFARX1 I_1168 (I20967,I251,I21255,I21300,);
not I_1169 (I21309,I21300);
not I_1170 (I21327,I20967);
nor I_1171 (I21345,I21327,I21075);
not I_1172 (I21363,I20814);
nor I_1173 (I21381,I21345,I20949);
nor I_1174 (I21399,I21300,I21381);
DFFARX1 I_1175 (I21399,I251,I21255,I21426,);
nor I_1176 (I21435,I20949,I21075);
nand I_1177 (I21453,I21435,I20967);
DFFARX1 I_1178 (I21453,I251,I21255,I21480,);
nor I_1179 (I21489,I21363,I20949);
nand I_1180 (I21507,I21489,I21192);
nor I_1181 (I21525,I21282,I21507);
DFFARX1 I_1182 (I21525,I251,I21255,I21552,);
not I_1183 (I21561,I21507);
nand I_1184 (I21579,I21300,I21561);
DFFARX1 I_1185 (I21507,I251,I21255,I21606,);
not I_1186 (I21615,I21606);
not I_1187 (I21633,I20949);
not I_1188 (I21651,I21237);
nor I_1189 (I21669,I21651,I20814);
nor I_1190 (I21687,I21615,I21669);
nor I_1191 (I21705,I21651,I21156);
and I_1192 (I21723,I21705,I20913);
or I_1193 (I21741,I21723,I21192);
DFFARX1 I_1194 (I21741,I251,I21255,I21768,);
nor I_1195 (I21777,I21768,I21282);
not I_1196 (I21795,I21768);
and I_1197 (I21813,I21795,I21282);
nor I_1198 (I21831,I21309,I21813);
nand I_1199 (I21849,I21795,I21363);
nor I_1200 (I21867,I21651,I21849);
nand I_1201 (I21885,I21795,I21561);
nand I_1202 (I21903,I21363,I21237);
nor I_1203 (I21921,I21633,I21903);
not I_1204 (I21939,I258);
DFFARX1 I_1205 (I21885,I251,I21939,I21966,);
DFFARX1 I_1206 (I21480,I251,I21939,I21984,);
not I_1207 (I21993,I21984);
nor I_1208 (I22011,I21966,I21993);
DFFARX1 I_1209 (I21993,I251,I21939,I22038,);
nor I_1210 (I22047,I21867,I21777);
and I_1211 (I22065,I22047,I21552);
nor I_1212 (I22083,I22065,I21867);
not I_1213 (I22101,I21867);
and I_1214 (I22119,I22101,I21831);
nand I_1215 (I22137,I22119,I21426);
nor I_1216 (I22155,I22101,I22137);
DFFARX1 I_1217 (I22155,I251,I21939,I22182,);
not I_1218 (I22191,I22137);
nand I_1219 (I22209,I21993,I22191);
nand I_1220 (I22227,I22065,I22191);
DFFARX1 I_1221 (I22101,I251,I21939,I22254,);
not I_1222 (I22263,I21579);
nor I_1223 (I22281,I22263,I21831);
nor I_1224 (I22299,I22281,I22083);
DFFARX1 I_1225 (I22299,I251,I21939,I22326,);
not I_1226 (I22335,I22281);
DFFARX1 I_1227 (I22335,I251,I21939,I22362,);
not I_1228 (I22371,I22362);
nor I_1229 (I22389,I22371,I22281);
nor I_1230 (I22407,I22263,I21552);
and I_1231 (I22425,I22407,I21687);
or I_1232 (I22443,I22425,I21921);
DFFARX1 I_1233 (I22443,I251,I21939,I22470,);
not I_1234 (I22479,I22470);
nand I_1235 (I22497,I22479,I22191);
not I_1236 (I22515,I22497);
nand I_1237 (I22533,I22497,I22209);
nand I_1238 (I22551,I22479,I22065);
not I_1239 (I22569,I258);
DFFARX1 I_1240 (I22254,I251,I22569,I22596,);
not I_1241 (I22605,I22596);
nand I_1242 (I22623,I22227,I22182);
and I_1243 (I22641,I22623,I22515);
DFFARX1 I_1244 (I22641,I251,I22569,I22668,);
not I_1245 (I22677,I22182);
DFFARX1 I_1246 (I22038,I251,I22569,I22704,);
not I_1247 (I22713,I22704);
nor I_1248 (I22731,I22713,I22605);
and I_1249 (I22749,I22731,I22182);
nor I_1250 (I22767,I22713,I22677);
nor I_1251 (I22785,I22668,I22767);
DFFARX1 I_1252 (I22551,I251,I22569,I22812,);
nor I_1253 (I22821,I22812,I22668);
not I_1254 (I22839,I22821);
not I_1255 (I22857,I22812);
nor I_1256 (I22875,I22857,I22749);
DFFARX1 I_1257 (I22875,I251,I22569,I22902,);
nand I_1258 (I22911,I22011,I22533);
and I_1259 (I22929,I22911,I22326);
DFFARX1 I_1260 (I22929,I251,I22569,I22956,);
nor I_1261 (I22965,I22956,I22812);
DFFARX1 I_1262 (I22965,I251,I22569,I22992,);
nand I_1263 (I23001,I22956,I22857);
nand I_1264 (I23019,I22839,I23001);
not I_1265 (I23037,I22956);
nor I_1266 (I23055,I23037,I22749);
DFFARX1 I_1267 (I23055,I251,I22569,I23082,);
nor I_1268 (I23091,I22389,I22533);
or I_1269 (I23109,I22812,I23091);
nor I_1270 (I23127,I22956,I23091);
or I_1271 (I23145,I22668,I23091);
DFFARX1 I_1272 (I23091,I251,I22569,I23172,);
endmodule


