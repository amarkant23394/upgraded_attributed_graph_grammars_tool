module test_final(IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_4_2_l_10,IN_5_2_l_10,IN_1_6_l_10,IN_2_6_l_10,IN_3_6_l_10,IN_4_6_l_10,IN_5_6_l_10,IN_1_9_l_10,IN_2_9_l_10,IN_3_9_l_10,IN_4_9_l_10,IN_5_9_l_10,blif_clk_net_5_r_13,blif_reset_net_5_r_13,N1371_0_r_13,N1508_0_r_13,n_429_or_0_5_r_13,G78_5_r_13,n_576_5_r_13,n_547_5_r_13,G42_7_r_13,n_572_7_r_13,n_573_7_r_13,n_549_7_r_13,n_569_7_r_13,n_452_7_r_13);
input IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_4_2_l_10,IN_5_2_l_10,IN_1_6_l_10,IN_2_6_l_10,IN_3_6_l_10,IN_4_6_l_10,IN_5_6_l_10,IN_1_9_l_10,IN_2_9_l_10,IN_3_9_l_10,IN_4_9_l_10,IN_5_9_l_10,blif_clk_net_5_r_13,blif_reset_net_5_r_13;
output N1371_0_r_13,N1508_0_r_13,n_429_or_0_5_r_13,G78_5_r_13,n_576_5_r_13,n_547_5_r_13,G42_7_r_13,n_572_7_r_13,n_573_7_r_13,n_549_7_r_13,n_569_7_r_13,n_452_7_r_13;
wire N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1372_4_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10,I_BUFF_1_9_r_10,N3_8_r_10,n35_10,n36_10,n37_10,n38_10,n39_10,n40_10,n41_10,n42_10,n43_10,n44_10,n45_10,n46_10,n47_10,n48_10,n49_10,n50_10,n51_10,n52_10,n53_10,n54_10,n55_10,n56_10,n57_10,n58_10,n59_10,n60_10,n61_10,n62_10,n63_10,n64_10,n_102_5_r_13,n4_7_l_13,n9_13,n62_13,n33_13,n_431_5_r_13,n1_13,n34_13,n35_13,n36_13,n37_13,n38_13,n39_13,n40_13,n41_13,n42_13,n43_13,n44_13,n45_13,n46_13,n47_13,n48_13,n49_13,n50_13,n51_13,n52_13,n53_13,n54_13,n55_13,n56_13,n57_13,n58_13,n59_13,n60_13,n61_13;
nor I_0(N1371_0_r_10,n37_10,n38_10);
nor I_1(N1508_0_r_10,n37_10,n58_10);
nand I_2(N6147_2_r_10,n39_10,n40_10);
not I_3(N6147_3_r_10,n39_10);
nor I_4(N1372_4_r_10,n46_10,n49_10);
nor I_5(N1508_4_r_10,n51_10,n52_10);
nor I_6(N1507_6_r_10,n49_10,n60_10);
nor I_7(N1508_6_r_10,n49_10,n50_10);
nor I_8(n_42_8_r_10,I_BUFF_1_9_r_10,n35_10);
DFFARX1 I_9(N3_8_r_10,blif_clk_net_5_r_13,n9_13,G199_8_r_10,);
nor I_10(N6147_9_r_10,n36_10,n37_10);
nor I_11(N6134_9_r_10,I_BUFF_1_9_r_10,n46_10);
not I_12(I_BUFF_1_9_r_10,n48_10);
nor I_13(N3_8_r_10,n44_10,n47_10);
not I_14(n35_10,n49_10);
nor I_15(n36_10,I_BUFF_1_9_r_10,n38_10);
not I_16(n37_10,IN_1_9_l_10);
not I_17(n38_10,n46_10);
nand I_18(n39_10,n43_10,n44_10);
nand I_19(n40_10,I_BUFF_1_9_r_10,n41_10);
nor I_20(n41_10,IN_1_9_l_10,n42_10);
not I_21(n42_10,n44_10);
nor I_22(n43_10,IN_1_9_l_10,n45_10);
nand I_23(n44_10,IN_2_6_l_10,n54_10);
nor I_24(n45_10,IN_5_9_l_10,n59_10);
nand I_25(n46_10,IN_2_9_l_10,n61_10);
nor I_26(n47_10,n46_10,n48_10);
nand I_27(n48_10,n62_10,n63_10);
nand I_28(n49_10,IN_5_6_l_10,n56_10);
not I_29(n50_10,n45_10);
nor I_30(n51_10,n42_10,n53_10);
not I_31(n52_10,N1372_4_r_10);
nor I_32(n53_10,n48_10,n50_10);
and I_33(n54_10,IN_1_6_l_10,n55_10);
nand I_34(n55_10,n56_10,n57_10);
nand I_35(n56_10,IN_3_6_l_10,IN_4_6_l_10);
not I_36(n57_10,IN_5_6_l_10);
nor I_37(n58_10,n35_10,n45_10);
nor I_38(n59_10,IN_3_9_l_10,IN_4_9_l_10);
nor I_39(n60_10,n37_10,n46_10);
or I_40(n61_10,IN_3_9_l_10,IN_4_9_l_10);
nor I_41(n62_10,IN_1_2_l_10,IN_2_2_l_10);
or I_42(n63_10,IN_5_2_l_10,n64_10);
nor I_43(n64_10,IN_3_2_l_10,IN_4_2_l_10);
nor I_44(N1371_0_r_13,n59_13,n61_13);
nor I_45(N1508_0_r_13,n59_13,n60_13);
not I_46(n_429_or_0_5_r_13,n46_13);
DFFARX1 I_47(n_431_5_r_13,blif_clk_net_5_r_13,n9_13,G78_5_r_13,);
nand I_48(n_576_5_r_13,n_102_5_r_13,n34_13);
nor I_49(n_102_5_r_13,N1508_0_r_10,N1508_4_r_10);
nand I_50(n_547_5_r_13,n48_13,n49_13);
DFFARX1 I_51(n1_13,blif_clk_net_5_r_13,n9_13,G42_7_r_13,);
nor I_52(n_572_7_r_13,n40_13,n41_13);
nand I_53(n_573_7_r_13,n37_13,n38_13);
nor I_54(n_549_7_r_13,n46_13,n47_13);
nand I_55(n_569_7_r_13,n37_13,n43_13);
nand I_56(n_452_7_r_13,n52_13,n53_13);
nor I_57(n4_7_l_13,N6147_3_r_10,N1507_6_r_10);
not I_58(n9_13,blif_reset_net_5_r_13);
DFFARX1 I_59(n4_7_l_13,blif_clk_net_5_r_13,n9_13,n62_13,);
not I_60(n33_13,n62_13);
nand I_61(n_431_5_r_13,n54_13,n55_13);
not I_62(n1_13,n52_13);
nor I_63(n34_13,n35_13,n36_13);
nor I_64(n35_13,n42_13,N6147_9_r_10);
nand I_65(n36_13,n50_13,n58_13);
nand I_66(n37_13,n44_13,n45_13);
or I_67(n38_13,n39_13,G199_8_r_10);
nand I_68(n39_13,N1371_0_r_10,N1508_0_r_10);
not I_69(n40_13,n36_13);
nor I_70(n41_13,n35_13,N1508_0_r_10);
not I_71(n42_13,N6147_2_r_10);
or I_72(n43_13,N6147_3_r_10,N6134_9_r_10);
not I_73(n44_13,N6147_9_r_10);
not I_74(n45_13,N1371_0_r_10);
nor I_75(n46_13,n39_13,n40_13);
nor I_76(n47_13,N6147_3_r_10,N6134_9_r_10);
nor I_77(n48_13,n50_13,n51_13);
nor I_78(n49_13,N1371_0_r_10,N6147_9_r_10);
not I_79(n50_13,n59_13);
not I_80(n51_13,n_102_5_r_13);
nand I_81(n52_13,n33_13,n39_13);
nand I_82(n53_13,n33_13,G199_8_r_10);
nor I_83(n54_13,N1508_4_r_10,N6134_9_r_10);
nand I_84(n55_13,n62_13,n56_13);
nor I_85(n56_13,n39_13,n57_13);
not I_86(n57_13,N6147_3_r_10);
or I_87(n58_13,N1508_6_r_10,N6147_3_r_10);
nand I_88(n59_13,n_42_8_r_10,N6147_2_r_10);
nor I_89(n60_13,n51_13,N6134_9_r_10);
nor I_90(n61_13,n39_13,G199_8_r_10);
endmodule


