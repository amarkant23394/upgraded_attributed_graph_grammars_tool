module test_I12608(I9465,I9477,I1477,I1470,I11088,I12608);
input I9465,I9477,I1477,I1470,I11088;
output I12608;
wire I12619,I10647,I11105,I12913,I13023,I12930,I10715,I10633,I10766,I10896,I10636,I10732,I11026,I10609;
not I_0(I12619,I1477);
not I_1(I10647,I1477);
and I_2(I11105,I10766,I11088);
DFFARX1 I_3(I10633,I1470,I12619,,,I12913,);
DFFARX1 I_4(I10636,I1470,I12619,,,I13023,);
and I_5(I12930,I12913,I10609);
nor I_6(I12608,I13023,I12930);
nor I_7(I10715,I9477);
nand I_8(I10633,I10896,I11026);
not I_9(I10766,I9477);
DFFARX1 I_10(I1470,I10647,,,I10896,);
nor I_11(I10636,I10732,I10766);
nand I_12(I10732,I10715,I9465);
nor I_13(I11026,I10732);
DFFARX1 I_14(I11105,I1470,I10647,,,I10609,);
endmodule


