module test_I3620(I1383,I1477,I1215,I1423,I1470,I1535,I3620);
input I1383,I1477,I1215,I1423,I1470,I1535;
output I3620;
wire I1518,I1668,I1637,I1880,I1586,I1603,I1492,I1483;
not I_0(I1518,I1477);
not I_1(I1668,I1637);
not I_2(I1637,I1215);
nor I_3(I3620,I1492,I1483);
DFFARX1 I_4(I1383,I1470,I1518,,,I1880,);
nor I_5(I1586,I1535,I1215);
nand I_6(I1603,I1586,I1423);
nand I_7(I1492,I1603,I1668);
DFFARX1 I_8(I1880,I1470,I1518,,,I1483,);
endmodule


