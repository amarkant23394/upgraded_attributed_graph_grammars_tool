module test_I2600(I1342,I1294,I1577,I2600);
input I1342,I1294,I1577;
output I2600;
wire I1911,I2406,I2070,I2389,I1310,I2488;
not I_0(I2600,I1911);
nand I_1(I1911,I2070,I2488);
not I_2(I2406,I2389);
not I_3(I2070,I1310);
DFFARX1 I_4(I1294,,,I2389,);
DFFARX1 I_5(I1577,I1294,I1342,,,I1310,);
not I_6(I2488,I2406);
endmodule


