module test_final(IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_6_2_l_6,IN_1_3_l_6,IN_2_3_l_6,IN_4_3_l_6,IN_1_4_l_6,IN_2_4_l_6,IN_3_4_l_6,IN_6_4_l_6,blif_clk_net_1_r_1,blif_reset_net_1_r_1,G42_1_r_1,n_572_1_r_1,n_573_1_r_1,n_549_1_r_1,n_452_1_r_1,ACVQN2_3_r_1,n_266_and_0_3_r_1,G199_4_r_1,G214_4_r_1);
input IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_6_2_l_6,IN_1_3_l_6,IN_2_3_l_6,IN_4_3_l_6,IN_1_4_l_6,IN_2_4_l_6,IN_3_4_l_6,IN_6_4_l_6,blif_clk_net_1_r_1,blif_reset_net_1_r_1;
output G42_1_r_1,n_572_1_r_1,n_573_1_r_1,n_549_1_r_1,n_452_1_r_1,ACVQN2_3_r_1,n_266_and_0_3_r_1,G199_4_r_1,G214_4_r_1;
wire G42_1_r_6,n_572_1_r_6,n_573_1_r_6,n_549_1_r_6,n_569_1_r_6,n_452_1_r_6,G199_4_r_6,G214_4_r_6,ACVQN1_5_r_6,P6_5_r_6,N3_2_l_6,n27_6,n17_6,n28_6,n26_6,N1_4_l_6,n29_6,n18_6,G214_4_l_6,n12_6,n4_1_r_6,N1_4_r_6,n_42_2_l_6,P6_5_r_internal_6,n19_6,n20_6,n21_6,n22_6,n23_6,n24_6,n25_6,N3_2_l_1,n5_1,n26_1,n17_1,n16_internal_1,n16_1,ACVQN1_3_l_1,N1_4_l_1,G199_4_l_1,G214_4_l_1,n4_1_r_1,n14_internal_1,n14_1,N1_4_r_1,n18_1,n19_1,n20_1,n21_1,n22_1,n23_1,n24_1,n25_1;
DFFARX1 I_0(n4_1_r_6,blif_clk_net_1_r_1,n5_1,G42_1_r_6,);
nor I_1(n_572_1_r_6,n27_6,n28_6);
nand I_2(n_573_1_r_6,n18_6,n19_6);
nor I_3(n_549_1_r_6,n_42_2_l_6,n21_6);
nand I_4(n_569_1_r_6,n19_6,n20_6);
nor I_5(n_452_1_r_6,n28_6,n29_6);
DFFARX1 I_6(N1_4_r_6,blif_clk_net_1_r_1,n5_1,G199_4_r_6,);
DFFARX1 I_7(n_42_2_l_6,blif_clk_net_1_r_1,n5_1,G214_4_r_6,);
DFFARX1 I_8(n_42_2_l_6,blif_clk_net_1_r_1,n5_1,ACVQN1_5_r_6,);
not I_9(P6_5_r_6,P6_5_r_internal_6);
and I_10(N3_2_l_6,IN_6_2_l_6,n23_6);
DFFARX1 I_11(N3_2_l_6,blif_clk_net_1_r_1,n5_1,n27_6,);
not I_12(n17_6,n27_6);
DFFARX1 I_13(IN_1_3_l_6,blif_clk_net_1_r_1,n5_1,n28_6,);
DFFARX1 I_14(IN_2_3_l_6,blif_clk_net_1_r_1,n5_1,n26_6,);
and I_15(N1_4_l_6,IN_6_4_l_6,n25_6);
DFFARX1 I_16(N1_4_l_6,blif_clk_net_1_r_1,n5_1,n29_6,);
not I_17(n18_6,n29_6);
DFFARX1 I_18(IN_3_4_l_6,blif_clk_net_1_r_1,n5_1,G214_4_l_6,);
not I_19(n12_6,G214_4_l_6);
nor I_20(n4_1_r_6,n28_6,n22_6);
nor I_21(N1_4_r_6,n12_6,n24_6);
nor I_22(n_42_2_l_6,IN_1_2_l_6,IN_3_2_l_6);
DFFARX1 I_23(G214_4_l_6,blif_clk_net_1_r_1,n5_1,P6_5_r_internal_6,);
nand I_24(n19_6,IN_4_3_l_6,n26_6);
not I_25(n20_6,n_42_2_l_6);
nor I_26(n21_6,n17_6,n28_6);
and I_27(n22_6,IN_4_3_l_6,n26_6);
nand I_28(n23_6,IN_2_2_l_6,IN_3_2_l_6);
nor I_29(n24_6,n17_6,n18_6);
nand I_30(n25_6,IN_1_4_l_6,IN_2_4_l_6);
DFFARX1 I_31(n4_1_r_1,blif_clk_net_1_r_1,n5_1,G42_1_r_1,);
nor I_32(n_572_1_r_1,n26_1,n19_1);
nand I_33(n_573_1_r_1,n16_1,n18_1);
nor I_34(n_549_1_r_1,n20_1,n21_1);
nor I_35(n_452_1_r_1,G214_4_l_1,n20_1);
DFFARX1 I_36(G199_4_l_1,blif_clk_net_1_r_1,n5_1,ACVQN2_3_r_1,);
nor I_37(n_266_and_0_3_r_1,n16_1,n14_1);
DFFARX1 I_38(N1_4_r_1,blif_clk_net_1_r_1,n5_1,G199_4_r_1,);
DFFARX1 I_39(G199_4_l_1,blif_clk_net_1_r_1,n5_1,G214_4_r_1,);
and I_40(N3_2_l_1,n23_1,n_549_1_r_6);
not I_41(n5_1,blif_reset_net_1_r_1);
DFFARX1 I_42(N3_2_l_1,blif_clk_net_1_r_1,n5_1,n26_1,);
not I_43(n17_1,n26_1);
DFFARX1 I_44(G214_4_r_6,blif_clk_net_1_r_1,n5_1,n16_internal_1,);
not I_45(n16_1,n16_internal_1);
DFFARX1 I_46(n_569_1_r_6,blif_clk_net_1_r_1,n5_1,ACVQN1_3_l_1,);
and I_47(N1_4_l_1,n25_1,ACVQN1_5_r_6);
DFFARX1 I_48(N1_4_l_1,blif_clk_net_1_r_1,n5_1,G199_4_l_1,);
DFFARX1 I_49(G42_1_r_6,blif_clk_net_1_r_1,n5_1,G214_4_l_1,);
nor I_50(n4_1_r_1,n26_1,G214_4_l_1);
DFFARX1 I_51(G214_4_l_1,blif_clk_net_1_r_1,n5_1,n14_internal_1,);
not I_52(n14_1,n14_internal_1);
nor I_53(N1_4_r_1,n17_1,n24_1);
nand I_54(n18_1,ACVQN1_3_l_1,n_452_1_r_6);
nor I_55(n19_1,n_573_1_r_6,P6_5_r_6);
not I_56(n20_1,n18_1);
nor I_57(n21_1,n26_1,n22_1);
not I_58(n22_1,n19_1);
nand I_59(n23_1,n_573_1_r_6,G199_4_r_6);
nor I_60(n24_1,n18_1,n22_1);
nand I_61(n25_1,n_572_1_r_6,G42_1_r_6);
endmodule


