module Benchmark_testing25000(I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1295,I1303,I1311,I1319,I1327,I1335,I1343,I1351,I1359,I1367,I1375,I1383,I1391,I1399,I1407,I1415,I1423,I1431,I1439,I1447,I1455,I1463,I1471,I1479,I1487,I1495,I1503,I1511,I1519,I1527,I1535,I1543,I1551,I1559,I1567,I1575,I1583,I1591,I1599,I1607,I1615,I1623,I1631,I1639,I1647,I1655,I1663,I1671,I1679,I1687,I1695,I1703,I1711,I1719,I1727,I1735,I1743,I1751,I1759,I1767,I1775,I1783,I1791,I1799,I1807,I1815,I1823,I1831,I1839,I1847,I1855,I1863,I1871,I1879,I1887,I1895,I1903,I1911,I1919,I1927,I1935,I1943,I1951,I1959,I1967,I1975,I1983,I1991,I1999,I2007,I2015,I2023,I2031,I2039,I2047,I2055,I2063,I2071,I2079,I2087,I2095,I2103,I2111,I2119,I2127,I2135,I2143,I2151,I2159,I2167,I2175,I2183,I2191,I2199,I2207,I2215,I2223,I2231,I2239,I2247,I2255,I2263,I2271,I2279,I2287,I2295,I2303,I2311,I2319,I2327,I2335,I2343,I2350,I2357,I12479,I12467,I12476,I12485,I12464,I12482,I12473,I12488,I12461,I12470,I12458,I25382,I25370,I25379,I25388,I25367,I25385,I25376,I25391,I25364,I25373,I25361,I71800,I71815,I71797,I71812,I71794,I71791,I71806,I71803,I71809,I71818,I71788,I139033,I139018,I139015,I139012,I139030,I139027,I139006,I139009,I139036,I139021,I139024,I149641,I149626,I149623,I149620,I149638,I149635,I149614,I149617,I149644,I149629,I149632,I248135,I248138,I248132,I248141,I248147,I248150,I248129,I248159,I248156,I248144,I248153,I255071,I255074,I255068,I255077,I255083,I255086,I255065,I255095,I255092,I255080,I255089,I283833,I283836,I283818,I283839,I283830,I283821,I283812,I283842,I283827,I283824,I283815,I292163,I292166,I292148,I292169,I292160,I292151,I292142,I292172,I292157,I292154,I292145,I318331,I318328,I318322,I318349,I318340,I318334,I318337,I318352,I318346,I318343,I318325,I351499,I351472,I351493,I351478,I351475,I351481,I351487,I351502,I351490,I351496,I351484,I379804,I379777,I379798,I379783,I379780,I379786,I379792,I379807,I379795,I379801,I379789,I383952,I383940,I383943,I383928,I383934,I383946,I383955,I383925,I383949,I383937,I383931);
input I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1295,I1303,I1311,I1319,I1327,I1335,I1343,I1351,I1359,I1367,I1375,I1383,I1391,I1399,I1407,I1415,I1423,I1431,I1439,I1447,I1455,I1463,I1471,I1479,I1487,I1495,I1503,I1511,I1519,I1527,I1535,I1543,I1551,I1559,I1567,I1575,I1583,I1591,I1599,I1607,I1615,I1623,I1631,I1639,I1647,I1655,I1663,I1671,I1679,I1687,I1695,I1703,I1711,I1719,I1727,I1735,I1743,I1751,I1759,I1767,I1775,I1783,I1791,I1799,I1807,I1815,I1823,I1831,I1839,I1847,I1855,I1863,I1871,I1879,I1887,I1895,I1903,I1911,I1919,I1927,I1935,I1943,I1951,I1959,I1967,I1975,I1983,I1991,I1999,I2007,I2015,I2023,I2031,I2039,I2047,I2055,I2063,I2071,I2079,I2087,I2095,I2103,I2111,I2119,I2127,I2135,I2143,I2151,I2159,I2167,I2175,I2183,I2191,I2199,I2207,I2215,I2223,I2231,I2239,I2247,I2255,I2263,I2271,I2279,I2287,I2295,I2303,I2311,I2319,I2327,I2335,I2343,I2350,I2357;
output I12479,I12467,I12476,I12485,I12464,I12482,I12473,I12488,I12461,I12470,I12458,I25382,I25370,I25379,I25388,I25367,I25385,I25376,I25391,I25364,I25373,I25361,I71800,I71815,I71797,I71812,I71794,I71791,I71806,I71803,I71809,I71818,I71788,I139033,I139018,I139015,I139012,I139030,I139027,I139006,I139009,I139036,I139021,I139024,I149641,I149626,I149623,I149620,I149638,I149635,I149614,I149617,I149644,I149629,I149632,I248135,I248138,I248132,I248141,I248147,I248150,I248129,I248159,I248156,I248144,I248153,I255071,I255074,I255068,I255077,I255083,I255086,I255065,I255095,I255092,I255080,I255089,I283833,I283836,I283818,I283839,I283830,I283821,I283812,I283842,I283827,I283824,I283815,I292163,I292166,I292148,I292169,I292160,I292151,I292142,I292172,I292157,I292154,I292145,I318331,I318328,I318322,I318349,I318340,I318334,I318337,I318352,I318346,I318343,I318325,I351499,I351472,I351493,I351478,I351475,I351481,I351487,I351502,I351490,I351496,I351484,I379804,I379777,I379798,I379783,I379780,I379786,I379792,I379807,I379795,I379801,I379789,I383952,I383940,I383943,I383928,I383934,I383946,I383955,I383925,I383949,I383937,I383931;
wire I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1295,I1303,I1311,I1319,I1327,I1335,I1343,I1351,I1359,I1367,I1375,I1383,I1391,I1399,I1407,I1415,I1423,I1431,I1439,I1447,I1455,I1463,I1471,I1479,I1487,I1495,I1503,I1511,I1519,I1527,I1535,I1543,I1551,I1559,I1567,I1575,I1583,I1591,I1599,I1607,I1615,I1623,I1631,I1639,I1647,I1655,I1663,I1671,I1679,I1687,I1695,I1703,I1711,I1719,I1727,I1735,I1743,I1751,I1759,I1767,I1775,I1783,I1791,I1799,I1807,I1815,I1823,I1831,I1839,I1847,I1855,I1863,I1871,I1879,I1887,I1895,I1903,I1911,I1919,I1927,I1935,I1943,I1951,I1959,I1967,I1975,I1983,I1991,I1999,I2007,I2015,I2023,I2031,I2039,I2047,I2055,I2063,I2071,I2079,I2087,I2095,I2103,I2111,I2119,I2127,I2135,I2143,I2151,I2159,I2167,I2175,I2183,I2191,I2199,I2207,I2215,I2223,I2231,I2239,I2247,I2255,I2263,I2271,I2279,I2287,I2295,I2303,I2311,I2319,I2327,I2335,I2343,I2350,I2357,I2398,I2415,I363423,I363426,I2432,I363432,I2449,I2466,I2483,I363444,I2381,I2369,I2528,I363453,I2545,I2562,I363441,I363438,I2579,I363450,I2596,I2378,I2627,I2644,I2661,I363447,I2678,I363435,I2387,I2366,I2723,I363429,I2740,I2384,I2771,I2375,I2390,I2816,I2833,I2850,I2867,I2363,I2372,I2360,I2959,I2976,I226977,I226968,I2993,I226971,I3010,I3027,I3044,I226947,I2942,I2930,I3089,I226962,I3106,I3123,I226950,I226965,I3140,I226959,I3157,I2939,I3188,I3205,I3222,I226974,I3239,I226953,I2948,I2927,I3284,I226956,I3301,I2945,I3332,I2936,I2951,I3377,I3394,I3411,I3428,I2924,I2933,I2921,I3520,I3537,I362794,I362797,I3554,I362803,I3571,I3588,I3605,I362815,I3503,I3491,I3650,I362824,I3667,I3684,I362812,I362809,I3701,I362821,I3718,I3500,I3749,I3766,I3783,I362818,I3800,I362806,I3509,I3488,I3845,I362800,I3862,I3506,I3893,I3497,I3512,I3938,I3955,I3972,I3989,I3485,I3494,I3482,I4081,I4098,I333860,I333863,I4115,I333869,I4132,I4149,I4166,I333881,I4064,I4052,I4211,I333890,I4228,I4245,I333878,I333875,I4262,I333887,I4279,I4061,I4310,I4327,I4344,I333884,I4361,I333872,I4070,I4049,I4406,I333866,I4423,I4067,I4454,I4058,I4073,I4499,I4516,I4533,I4550,I4046,I4055,I4043,I4642,I4659,I125804,I125807,I4676,I125801,I4693,I4710,I4727,I125792,I4625,I4613,I4772,I125780,I4789,I4806,I125789,I125783,I4823,I125795,I4840,I4622,I4871,I4888,I4905,I125810,I4922,I125798,I4631,I4610,I4967,I125786,I4984,I4628,I5015,I4619,I4634,I5060,I5077,I5094,I5111,I4607,I4616,I4604,I5203,I5220,I169528,I169519,I5237,I169534,I5254,I5271,I5288,I169504,I5186,I5174,I5333,I169507,I5350,I5367,I169525,I169522,I5384,I169510,I5401,I5183,I5432,I5449,I5466,I169531,I5483,I169516,I5192,I5171,I5528,I169513,I5545,I5189,I5576,I5180,I5195,I5621,I5638,I5655,I5672,I5168,I5177,I5165,I5764,I5781,I221809,I221800,I5798,I221803,I5815,I5832,I5849,I221779,I5747,I5735,I5894,I221794,I5911,I5928,I221782,I221797,I5945,I221791,I5962,I5744,I5993,I6010,I6027,I221806,I6044,I221785,I5753,I5732,I6089,I221788,I6106,I5750,I6137,I5741,I5756,I6182,I6199,I6216,I6233,I5729,I5738,I5726,I6325,I6342,I319533,I319521,I6359,I319518,I6376,I6393,I6410,I319539,I6308,I6296,I6455,I319542,I6472,I6489,I319512,I319530,I6506,I319527,I6523,I6305,I6554,I6571,I6588,I319536,I6605,I319524,I6314,I6293,I6650,I319515,I6667,I6311,I6698,I6302,I6317,I6743,I6760,I6777,I6794,I6290,I6299,I6287,I6886,I6903,I215349,I215340,I6920,I215343,I6937,I6954,I6971,I215319,I6869,I6857,I7016,I215334,I7033,I7050,I215322,I215337,I7067,I215331,I7084,I6866,I7115,I7132,I7149,I215346,I7166,I215325,I6875,I6854,I7211,I215328,I7228,I6872,I7259,I6863,I6878,I7304,I7321,I7338,I7355,I6851,I6860,I6848,I7447,I7464,I36925,I36928,I7481,I36910,I7498,I7515,I7532,I36907,I7430,I7418,I7577,I36931,I7594,I7611,I36916,I36922,I7628,I36934,I7645,I7427,I7676,I7693,I7710,I36913,I7727,I36904,I7436,I7415,I7772,I36919,I7789,I7433,I7820,I7424,I7439,I7865,I7882,I7899,I7916,I7412,I7421,I7409,I8008,I8025,I45323,I45326,I8042,I45308,I8059,I8076,I8093,I45305,I7991,I7979,I8138,I45329,I8155,I8172,I45314,I45320,I8189,I45332,I8206,I7988,I8237,I8254,I8271,I45311,I8288,I45302,I7997,I7976,I8333,I45317,I8350,I7994,I8381,I7985,I8000,I8426,I8443,I8460,I8477,I7973,I7982,I7970,I8569,I8586,I111900,I111897,I8603,I111894,I8620,I8637,I8654,I111918,I8552,I8540,I8699,I111912,I8716,I8733,I111891,I111903,I8750,I111906,I8767,I8549,I8798,I8815,I8832,I111915,I8849,I111921,I8558,I8537,I8894,I111909,I8911,I8555,I8942,I8546,I8561,I8987,I9004,I9021,I9038,I8534,I8543,I8531,I9130,I9147,I345182,I345185,I9164,I345191,I9181,I9198,I9215,I345203,I9113,I9101,I9260,I345212,I9277,I9294,I345200,I345197,I9311,I345209,I9328,I9110,I9359,I9376,I9393,I345206,I9410,I345194,I9119,I9098,I9455,I345188,I9472,I9116,I9503,I9107,I9122,I9548,I9565,I9582,I9599,I9095,I9104,I9092,I9691,I9708,I119259,I119262,I9725,I119256,I9742,I9759,I9776,I119247,I9674,I9662,I9821,I119235,I9838,I9855,I119244,I119238,I9872,I119250,I9889,I9671,I9920,I9937,I9954,I119265,I9971,I119253,I9680,I9659,I10016,I119241,I10033,I9677,I10064,I9668,I9683,I10109,I10126,I10143,I10160,I9656,I9665,I9653,I10252,I10269,I78269,I78272,I10286,I78254,I10303,I10320,I10337,I78251,I10235,I10223,I10382,I78275,I10399,I10416,I78260,I78266,I10433,I78278,I10450,I10232,I10481,I10498,I10515,I78257,I10532,I78248,I10241,I10220,I10577,I78263,I10594,I10238,I10625,I10229,I10244,I10670,I10687,I10704,I10721,I10217,I10226,I10214,I10813,I10830,I242939,I242936,I10847,I242930,I10864,I10881,I10898,I242942,I10796,I10784,I10943,I242954,I10960,I10977,I242945,I242927,I10994,I242957,I11011,I10793,I11042,I11059,I11076,I242933,I11093,I242951,I10802,I10781,I11138,I242948,I11155,I10799,I11186,I10790,I10805,I11231,I11248,I11265,I11282,I10778,I10787,I10775,I11374,I11391,I175495,I175486,I11408,I175501,I11425,I11442,I11459,I175471,I11357,I11345,I11504,I175474,I11521,I11538,I175492,I175489,I11555,I175477,I11572,I11354,I11603,I11620,I11637,I175498,I11654,I175483,I11363,I11342,I11699,I175480,I11716,I11360,I11747,I11351,I11366,I11792,I11809,I11826,I11843,I11339,I11348,I11336,I11935,I11952,I157594,I157585,I11969,I157600,I11986,I12003,I12020,I157570,I11918,I11906,I12065,I157573,I12082,I12099,I157591,I157588,I12116,I157576,I12133,I11915,I12164,I12181,I12198,I157597,I12215,I157582,I11924,I11903,I12260,I157579,I12277,I11921,I12308,I11912,I11927,I12353,I12370,I12387,I12404,I11900,I11909,I11897,I12496,I12513,I311780,I311783,I12530,I311795,I12547,I12564,I12581,I311789,I12626,I311792,I12643,I12660,I311786,I311804,I12677,I311807,I12694,I12725,I12742,I12759,I311777,I12776,I311798,I12821,I311801,I12838,I12869,I12914,I12931,I12948,I12965,I13057,I13074,I128779,I128782,I13091,I128776,I13108,I13125,I13142,I128767,I13040,I13028,I13187,I128755,I13204,I13221,I128764,I128758,I13238,I128770,I13255,I13037,I13286,I13303,I13320,I128785,I13337,I128773,I13046,I13025,I13382,I128761,I13399,I13043,I13430,I13034,I13049,I13475,I13492,I13509,I13526,I13022,I13031,I13019,I13618,I13635,I336376,I336379,I13652,I336385,I13669,I13686,I13703,I336397,I13601,I13589,I13748,I336406,I13765,I13782,I336394,I336391,I13799,I336403,I13816,I13598,I13847,I13864,I13881,I336400,I13898,I336388,I13607,I13586,I13943,I336382,I13960,I13604,I13991,I13595,I13610,I14036,I14053,I14070,I14087,I13583,I13592,I13580,I14179,I14196,I195969,I195960,I14213,I195963,I14230,I14247,I14264,I195939,I14162,I14150,I14309,I195954,I14326,I14343,I195942,I195957,I14360,I195951,I14377,I14159,I14408,I14425,I14442,I195966,I14459,I195945,I14168,I14147,I14504,I195948,I14521,I14165,I14552,I14156,I14171,I14597,I14614,I14631,I14648,I14144,I14153,I14141,I14740,I14757,I244673,I244670,I14774,I244664,I14791,I14808,I14825,I244676,I14723,I14711,I14870,I244688,I14887,I14904,I244679,I244661,I14921,I244691,I14938,I14720,I14969,I14986,I15003,I244667,I15020,I244685,I14729,I14708,I15065,I244682,I15082,I14726,I15113,I14717,I14732,I15158,I15175,I15192,I15209,I14705,I14714,I14702,I15301,I15318,I390870,I390891,I15335,I390879,I15352,I15369,I15386,I390885,I15284,I15272,I15431,I390873,I15448,I15465,I390864,I390882,I15482,I390876,I15499,I15281,I15530,I15547,I15564,I390888,I15581,I390861,I15290,I15269,I15626,I390867,I15643,I15287,I15674,I15278,I15293,I15719,I15736,I15753,I15770,I15266,I15275,I15263,I15862,I15879,I326673,I326661,I15896,I326658,I15913,I15930,I15947,I326679,I15845,I15833,I15992,I326682,I16009,I16026,I326652,I326670,I16043,I326667,I16060,I15842,I16091,I16108,I16125,I326676,I16142,I326664,I15851,I15830,I16187,I326655,I16204,I15848,I16235,I15839,I15854,I16280,I16297,I16314,I16331,I15827,I15836,I15824,I16423,I16440,I224393,I224384,I16457,I224387,I16474,I16491,I16508,I224363,I16406,I16394,I16553,I224378,I16570,I16587,I224366,I224381,I16604,I224375,I16621,I16403,I16652,I16669,I16686,I224390,I16703,I224369,I16412,I16391,I16748,I224372,I16765,I16409,I16796,I16400,I16415,I16841,I16858,I16875,I16892,I16388,I16397,I16385,I16984,I17001,I78915,I78918,I17018,I78900,I17035,I17052,I17069,I78897,I16967,I16955,I17114,I78921,I17131,I17148,I78906,I78912,I17165,I78924,I17182,I16964,I17213,I17230,I17247,I78903,I17264,I78894,I16973,I16952,I17309,I78909,I17326,I16970,I17357,I16961,I16976,I17402,I17419,I17436,I17453,I16949,I16958,I16946,I17545,I17562,I197907,I197898,I17579,I197901,I17596,I17613,I17630,I197877,I17528,I17516,I17675,I197892,I17692,I17709,I197880,I197895,I17726,I197889,I17743,I17525,I17774,I17791,I17808,I197904,I17825,I197883,I17534,I17513,I17870,I197886,I17887,I17531,I17918,I17522,I17537,I17963,I17980,I17997,I18014,I17510,I17519,I17507,I18106,I18123,I306425,I306428,I18140,I306440,I18157,I18174,I18191,I306434,I18089,I18077,I18236,I306437,I18253,I18270,I306431,I306449,I18287,I306452,I18304,I18086,I18335,I18352,I18369,I306422,I18386,I306443,I18095,I18074,I18431,I306446,I18448,I18092,I18479,I18083,I18098,I18524,I18541,I18558,I18575,I18071,I18080,I18068,I18667,I18684,I278460,I278463,I18701,I278475,I18718,I18735,I18752,I278469,I18650,I18638,I18797,I278472,I18814,I18831,I278466,I278484,I18848,I278487,I18865,I18647,I18896,I18913,I18930,I278457,I18947,I278478,I18656,I18635,I18992,I278481,I19009,I18653,I19040,I18644,I18659,I19085,I19102,I19119,I19136,I18632,I18641,I18629,I19228,I19245,I382200,I382221,I19262,I382209,I19279,I19296,I19313,I382215,I19211,I19199,I19358,I382203,I19375,I19392,I382194,I382212,I19409,I382206,I19426,I19208,I19457,I19474,I19491,I382218,I19508,I382191,I19217,I19196,I19553,I382197,I19570,I19214,I19601,I19205,I19220,I19646,I19663,I19680,I19697,I19193,I19202,I19190,I19789,I19806,I109911,I109908,I19823,I109905,I19840,I19857,I19874,I109929,I19772,I19760,I19919,I109923,I19936,I19953,I109902,I109914,I19970,I109917,I19987,I19769,I20018,I20035,I20052,I109926,I20069,I109932,I19778,I19757,I20114,I109920,I20131,I19775,I20162,I19766,I19781,I20207,I20224,I20241,I20258,I19754,I19763,I19751,I20350,I20367,I226331,I226322,I20384,I226325,I20401,I20418,I20435,I226301,I20333,I20321,I20480,I226316,I20497,I20514,I226304,I226319,I20531,I226313,I20548,I20330,I20579,I20596,I20613,I226328,I20630,I226307,I20339,I20318,I20675,I226310,I20692,I20336,I20723,I20327,I20342,I20768,I20785,I20802,I20819,I20315,I20324,I20312,I20911,I20928,I353359,I353362,I20945,I353368,I20962,I20979,I20996,I353380,I20894,I20882,I21041,I353389,I21058,I21075,I353377,I353374,I21092,I353386,I21109,I20891,I21140,I21157,I21174,I353383,I21191,I353371,I20900,I20879,I21236,I353365,I21253,I20897,I21284,I20888,I20903,I21329,I21346,I21363,I21380,I20876,I20885,I20873,I21472,I21489,I280245,I280248,I21506,I280260,I21523,I21540,I21557,I280254,I21455,I21443,I21602,I280257,I21619,I21636,I280251,I280269,I21653,I280272,I21670,I21452,I21701,I21718,I21735,I280242,I21752,I280263,I21461,I21440,I21797,I280266,I21814,I21458,I21845,I21449,I21464,I21890,I21907,I21924,I21941,I21437,I21446,I21434,I22033,I22050,I237066,I237060,I22067,I237072,I22084,I22101,I22118,I237069,I22016,I22004,I22163,I237048,I22180,I22197,I237054,I237063,I22214,I237051,I22231,I22013,I22262,I22279,I22296,I237075,I22313,I237045,I22022,I22001,I22358,I237057,I22375,I22019,I22406,I22010,I22025,I22451,I22468,I22485,I22502,I21998,I22007,I21995,I22594,I22611,I249297,I249294,I22628,I249288,I22645,I22662,I22679,I249300,I22577,I22565,I22724,I249312,I22741,I22758,I249303,I249285,I22775,I249315,I22792,I22574,I22823,I22840,I22857,I249291,I22874,I249309,I22583,I22562,I22919,I249306,I22936,I22580,I22967,I22571,I22586,I23012,I23029,I23046,I23063,I22559,I22568,I22556,I23155,I23172,I231499,I231490,I23189,I231493,I23206,I23223,I23240,I231469,I23138,I23126,I23285,I231484,I23302,I23319,I231472,I231487,I23336,I231481,I23353,I23135,I23384,I23401,I23418,I231496,I23435,I231475,I23144,I23123,I23480,I231478,I23497,I23141,I23528,I23132,I23147,I23573,I23590,I23607,I23624,I23120,I23129,I23117,I23716,I23733,I338892,I338895,I23750,I338901,I23767,I23784,I23801,I338913,I23699,I23687,I23846,I338922,I23863,I23880,I338910,I338907,I23897,I338919,I23914,I23696,I23945,I23962,I23979,I338916,I23996,I338904,I23705,I23684,I24041,I338898,I24058,I23702,I24089,I23693,I23708,I24134,I24151,I24168,I24185,I23681,I23690,I23678,I24277,I24294,I192070,I192061,I24311,I192076,I24328,I24345,I24362,I192046,I24260,I24248,I24407,I192049,I24424,I24441,I192067,I192064,I24458,I192052,I24475,I24257,I24506,I24523,I24540,I192073,I24557,I192058,I24266,I24245,I24602,I192055,I24619,I24263,I24650,I24254,I24269,I24695,I24712,I24729,I24746,I24242,I24251,I24239,I24838,I24855,I113226,I113223,I24872,I113220,I24889,I24906,I24923,I113244,I24821,I24809,I24968,I113238,I24985,I25002,I113217,I113229,I25019,I113232,I25036,I24818,I25067,I25084,I25101,I113241,I25118,I113247,I24827,I24806,I25163,I113235,I25180,I24824,I25211,I24815,I24830,I25256,I25273,I25290,I25307,I24803,I24812,I24800,I25399,I25416,I156931,I156922,I25433,I156937,I25450,I25467,I25484,I156907,I25529,I156910,I25546,I25563,I156928,I156925,I25580,I156913,I25597,I25628,I25645,I25662,I156934,I25679,I156919,I25724,I156916,I25741,I25772,I25817,I25834,I25851,I25868,I25960,I25977,I241208,I25994,I241196,I241202,I26011,I241193,I25934,I26042,I26059,I241199,I25949,I25931,I26104,I26121,I26138,I241211,I26155,I241223,I26172,I241205,I26189,I241220,I26206,I26223,I26240,I25946,I26271,I26288,I26305,I25928,I26336,I25925,I26367,I241214,I26384,I26401,I26418,I25940,I26449,I25937,I26480,I241217,I26497,I26514,I25943,I25952,I25922,I26606,I26623,I163555,I26640,I163552,I163540,I26657,I163543,I26580,I26688,I26705,I163549,I26595,I26577,I26750,I26767,I26784,I163561,I26801,I163537,I26818,I163558,I26835,I163546,I26852,I26869,I26886,I26592,I26917,I26934,I26951,I26574,I26982,I26571,I27013,I163567,I27030,I27047,I27064,I26586,I27095,I26583,I27126,I163564,I27143,I27160,I26589,I26598,I26568,I27252,I27269,I154936,I27286,I154933,I154921,I27303,I154924,I27226,I27334,I27351,I154930,I27241,I27223,I27396,I27413,I27430,I154942,I27447,I154918,I27464,I154939,I27481,I154927,I27498,I27515,I27532,I27238,I27563,I27580,I27597,I27220,I27628,I27217,I27659,I154948,I27676,I27693,I27710,I27232,I27741,I27229,I27772,I154945,I27789,I27806,I27235,I27244,I27214,I27898,I27915,I312399,I27932,I312375,I312381,I27949,I312384,I27872,I27980,I27997,I312393,I27887,I27869,I28042,I28059,I28076,I312372,I28093,I312387,I28110,I312378,I28127,I312390,I28144,I28161,I28178,I27884,I28209,I28226,I28243,I27866,I28274,I27863,I28305,I312402,I28322,I28339,I28356,I27878,I28387,I27875,I28418,I312396,I28435,I28452,I27881,I27890,I27860,I28544,I28561,I335118,I28578,I335133,I335148,I28595,I335136,I28518,I28626,I28643,I335139,I28533,I28515,I28688,I28705,I28722,I335145,I28739,I335142,I28756,I335121,I28773,I335130,I28790,I28807,I28824,I28530,I28855,I28872,I28889,I28512,I28920,I28509,I28951,I335127,I28968,I28985,I29002,I28524,I29033,I28521,I29064,I335124,I29081,I29098,I28527,I28536,I28506,I29190,I29207,I292764,I29224,I292740,I292746,I29241,I292749,I29164,I29272,I29289,I292758,I29179,I29161,I29334,I29351,I29368,I292737,I29385,I292752,I29402,I292743,I29419,I292755,I29436,I29453,I29470,I29176,I29501,I29518,I29535,I29158,I29566,I29155,I29597,I292767,I29614,I29631,I29648,I29170,I29679,I29167,I29710,I292761,I29727,I29744,I29173,I29182,I29152,I29836,I29853,I287409,I29870,I287385,I287391,I29887,I287394,I29810,I29918,I29935,I287403,I29825,I29807,I29980,I29997,I30014,I287382,I30031,I287397,I30048,I287388,I30065,I287400,I30082,I30099,I30116,I29822,I30147,I30164,I30181,I29804,I30212,I29801,I30243,I287412,I30260,I30277,I30294,I29816,I30325,I29813,I30356,I287406,I30373,I30390,I29819,I29828,I29798,I30482,I30499,I263172,I30516,I263160,I263166,I30533,I263157,I30456,I30564,I30581,I263163,I30471,I30453,I30626,I30643,I30660,I263175,I30677,I263187,I30694,I263169,I30711,I263184,I30728,I30745,I30762,I30468,I30793,I30810,I30827,I30450,I30858,I30447,I30889,I263178,I30906,I30923,I30940,I30462,I30971,I30459,I31002,I263181,I31019,I31036,I30465,I30474,I30444,I31128,I31145,I123400,I31162,I123430,I123409,I31179,I123421,I31102,I31210,I31227,I123403,I31117,I31099,I31272,I31289,I31306,I123406,I31323,I123424,I31340,I123415,I31357,I123412,I31374,I31391,I31408,I31114,I31439,I31456,I31473,I31096,I31504,I31093,I31535,I123418,I31552,I31569,I31586,I31108,I31617,I31105,I31648,I123427,I31665,I31682,I31111,I31120,I31090,I31774,I31791,I356504,I31808,I356519,I356534,I31825,I356522,I31748,I31856,I31873,I356525,I31763,I31745,I31918,I31935,I31952,I356531,I31969,I356528,I31986,I356507,I32003,I356516,I32020,I32037,I32054,I31760,I32085,I32102,I32119,I31742,I32150,I31739,I32181,I356513,I32198,I32215,I32232,I31754,I32263,I31751,I32294,I356510,I32311,I32328,I31757,I31766,I31736,I32420,I32437,I236451,I32454,I236433,I236448,I32471,I236457,I32394,I32502,I32519,I236460,I32409,I32391,I32564,I32581,I32598,I236463,I32615,I236439,I32632,I236442,I32649,I236436,I32666,I32683,I32700,I32406,I32731,I32748,I32765,I32388,I32796,I32385,I32827,I236445,I32844,I32861,I32878,I32400,I32909,I32397,I32940,I236454,I32957,I32974,I32403,I32412,I32382,I33066,I33083,I116260,I33100,I116290,I116269,I33117,I116281,I33040,I33148,I33165,I116263,I33055,I33037,I33210,I33227,I33244,I116266,I33261,I116284,I33278,I116275,I33295,I116272,I33312,I33329,I33346,I33052,I33377,I33394,I33411,I33034,I33442,I33031,I33473,I116278,I33490,I33507,I33524,I33046,I33555,I33043,I33586,I116287,I33603,I33620,I33049,I33058,I33028,I33712,I33729,I323692,I33746,I323677,I323704,I33763,I323680,I33686,I33794,I33811,I323695,I33701,I33683,I33856,I33873,I33890,I323707,I33907,I323689,I33924,I323698,I33941,I323683,I33958,I33975,I33992,I33698,I34023,I34040,I34057,I33680,I34088,I33677,I34119,I323686,I34136,I34153,I34170,I33692,I34201,I33689,I34232,I323701,I34249,I34266,I33695,I33704,I33674,I34358,I34375,I34392,I34409,I34332,I34440,I34457,I34347,I34329,I34502,I34519,I34536,I34553,I34570,I34587,I34604,I34621,I34638,I34344,I34669,I34686,I34703,I34326,I34734,I34323,I34765,I34782,I34799,I34816,I34338,I34847,I34335,I34878,I34895,I34912,I34341,I34350,I34320,I35004,I35021,I251034,I35038,I251022,I251028,I35055,I251019,I34978,I35086,I35103,I251025,I34993,I34975,I35148,I35165,I35182,I251037,I35199,I251049,I35216,I251031,I35233,I251046,I35250,I35267,I35284,I34990,I35315,I35332,I35349,I34972,I35380,I34969,I35411,I251040,I35428,I35445,I35462,I34984,I35493,I34981,I35524,I251043,I35541,I35558,I34987,I34996,I34966,I35650,I35667,I35684,I35701,I35624,I35732,I35749,I35639,I35621,I35794,I35811,I35828,I35845,I35862,I35879,I35896,I35913,I35930,I35636,I35961,I35978,I35995,I35618,I36026,I35615,I36057,I36074,I36091,I36108,I35630,I36139,I35627,I36170,I36187,I36204,I35633,I35642,I35612,I36296,I36313,I93345,I36330,I93333,I93339,I36347,I93348,I36270,I36378,I36395,I93336,I36285,I36267,I36440,I36457,I36474,I93357,I36491,I93330,I36508,I93351,I36525,I93342,I36542,I36559,I36576,I36282,I36607,I36624,I36641,I36264,I36672,I36261,I36703,I93327,I36720,I36737,I36754,I36276,I36785,I36273,I36816,I93354,I36833,I36850,I36279,I36288,I36258,I36942,I36959,I166207,I36976,I166204,I166192,I36993,I166195,I37024,I37041,I166201,I37086,I37103,I37120,I166213,I37137,I166189,I37154,I166210,I37171,I166198,I37188,I37205,I37222,I37253,I37270,I37287,I37318,I37349,I166219,I37366,I37383,I37400,I37431,I37462,I166216,I37479,I37496,I37588,I37605,I202417,I37622,I202429,I202411,I37639,I202426,I37562,I37670,I37687,I202414,I37577,I37559,I37732,I37749,I37766,I202423,I37783,I202402,I37800,I202405,I37817,I202408,I37834,I37851,I37868,I37574,I37899,I37916,I37933,I37556,I37964,I37553,I37995,I202399,I38012,I38029,I38046,I37568,I38077,I37565,I38108,I202420,I38125,I38142,I37571,I37580,I37550,I38234,I38251,I216629,I38268,I216641,I216623,I38285,I216638,I38208,I38316,I38333,I216626,I38223,I38205,I38378,I38395,I38412,I216635,I38429,I216614,I38446,I216617,I38463,I216620,I38480,I38497,I38514,I38220,I38545,I38562,I38579,I38202,I38610,I38199,I38641,I216611,I38658,I38675,I38692,I38214,I38723,I38211,I38754,I216632,I38771,I38788,I38217,I38226,I38196,I38880,I38897,I381044,I38914,I381041,I381038,I38931,I381059,I38854,I38962,I38979,I381062,I38869,I38851,I39024,I39041,I39058,I381035,I39075,I381047,I39092,I381056,I39109,I381050,I39126,I39143,I39160,I38866,I39191,I39208,I39225,I38848,I39256,I38845,I39287,I381065,I39304,I39321,I39338,I38860,I39369,I38857,I39400,I381053,I39417,I39434,I38863,I38872,I38842,I39526,I39543,I310614,I39560,I310590,I310596,I39577,I310599,I39500,I39608,I39625,I310608,I39515,I39497,I39670,I39687,I39704,I310587,I39721,I310602,I39738,I310593,I39755,I310605,I39772,I39789,I39806,I39512,I39837,I39854,I39871,I39494,I39902,I39491,I39933,I310617,I39950,I39967,I39984,I39506,I40015,I39503,I40046,I310611,I40063,I40080,I39509,I39518,I39488,I40172,I40189,I256236,I40206,I256224,I256230,I40223,I256221,I40146,I40254,I40271,I256227,I40161,I40143,I40316,I40333,I40350,I256239,I40367,I256251,I40384,I256233,I40401,I256248,I40418,I40435,I40452,I40158,I40483,I40500,I40517,I40140,I40548,I40137,I40579,I256242,I40596,I40613,I40630,I40152,I40661,I40149,I40692,I256245,I40709,I40726,I40155,I40164,I40134,I40818,I40835,I383356,I40852,I383353,I383350,I40869,I383371,I40792,I40900,I40917,I383374,I40807,I40789,I40962,I40979,I40996,I383347,I41013,I383359,I41030,I383368,I41047,I383362,I41064,I41081,I41098,I40804,I41129,I41146,I41163,I40786,I41194,I40783,I41225,I383377,I41242,I41259,I41276,I40798,I41307,I40795,I41338,I383365,I41355,I41372,I40801,I40810,I40780,I41464,I41481,I308829,I41498,I308805,I308811,I41515,I308814,I41438,I41546,I41563,I308823,I41453,I41435,I41608,I41625,I41642,I308802,I41659,I308817,I41676,I308808,I41693,I308820,I41710,I41727,I41744,I41450,I41775,I41792,I41809,I41432,I41840,I41429,I41871,I308832,I41888,I41905,I41922,I41444,I41953,I41441,I41984,I308826,I42001,I42018,I41447,I41456,I41426,I42110,I42127,I288599,I42144,I288575,I288581,I42161,I288584,I42084,I42192,I42209,I288593,I42099,I42081,I42254,I42271,I42288,I288572,I42305,I288587,I42322,I288578,I42339,I288590,I42356,I42373,I42390,I42096,I42421,I42438,I42455,I42078,I42486,I42075,I42517,I288602,I42534,I42551,I42568,I42090,I42599,I42087,I42630,I288596,I42647,I42664,I42093,I42102,I42072,I42756,I42773,I42790,I42807,I42730,I42838,I42855,I42745,I42727,I42900,I42917,I42934,I42951,I42968,I42985,I43002,I43019,I43036,I42742,I43067,I43084,I43101,I42724,I43132,I42721,I43163,I43180,I43197,I43214,I42736,I43245,I42733,I43276,I43293,I43310,I42739,I42748,I42718,I43402,I43419,I364052,I43436,I364067,I364082,I43453,I364070,I43376,I43484,I43501,I364073,I43391,I43373,I43546,I43563,I43580,I364079,I43597,I364076,I43614,I364055,I43631,I364064,I43648,I43665,I43682,I43388,I43713,I43730,I43747,I43370,I43778,I43367,I43809,I364061,I43826,I43843,I43860,I43382,I43891,I43379,I43922,I364058,I43939,I43956,I43385,I43394,I43364,I44048,I44065,I203063,I44082,I203075,I203057,I44099,I203072,I44022,I44130,I44147,I203060,I44037,I44019,I44192,I44209,I44226,I203069,I44243,I203048,I44260,I203051,I44277,I203054,I44294,I44311,I44328,I44034,I44359,I44376,I44393,I44016,I44424,I44013,I44455,I203045,I44472,I44489,I44506,I44028,I44537,I44025,I44568,I203066,I44585,I44602,I44031,I44040,I44010,I44694,I44711,I135306,I44728,I135327,I135300,I44745,I135315,I44668,I44776,I44793,I135330,I44683,I44665,I44838,I44855,I44872,I135303,I44889,I135321,I44906,I135309,I44923,I135312,I44940,I44957,I44974,I44680,I45005,I45022,I45039,I44662,I45070,I44659,I45101,I135324,I45118,I45135,I45152,I44674,I45183,I44671,I45214,I135318,I45231,I45248,I44677,I44686,I44656,I45340,I45357,I256814,I45374,I256802,I256808,I45391,I256799,I45422,I45439,I256805,I45484,I45501,I45518,I256817,I45535,I256829,I45552,I256811,I45569,I256826,I45586,I45603,I45620,I45651,I45668,I45685,I45716,I45747,I256820,I45764,I45781,I45798,I45829,I45860,I256823,I45877,I45894,I45986,I46003,I326072,I46020,I326057,I326084,I46037,I326060,I45960,I46068,I46085,I326075,I45975,I45957,I46130,I46147,I46164,I326087,I46181,I326069,I46198,I326078,I46215,I326063,I46232,I46249,I46266,I45972,I46297,I46314,I46331,I45954,I46362,I45951,I46393,I326066,I46410,I46427,I46444,I45966,I46475,I45963,I46506,I326081,I46523,I46540,I45969,I45978,I45948,I46632,I46649,I385668,I46666,I385665,I385662,I46683,I385683,I46606,I46714,I46731,I385686,I46621,I46603,I46776,I46793,I46810,I385659,I46827,I385671,I46844,I385680,I46861,I385674,I46878,I46895,I46912,I46618,I46943,I46960,I46977,I46600,I47008,I46597,I47039,I385689,I47056,I47073,I47090,I46612,I47121,I46609,I47152,I385677,I47169,I47186,I46615,I46624,I46594,I47278,I47295,I144328,I47312,I144325,I144313,I47329,I144316,I47252,I47360,I47377,I144322,I47267,I47249,I47422,I47439,I47456,I144334,I47473,I144310,I47490,I144331,I47507,I144319,I47524,I47541,I47558,I47264,I47589,I47606,I47623,I47246,I47654,I47243,I47685,I144340,I47702,I47719,I47736,I47258,I47767,I47255,I47798,I144337,I47815,I47832,I47261,I47270,I47240,I47924,I47941,I359649,I47958,I359664,I359679,I47975,I359667,I47898,I48006,I48023,I359670,I47913,I47895,I48068,I48085,I48102,I359676,I48119,I359673,I48136,I359652,I48153,I359661,I48170,I48187,I48204,I47910,I48235,I48252,I48269,I47892,I48300,I47889,I48331,I359658,I48348,I48365,I48382,I47904,I48413,I47901,I48444,I359655,I48461,I48478,I47907,I47916,I47886,I48570,I48587,I184108,I48604,I184105,I184093,I48621,I184096,I48544,I48652,I48669,I184102,I48559,I48541,I48714,I48731,I48748,I184114,I48765,I184090,I48782,I184111,I48799,I184099,I48816,I48833,I48850,I48556,I48881,I48898,I48915,I48538,I48946,I48535,I48977,I184120,I48994,I49011,I49028,I48550,I49059,I48547,I49090,I184117,I49107,I49124,I48553,I48562,I48532,I49216,I49233,I89367,I49250,I89355,I89361,I49267,I89370,I49190,I49298,I49315,I89358,I49205,I49187,I49360,I49377,I49394,I89379,I49411,I89352,I49428,I89373,I49445,I89364,I49462,I49479,I49496,I49202,I49527,I49544,I49561,I49184,I49592,I49181,I49623,I89349,I49640,I49657,I49674,I49196,I49705,I49193,I49736,I89376,I49753,I49770,I49199,I49208,I49178,I49862,I49879,I247566,I49896,I247554,I247560,I49913,I247551,I49836,I49944,I49961,I247557,I49851,I49833,I50006,I50023,I50040,I247569,I50057,I247581,I50074,I247563,I50091,I247578,I50108,I50125,I50142,I49848,I50173,I50190,I50207,I49830,I50238,I49827,I50269,I247572,I50286,I50303,I50320,I49842,I50351,I49839,I50382,I247575,I50399,I50416,I49845,I49854,I49824,I50508,I50525,I244098,I50542,I244086,I244092,I50559,I244083,I50482,I50590,I50607,I244089,I50497,I50479,I50652,I50669,I50686,I244101,I50703,I244113,I50720,I244095,I50737,I244110,I50754,I50771,I50788,I50494,I50819,I50836,I50853,I50476,I50884,I50473,I50915,I244104,I50932,I50949,I50966,I50488,I50997,I50485,I51028,I244107,I51045,I51062,I50491,I50500,I50470,I51154,I51171,I396072,I51188,I396069,I396066,I51205,I396087,I51128,I51236,I51253,I396090,I51143,I51125,I51298,I51315,I51332,I396063,I51349,I396075,I51366,I396084,I51383,I396078,I51400,I51417,I51434,I51140,I51465,I51482,I51499,I51122,I51530,I51119,I51561,I396093,I51578,I51595,I51612,I51134,I51643,I51131,I51674,I396081,I51691,I51708,I51137,I51146,I51116,I51800,I51817,I144991,I51834,I144988,I144976,I51851,I144979,I51774,I51882,I51899,I144985,I51789,I51771,I51944,I51961,I51978,I144997,I51995,I144973,I52012,I144994,I52029,I144982,I52046,I52063,I52080,I51786,I52111,I52128,I52145,I51768,I52176,I51765,I52207,I145003,I52224,I52241,I52258,I51780,I52289,I51777,I52320,I145000,I52337,I52354,I51783,I51792,I51762,I52446,I52463,I248722,I52480,I248710,I248716,I52497,I248707,I52420,I52528,I52545,I248713,I52435,I52417,I52590,I52607,I52624,I248725,I52641,I248737,I52658,I248719,I52675,I248734,I52692,I52709,I52726,I52432,I52757,I52774,I52791,I52414,I52822,I52411,I52853,I248728,I52870,I52887,I52904,I52426,I52935,I52423,I52966,I248731,I52983,I53000,I52429,I52438,I52408,I53092,I53109,I271539,I53126,I271551,I271533,I53143,I271542,I53066,I53174,I53191,I271548,I53081,I53063,I53236,I53253,I53270,I271521,I53287,I271524,I53304,I271530,I53321,I271545,I53338,I53355,I53372,I53078,I53403,I53420,I53437,I53060,I53468,I53057,I53499,I271527,I53516,I53533,I53550,I53072,I53581,I53069,I53612,I271536,I53629,I53646,I53075,I53084,I53054,I53738,I53755,I240630,I53772,I240618,I240624,I53789,I240615,I53712,I53820,I53837,I240621,I53727,I53709,I53882,I53899,I53916,I240633,I53933,I240645,I53950,I240627,I53967,I240642,I53984,I54001,I54018,I53724,I54049,I54066,I54083,I53706,I54114,I53703,I54145,I240636,I54162,I54179,I54196,I53718,I54227,I53715,I54258,I240639,I54275,I54292,I53721,I53730,I53700,I54384,I54401,I54418,I54435,I54358,I54466,I54483,I54373,I54355,I54528,I54545,I54562,I54579,I54596,I54613,I54630,I54647,I54664,I54370,I54695,I54712,I54729,I54352,I54760,I54349,I54791,I54808,I54825,I54842,I54364,I54873,I54361,I54904,I54921,I54938,I54367,I54376,I54346,I55030,I55047,I252768,I55064,I252756,I252762,I55081,I252753,I55004,I55112,I55129,I252759,I55019,I55001,I55174,I55191,I55208,I252771,I55225,I252783,I55242,I252765,I55259,I252780,I55276,I55293,I55310,I55016,I55341,I55358,I55375,I54998,I55406,I54995,I55437,I252774,I55454,I55471,I55488,I55010,I55519,I55007,I55550,I252777,I55567,I55584,I55013,I55022,I54992,I55676,I55693,I340150,I55710,I340165,I340180,I55727,I340168,I55650,I55758,I55775,I340171,I55665,I55647,I55820,I55837,I55854,I340177,I55871,I340174,I55888,I340153,I55905,I340162,I55922,I55939,I55956,I55662,I55987,I56004,I56021,I55644,I56052,I55641,I56083,I340159,I56100,I56117,I56134,I55656,I56165,I55653,I56196,I340156,I56213,I56230,I55659,I55668,I55638,I56322,I56339,I267261,I56356,I267243,I267252,I56373,I267264,I56296,I56404,I56421,I267249,I56311,I56293,I56466,I56483,I56500,I267240,I56517,I267258,I56534,I267246,I56551,I267267,I56568,I56585,I56602,I56308,I56633,I56650,I56667,I56290,I56698,I56287,I56729,I267255,I56746,I56763,I56780,I56302,I56811,I56299,I56842,I267237,I56859,I56876,I56305,I56314,I56284,I56968,I56985,I103290,I57002,I103278,I103284,I57019,I103293,I56942,I57050,I57067,I103281,I56957,I56939,I57112,I57129,I57146,I103302,I57163,I103275,I57180,I103296,I57197,I103287,I57214,I57231,I57248,I56954,I57279,I57296,I57313,I56936,I57344,I56933,I57375,I103272,I57392,I57409,I57426,I56948,I57457,I56945,I57488,I103299,I57505,I57522,I56951,I56960,I56930,I57614,I57631,I329047,I57648,I329032,I329059,I57665,I329035,I57588,I57696,I57713,I329050,I57603,I57585,I57758,I57775,I57792,I329062,I57809,I329044,I57826,I329053,I57843,I329038,I57860,I57877,I57894,I57600,I57925,I57942,I57959,I57582,I57990,I57579,I58021,I329041,I58038,I58055,I58072,I57594,I58103,I57591,I58134,I329056,I58151,I58168,I57597,I57606,I57576,I58260,I58277,I99312,I58294,I99300,I99306,I58311,I99315,I58234,I58342,I58359,I99303,I58249,I58231,I58404,I58421,I58438,I99324,I58455,I99297,I58472,I99318,I58489,I99309,I58506,I58523,I58540,I58246,I58571,I58588,I58605,I58228,I58636,I58225,I58667,I99294,I58684,I58701,I58718,I58240,I58749,I58237,I58780,I99321,I58797,I58814,I58243,I58252,I58222,I58906,I58923,I370971,I58940,I370986,I371001,I58957,I370989,I58880,I58988,I59005,I370992,I58895,I58877,I59050,I59067,I59084,I370998,I59101,I370995,I59118,I370974,I59135,I370983,I59152,I59169,I59186,I58892,I59217,I59234,I59251,I58874,I59282,I58871,I59313,I370980,I59330,I59347,I59364,I58886,I59395,I58883,I59426,I370977,I59443,I59460,I58889,I58898,I58868,I59552,I59569,I387980,I59586,I387977,I387974,I59603,I387995,I59526,I59634,I59651,I387998,I59541,I59523,I59696,I59713,I59730,I387971,I59747,I387983,I59764,I387992,I59781,I387986,I59798,I59815,I59832,I59538,I59863,I59880,I59897,I59520,I59928,I59517,I59959,I388001,I59976,I59993,I60010,I59532,I60041,I59529,I60072,I387989,I60089,I60106,I59535,I59544,I59514,I60198,I60215,I251612,I60232,I251600,I251606,I60249,I251597,I60172,I60280,I60297,I251603,I60187,I60169,I60342,I60359,I60376,I251615,I60393,I251627,I60410,I251609,I60427,I251624,I60444,I60461,I60478,I60184,I60509,I60526,I60543,I60166,I60574,I60163,I60605,I251618,I60622,I60639,I60656,I60178,I60687,I60175,I60718,I251621,I60735,I60752,I60181,I60190,I60160,I60844,I60861,I60878,I60895,I60818,I60926,I60943,I60833,I60815,I60988,I61005,I61022,I61039,I61056,I61073,I61090,I61107,I61124,I60830,I61155,I61172,I61189,I60812,I61220,I60809,I61251,I61268,I61285,I61302,I60824,I61333,I60821,I61364,I61381,I61398,I60827,I60836,I60806,I61490,I61507,I172837,I61524,I172834,I172822,I61541,I172825,I61464,I61572,I61589,I172831,I61479,I61461,I61634,I61651,I61668,I172843,I61685,I172819,I61702,I172840,I61719,I172828,I61736,I61753,I61770,I61476,I61801,I61818,I61835,I61458,I61866,I61455,I61897,I172849,I61914,I61931,I61948,I61470,I61979,I61467,I62010,I172846,I62027,I62044,I61473,I61482,I61452,I62136,I62153,I206293,I62170,I206305,I206287,I62187,I206302,I62110,I62218,I62235,I206290,I62125,I62107,I62280,I62297,I62314,I206299,I62331,I206278,I62348,I206281,I62365,I206284,I62382,I62399,I62416,I62122,I62447,I62464,I62481,I62104,I62512,I62101,I62543,I206275,I62560,I62577,I62594,I62116,I62625,I62113,I62656,I206296,I62673,I62690,I62119,I62128,I62098,I62782,I62799,I239474,I62816,I239462,I239468,I62833,I239459,I62756,I62864,I62881,I239465,I62771,I62753,I62926,I62943,I62960,I239477,I62977,I239489,I62994,I239471,I63011,I239486,I63028,I63045,I63062,I62768,I63093,I63110,I63127,I62750,I63158,I62747,I63189,I239480,I63206,I63223,I63240,I62762,I63271,I62759,I63302,I239483,I63319,I63336,I62765,I62774,I62744,I63428,I63445,I241786,I63462,I241774,I241780,I63479,I241771,I63402,I63510,I63527,I241777,I63417,I63399,I63572,I63589,I63606,I241789,I63623,I241801,I63640,I241783,I63657,I241798,I63674,I63691,I63708,I63414,I63739,I63756,I63773,I63396,I63804,I63393,I63835,I241792,I63852,I63869,I63886,I63408,I63917,I63405,I63948,I241795,I63965,I63982,I63411,I63420,I63390,I64074,I64091,I296929,I64108,I296905,I296911,I64125,I296914,I64048,I64156,I64173,I296923,I64063,I64045,I64218,I64235,I64252,I296902,I64269,I296917,I64286,I296908,I64303,I296920,I64320,I64337,I64354,I64060,I64385,I64402,I64419,I64042,I64450,I64039,I64481,I296932,I64498,I64515,I64532,I64054,I64563,I64051,I64594,I296926,I64611,I64628,I64057,I64066,I64036,I64720,I64737,I392026,I64754,I392023,I392020,I64771,I392041,I64694,I64802,I64819,I392044,I64709,I64691,I64864,I64881,I64898,I392017,I64915,I392029,I64932,I392038,I64949,I392032,I64966,I64983,I65000,I64706,I65031,I65048,I65065,I64688,I65096,I64685,I65127,I392047,I65144,I65161,I65178,I64700,I65209,I64697,I65240,I392035,I65257,I65274,I64703,I64712,I64682,I65366,I65383,I233391,I65400,I233373,I233388,I65417,I233397,I65340,I65448,I65465,I233400,I65355,I65337,I65510,I65527,I65544,I233403,I65561,I233379,I65578,I233382,I65595,I233376,I65612,I65629,I65646,I65352,I65677,I65694,I65711,I65334,I65742,I65331,I65773,I233385,I65790,I65807,I65824,I65346,I65855,I65343,I65886,I233394,I65903,I65920,I65349,I65358,I65328,I66012,I66029,I66046,I66063,I65986,I66094,I66111,I66001,I65983,I66156,I66173,I66190,I66207,I66224,I66241,I66258,I66275,I66292,I65998,I66323,I66340,I66357,I65980,I66388,I65977,I66419,I66436,I66453,I66470,I65992,I66501,I65989,I66532,I66549,I66566,I65995,I66004,I65974,I66658,I66675,I211461,I66692,I211473,I211455,I66709,I211470,I66632,I66740,I66757,I211458,I66647,I66629,I66802,I66819,I66836,I211467,I66853,I211446,I66870,I211449,I66887,I211452,I66904,I66921,I66938,I66644,I66969,I66986,I67003,I66626,I67034,I66623,I67065,I211443,I67082,I67099,I67116,I66638,I67147,I66635,I67178,I211464,I67195,I67212,I66641,I66650,I66620,I67304,I67321,I160240,I67338,I160237,I160225,I67355,I160228,I67278,I67386,I67403,I160234,I67293,I67275,I67448,I67465,I67482,I160246,I67499,I160222,I67516,I160243,I67533,I160231,I67550,I67567,I67584,I67290,I67615,I67632,I67649,I67272,I67680,I67269,I67711,I160252,I67728,I67745,I67762,I67284,I67793,I67281,I67824,I160249,I67841,I67858,I67287,I67296,I67266,I67950,I67967,I86715,I67984,I86703,I86709,I68001,I86718,I67924,I68032,I68049,I86706,I67939,I67921,I68094,I68111,I68128,I86727,I68145,I86700,I68162,I86721,I68179,I86712,I68196,I68213,I68230,I67936,I68261,I68278,I68295,I67918,I68326,I67915,I68357,I86697,I68374,I68391,I68408,I67930,I68439,I67927,I68470,I86724,I68487,I68504,I67933,I67942,I67912,I68596,I68613,I290979,I68630,I290955,I290961,I68647,I290964,I68570,I68678,I68695,I290973,I68585,I68567,I68740,I68757,I68774,I290952,I68791,I290967,I68808,I290958,I68825,I290970,I68842,I68859,I68876,I68582,I68907,I68924,I68941,I68564,I68972,I68561,I69003,I290982,I69020,I69037,I69054,I68576,I69085,I68573,I69116,I290976,I69133,I69150,I68579,I68588,I68558,I69242,I69259,I355246,I69276,I355261,I355276,I69293,I355264,I69216,I69324,I69341,I355267,I69231,I69213,I69386,I69403,I69420,I355273,I69437,I355270,I69454,I355249,I69471,I355258,I69488,I69505,I69522,I69228,I69553,I69570,I69587,I69210,I69618,I69207,I69649,I355255,I69666,I69683,I69700,I69222,I69731,I69219,I69762,I355252,I69779,I69796,I69225,I69234,I69204,I69888,I69905,I294549,I69922,I294525,I294531,I69939,I294534,I69862,I69970,I69987,I294543,I69877,I69859,I70032,I70049,I70066,I294522,I70083,I294537,I70100,I294528,I70117,I294540,I70134,I70151,I70168,I69874,I70199,I70216,I70233,I69856,I70264,I69853,I70295,I294552,I70312,I70329,I70346,I69868,I70377,I69865,I70408,I294546,I70425,I70442,I69871,I69880,I69850,I70534,I70551,I328452,I70568,I328437,I328464,I70585,I328440,I70508,I70616,I70633,I328455,I70523,I70505,I70678,I70695,I70712,I328467,I70729,I328449,I70746,I328458,I70763,I328443,I70780,I70797,I70814,I70520,I70845,I70862,I70879,I70502,I70910,I70499,I70941,I328446,I70958,I70975,I70992,I70514,I71023,I70511,I71054,I328461,I71071,I71088,I70517,I70526,I70496,I71180,I71197,I71214,I71231,I71154,I71262,I71279,I71169,I71151,I71324,I71341,I71358,I71375,I71392,I71409,I71426,I71443,I71460,I71166,I71491,I71508,I71525,I71148,I71556,I71145,I71587,I71604,I71621,I71638,I71160,I71669,I71157,I71700,I71717,I71734,I71163,I71172,I71142,I71826,I71843,I352730,I71860,I352745,I352760,I71877,I352748,I71908,I71925,I352751,I71970,I71987,I72004,I352757,I72021,I352754,I72038,I352733,I72055,I352742,I72072,I72089,I72106,I72137,I72154,I72171,I72202,I72233,I352739,I72250,I72267,I72284,I72315,I72346,I352736,I72363,I72380,I72472,I72489,I298714,I72506,I298690,I298696,I72523,I298699,I72446,I72554,I72571,I298708,I72461,I72443,I72616,I72633,I72650,I298687,I72667,I298702,I72684,I298693,I72701,I298705,I72718,I72735,I72752,I72458,I72783,I72800,I72817,I72440,I72848,I72437,I72879,I298717,I72896,I72913,I72930,I72452,I72961,I72449,I72992,I298711,I73009,I73026,I72455,I72464,I72434,I73118,I73135,I257392,I73152,I257380,I257386,I73169,I257377,I73092,I73200,I73217,I257383,I73107,I73089,I73262,I73279,I73296,I257395,I73313,I257407,I73330,I257389,I73347,I257404,I73364,I73381,I73398,I73104,I73429,I73446,I73463,I73086,I73494,I73083,I73525,I257398,I73542,I73559,I73576,I73098,I73607,I73095,I73638,I257401,I73655,I73672,I73101,I73110,I73080,I73764,I73781,I180793,I73798,I180790,I180778,I73815,I180781,I73738,I73846,I73863,I180787,I73753,I73735,I73908,I73925,I73942,I180799,I73959,I180775,I73976,I180796,I73993,I180784,I74010,I74027,I74044,I73750,I74075,I74092,I74109,I73732,I74140,I73729,I74171,I180805,I74188,I74205,I74222,I73744,I74253,I73741,I74284,I180802,I74301,I74318,I73747,I73756,I73726,I74410,I74427,I178804,I74444,I178801,I178789,I74461,I178792,I74384,I74492,I74509,I178798,I74399,I74381,I74554,I74571,I74588,I178810,I74605,I178786,I74622,I178807,I74639,I178795,I74656,I74673,I74690,I74396,I74721,I74738,I74755,I74378,I74786,I74375,I74817,I178816,I74834,I74851,I74868,I74390,I74899,I74387,I74930,I178813,I74947,I74964,I74393,I74402,I74372,I75056,I75073,I150958,I75090,I150955,I150943,I75107,I150946,I75030,I75138,I75155,I150952,I75045,I75027,I75200,I75217,I75234,I150964,I75251,I150940,I75268,I150961,I75285,I150949,I75302,I75319,I75336,I75042,I75367,I75384,I75401,I75024,I75432,I75021,I75463,I150970,I75480,I75497,I75514,I75036,I75545,I75033,I75576,I150967,I75593,I75610,I75039,I75048,I75018,I75702,I75719,I305259,I75736,I305235,I305241,I75753,I305244,I75676,I75784,I75801,I305253,I75691,I75673,I75846,I75863,I75880,I305232,I75897,I305247,I75914,I305238,I75931,I305250,I75948,I75965,I75982,I75688,I76013,I76030,I76047,I75670,I76078,I75667,I76109,I305262,I76126,I76143,I76160,I75682,I76191,I75679,I76222,I305256,I76239,I76256,I75685,I75694,I75664,I76348,I76365,I145654,I76382,I145651,I145639,I76399,I145642,I76322,I76430,I76447,I145648,I76337,I76319,I76492,I76509,I76526,I145660,I76543,I145636,I76560,I145657,I76577,I145645,I76594,I76611,I76628,I76334,I76659,I76676,I76693,I76316,I76724,I76313,I76755,I145666,I76772,I76789,I76806,I76328,I76837,I76325,I76868,I145663,I76885,I76902,I76331,I76340,I76310,I76994,I77011,I295739,I77028,I295715,I295721,I77045,I295724,I76968,I77076,I77093,I295733,I76983,I76965,I77138,I77155,I77172,I295712,I77189,I295727,I77206,I295718,I77223,I295730,I77240,I77257,I77274,I76980,I77305,I77322,I77339,I76962,I77370,I76959,I77401,I295742,I77418,I77435,I77452,I76974,I77483,I76971,I77514,I295736,I77531,I77548,I76977,I76986,I76956,I77640,I77657,I77674,I77691,I77614,I77722,I77739,I77629,I77611,I77784,I77801,I77818,I77835,I77852,I77869,I77886,I77903,I77920,I77626,I77951,I77968,I77985,I77608,I78016,I77605,I78047,I78064,I78081,I78098,I77620,I78129,I77617,I78160,I78177,I78194,I77623,I77632,I77602,I78286,I78303,I78320,I78337,I78368,I78385,I78430,I78447,I78464,I78481,I78498,I78515,I78532,I78549,I78566,I78597,I78614,I78631,I78662,I78693,I78710,I78727,I78744,I78775,I78806,I78823,I78840,I78932,I78949,I122210,I78966,I122240,I122219,I78983,I122231,I79014,I79031,I122213,I79076,I79093,I79110,I122216,I79127,I122234,I79144,I122225,I79161,I122222,I79178,I79195,I79212,I79243,I79260,I79277,I79308,I79339,I122228,I79356,I79373,I79390,I79421,I79452,I122237,I79469,I79486,I79578,I79595,I194665,I79612,I194677,I194659,I79629,I194674,I79552,I79660,I79677,I194662,I79567,I79549,I79722,I79739,I79756,I194671,I79773,I194650,I79790,I194653,I79807,I194656,I79824,I79841,I79858,I79564,I79889,I79906,I79923,I79546,I79954,I79543,I79985,I194647,I80002,I80019,I80036,I79558,I80067,I79555,I80098,I194668,I80115,I80132,I79561,I79570,I79540,I80224,I80241,I258548,I80258,I258536,I258542,I80275,I258533,I80198,I80306,I80323,I258539,I80213,I80195,I80368,I80385,I80402,I258551,I80419,I258563,I80436,I258545,I80453,I258560,I80470,I80487,I80504,I80210,I80535,I80552,I80569,I80192,I80600,I80189,I80631,I258554,I80648,I80665,I80682,I80204,I80713,I80201,I80744,I258557,I80761,I80778,I80207,I80216,I80186,I80870,I80887,I299309,I80904,I299285,I299291,I80921,I299294,I80844,I80952,I80969,I299303,I80859,I80841,I81014,I81031,I81048,I299282,I81065,I299297,I81082,I299288,I81099,I299300,I81116,I81133,I81150,I80856,I81181,I81198,I81215,I80838,I81246,I80835,I81277,I299312,I81294,I81311,I81328,I80850,I81359,I80847,I81390,I299306,I81407,I81424,I80853,I80862,I80832,I81516,I81533,I146317,I81550,I146314,I146302,I81567,I146305,I81490,I81598,I81615,I146311,I81505,I81487,I81660,I81677,I81694,I146323,I81711,I146299,I81728,I146320,I81745,I146308,I81762,I81779,I81796,I81502,I81827,I81844,I81861,I81484,I81892,I81481,I81923,I146329,I81940,I81957,I81974,I81496,I82005,I81493,I82036,I146326,I82053,I82070,I81499,I81508,I81478,I82162,I82179,I312994,I82196,I312970,I312976,I82213,I312979,I82136,I82244,I82261,I312988,I82151,I82133,I82306,I82323,I82340,I312967,I82357,I312982,I82374,I312973,I82391,I312985,I82408,I82425,I82442,I82148,I82473,I82490,I82507,I82130,I82538,I82127,I82569,I312997,I82586,I82603,I82620,I82142,I82651,I82139,I82682,I312991,I82699,I82716,I82145,I82154,I82124,I82808,I82825,I214691,I82842,I214703,I214685,I82859,I214700,I82782,I82890,I82907,I214688,I82797,I82779,I82952,I82969,I82986,I214697,I83003,I214676,I83020,I214679,I83037,I214682,I83054,I83071,I83088,I82794,I83119,I83136,I83153,I82776,I83184,I82773,I83215,I214673,I83232,I83249,I83266,I82788,I83297,I82785,I83328,I214694,I83345,I83362,I82791,I82800,I82770,I83454,I83471,I323097,I83488,I323082,I323109,I83505,I323085,I83428,I83536,I83553,I323100,I83443,I83425,I83598,I83615,I83632,I323112,I83649,I323094,I83666,I323103,I83683,I323088,I83700,I83717,I83734,I83440,I83765,I83782,I83799,I83422,I83830,I83419,I83861,I323091,I83878,I83895,I83912,I83434,I83943,I83431,I83974,I323106,I83991,I84008,I83437,I83446,I83416,I84100,I84117,I186760,I84134,I186757,I186745,I84151,I186748,I84074,I84182,I84199,I186754,I84089,I84071,I84244,I84261,I84278,I186766,I84295,I186742,I84312,I186763,I84329,I186751,I84346,I84363,I84380,I84086,I84411,I84428,I84445,I84068,I84476,I84065,I84507,I186772,I84524,I84541,I84558,I84080,I84589,I84077,I84620,I186769,I84637,I84654,I84083,I84092,I84062,I84746,I84763,I345823,I84780,I345829,I345841,I84797,I345832,I84717,I84828,I84845,I345811,I84862,I84879,I84896,I345826,I84913,I345814,I84930,I345835,I84947,I345817,I84964,I84981,I84732,I84729,I85026,I84714,I85057,I84711,I85088,I85105,I85122,I85139,I345838,I85156,I85173,I84738,I85204,I84726,I84720,I85249,I345820,I85266,I84735,I85297,I85314,I85331,I84723,I84708,I85409,I85426,I165526,I85443,I165535,I165547,I85460,I165538,I85380,I85491,I85508,I165550,I85525,I85542,I85559,I165556,I85576,I165532,I85593,I165541,I85610,I165529,I85627,I85644,I85395,I85392,I85689,I85377,I85720,I85374,I85751,I85768,I85785,I85802,I165553,I85819,I85836,I85401,I85867,I85389,I85383,I85912,I165544,I85929,I85398,I85960,I85977,I85994,I85386,I85371,I86072,I86089,I190720,I86106,I190729,I190741,I86123,I190732,I86043,I86154,I86171,I190744,I86188,I86205,I86222,I190750,I86239,I190726,I86256,I190735,I86273,I190723,I86290,I86307,I86058,I86055,I86352,I86040,I86383,I86037,I86414,I86431,I86448,I86465,I190747,I86482,I86499,I86064,I86530,I86052,I86046,I86575,I190738,I86592,I86061,I86623,I86640,I86657,I86049,I86034,I86735,I86752,I199187,I86769,I199196,I199169,I86786,I199181,I86817,I86834,I199193,I86851,I86868,I86885,I199172,I86902,I199178,I86919,I199190,I86936,I199175,I86953,I86970,I87015,I87046,I87077,I87094,I87111,I87128,I199199,I87145,I87162,I87193,I87238,I199184,I87255,I87286,I87303,I87320,I87398,I87415,I230195,I87432,I230204,I230177,I87449,I230189,I87369,I87480,I87497,I230201,I87514,I87531,I87548,I230180,I87565,I230186,I87582,I230198,I87599,I230183,I87616,I87633,I87384,I87381,I87678,I87366,I87709,I87363,I87740,I87757,I87774,I87791,I230207,I87808,I87825,I87390,I87856,I87378,I87372,I87901,I230192,I87918,I87387,I87949,I87966,I87983,I87375,I87360,I88061,I88078,I266047,I88095,I266053,I266050,I88112,I266068,I88032,I88143,I88160,I266077,I88177,I88194,I88211,I266071,I88228,I266062,I88245,I266065,I88262,I266056,I88279,I88296,I88047,I88044,I88341,I88029,I88372,I88026,I88403,I88420,I88437,I88454,I266074,I88471,I88488,I88053,I88519,I88041,I88035,I88564,I266059,I88581,I88050,I88612,I88629,I88646,I88038,I88023,I88724,I88741,I352113,I88758,I352119,I352131,I88775,I352122,I88695,I88806,I88823,I352101,I88840,I88857,I88874,I352116,I88891,I352104,I88908,I352125,I88925,I352107,I88942,I88959,I88710,I88707,I89004,I88692,I89035,I88689,I89066,I89083,I89100,I89117,I352128,I89134,I89151,I88716,I89182,I88704,I88698,I89227,I352110,I89244,I88713,I89275,I89292,I89309,I88701,I88686,I89387,I89404,I338275,I89421,I338281,I338293,I89438,I338284,I89469,I89486,I338263,I89503,I89520,I89537,I338278,I89554,I338266,I89571,I338287,I89588,I338269,I89605,I89622,I89667,I89698,I89729,I89746,I89763,I89780,I338290,I89797,I89814,I89845,I89890,I338272,I89907,I89938,I89955,I89972,I90050,I90067,I90084,I90101,I90021,I90132,I90149,I90166,I90183,I90200,I90217,I90234,I90251,I90268,I90285,I90036,I90033,I90330,I90018,I90361,I90015,I90392,I90409,I90426,I90443,I90460,I90477,I90042,I90508,I90030,I90024,I90553,I90570,I90039,I90601,I90618,I90635,I90027,I90012,I90713,I90730,I127589,I90747,I127571,I127565,I90764,I127568,I90684,I90795,I90812,I127577,I90829,I90846,I90863,I127586,I90880,I127574,I90897,I127580,I90914,I127595,I90931,I90948,I90699,I90696,I90993,I90681,I91024,I90678,I91055,I91072,I91089,I91106,I127583,I91123,I91140,I90705,I91171,I90693,I90687,I91216,I127592,I91233,I90702,I91264,I91281,I91298,I90690,I90675,I91376,I91393,I146962,I91410,I146971,I146983,I91427,I146974,I91347,I91458,I91475,I146986,I91492,I91509,I91526,I146992,I91543,I146968,I91560,I146977,I91577,I146965,I91594,I91611,I91362,I91359,I91656,I91344,I91687,I91341,I91718,I91735,I91752,I91769,I146989,I91786,I91803,I91368,I91834,I91356,I91350,I91879,I146980,I91896,I91365,I91927,I91944,I91961,I91353,I91338,I92039,I92056,I333243,I92073,I333249,I333261,I92090,I333252,I92010,I92121,I92138,I333231,I92155,I92172,I92189,I333246,I92206,I333234,I92223,I333255,I92240,I333237,I92257,I92274,I92025,I92022,I92319,I92007,I92350,I92004,I92381,I92398,I92415,I92432,I333258,I92449,I92466,I92031,I92497,I92019,I92013,I92542,I333240,I92559,I92028,I92590,I92607,I92624,I92016,I92001,I92702,I92719,I343936,I92736,I343942,I343954,I92753,I343945,I92673,I92784,I92801,I343924,I92818,I92835,I92852,I343939,I92869,I343927,I92886,I343948,I92903,I343930,I92920,I92937,I92688,I92685,I92982,I92670,I93013,I92667,I93044,I93061,I93078,I93095,I343951,I93112,I93129,I92694,I93160,I92682,I92676,I93205,I343933,I93222,I92691,I93253,I93270,I93287,I92679,I92664,I93365,I93382,I259111,I93399,I259117,I259114,I93416,I259132,I93447,I93464,I259141,I93481,I93498,I93515,I259135,I93532,I259126,I93549,I259129,I93566,I259120,I93583,I93600,I93645,I93676,I93707,I93724,I93741,I93758,I259138,I93775,I93792,I93823,I93868,I259123,I93885,I93916,I93933,I93950,I94028,I94045,I354629,I94062,I354635,I354647,I94079,I354638,I93999,I94110,I94127,I354617,I94144,I94161,I94178,I354632,I94195,I354620,I94212,I354641,I94229,I354623,I94246,I94263,I94014,I94011,I94308,I93996,I94339,I93993,I94370,I94387,I94404,I94421,I354644,I94438,I94455,I94020,I94486,I94008,I94002,I94531,I354626,I94548,I94017,I94579,I94596,I94613,I94005,I93990,I94691,I94708,I94725,I94742,I94662,I94773,I94790,I94807,I94824,I94841,I94858,I94875,I94892,I94909,I94926,I94677,I94674,I94971,I94659,I95002,I94656,I95033,I95050,I95067,I95084,I95101,I95118,I94683,I95149,I94671,I94665,I95194,I95211,I94680,I95242,I95259,I95276,I94668,I94653,I95354,I95371,I273255,I95388,I273267,I273270,I95405,I273276,I95325,I95436,I95453,I273279,I95470,I95487,I95504,I273258,I95521,I273273,I95538,I273282,I95555,I273285,I95572,I95589,I95340,I95337,I95634,I95322,I95665,I95319,I95696,I95713,I95730,I95747,I273261,I95764,I95781,I95346,I95812,I95334,I95328,I95857,I273264,I95874,I95343,I95905,I95922,I95939,I95331,I95316,I96017,I96034,I96051,I96068,I95988,I96099,I96116,I96133,I96150,I96167,I96184,I96201,I96218,I96235,I96252,I96003,I96000,I96297,I95985,I96328,I95982,I96359,I96376,I96393,I96410,I96427,I96444,I96009,I96475,I95997,I95991,I96520,I96537,I96006,I96568,I96585,I96602,I95994,I95979,I96680,I96697,I324278,I96714,I324293,I324275,I96731,I324287,I96651,I96762,I96779,I324284,I96796,I96813,I96830,I324302,I96847,I324272,I96864,I324281,I96881,I324299,I96898,I96915,I96666,I96663,I96960,I96648,I96991,I96645,I97022,I97039,I97056,I97073,I324290,I97090,I97107,I96672,I97138,I96660,I96654,I97183,I324296,I97200,I96669,I97231,I97248,I97265,I96657,I96642,I97343,I97360,I97377,I97394,I97314,I97425,I97442,I97459,I97476,I97493,I97510,I97527,I97544,I97561,I97578,I97329,I97326,I97623,I97311,I97654,I97308,I97685,I97702,I97719,I97736,I97753,I97770,I97335,I97801,I97323,I97317,I97846,I97863,I97332,I97894,I97911,I97928,I97320,I97305,I98006,I98023,I209523,I98040,I209532,I209505,I98057,I209517,I97977,I98088,I98105,I209529,I98122,I98139,I98156,I209508,I98173,I209514,I98190,I209526,I98207,I209511,I98224,I98241,I97992,I97989,I98286,I97974,I98317,I97971,I98348,I98365,I98382,I98399,I209535,I98416,I98433,I97998,I98464,I97986,I97980,I98509,I209520,I98526,I97995,I98557,I98574,I98591,I97983,I97968,I98669,I98686,I233997,I98703,I234015,I234003,I98720,I234009,I98640,I98751,I98768,I234012,I98785,I98802,I98819,I233991,I98836,I233985,I98853,I233994,I98870,I234006,I98887,I98904,I98655,I98652,I98949,I98637,I98980,I98634,I99011,I99028,I99045,I99062,I234000,I99079,I99096,I98661,I99127,I98649,I98643,I99172,I233988,I99189,I98658,I99220,I99237,I99254,I98646,I98631,I99332,I99349,I301082,I99366,I301094,I301097,I99383,I301085,I99414,I99431,I301070,I99448,I99465,I99482,I301073,I99499,I301076,I99516,I301079,I99533,I301088,I99550,I99567,I99612,I99643,I99674,I99691,I99708,I99725,I301091,I99742,I99759,I99790,I99835,I301067,I99852,I99883,I99900,I99917,I99995,I100012,I253909,I100029,I253915,I253912,I100046,I253930,I99966,I100077,I100094,I253939,I100111,I100128,I100145,I253933,I100162,I253924,I100179,I253927,I100196,I253918,I100213,I100230,I99981,I99978,I100275,I99963,I100306,I99960,I100337,I100354,I100371,I100388,I253936,I100405,I100422,I99987,I100453,I99975,I99969,I100498,I253921,I100515,I99984,I100546,I100563,I100580,I99972,I99957,I100658,I100675,I100692,I100709,I100629,I100740,I100757,I100774,I100791,I100808,I100825,I100842,I100859,I100876,I100893,I100644,I100641,I100938,I100626,I100969,I100623,I101000,I101017,I101034,I101051,I101068,I101085,I100650,I101116,I100638,I100632,I101161,I101178,I100647,I101209,I101226,I101243,I100635,I100620,I101321,I101338,I101355,I101372,I101292,I101403,I101420,I101437,I101454,I101471,I101488,I101505,I101522,I101539,I101556,I101307,I101304,I101601,I101289,I101632,I101286,I101663,I101680,I101697,I101714,I101731,I101748,I101313,I101779,I101301,I101295,I101824,I101841,I101310,I101872,I101889,I101906,I101298,I101283,I101984,I102001,I385105,I102018,I385084,I385096,I102035,I385090,I101955,I102066,I102083,I385111,I102100,I102117,I102134,I385087,I102151,I385099,I102168,I385102,I102185,I385108,I102202,I102219,I101970,I101967,I102264,I101952,I102295,I101949,I102326,I102343,I102360,I102377,I385081,I102394,I102411,I101976,I102442,I101964,I101958,I102487,I385093,I102504,I101973,I102535,I102552,I102569,I101961,I101946,I102647,I102664,I161548,I102681,I161557,I161569,I102698,I161560,I102618,I102729,I102746,I161572,I102763,I102780,I102797,I161578,I102814,I161554,I102831,I161563,I102848,I161551,I102865,I102882,I102633,I102630,I102927,I102615,I102958,I102612,I102989,I103006,I103023,I103040,I161575,I103057,I103074,I102639,I103105,I102627,I102621,I103150,I161566,I103167,I102636,I103198,I103215,I103232,I102624,I102609,I103310,I103327,I254487,I103344,I254493,I254490,I103361,I254508,I103392,I103409,I254517,I103426,I103443,I103460,I254511,I103477,I254502,I103494,I254505,I103511,I254496,I103528,I103545,I103590,I103621,I103652,I103669,I103686,I103703,I254514,I103720,I103737,I103768,I103813,I254499,I103830,I103861,I103878,I103895,I103973,I103990,I316543,I104007,I316558,I316540,I104024,I316552,I103944,I104055,I104072,I316549,I104089,I104106,I104123,I316567,I104140,I316537,I104157,I316546,I104174,I316564,I104191,I104208,I103959,I103956,I104253,I103941,I104284,I103938,I104315,I104332,I104349,I104366,I316555,I104383,I104400,I103965,I104431,I103953,I103947,I104476,I316561,I104493,I103962,I104524,I104541,I104558,I103950,I103935,I104636,I104653,I266631,I104670,I266637,I266628,I104687,I266646,I104607,I104718,I104735,I266625,I104752,I104769,I104786,I266655,I104803,I266634,I104820,I266643,I104837,I266649,I104854,I104871,I104622,I104619,I104916,I104604,I104947,I104601,I104978,I104995,I105012,I105029,I266640,I105046,I105063,I104628,I105094,I104616,I104610,I105139,I266652,I105156,I104625,I105187,I105204,I105221,I104613,I104598,I105299,I105316,I105333,I105350,I105270,I105381,I105398,I105415,I105432,I105449,I105466,I105483,I105500,I105517,I105534,I105285,I105282,I105579,I105267,I105610,I105264,I105641,I105658,I105675,I105692,I105709,I105726,I105291,I105757,I105279,I105273,I105802,I105819,I105288,I105850,I105867,I105884,I105276,I105261,I105962,I105979,I320708,I105996,I320723,I320705,I106013,I320717,I105933,I106044,I106061,I320714,I106078,I106095,I106112,I320732,I106129,I320702,I106146,I320711,I106163,I320729,I106180,I106197,I105948,I105945,I106242,I105930,I106273,I105927,I106304,I106321,I106338,I106355,I320720,I106372,I106389,I105954,I106420,I105942,I105936,I106465,I320726,I106482,I105951,I106513,I106530,I106547,I105939,I105924,I106625,I106642,I106659,I106676,I106596,I106707,I106724,I106741,I106758,I106775,I106792,I106809,I106826,I106843,I106860,I106611,I106608,I106905,I106593,I106936,I106590,I106967,I106984,I107001,I107018,I107035,I107052,I106617,I107083,I106605,I106599,I107128,I107145,I106614,I107176,I107193,I107210,I106602,I106587,I107288,I107305,I107322,I107339,I107259,I107370,I107387,I107404,I107421,I107438,I107455,I107472,I107489,I107506,I107523,I107274,I107271,I107568,I107256,I107599,I107253,I107630,I107647,I107664,I107681,I107698,I107715,I107280,I107746,I107268,I107262,I107791,I107808,I107277,I107839,I107856,I107873,I107265,I107250,I107951,I107968,I107985,I108002,I107922,I108033,I108050,I108067,I108084,I108101,I108118,I108135,I108152,I108169,I108186,I107937,I107934,I108231,I107919,I108262,I107916,I108293,I108310,I108327,I108344,I108361,I108378,I107943,I108409,I107931,I107925,I108454,I108471,I107940,I108502,I108519,I108536,I107928,I107913,I108614,I108631,I108648,I108665,I108585,I108696,I108713,I108730,I108747,I108764,I108781,I108798,I108815,I108832,I108849,I108600,I108597,I108894,I108582,I108925,I108579,I108956,I108973,I108990,I109007,I109024,I109041,I108606,I109072,I108594,I108588,I109117,I109134,I108603,I109165,I109182,I109199,I108591,I108576,I109277,I109294,I310007,I109311,I310019,I310022,I109328,I310010,I109248,I109359,I109376,I309995,I109393,I109410,I109427,I309998,I109444,I310001,I109461,I310004,I109478,I310013,I109495,I109512,I109263,I109260,I109557,I109245,I109588,I109242,I109619,I109636,I109653,I109670,I310016,I109687,I109704,I109269,I109735,I109257,I109251,I109780,I309992,I109797,I109266,I109828,I109845,I109862,I109254,I109239,I109940,I109957,I393197,I109974,I393176,I393188,I109991,I393182,I110022,I110039,I393203,I110056,I110073,I110090,I393179,I110107,I393191,I110124,I393194,I110141,I393200,I110158,I110175,I110220,I110251,I110282,I110299,I110316,I110333,I393173,I110350,I110367,I110398,I110443,I393185,I110460,I110491,I110508,I110525,I110603,I110620,I286207,I110637,I286219,I286222,I110654,I286210,I110574,I110685,I110702,I286195,I110719,I110736,I110753,I286198,I110770,I286201,I110787,I286204,I110804,I286213,I110821,I110838,I110589,I110586,I110883,I110571,I110914,I110568,I110945,I110962,I110979,I110996,I286216,I111013,I111030,I110595,I111061,I110583,I110577,I111106,I286192,I111123,I110592,I111154,I111171,I111188,I110580,I110565,I111266,I111283,I111300,I111317,I111237,I111348,I111365,I111382,I111399,I111416,I111433,I111450,I111467,I111484,I111501,I111252,I111249,I111546,I111234,I111577,I111231,I111608,I111625,I111642,I111659,I111676,I111693,I111258,I111724,I111246,I111240,I111769,I111786,I111255,I111817,I111834,I111851,I111243,I111228,I111929,I111946,I126994,I111963,I126976,I126970,I111980,I126973,I112011,I112028,I126982,I112045,I112062,I112079,I126991,I112096,I126979,I112113,I126985,I112130,I127000,I112147,I112164,I112209,I112240,I112271,I112288,I112305,I112322,I126988,I112339,I112356,I112387,I112432,I126997,I112449,I112480,I112497,I112514,I112592,I112609,I112626,I112643,I112563,I112674,I112691,I112708,I112725,I112742,I112759,I112776,I112793,I112810,I112827,I112578,I112575,I112872,I112560,I112903,I112557,I112934,I112951,I112968,I112985,I113002,I113019,I112584,I113050,I112572,I112566,I113095,I113112,I112581,I113143,I113160,I113177,I112569,I112554,I113255,I113272,I113289,I113306,I113337,I113354,I113371,I113388,I113405,I113422,I113439,I113456,I113473,I113490,I113535,I113566,I113597,I113614,I113631,I113648,I113665,I113682,I113713,I113758,I113775,I113806,I113823,I113840,I113918,I113935,I217275,I217272,I113952,I217257,I113892,I113983,I217266,I217269,I114000,I114017,I114034,I217281,I114051,I114068,I217287,I217263,I114085,I114102,I114119,I113886,I114150,I114167,I113883,I114198,I217278,I114215,I217284,I114232,I113895,I113880,I114277,I217260,I114294,I114311,I114328,I114345,I113901,I114376,I113910,I114407,I113904,I113907,I113898,I113889,I114513,I114530,I114547,I114487,I114578,I114595,I114612,I114629,I114646,I114663,I114680,I114697,I114714,I114481,I114745,I114762,I114478,I114793,I114810,I114827,I114490,I114475,I114872,I114889,I114906,I114923,I114940,I114496,I114971,I114505,I115002,I114499,I114502,I114493,I114484,I115108,I115125,I115142,I115082,I115173,I115190,I115207,I115224,I115241,I115258,I115275,I115292,I115309,I115076,I115340,I115357,I115073,I115388,I115405,I115422,I115085,I115070,I115467,I115484,I115501,I115518,I115535,I115091,I115566,I115100,I115597,I115094,I115097,I115088,I115079,I115703,I115720,I143647,I143662,I115737,I143650,I115677,I115768,I143653,I143668,I115785,I115802,I115819,I143656,I115836,I115853,I143659,I143677,I115870,I115887,I115904,I115671,I115935,I115952,I115668,I115983,I143674,I116000,I143665,I116017,I115680,I115665,I116062,I143671,I116079,I116096,I116113,I116130,I115686,I116161,I115695,I116192,I115689,I115692,I115683,I115674,I116298,I116315,I253361,I253346,I116332,I253358,I116363,I253340,I253331,I116380,I116397,I116414,I253355,I116431,I116448,I253334,I253352,I116465,I116482,I116499,I116530,I116547,I116578,I253343,I116595,I253337,I116612,I116657,I253349,I116674,I116691,I116708,I116725,I116756,I116787,I116893,I116910,I116927,I116867,I116958,I116975,I116992,I117009,I117026,I117043,I117060,I117077,I117094,I116861,I117125,I117142,I116858,I117173,I117190,I117207,I116870,I116855,I117252,I117269,I117286,I117303,I117320,I116876,I117351,I116885,I117382,I116879,I116882,I116873,I116864,I117488,I117505,I117522,I117462,I117553,I117570,I117587,I117604,I117621,I117638,I117655,I117672,I117689,I117456,I117720,I117737,I117453,I117768,I117785,I117802,I117465,I117450,I117847,I117864,I117881,I117898,I117915,I117471,I117946,I117480,I117977,I117474,I117477,I117468,I117459,I118083,I118100,I315359,I315353,I118117,I315347,I118057,I118148,I315350,I315356,I118165,I118182,I118199,I315374,I118216,I118233,I315377,I315368,I118250,I118267,I118284,I118051,I118315,I118332,I118048,I118363,I315365,I118380,I315362,I118397,I118060,I118045,I118442,I315371,I118459,I118476,I118493,I118510,I118066,I118541,I118075,I118572,I118069,I118072,I118063,I118054,I118678,I118695,I222443,I222440,I118712,I222425,I118652,I118743,I222434,I222437,I118760,I118777,I118794,I222449,I118811,I118828,I222455,I222431,I118845,I118862,I118879,I118646,I118910,I118927,I118643,I118958,I222446,I118975,I222452,I118992,I118655,I118640,I119037,I222428,I119054,I119071,I119088,I119105,I118661,I119136,I118670,I119167,I118664,I118667,I118658,I118649,I119273,I119290,I119307,I119338,I119355,I119372,I119389,I119406,I119423,I119440,I119457,I119474,I119505,I119522,I119553,I119570,I119587,I119632,I119649,I119666,I119683,I119700,I119731,I119762,I119868,I119885,I119902,I119842,I119933,I119950,I119967,I119984,I120001,I120018,I120035,I120052,I120069,I119836,I120100,I120117,I119833,I120148,I120165,I120182,I119845,I119830,I120227,I120244,I120261,I120278,I120295,I119851,I120326,I119860,I120357,I119854,I119857,I119848,I119839,I120463,I120480,I152266,I152281,I120497,I152269,I120437,I120528,I152272,I152287,I120545,I120562,I120579,I152275,I120596,I120613,I152278,I152296,I120630,I120647,I120664,I120431,I120695,I120712,I120428,I120743,I152293,I120760,I152284,I120777,I120440,I120425,I120822,I152290,I120839,I120856,I120873,I120890,I120446,I120921,I120455,I120952,I120449,I120452,I120443,I120434,I121058,I121075,I347701,I347698,I121092,I347728,I121032,I121123,I347707,I347713,I121140,I121157,I121174,I347704,I121191,I121208,I347716,I347725,I121225,I121242,I121259,I121026,I121290,I121307,I121023,I121338,I347719,I121355,I347710,I121372,I121035,I121020,I121417,I347722,I121434,I121451,I121468,I121485,I121041,I121516,I121050,I121547,I121044,I121047,I121038,I121029,I121653,I121670,I327854,I327848,I121687,I327842,I121627,I121718,I327845,I327851,I121735,I121752,I121769,I327869,I121786,I121803,I327872,I327863,I121820,I121837,I121854,I121621,I121885,I121902,I121618,I121933,I327860,I121950,I327857,I121967,I121630,I121615,I122012,I327866,I122029,I122046,I122063,I122080,I121636,I122111,I121645,I122142,I121639,I121642,I121633,I121624,I122248,I122265,I122282,I122313,I122330,I122347,I122364,I122381,I122398,I122415,I122432,I122449,I122480,I122497,I122528,I122545,I122562,I122607,I122624,I122641,I122658,I122675,I122706,I122737,I122843,I122860,I225027,I225024,I122877,I225009,I122817,I122908,I225018,I225021,I122925,I122942,I122959,I225033,I122976,I122993,I225039,I225015,I123010,I123027,I123044,I122811,I123075,I123092,I122808,I123123,I225030,I123140,I225036,I123157,I122820,I122805,I123202,I225012,I123219,I123236,I123253,I123270,I122826,I123301,I122835,I123332,I122829,I122832,I122823,I122814,I123438,I123455,I123472,I123503,I123520,I123537,I123554,I123571,I123588,I123605,I123622,I123639,I123670,I123687,I123718,I123735,I123752,I123797,I123814,I123831,I123848,I123865,I123896,I123927,I124033,I124050,I124067,I124007,I124098,I124115,I124132,I124149,I124166,I124183,I124200,I124217,I124234,I124001,I124265,I124282,I123998,I124313,I124330,I124347,I124010,I123995,I124392,I124409,I124426,I124443,I124460,I124016,I124491,I124025,I124522,I124019,I124022,I124013,I124004,I124628,I124645,I124662,I124602,I124693,I124710,I124727,I124744,I124761,I124778,I124795,I124812,I124829,I124596,I124860,I124877,I124593,I124908,I124925,I124942,I124605,I124590,I124987,I125004,I125021,I125038,I125055,I124611,I125086,I124620,I125117,I124614,I124617,I124608,I124599,I125223,I125240,I380409,I380406,I125257,I380436,I125197,I125288,I380415,I380421,I125305,I125322,I125339,I380412,I125356,I125373,I380424,I380433,I125390,I125407,I125424,I125191,I125455,I125472,I125188,I125503,I380427,I125520,I380418,I125537,I125200,I125185,I125582,I380430,I125599,I125616,I125633,I125650,I125206,I125681,I125215,I125712,I125209,I125212,I125203,I125194,I125818,I125835,I166852,I166867,I125852,I166855,I125883,I166858,I166873,I125900,I125917,I125934,I166861,I125951,I125968,I166864,I166882,I125985,I126002,I126019,I126050,I126067,I126098,I166879,I126115,I166870,I126132,I126177,I166876,I126194,I126211,I126228,I126245,I126276,I126307,I126413,I126430,I377893,I377890,I126447,I377920,I126387,I126478,I377899,I377905,I126495,I126512,I126529,I377896,I126546,I126563,I377908,I377917,I126580,I126597,I126614,I126381,I126645,I126662,I126378,I126693,I377911,I126710,I377902,I126727,I126390,I126375,I126772,I377914,I126789,I126806,I126823,I126840,I126396,I126871,I126405,I126902,I126399,I126402,I126393,I126384,I127008,I127025,I368458,I368455,I127042,I368485,I127073,I368464,I368470,I127090,I127107,I127124,I368461,I127141,I127158,I368473,I368482,I127175,I127192,I127209,I127240,I127257,I127288,I368476,I127305,I368467,I127322,I127367,I368479,I127384,I127401,I127418,I127435,I127466,I127497,I127603,I127620,I177460,I177475,I127637,I177463,I127668,I177466,I177481,I127685,I127702,I127719,I177469,I127736,I127753,I177472,I177490,I127770,I127787,I127804,I127835,I127852,I127883,I177487,I127900,I177478,I127917,I127962,I177484,I127979,I127996,I128013,I128030,I128061,I128092,I128198,I128215,I301677,I301662,I128232,I301683,I128172,I128263,I301689,I301671,I128280,I128297,I128314,I301668,I128331,I128348,I301665,I301674,I128365,I128382,I128399,I128166,I128430,I128447,I128163,I128478,I301692,I128495,I301680,I128512,I128175,I128160,I128557,I301686,I128574,I128591,I128608,I128625,I128181,I128656,I128190,I128687,I128184,I128187,I128178,I128169,I128793,I128810,I314169,I314163,I128827,I314157,I128858,I314160,I314166,I128875,I128892,I128909,I314184,I128926,I128943,I314187,I314178,I128960,I128977,I128994,I129025,I129042,I129073,I314175,I129090,I314172,I129107,I129152,I314181,I129169,I129186,I129203,I129220,I129251,I129282,I129388,I129405,I269706,I269715,I129422,I269709,I129362,I129453,I269694,I269685,I129470,I129487,I129504,I269712,I129521,I129538,I269688,I269697,I129555,I129572,I129589,I129356,I129620,I129637,I129353,I129668,I269691,I129685,I269703,I129702,I129365,I129350,I129747,I269700,I129764,I129781,I129798,I129815,I129371,I129846,I129380,I129877,I129374,I129377,I129368,I129359,I129983,I130000,I170845,I170833,I129966,I129945,I130045,I170830,I130062,I170860,I170851,I130079,I130096,I130113,I170839,I130130,I130147,I130164,I170842,I170836,I130181,I129972,I130212,I130229,I130246,I130263,I129975,I130294,I170857,I130311,I170854,I130328,I130345,I130362,I129960,I130393,I130410,I129963,I129957,I129951,I130469,I170848,I129969,I130500,I129954,I129948,I130578,I130595,I130561,I130540,I130640,I130657,I130674,I130691,I130708,I130725,I130742,I130759,I130776,I130567,I130807,I130824,I130841,I130858,I130570,I130889,I130906,I130923,I130940,I130957,I130555,I130988,I131005,I130558,I130552,I130546,I131064,I130564,I131095,I130549,I130543,I131173,I131190,I131156,I131135,I131235,I131252,I131269,I131286,I131303,I131320,I131337,I131354,I131371,I131162,I131402,I131419,I131436,I131453,I131165,I131484,I131501,I131518,I131535,I131552,I131150,I131583,I131600,I131153,I131147,I131141,I131659,I131159,I131690,I131144,I131138,I131768,I131785,I183442,I183430,I131751,I131730,I131830,I183427,I131847,I183457,I183448,I131864,I131881,I131898,I183436,I131915,I131932,I131949,I183439,I183433,I131966,I131757,I131997,I132014,I132031,I132048,I131760,I132079,I183454,I132096,I183451,I132113,I132130,I132147,I131745,I132178,I132195,I131748,I131742,I131736,I132254,I183445,I131754,I132285,I131739,I131733,I132363,I132380,I132346,I132325,I132425,I132442,I132459,I132476,I132493,I132510,I132527,I132544,I132561,I132352,I132592,I132609,I132626,I132643,I132355,I132674,I132691,I132708,I132725,I132742,I132340,I132773,I132790,I132343,I132337,I132331,I132849,I132349,I132880,I132334,I132328,I132958,I132975,I245817,I245847,I132941,I132920,I133020,I245826,I133037,I245832,I245829,I133054,I133071,I133088,I245838,I133105,I133122,I133139,I245823,I245841,I133156,I132947,I133187,I133204,I133221,I133238,I132950,I133269,I245844,I133286,I245835,I133303,I133320,I133337,I132935,I133368,I133385,I132938,I132932,I132926,I133444,I245820,I132944,I133475,I132929,I132923,I133553,I133570,I133536,I133515,I133615,I133632,I133649,I133666,I133683,I133700,I133717,I133734,I133751,I133542,I133782,I133799,I133816,I133833,I133545,I133864,I133881,I133898,I133915,I133932,I133530,I133963,I133980,I133533,I133527,I133521,I134039,I133539,I134070,I133524,I133518,I134148,I134165,I152944,I152932,I134131,I134110,I134210,I152929,I134227,I152959,I152950,I134244,I134261,I134278,I152938,I134295,I134312,I134329,I152941,I152935,I134346,I134137,I134377,I134394,I134411,I134428,I134140,I134459,I152956,I134476,I152953,I134493,I134510,I134527,I134125,I134558,I134575,I134128,I134122,I134116,I134634,I152947,I134134,I134665,I134119,I134113,I134743,I134760,I348333,I348342,I134726,I134705,I134805,I348351,I134822,I348345,I348339,I134839,I134856,I134873,I348348,I134890,I134907,I134924,I348336,I348354,I134941,I134732,I134972,I134989,I135006,I135023,I134735,I135054,I348357,I135071,I348330,I135088,I135105,I135122,I134720,I135153,I135170,I134723,I134717,I134711,I135229,I348327,I134729,I135260,I134714,I134708,I135338,I135355,I135400,I135417,I135434,I135451,I135468,I135485,I135502,I135519,I135536,I135567,I135584,I135601,I135618,I135649,I135666,I135683,I135700,I135717,I135748,I135765,I135824,I135855,I135933,I135950,I135916,I135895,I135995,I136012,I136029,I136046,I136063,I136080,I136097,I136114,I136131,I135922,I136162,I136179,I136196,I136213,I135925,I136244,I136261,I136278,I136295,I136312,I135910,I136343,I136360,I135913,I135907,I135901,I136419,I135919,I136450,I135904,I135898,I136528,I136545,I136511,I136490,I136590,I136607,I136624,I136641,I136658,I136675,I136692,I136709,I136726,I136517,I136757,I136774,I136791,I136808,I136520,I136839,I136856,I136873,I136890,I136907,I136505,I136938,I136955,I136508,I136502,I136496,I137014,I136514,I137045,I136499,I136493,I137123,I137140,I137106,I137085,I137185,I137202,I137219,I137236,I137253,I137270,I137287,I137304,I137321,I137112,I137352,I137369,I137386,I137403,I137115,I137434,I137451,I137468,I137485,I137502,I137100,I137533,I137550,I137103,I137097,I137091,I137609,I137109,I137640,I137094,I137088,I137718,I137735,I317150,I137752,I317147,I317138,I137769,I317141,I137786,I137803,I317135,I137820,I137837,I137707,I137868,I137692,I137899,I317156,I137916,I317159,I137933,I317144,I137950,I317132,I137967,I137984,I138001,I137689,I138032,I138049,I137686,I138080,I317153,I138097,I137704,I138128,I137701,I138159,I138176,I137680,I137683,I138221,I317162,I138238,I138255,I138272,I137710,I138303,I137695,I137698,I138381,I138398,I138415,I138432,I138449,I138466,I138483,I138500,I138370,I138531,I138355,I138562,I138579,I138596,I138613,I138630,I138647,I138664,I138352,I138695,I138712,I138349,I138743,I138760,I138367,I138791,I138364,I138822,I138839,I138343,I138346,I138884,I138901,I138918,I138935,I138373,I138966,I138358,I138361,I139044,I139061,I332608,I139078,I332626,I332617,I139095,I332623,I139112,I139129,I332629,I139146,I139163,I139194,I139225,I332605,I139242,I332620,I139259,I332602,I139276,I332611,I139293,I139310,I139327,I139358,I139375,I139406,I332614,I139423,I139454,I139485,I139502,I139547,I332632,I139564,I139581,I139598,I139629,I139707,I139724,I208871,I139741,I208868,I208886,I139758,I208889,I139775,I139792,I208874,I139809,I139826,I139696,I139857,I139681,I139888,I208883,I139905,I208865,I139922,I208859,I139939,I208877,I139956,I139973,I139990,I139678,I140021,I140038,I139675,I140069,I208862,I140086,I139693,I140117,I139690,I140148,I140165,I139669,I139672,I140210,I208880,I140227,I140244,I140261,I139699,I140292,I139684,I139687,I140370,I140387,I313580,I140404,I313577,I313568,I140421,I313571,I140438,I140455,I313565,I140472,I140489,I140359,I140520,I140344,I140551,I313586,I140568,I313589,I140585,I313574,I140602,I313562,I140619,I140636,I140653,I140341,I140684,I140701,I140338,I140732,I313583,I140749,I140356,I140780,I140353,I140811,I140828,I140332,I140335,I140873,I313592,I140890,I140907,I140924,I140362,I140955,I140347,I140350,I141033,I141050,I274992,I141067,I275013,I275019,I141084,I275007,I141101,I141118,I274989,I141135,I141152,I141022,I141183,I141007,I141214,I274995,I141231,I275016,I141248,I275004,I141265,I275010,I141282,I141299,I141316,I141004,I141347,I141364,I141001,I141395,I275001,I141412,I141019,I141443,I141016,I141474,I141491,I140995,I140998,I141536,I274998,I141553,I141570,I141587,I141025,I141618,I141010,I141013,I141696,I141713,I141730,I141747,I141764,I141781,I141798,I141815,I141685,I141846,I141670,I141877,I141894,I141911,I141928,I141945,I141962,I141979,I141667,I142010,I142027,I141664,I142058,I142075,I141682,I142106,I141679,I142137,I142154,I141658,I141661,I142199,I142216,I142233,I142250,I141688,I142281,I141673,I141676,I142359,I142376,I357768,I142393,I357786,I357777,I142410,I357783,I142427,I142444,I357789,I142461,I142478,I142348,I142509,I142333,I142540,I357765,I142557,I357780,I142574,I357762,I142591,I357771,I142608,I142625,I142642,I142330,I142673,I142690,I142327,I142721,I357774,I142738,I142345,I142769,I142342,I142800,I142817,I142321,I142324,I142862,I357792,I142879,I142896,I142913,I142351,I142944,I142336,I142339,I143022,I143039,I143056,I143073,I143090,I143107,I143124,I143141,I143011,I143172,I142996,I143203,I143220,I143237,I143254,I143271,I143288,I143305,I142993,I143336,I143353,I142990,I143384,I143401,I143008,I143432,I143005,I143463,I143480,I142984,I142987,I143525,I143542,I143559,I143576,I143014,I143607,I142999,I143002,I143685,I143702,I201119,I143719,I201116,I201134,I143736,I201137,I143753,I143770,I201122,I143787,I143804,I143835,I143866,I201131,I143883,I201113,I143900,I201107,I143917,I201125,I143934,I143951,I143968,I143999,I144016,I144047,I201110,I144064,I144095,I144126,I144143,I144188,I201128,I144205,I144222,I144239,I144270,I144348,I144365,I262594,I144382,I262606,I262588,I144399,I262609,I144416,I144433,I262600,I144450,I144467,I144498,I144529,I262591,I144546,I262585,I144563,I262597,I144580,I262582,I144597,I144614,I144631,I144662,I144679,I144710,I262579,I144727,I144758,I144789,I144806,I144851,I262603,I144868,I144885,I144902,I144933,I145011,I145028,I145045,I145062,I145079,I145096,I145113,I145130,I145161,I145192,I145209,I145226,I145243,I145260,I145277,I145294,I145325,I145342,I145373,I145390,I145421,I145452,I145469,I145514,I145531,I145548,I145565,I145596,I145674,I145691,I382781,I145708,I382772,I382778,I145725,I382790,I145742,I145759,I382775,I145776,I145793,I145824,I145855,I382799,I145872,I382793,I145889,I382784,I145906,I382769,I145923,I145940,I145957,I145988,I146005,I146036,I382787,I146053,I146084,I146115,I146132,I146177,I382796,I146194,I146211,I146228,I146259,I146337,I146354,I199827,I146371,I199824,I199842,I146388,I199845,I146405,I146422,I199830,I146439,I146456,I146487,I146518,I199839,I146535,I199821,I146552,I199815,I146569,I199833,I146586,I146603,I146620,I146651,I146668,I146699,I199818,I146716,I146747,I146778,I146795,I146840,I199836,I146857,I146874,I146891,I146922,I147000,I147017,I147034,I147051,I147068,I147085,I147102,I147119,I147150,I147181,I147198,I147215,I147232,I147249,I147266,I147283,I147314,I147331,I147362,I147379,I147410,I147441,I147458,I147503,I147520,I147537,I147554,I147585,I147663,I147680,I147697,I147714,I147731,I147748,I147765,I147782,I147652,I147813,I147637,I147844,I147861,I147878,I147895,I147912,I147929,I147946,I147634,I147977,I147994,I147631,I148025,I148042,I147649,I148073,I147646,I148104,I148121,I147625,I147628,I148166,I148183,I148200,I148217,I147655,I148248,I147640,I147643,I148326,I148343,I379154,I148360,I379172,I379163,I148377,I379169,I148394,I148411,I379175,I148428,I148445,I148315,I148476,I148300,I148507,I379151,I148524,I379166,I148541,I379148,I148558,I379157,I148575,I148592,I148609,I148297,I148640,I148657,I148294,I148688,I379160,I148705,I148312,I148736,I148309,I148767,I148784,I148288,I148291,I148829,I379178,I148846,I148863,I148880,I148318,I148911,I148303,I148306,I148989,I149006,I149023,I149040,I149057,I149074,I149091,I149108,I148978,I149139,I148963,I149170,I149187,I149204,I149221,I149238,I149255,I149272,I148960,I149303,I149320,I148957,I149351,I149368,I148975,I149399,I148972,I149430,I149447,I148951,I148954,I149492,I149509,I149526,I149543,I148981,I149574,I148966,I148969,I149652,I149669,I305845,I149686,I305854,I305836,I149703,I305857,I149720,I149737,I305848,I149754,I149771,I149802,I149833,I305842,I149850,I305833,I149867,I305830,I149884,I305827,I149901,I149918,I149935,I149966,I149983,I150014,I305851,I150031,I150062,I150093,I150110,I150155,I305839,I150172,I150189,I150206,I150237,I150315,I150332,I150349,I150366,I150383,I150400,I150417,I150434,I150304,I150465,I150289,I150496,I150513,I150530,I150547,I150564,I150581,I150598,I150286,I150629,I150646,I150283,I150677,I150694,I150301,I150725,I150298,I150756,I150773,I150277,I150280,I150818,I150835,I150852,I150869,I150307,I150900,I150292,I150295,I150978,I150995,I151012,I151029,I151046,I151063,I151080,I151097,I151128,I151159,I151176,I151193,I151210,I151227,I151244,I151261,I151292,I151309,I151340,I151357,I151388,I151419,I151436,I151481,I151498,I151515,I151532,I151563,I151641,I151658,I151675,I151692,I151709,I151726,I151743,I151760,I151630,I151791,I151615,I151822,I151839,I151856,I151873,I151890,I151907,I151924,I151612,I151955,I151972,I151609,I152003,I152020,I151627,I152051,I151624,I152082,I152099,I151603,I151606,I152144,I152161,I152178,I152195,I151633,I152226,I151618,I151621,I152304,I152321,I201765,I152338,I201762,I201780,I152355,I201783,I152372,I152389,I201768,I152406,I152423,I152454,I152485,I201777,I152502,I201759,I152519,I201753,I152536,I201771,I152553,I152570,I152587,I152618,I152635,I152666,I201756,I152683,I152714,I152745,I152762,I152807,I201774,I152824,I152841,I152858,I152889,I152967,I152984,I302275,I153001,I302284,I302266,I153018,I302287,I153035,I153052,I302278,I153069,I153086,I153117,I153148,I302272,I153165,I302263,I153182,I302260,I153199,I302257,I153216,I153233,I153250,I153281,I153298,I153329,I302281,I153346,I153377,I153408,I153425,I153470,I302269,I153487,I153504,I153521,I153552,I153630,I153647,I273836,I153664,I273857,I273863,I153681,I273851,I153698,I153715,I273833,I153732,I153749,I153619,I153780,I153604,I153811,I273839,I153828,I273860,I153845,I273848,I153862,I273854,I153879,I153896,I153913,I153601,I153944,I153961,I153598,I153992,I273845,I154009,I153616,I154040,I153613,I154071,I154088,I153592,I153595,I154133,I273842,I154150,I154167,I154184,I153622,I154215,I153607,I153610,I154293,I154310,I154327,I154344,I154361,I154378,I154395,I154412,I154282,I154443,I154267,I154474,I154491,I154508,I154525,I154542,I154559,I154576,I154264,I154607,I154624,I154261,I154655,I154672,I154279,I154703,I154276,I154734,I154751,I154255,I154258,I154796,I154813,I154830,I154847,I154285,I154878,I154270,I154273,I154956,I154973,I279665,I154990,I279674,I279656,I155007,I279677,I155024,I155041,I279668,I155058,I155075,I155106,I155137,I279662,I155154,I279653,I155171,I279650,I155188,I279647,I155205,I155222,I155239,I155270,I155287,I155318,I279671,I155335,I155366,I155397,I155414,I155459,I279659,I155476,I155493,I155510,I155541,I155619,I155636,I204349,I155653,I204346,I204364,I155670,I204367,I155687,I155704,I204352,I155721,I155738,I155608,I155769,I155593,I155800,I204361,I155817,I204343,I155834,I204337,I155851,I204355,I155868,I155885,I155902,I155590,I155933,I155950,I155587,I155981,I204340,I155998,I155605,I156029,I155602,I156060,I156077,I155581,I155584,I156122,I204358,I156139,I156156,I156173,I155611,I156204,I155596,I155599,I156282,I156299,I377267,I156316,I377285,I377276,I156333,I377282,I156350,I156367,I377288,I156384,I156401,I156271,I156432,I156256,I156463,I377264,I156480,I377279,I156497,I377261,I156514,I377270,I156531,I156548,I156565,I156253,I156596,I156613,I156250,I156644,I377273,I156661,I156268,I156692,I156265,I156723,I156740,I156244,I156247,I156785,I377291,I156802,I156819,I156836,I156274,I156867,I156259,I156262,I156945,I156962,I156979,I156996,I157013,I157030,I157047,I157064,I157095,I157126,I157143,I157160,I157177,I157194,I157211,I157228,I157259,I157276,I157307,I157324,I157355,I157386,I157403,I157448,I157465,I157482,I157499,I157530,I157608,I157625,I157642,I157659,I157676,I157693,I157710,I157727,I157758,I157789,I157806,I157823,I157840,I157857,I157874,I157891,I157922,I157939,I157970,I157987,I158018,I158049,I158066,I158111,I158128,I158145,I158162,I158193,I158271,I158288,I158305,I158322,I158339,I158356,I158373,I158390,I158260,I158421,I158245,I158452,I158469,I158486,I158503,I158520,I158537,I158554,I158242,I158585,I158602,I158239,I158633,I158650,I158257,I158681,I158254,I158712,I158729,I158233,I158236,I158774,I158791,I158808,I158825,I158263,I158856,I158248,I158251,I158934,I158951,I277882,I158968,I277903,I277909,I158985,I277897,I159002,I159019,I277879,I159036,I159053,I158923,I159084,I158908,I159115,I277885,I159132,I277906,I159149,I277894,I159166,I277900,I159183,I159200,I159217,I158905,I159248,I159265,I158902,I159296,I277891,I159313,I158920,I159344,I158917,I159375,I159392,I158896,I158899,I159437,I277888,I159454,I159471,I159488,I158926,I159519,I158911,I158914,I159597,I159614,I272680,I159631,I272701,I272707,I159648,I272695,I159665,I159682,I272677,I159699,I159716,I159586,I159747,I159571,I159778,I272683,I159795,I272704,I159812,I272692,I159829,I272698,I159846,I159863,I159880,I159568,I159911,I159928,I159565,I159959,I272689,I159976,I159583,I160007,I159580,I160038,I160055,I159559,I159562,I160100,I272686,I160117,I160134,I160151,I159589,I160182,I159574,I159577,I160260,I160277,I330240,I160294,I330237,I330228,I160311,I330231,I160328,I160345,I330225,I160362,I160379,I160410,I160441,I330246,I160458,I330249,I160475,I330234,I160492,I330222,I160509,I160526,I160543,I160574,I160591,I160622,I330243,I160639,I160670,I160701,I160718,I160763,I330252,I160780,I160797,I160814,I160845,I160923,I160940,I160957,I160974,I160991,I161008,I161025,I161042,I160912,I161073,I160897,I161104,I161121,I161138,I161155,I161172,I161189,I161206,I160894,I161237,I161254,I160891,I161285,I161302,I160909,I161333,I160906,I161364,I161381,I160885,I160888,I161426,I161443,I161460,I161477,I160915,I161508,I160900,I160903,I161586,I161603,I161620,I161637,I161654,I161671,I161688,I161705,I161736,I161767,I161784,I161801,I161818,I161835,I161852,I161869,I161900,I161917,I161948,I161965,I161996,I162027,I162044,I162089,I162106,I162123,I162140,I162171,I162249,I162266,I392607,I162283,I392598,I392604,I162300,I392616,I162317,I162334,I392601,I162351,I162368,I162238,I162399,I162223,I162430,I392625,I162447,I392619,I162464,I392610,I162481,I392595,I162498,I162515,I162532,I162220,I162563,I162580,I162217,I162611,I392613,I162628,I162235,I162659,I162232,I162690,I162707,I162211,I162214,I162752,I392622,I162769,I162786,I162803,I162241,I162834,I162226,I162229,I162912,I162929,I162946,I162963,I162980,I162997,I163014,I163031,I162901,I163062,I162886,I163093,I163110,I163127,I163144,I163161,I163178,I163195,I162883,I163226,I163243,I162880,I163274,I163291,I162898,I163322,I162895,I163353,I163370,I162874,I162877,I163415,I163432,I163449,I163466,I162904,I163497,I162889,I162892,I163575,I163592,I163609,I163626,I163643,I163660,I163677,I163694,I163725,I163756,I163773,I163790,I163807,I163824,I163841,I163858,I163889,I163906,I163937,I163954,I163985,I164016,I164033,I164078,I164095,I164112,I164129,I164160,I164238,I164255,I164272,I164289,I164306,I164323,I164340,I164357,I164227,I164388,I164212,I164419,I164436,I164453,I164470,I164487,I164504,I164521,I164209,I164552,I164569,I164206,I164600,I164617,I164224,I164648,I164221,I164679,I164696,I164200,I164203,I164741,I164758,I164775,I164792,I164230,I164823,I164215,I164218,I164901,I164918,I320125,I164935,I320122,I320113,I164952,I320116,I164969,I164986,I320110,I165003,I165020,I164890,I165051,I164875,I165082,I320131,I165099,I320134,I165116,I320119,I165133,I320107,I165150,I165167,I165184,I164872,I165215,I165232,I164869,I165263,I320128,I165280,I164887,I165311,I164884,I165342,I165359,I164863,I164866,I165404,I320137,I165421,I165438,I165455,I164893,I165486,I164878,I164881,I165564,I165581,I371606,I165598,I371624,I371615,I165615,I371621,I165632,I165649,I371627,I165666,I165683,I165714,I165745,I371603,I165762,I371618,I165779,I371600,I165796,I371609,I165813,I165830,I165847,I165878,I165895,I165926,I371612,I165943,I165974,I166005,I166022,I166067,I371630,I166084,I166101,I166118,I166149,I166227,I166244,I366574,I166261,I366592,I366583,I166278,I366589,I166295,I166312,I366595,I166329,I166346,I166377,I166408,I366571,I166425,I366586,I166442,I366568,I166459,I366577,I166476,I166493,I166510,I166541,I166558,I166589,I366580,I166606,I166637,I166668,I166685,I166730,I366598,I166747,I166764,I166781,I166812,I166890,I166907,I166924,I166941,I166958,I166975,I166992,I167009,I167040,I167071,I167088,I167105,I167122,I167139,I167156,I167173,I167204,I167221,I167252,I167269,I167300,I167331,I167348,I167393,I167410,I167427,I167444,I167475,I167553,I167570,I210809,I167587,I210806,I210824,I167604,I210827,I167621,I167638,I210812,I167655,I167672,I167542,I167703,I167527,I167734,I210821,I167751,I210803,I167768,I210797,I167785,I210815,I167802,I167819,I167836,I167524,I167867,I167884,I167521,I167915,I210800,I167932,I167539,I167963,I167536,I167994,I168011,I167515,I167518,I168056,I210818,I168073,I168090,I168107,I167545,I168138,I167530,I167533,I168216,I168233,I168250,I168267,I168284,I168301,I168318,I168335,I168205,I168366,I168190,I168397,I168414,I168431,I168448,I168465,I168482,I168499,I168187,I168530,I168547,I168184,I168578,I168595,I168202,I168626,I168199,I168657,I168674,I168178,I168181,I168719,I168736,I168753,I168770,I168208,I168801,I168193,I168196,I168879,I168896,I290375,I168913,I290384,I290366,I168930,I290387,I168947,I168964,I290378,I168981,I168998,I168868,I169029,I168853,I169060,I290372,I169077,I290363,I169094,I290360,I169111,I290357,I169128,I169145,I169162,I168850,I169193,I169210,I168847,I169241,I290381,I169258,I168865,I169289,I168862,I169320,I169337,I168841,I168844,I169382,I290369,I169399,I169416,I169433,I168871,I169464,I168856,I168859,I169542,I169559,I317745,I169576,I317742,I317733,I169593,I317736,I169610,I169627,I317730,I169644,I169661,I169692,I169723,I317751,I169740,I317754,I169757,I317739,I169774,I317727,I169791,I169808,I169825,I169856,I169873,I169904,I317748,I169921,I169952,I169983,I170000,I170045,I317757,I170062,I170079,I170096,I170127,I170205,I170222,I170239,I170256,I170273,I170290,I170307,I170324,I170194,I170355,I170179,I170386,I170403,I170420,I170437,I170454,I170471,I170488,I170176,I170519,I170536,I170173,I170567,I170584,I170191,I170615,I170188,I170646,I170663,I170167,I170170,I170708,I170725,I170742,I170759,I170197,I170790,I170182,I170185,I170868,I170885,I270927,I170902,I270924,I270921,I170919,I270909,I170936,I170953,I270930,I170970,I170987,I171018,I171049,I270912,I171066,I270918,I171083,I270915,I171100,I270939,I171117,I171134,I171151,I171182,I171199,I171230,I270936,I171247,I171278,I171309,I171326,I171371,I270933,I171388,I171405,I171422,I171453,I171531,I171548,I208225,I171565,I208222,I208240,I171582,I208243,I171599,I171616,I208228,I171633,I171650,I171520,I171681,I171505,I171712,I208237,I171729,I208219,I171746,I208213,I171763,I208231,I171780,I171797,I171814,I171502,I171845,I171862,I171499,I171893,I208216,I171910,I171517,I171941,I171514,I171972,I171989,I171493,I171496,I172034,I208234,I172051,I172068,I172085,I171523,I172116,I171508,I171511,I172194,I172211,I252190,I172228,I252202,I252184,I172245,I252205,I172262,I172279,I252196,I172296,I172313,I172183,I172344,I172168,I172375,I252187,I172392,I252181,I172409,I252193,I172426,I252178,I172443,I172460,I172477,I172165,I172508,I172525,I172162,I172556,I252175,I172573,I172180,I172604,I172177,I172635,I172652,I172156,I172159,I172697,I252199,I172714,I172731,I172748,I172186,I172779,I172171,I172174,I172857,I172874,I172891,I172908,I172925,I172942,I172959,I172976,I173007,I173038,I173055,I173072,I173089,I173106,I173123,I173140,I173171,I173188,I173219,I173236,I173267,I173298,I173315,I173360,I173377,I173394,I173411,I173442,I173520,I173537,I360913,I173554,I360931,I360922,I173571,I360928,I173588,I173605,I360934,I173622,I173639,I173509,I173670,I173494,I173701,I360910,I173718,I360925,I173735,I360907,I173752,I360916,I173769,I173786,I173803,I173491,I173834,I173851,I173488,I173882,I360919,I173899,I173506,I173930,I173503,I173961,I173978,I173482,I173485,I174023,I360937,I174040,I174057,I174074,I173512,I174105,I173497,I173500,I174183,I174200,I229543,I174217,I229540,I229558,I174234,I229561,I174251,I174268,I229546,I174285,I174302,I174172,I174333,I174157,I174364,I229555,I174381,I229537,I174398,I229531,I174415,I229549,I174432,I174449,I174466,I174154,I174497,I174514,I174151,I174545,I229534,I174562,I174169,I174593,I174166,I174624,I174641,I174145,I174148,I174686,I229552,I174703,I174720,I174737,I174175,I174768,I174160,I174163,I174846,I174863,I235215,I174880,I235218,I235224,I174897,I235230,I174914,I174931,I235209,I174948,I174965,I174835,I174996,I174820,I175027,I235221,I175044,I235236,I175061,I235239,I175078,I235212,I175095,I175112,I175129,I174817,I175160,I175177,I174814,I175208,I235233,I175225,I174832,I175256,I174829,I175287,I175304,I174808,I174811,I175349,I235227,I175366,I175383,I175400,I174838,I175431,I174823,I174826,I175509,I175526,I372235,I175543,I372253,I372244,I175560,I372250,I175577,I175594,I372256,I175611,I175628,I175659,I175690,I372232,I175707,I372247,I175724,I372229,I175741,I372238,I175758,I175775,I175792,I175823,I175840,I175871,I372241,I175888,I175919,I175950,I175967,I176012,I372259,I176029,I176046,I176063,I176094,I176172,I176189,I365945,I176206,I365963,I365954,I176223,I365960,I176240,I176257,I365966,I176274,I176291,I176161,I176322,I176146,I176353,I365942,I176370,I365957,I176387,I365939,I176404,I365948,I176421,I176438,I176455,I176143,I176486,I176503,I176140,I176534,I365951,I176551,I176158,I176582,I176155,I176613,I176630,I176134,I176137,I176675,I365969,I176692,I176709,I176726,I176164,I176757,I176149,I176152,I176835,I176852,I277304,I176869,I277325,I277331,I176886,I277319,I176903,I176920,I277301,I176937,I176954,I176824,I176985,I176809,I177016,I277307,I177033,I277328,I177050,I277316,I177067,I277322,I177084,I177101,I177118,I176806,I177149,I177166,I176803,I177197,I277313,I177214,I176821,I177245,I176818,I177276,I177293,I176797,I176800,I177338,I277310,I177355,I177372,I177389,I176827,I177420,I176812,I176815,I177498,I177515,I362171,I177532,I362189,I362180,I177549,I362186,I177566,I177583,I362192,I177600,I177617,I177648,I177679,I362168,I177696,I362183,I177713,I362165,I177730,I362174,I177747,I177764,I177781,I177812,I177829,I177860,I362177,I177877,I177908,I177939,I177956,I178001,I362195,I178018,I178035,I178052,I178083,I178161,I178178,I178195,I178212,I178229,I178246,I178263,I178280,I178150,I178311,I178135,I178342,I178359,I178376,I178393,I178410,I178427,I178444,I178132,I178475,I178492,I178129,I178523,I178540,I178147,I178571,I178144,I178602,I178619,I178123,I178126,I178664,I178681,I178698,I178715,I178153,I178746,I178138,I178141,I178824,I178841,I178858,I178875,I178892,I178909,I178926,I178943,I178974,I179005,I179022,I179039,I179056,I179073,I179090,I179107,I179138,I179155,I179186,I179203,I179234,I179265,I179282,I179327,I179344,I179361,I179378,I179409,I179487,I179504,I374122,I179521,I374140,I374131,I179538,I374137,I179555,I179572,I374143,I179589,I179606,I179476,I179637,I179461,I179668,I374119,I179685,I374134,I179702,I374116,I179719,I374125,I179736,I179753,I179770,I179458,I179801,I179818,I179455,I179849,I374128,I179866,I179473,I179897,I179470,I179928,I179945,I179449,I179452,I179990,I374146,I180007,I180024,I180041,I179479,I180072,I179464,I179467,I180150,I180167,I367203,I180184,I367221,I367212,I180201,I367218,I180218,I180235,I367224,I180252,I180269,I180139,I180300,I180124,I180331,I367200,I180348,I367215,I180365,I367197,I180382,I367206,I180399,I180416,I180433,I180121,I180464,I180481,I180118,I180512,I367209,I180529,I180136,I180560,I180133,I180591,I180608,I180112,I180115,I180653,I367227,I180670,I180687,I180704,I180142,I180735,I180127,I180130,I180813,I180830,I249878,I180847,I249890,I249872,I180864,I249893,I180881,I180898,I249884,I180915,I180932,I180963,I180994,I249875,I181011,I249869,I181028,I249881,I181045,I249866,I181062,I181079,I181096,I181127,I181144,I181175,I249863,I181192,I181223,I181254,I181271,I181316,I249887,I181333,I181350,I181367,I181398,I181476,I181493,I264328,I181510,I264340,I264322,I181527,I264343,I181544,I181561,I264334,I181578,I181595,I181465,I181626,I181450,I181657,I264325,I181674,I264319,I181691,I264331,I181708,I264316,I181725,I181742,I181759,I181447,I181790,I181807,I181444,I181838,I264313,I181855,I181462,I181886,I181459,I181917,I181934,I181438,I181441,I181979,I264337,I181996,I182013,I182030,I181468,I182061,I181453,I181456,I182139,I182156,I182173,I182190,I182207,I182224,I182241,I182258,I182128,I182289,I182113,I182320,I182337,I182354,I182371,I182388,I182405,I182422,I182110,I182453,I182470,I182107,I182501,I182518,I182125,I182549,I182122,I182580,I182597,I182101,I182104,I182642,I182659,I182676,I182693,I182131,I182724,I182116,I182119,I182802,I182819,I365316,I182836,I365334,I365325,I182853,I365331,I182870,I182887,I365337,I182904,I182921,I182791,I182952,I182776,I182983,I365313,I183000,I365328,I183017,I365310,I183034,I365319,I183051,I183068,I183085,I182773,I183116,I183133,I182770,I183164,I365322,I183181,I182788,I183212,I182785,I183243,I183260,I182764,I182767,I183305,I365340,I183322,I183339,I183356,I182794,I183387,I182779,I182782,I183465,I183482,I289780,I183499,I289789,I289771,I183516,I289792,I183533,I183550,I289783,I183567,I183584,I183615,I183646,I289777,I183663,I289768,I183680,I289765,I183697,I289762,I183714,I183731,I183748,I183779,I183796,I183827,I289786,I183844,I183875,I183906,I183923,I183968,I289774,I183985,I184002,I184019,I184050,I184128,I184145,I184162,I184179,I184196,I184213,I184230,I184247,I184278,I184309,I184326,I184343,I184360,I184377,I184394,I184411,I184442,I184459,I184490,I184507,I184538,I184569,I184586,I184631,I184648,I184665,I184682,I184713,I184791,I184808,I255658,I184825,I255670,I255652,I184842,I255673,I184859,I184876,I255664,I184893,I184910,I184780,I184941,I184765,I184972,I255655,I184989,I255649,I185006,I255661,I185023,I255646,I185040,I185057,I185074,I184762,I185105,I185122,I184759,I185153,I255643,I185170,I184777,I185201,I184774,I185232,I185249,I184753,I184756,I185294,I255667,I185311,I185328,I185345,I184783,I185376,I184768,I184771,I185454,I185471,I358397,I185488,I358415,I358406,I185505,I358412,I185522,I185539,I358418,I185556,I185573,I185443,I185604,I185428,I185635,I358394,I185652,I358409,I185669,I358391,I185686,I358400,I185703,I185720,I185737,I185425,I185768,I185785,I185422,I185816,I358403,I185833,I185440,I185864,I185437,I185895,I185912,I185416,I185419,I185957,I358421,I185974,I185991,I186008,I185446,I186039,I185431,I185434,I186117,I186134,I245254,I186151,I245266,I245248,I186168,I245269,I186185,I186202,I245260,I186219,I186236,I186106,I186267,I186091,I186298,I245251,I186315,I245245,I186332,I245257,I186349,I245242,I186366,I186383,I186400,I186088,I186431,I186448,I186085,I186479,I245239,I186496,I186103,I186527,I186100,I186558,I186575,I186079,I186082,I186620,I245263,I186637,I186654,I186671,I186109,I186702,I186094,I186097,I186780,I186797,I308225,I186814,I308234,I308216,I186831,I308237,I186848,I186865,I308228,I186882,I186899,I186930,I186961,I308222,I186978,I308213,I186995,I308210,I187012,I308207,I187029,I187046,I187063,I187094,I187111,I187142,I308231,I187159,I187190,I187221,I187238,I187283,I308219,I187300,I187317,I187334,I187365,I187443,I187460,I285615,I187477,I285624,I285606,I187494,I285627,I187511,I187528,I285618,I187545,I187562,I187432,I187593,I187417,I187624,I285612,I187641,I285603,I187658,I285600,I187675,I285597,I187692,I187709,I187726,I187414,I187757,I187774,I187411,I187805,I285621,I187822,I187429,I187853,I187426,I187884,I187901,I187405,I187408,I187946,I285609,I187963,I187980,I187997,I187435,I188028,I187420,I187423,I188106,I188123,I188140,I188157,I188174,I188191,I188208,I188225,I188095,I188256,I188080,I188287,I188304,I188321,I188338,I188355,I188372,I188389,I188077,I188420,I188437,I188074,I188468,I188485,I188092,I188516,I188089,I188547,I188564,I188068,I188071,I188609,I188626,I188643,I188660,I188098,I188691,I188083,I188086,I188769,I188786,I188803,I188820,I188837,I188854,I188871,I188888,I188758,I188919,I188743,I188950,I188967,I188984,I189001,I189018,I189035,I189052,I188740,I189083,I189100,I188737,I189131,I189148,I188755,I189179,I188752,I189210,I189227,I188731,I188734,I189272,I189289,I189306,I189323,I188761,I189354,I188746,I188749,I189432,I189449,I227605,I189466,I227602,I227620,I189483,I227623,I189500,I189517,I227608,I189534,I189551,I189421,I189582,I189406,I189613,I227617,I189630,I227599,I189647,I227593,I189664,I227611,I189681,I189698,I189715,I189403,I189746,I189763,I189400,I189794,I227596,I189811,I189418,I189842,I189415,I189873,I189890,I189394,I189397,I189935,I227614,I189952,I189969,I189986,I189424,I190017,I189409,I189412,I190095,I190112,I355881,I190129,I355899,I355890,I190146,I355896,I190163,I190180,I355902,I190197,I190214,I190084,I190245,I190069,I190276,I355878,I190293,I355893,I190310,I355875,I190327,I355884,I190344,I190361,I190378,I190066,I190409,I190426,I190063,I190457,I355887,I190474,I190081,I190505,I190078,I190536,I190553,I190057,I190060,I190598,I355905,I190615,I190632,I190649,I190087,I190680,I190072,I190075,I190758,I190775,I190792,I190809,I190826,I190843,I190860,I190877,I190908,I190939,I190956,I190973,I190990,I191007,I191024,I191041,I191072,I191089,I191120,I191137,I191168,I191199,I191216,I191261,I191278,I191295,I191312,I191343,I191421,I191438,I390295,I191455,I390286,I390292,I191472,I390304,I191489,I191506,I390289,I191523,I191540,I191410,I191571,I191395,I191602,I390313,I191619,I390307,I191636,I390298,I191653,I390283,I191670,I191687,I191704,I191392,I191735,I191752,I191389,I191783,I390301,I191800,I191407,I191831,I191404,I191862,I191879,I191383,I191386,I191924,I390310,I191941,I191958,I191975,I191413,I192006,I191398,I191401,I192084,I192101,I192118,I192135,I192152,I192169,I192186,I192203,I192234,I192265,I192282,I192299,I192316,I192333,I192350,I192367,I192398,I192415,I192446,I192463,I192494,I192525,I192542,I192587,I192604,I192621,I192638,I192669,I192747,I192764,I192781,I192798,I192815,I192832,I192849,I192718,I192880,I192897,I192914,I192931,I192948,I192965,I192982,I192715,I193013,I192709,I193044,I193061,I193078,I192739,I192712,I193123,I192736,I193154,I192733,I192730,I193199,I193216,I193233,I193250,I193267,I192724,I193298,I193315,I192727,I192721,I193393,I193410,I193427,I193444,I193461,I193478,I193495,I193364,I193526,I193543,I193560,I193577,I193594,I193611,I193628,I193361,I193659,I193355,I193690,I193707,I193724,I193385,I193358,I193769,I193382,I193800,I193379,I193376,I193845,I193862,I193879,I193896,I193913,I193370,I193944,I193961,I193373,I193367,I194039,I194056,I321315,I194073,I321303,I321312,I194090,I321327,I194107,I194124,I321309,I194141,I194010,I194172,I194189,I194206,I321297,I194223,I321318,I194240,I321300,I194257,I321306,I194274,I194007,I194305,I194001,I194336,I194353,I194370,I194031,I194004,I194415,I321324,I194028,I194446,I194025,I194022,I194491,I321321,I194508,I194525,I194542,I194559,I194016,I194590,I194607,I194019,I194013,I194685,I194702,I194719,I194736,I194753,I194770,I194787,I194818,I194835,I194852,I194869,I194886,I194903,I194920,I194951,I194982,I194999,I195016,I195061,I195092,I195137,I195154,I195171,I195188,I195205,I195236,I195253,I195331,I195348,I304646,I195365,I304658,I304652,I195382,I304637,I195399,I195416,I304664,I195433,I195302,I195464,I195481,I195498,I304661,I195515,I304643,I195532,I304640,I195549,I304667,I195566,I195299,I195597,I195293,I195628,I195645,I195662,I195323,I195296,I195707,I304655,I195320,I195738,I195317,I195314,I195783,I304649,I195800,I195817,I195834,I195851,I195308,I195882,I195899,I195311,I195305,I195977,I195994,I196011,I196028,I196045,I196062,I196079,I196110,I196127,I196144,I196161,I196178,I196195,I196212,I196243,I196274,I196291,I196308,I196353,I196384,I196429,I196446,I196463,I196480,I196497,I196528,I196545,I196623,I196640,I196657,I196674,I196691,I196708,I196725,I196594,I196756,I196773,I196790,I196807,I196824,I196841,I196858,I196591,I196889,I196585,I196920,I196937,I196954,I196615,I196588,I196999,I196612,I197030,I196609,I196606,I197075,I197092,I197109,I197126,I197143,I196600,I197174,I197191,I196603,I196597,I197269,I197286,I261438,I197303,I261441,I261423,I197320,I261450,I197337,I197354,I261429,I197371,I197240,I197402,I197419,I197436,I261435,I197453,I261447,I197470,I261453,I197487,I261432,I197504,I197237,I197535,I197231,I197566,I197583,I197600,I197261,I197234,I197645,I261444,I197258,I197676,I197255,I197252,I197721,I261426,I197738,I197755,I197772,I197789,I197246,I197820,I197837,I197249,I197243,I197915,I197932,I197949,I197966,I197983,I198000,I198017,I198048,I198065,I198082,I198099,I198116,I198133,I198150,I198181,I198212,I198229,I198246,I198291,I198322,I198367,I198384,I198401,I198418,I198435,I198466,I198483,I198561,I198578,I369105,I198595,I369102,I369087,I198612,I369096,I198629,I198646,I369111,I198663,I198532,I198694,I198711,I198728,I369084,I198745,I369090,I198762,I369114,I198779,I369108,I198796,I198529,I198827,I198523,I198858,I198875,I198892,I198553,I198526,I198937,I369093,I198550,I198968,I198547,I198544,I199013,I369099,I199030,I199047,I199064,I199081,I198538,I199112,I199129,I198541,I198535,I199207,I199224,I199241,I199258,I199275,I199292,I199309,I199340,I199357,I199374,I199391,I199408,I199425,I199442,I199473,I199504,I199521,I199538,I199583,I199614,I199659,I199676,I199693,I199710,I199727,I199758,I199775,I199853,I199870,I324885,I199887,I324873,I324882,I199904,I324897,I199921,I199938,I324879,I199955,I199986,I200003,I200020,I324867,I200037,I324888,I200054,I324870,I200071,I324876,I200088,I200119,I200150,I200167,I200184,I200229,I324894,I200260,I200305,I324891,I200322,I200339,I200356,I200373,I200404,I200421,I200499,I200516,I200533,I200550,I200567,I200584,I200601,I200470,I200632,I200649,I200666,I200683,I200700,I200717,I200734,I200467,I200765,I200461,I200796,I200813,I200830,I200491,I200464,I200875,I200488,I200906,I200485,I200482,I200951,I200968,I200985,I201002,I201019,I200476,I201050,I201067,I200479,I200473,I201145,I201162,I201179,I201196,I201213,I201230,I201247,I201278,I201295,I201312,I201329,I201346,I201363,I201380,I201411,I201442,I201459,I201476,I201521,I201552,I201597,I201614,I201631,I201648,I201665,I201696,I201713,I201791,I201808,I373508,I201825,I373505,I373490,I201842,I373499,I201859,I201876,I373514,I201893,I201924,I201941,I201958,I373487,I201975,I373493,I201992,I373517,I202009,I373511,I202026,I202057,I202088,I202105,I202122,I202167,I373496,I202198,I202243,I373502,I202260,I202277,I202294,I202311,I202342,I202359,I202437,I202454,I202471,I202488,I202505,I202522,I202539,I202570,I202587,I202604,I202621,I202638,I202655,I202672,I202703,I202734,I202751,I202768,I202813,I202844,I202889,I202906,I202923,I202940,I202957,I202988,I203005,I203083,I203100,I203117,I203134,I203151,I203168,I203185,I203216,I203233,I203250,I203267,I203284,I203301,I203318,I203349,I203380,I203397,I203414,I203459,I203490,I203535,I203552,I203569,I203586,I203603,I203634,I203651,I203729,I203746,I203763,I203780,I203797,I203814,I203831,I203700,I203862,I203879,I203896,I203913,I203930,I203947,I203964,I203697,I203995,I203691,I204026,I204043,I204060,I203721,I203694,I204105,I203718,I204136,I203715,I203712,I204181,I204198,I204215,I204232,I204249,I203706,I204280,I204297,I203709,I203703,I204375,I204392,I246988,I204409,I246991,I246973,I204426,I247000,I204443,I204460,I246979,I204477,I204508,I204525,I204542,I246985,I204559,I246997,I204576,I247003,I204593,I246982,I204610,I204641,I204672,I204689,I204706,I204751,I246994,I204782,I204827,I246976,I204844,I204861,I204878,I204895,I204926,I204943,I205021,I205038,I276741,I205055,I276747,I276732,I205072,I276726,I205089,I205106,I276753,I205123,I204992,I205154,I205171,I205188,I276738,I205205,I276744,I205222,I276750,I205239,I276723,I205256,I204989,I205287,I204983,I205318,I205335,I205352,I205013,I204986,I205397,I276729,I205010,I205428,I205007,I205004,I205473,I276735,I205490,I205507,I205524,I205541,I204998,I205572,I205589,I205001,I204995,I205667,I205684,I205701,I205718,I205735,I205752,I205769,I205638,I205800,I205817,I205834,I205851,I205868,I205885,I205902,I205635,I205933,I205629,I205964,I205981,I205998,I205659,I205632,I206043,I205656,I206074,I205653,I205650,I206119,I206136,I206153,I206170,I206187,I205644,I206218,I206235,I205647,I205641,I206313,I206330,I206347,I206364,I206381,I206398,I206415,I206446,I206463,I206480,I206497,I206514,I206531,I206548,I206579,I206610,I206627,I206644,I206689,I206720,I206765,I206782,I206799,I206816,I206833,I206864,I206881,I206959,I206976,I206993,I207010,I207027,I207044,I207061,I206930,I207092,I207109,I207126,I207143,I207160,I207177,I207194,I206927,I207225,I206921,I207256,I207273,I207290,I206951,I206924,I207335,I206948,I207366,I206945,I206942,I207411,I207428,I207445,I207462,I207479,I206936,I207510,I207527,I206939,I206933,I207605,I207622,I207639,I207656,I207673,I207690,I207707,I207576,I207738,I207755,I207772,I207789,I207806,I207823,I207840,I207573,I207871,I207567,I207902,I207919,I207936,I207597,I207570,I207981,I207594,I208012,I207591,I207588,I208057,I208074,I208091,I208108,I208125,I207582,I208156,I208173,I207585,I207579,I208251,I208268,I342687,I208285,I342684,I342669,I208302,I342678,I208319,I208336,I342693,I208353,I208384,I208401,I208418,I342666,I208435,I342672,I208452,I342696,I208469,I342690,I208486,I208517,I208548,I208565,I208582,I208627,I342675,I208658,I208703,I342681,I208720,I208737,I208754,I208771,I208802,I208819,I208897,I208914,I361557,I208931,I361554,I361539,I208948,I361548,I208965,I208982,I361563,I208999,I209030,I209047,I209064,I361536,I209081,I361542,I209098,I361566,I209115,I361560,I209132,I209163,I209194,I209211,I209228,I209273,I361545,I209304,I209349,I361551,I209366,I209383,I209400,I209417,I209448,I209465,I209543,I209560,I376653,I209577,I376650,I376635,I209594,I376644,I209611,I209628,I376659,I209645,I209676,I209693,I209710,I376632,I209727,I376638,I209744,I376662,I209761,I376656,I209778,I209809,I209840,I209857,I209874,I209919,I376641,I209950,I209995,I376647,I210012,I210029,I210046,I210063,I210094,I210111,I210189,I210206,I393769,I210223,I393754,I393760,I210240,I393757,I210257,I210274,I393766,I210291,I210160,I210322,I210339,I210356,I393781,I210373,I393775,I210390,I393772,I210407,I393751,I210424,I210157,I210455,I210151,I210486,I210503,I210520,I210181,I210154,I210565,I393778,I210178,I210596,I210175,I210172,I210641,I393763,I210658,I210675,I210692,I210709,I210166,I210740,I210757,I210169,I210163,I210835,I210852,I291556,I210869,I291568,I291562,I210886,I291547,I210903,I210920,I291574,I210937,I210968,I210985,I211002,I291571,I211019,I291553,I211036,I291550,I211053,I291577,I211070,I211101,I211132,I211149,I211166,I211211,I291565,I211242,I211287,I291559,I211304,I211321,I211338,I211355,I211386,I211403,I211481,I211498,I211515,I211532,I211549,I211566,I211583,I211614,I211631,I211648,I211665,I211682,I211699,I211716,I211747,I211778,I211795,I211812,I211857,I211888,I211933,I211950,I211967,I211984,I212001,I212032,I212049,I212127,I212144,I321910,I212161,I321898,I321907,I212178,I321922,I212195,I212212,I321904,I212229,I212098,I212260,I212277,I212294,I321892,I212311,I321913,I212328,I321895,I212345,I321901,I212362,I212095,I212393,I212089,I212424,I212441,I212458,I212119,I212092,I212503,I321919,I212116,I212534,I212113,I212110,I212579,I321916,I212596,I212613,I212630,I212647,I212104,I212678,I212695,I212107,I212101,I212773,I212790,I212807,I212824,I212841,I212858,I212875,I212744,I212906,I212923,I212940,I212957,I212974,I212991,I213008,I212741,I213039,I212735,I213070,I213087,I213104,I212765,I212738,I213149,I212762,I213180,I212759,I212756,I213225,I213242,I213259,I213276,I213293,I212750,I213324,I213341,I212753,I212747,I213419,I213436,I348977,I213453,I348974,I348959,I213470,I348968,I213487,I213504,I348983,I213521,I213390,I213552,I213569,I213586,I348956,I213603,I348962,I213620,I348986,I213637,I348980,I213654,I213387,I213685,I213381,I213716,I213733,I213750,I213411,I213384,I213795,I348965,I213408,I213826,I213405,I213402,I213871,I348971,I213888,I213905,I213922,I213939,I213396,I213970,I213987,I213399,I213393,I214065,I214082,I214099,I214116,I214133,I214150,I214167,I214036,I214198,I214215,I214232,I214249,I214266,I214283,I214300,I214033,I214331,I214027,I214362,I214379,I214396,I214057,I214030,I214441,I214054,I214472,I214051,I214048,I214517,I214534,I214551,I214568,I214585,I214042,I214616,I214633,I214045,I214039,I214711,I214728,I214745,I214762,I214779,I214796,I214813,I214844,I214861,I214878,I214895,I214912,I214929,I214946,I214977,I215008,I215025,I215042,I215087,I215118,I215163,I215180,I215197,I215214,I215231,I215262,I215279,I215357,I215374,I360299,I215391,I360296,I360281,I215408,I360290,I215425,I215442,I360305,I215459,I215490,I215507,I215524,I360278,I215541,I360284,I215558,I360308,I215575,I360302,I215592,I215623,I215654,I215671,I215688,I215733,I360287,I215764,I215809,I360293,I215826,I215843,I215860,I215877,I215908,I215925,I216003,I216020,I364702,I216037,I364699,I364684,I216054,I364693,I216071,I216088,I364708,I216105,I215974,I216136,I216153,I216170,I364681,I216187,I364687,I216204,I364711,I216221,I364705,I216238,I215971,I216269,I215965,I216300,I216317,I216334,I215995,I215968,I216379,I364690,I215992,I216410,I215989,I215986,I216455,I364696,I216472,I216489,I216506,I216523,I215980,I216554,I216571,I215983,I215977,I216649,I216666,I295126,I216683,I295138,I295132,I216700,I295117,I216717,I216734,I295144,I216751,I216782,I216799,I216816,I295141,I216833,I295123,I216850,I295120,I216867,I295147,I216884,I216915,I216946,I216963,I216980,I217025,I295135,I217056,I217101,I295129,I217118,I217135,I217152,I217169,I217200,I217217,I217295,I217312,I217329,I217346,I217363,I217380,I217397,I217428,I217445,I217462,I217479,I217496,I217513,I217530,I217561,I217592,I217609,I217626,I217671,I217702,I217747,I217764,I217781,I217798,I217815,I217846,I217863,I217941,I217958,I389145,I217975,I389130,I389136,I217992,I389133,I218009,I218026,I389142,I218043,I217912,I218074,I218091,I218108,I389157,I218125,I389151,I218142,I389148,I218159,I389127,I218176,I217909,I218207,I217903,I218238,I218255,I218272,I217933,I217906,I218317,I389154,I217930,I218348,I217927,I217924,I218393,I389139,I218410,I218427,I218444,I218461,I217918,I218492,I218509,I217921,I217915,I218587,I218604,I218621,I218638,I218655,I218672,I218689,I218558,I218720,I218737,I218754,I218771,I218788,I218805,I218822,I218555,I218853,I218549,I218884,I218901,I218918,I218579,I218552,I218963,I218576,I218994,I218573,I218570,I219039,I219056,I219073,I219090,I219107,I218564,I219138,I219155,I218567,I218561,I219233,I219250,I219267,I219284,I219301,I219318,I219335,I219204,I219366,I219383,I219400,I219417,I219434,I219451,I219468,I219201,I219499,I219195,I219530,I219547,I219564,I219225,I219198,I219609,I219222,I219640,I219219,I219216,I219685,I219702,I219719,I219736,I219753,I219210,I219784,I219801,I219213,I219207,I219879,I219896,I342058,I219913,I342055,I342040,I219930,I342049,I219947,I219964,I342064,I219981,I219850,I220012,I220029,I220046,I342037,I220063,I342043,I220080,I342067,I220097,I342061,I220114,I219847,I220145,I219841,I220176,I220193,I220210,I219871,I219844,I220255,I342046,I219868,I220286,I219865,I219862,I220331,I342052,I220348,I220365,I220382,I220399,I219856,I220430,I220447,I219859,I219853,I220525,I220542,I220559,I220576,I220593,I220610,I220627,I220496,I220658,I220675,I220692,I220709,I220726,I220743,I220760,I220493,I220791,I220487,I220822,I220839,I220856,I220517,I220490,I220901,I220514,I220932,I220511,I220508,I220977,I220994,I221011,I221028,I221045,I220502,I221076,I221093,I220505,I220499,I221171,I221188,I221205,I221222,I221239,I221256,I221273,I221142,I221304,I221321,I221338,I221355,I221372,I221389,I221406,I221139,I221437,I221133,I221468,I221485,I221502,I221163,I221136,I221547,I221160,I221578,I221157,I221154,I221623,I221640,I221657,I221674,I221691,I221148,I221722,I221739,I221151,I221145,I221817,I221834,I221851,I221868,I221885,I221902,I221919,I221950,I221967,I221984,I222001,I222018,I222035,I222052,I222083,I222114,I222131,I222148,I222193,I222224,I222269,I222286,I222303,I222320,I222337,I222368,I222385,I222463,I222480,I222497,I222514,I222531,I222548,I222565,I222596,I222613,I222630,I222647,I222664,I222681,I222698,I222729,I222760,I222777,I222794,I222839,I222870,I222915,I222932,I222949,I222966,I222983,I223014,I223031,I223109,I223126,I346461,I223143,I346458,I346443,I223160,I346452,I223177,I223194,I346467,I223211,I223080,I223242,I223259,I223276,I346440,I223293,I346446,I223310,I346470,I223327,I346464,I223344,I223077,I223375,I223071,I223406,I223423,I223440,I223101,I223074,I223485,I346449,I223098,I223516,I223095,I223092,I223561,I346455,I223578,I223595,I223612,I223629,I223086,I223660,I223677,I223089,I223083,I223755,I223772,I223789,I223806,I223823,I223840,I223857,I223726,I223888,I223905,I223922,I223939,I223956,I223973,I223990,I223723,I224021,I223717,I224052,I224069,I224086,I223747,I223720,I224131,I223744,I224162,I223741,I223738,I224207,I224224,I224241,I224258,I224275,I223732,I224306,I224323,I223735,I223729,I224401,I224418,I234615,I224435,I234624,I234609,I224452,I234597,I224469,I224486,I234600,I224503,I224534,I224551,I224568,I234612,I224585,I234606,I224602,I234603,I224619,I234618,I224636,I224667,I224698,I224715,I224732,I224777,I234627,I224808,I224853,I234621,I224870,I224887,I224904,I224921,I224952,I224969,I225047,I225064,I225081,I225098,I225115,I225132,I225149,I225180,I225197,I225214,I225231,I225248,I225265,I225282,I225313,I225344,I225361,I225378,I225423,I225454,I225499,I225516,I225533,I225550,I225567,I225598,I225615,I225693,I225710,I225727,I225744,I225761,I225778,I225795,I225664,I225826,I225843,I225860,I225877,I225894,I225911,I225928,I225661,I225959,I225655,I225990,I226007,I226024,I225685,I225658,I226069,I225682,I226100,I225679,I225676,I226145,I226162,I226179,I226196,I226213,I225670,I226244,I226261,I225673,I225667,I226339,I226356,I226373,I226390,I226407,I226424,I226441,I226472,I226489,I226506,I226523,I226540,I226557,I226574,I226605,I226636,I226653,I226670,I226715,I226746,I226791,I226808,I226825,I226842,I226859,I226890,I226907,I226985,I227002,I227019,I227036,I227053,I227070,I227087,I227118,I227135,I227152,I227169,I227186,I227203,I227220,I227251,I227282,I227299,I227316,I227361,I227392,I227437,I227454,I227471,I227488,I227505,I227536,I227553,I227631,I227648,I376024,I227665,I376021,I376006,I227682,I376015,I227699,I227716,I376030,I227733,I227764,I227781,I227798,I376003,I227815,I376009,I227832,I376033,I227849,I376027,I227866,I227897,I227928,I227945,I227962,I228007,I376012,I228038,I228083,I376018,I228100,I228117,I228134,I228151,I228182,I228199,I228277,I228294,I343316,I228311,I343313,I343298,I228328,I343307,I228345,I228362,I343322,I228379,I228248,I228410,I228427,I228444,I343295,I228461,I343301,I228478,I343325,I228495,I343319,I228512,I228245,I228543,I228239,I228574,I228591,I228608,I228269,I228242,I228653,I343304,I228266,I228684,I228263,I228260,I228729,I343310,I228746,I228763,I228780,I228797,I228254,I228828,I228845,I228257,I228251,I228923,I228940,I228957,I228974,I228991,I229008,I229025,I228894,I229056,I229073,I229090,I229107,I229124,I229141,I229158,I228891,I229189,I228885,I229220,I229237,I229254,I228915,I228888,I229299,I228912,I229330,I228909,I228906,I229375,I229392,I229409,I229426,I229443,I228900,I229474,I229491,I228903,I228897,I229569,I229586,I264906,I229603,I264909,I264891,I229620,I264918,I229637,I229654,I264897,I229671,I229702,I229719,I229736,I264903,I229753,I264915,I229770,I264921,I229787,I264900,I229804,I229835,I229866,I229883,I229900,I229945,I264912,I229976,I230021,I264894,I230038,I230055,I230072,I230089,I230120,I230137,I230215,I230232,I232779,I230249,I232788,I232773,I230266,I232761,I230283,I230300,I232764,I230317,I230348,I230365,I230382,I232776,I230399,I232770,I230416,I232767,I230433,I232782,I230450,I230481,I230512,I230529,I230546,I230591,I232791,I230622,I230667,I232785,I230684,I230701,I230718,I230735,I230766,I230783,I230861,I230878,I237675,I230895,I237684,I237669,I230912,I237657,I230929,I230946,I237660,I230963,I230832,I230994,I231011,I231028,I237672,I231045,I237666,I231062,I237663,I231079,I237678,I231096,I230829,I231127,I230823,I231158,I231175,I231192,I230853,I230826,I231237,I237687,I230850,I231268,I230847,I230844,I231313,I237681,I231330,I231347,I231364,I231381,I230838,I231412,I231429,I230841,I230835,I231507,I231524,I231541,I231558,I231575,I231592,I231609,I231640,I231657,I231674,I231691,I231708,I231725,I231742,I231773,I231804,I231821,I231838,I231883,I231914,I231959,I231976,I231993,I232010,I232027,I232058,I232075,I232153,I232170,I232187,I232204,I232221,I232238,I232255,I232124,I232286,I232303,I232320,I232337,I232354,I232371,I232388,I232121,I232419,I232115,I232450,I232467,I232484,I232145,I232118,I232529,I232142,I232560,I232139,I232136,I232605,I232622,I232639,I232656,I232673,I232130,I232704,I232721,I232133,I232127,I232799,I232816,I232833,I232850,I232867,I232898,I232915,I232932,I232949,I232966,I232983,I233014,I233045,I233062,I233079,I233096,I233141,I233158,I233175,I233206,I233251,I233268,I233285,I233330,I233347,I233411,I233428,I233445,I233462,I233479,I233510,I233527,I233544,I233561,I233578,I233595,I233626,I233657,I233674,I233691,I233708,I233753,I233770,I233787,I233818,I233863,I233880,I233897,I233942,I233959,I234023,I234040,I344574,I344577,I234057,I344583,I234074,I344580,I344556,I234091,I234122,I234139,I344559,I234156,I234173,I344568,I344553,I234190,I234207,I234238,I234269,I344571,I234286,I344565,I234303,I234320,I234365,I234382,I234399,I234430,I234475,I344562,I234492,I234509,I234554,I234571,I234635,I234652,I234669,I234686,I234703,I234734,I234751,I234768,I234785,I234802,I234819,I234850,I234881,I234898,I234915,I234932,I234977,I234994,I235011,I235042,I235087,I235104,I235121,I235166,I235183,I235247,I235264,I235281,I235298,I235315,I235346,I235363,I235380,I235397,I235414,I235431,I235462,I235493,I235510,I235527,I235544,I235589,I235606,I235623,I235654,I235699,I235716,I235733,I235778,I235795,I235859,I235876,I235893,I235910,I235927,I235821,I235958,I235975,I235992,I236009,I236026,I236043,I235830,I236074,I235824,I236105,I236122,I236139,I236156,I235851,I235848,I236201,I236218,I236235,I235845,I236266,I235842,I235833,I236311,I236328,I236345,I235836,I235839,I236390,I236407,I235827,I236471,I236488,I236505,I236522,I236539,I236570,I236587,I236604,I236621,I236638,I236655,I236686,I236717,I236734,I236751,I236768,I236813,I236830,I236847,I236878,I236923,I236940,I236957,I237002,I237019,I237083,I237100,I237117,I237134,I237151,I237182,I237199,I237216,I237233,I237250,I237267,I237298,I237329,I237346,I237363,I237380,I237425,I237442,I237459,I237490,I237535,I237552,I237569,I237614,I237631,I237695,I237712,I237729,I237746,I237763,I237794,I237811,I237828,I237845,I237862,I237879,I237910,I237941,I237958,I237975,I237992,I238037,I238054,I238071,I238102,I238147,I238164,I238181,I238226,I238243,I238307,I238324,I238341,I238358,I238375,I238269,I238406,I238423,I238440,I238457,I238474,I238491,I238278,I238522,I238272,I238553,I238570,I238587,I238604,I238299,I238296,I238649,I238666,I238683,I238293,I238714,I238290,I238281,I238759,I238776,I238793,I238284,I238287,I238838,I238855,I238275,I238919,I238936,I238953,I238970,I238987,I238887,I239018,I239035,I239052,I238890,I239083,I238884,I239114,I239131,I239148,I239165,I239182,I238893,I239213,I239230,I239247,I239264,I238899,I238902,I238881,I239323,I239340,I239357,I238911,I238908,I239402,I239419,I238896,I238905,I239497,I239514,I354006,I354009,I239531,I354015,I239548,I239565,I239596,I354012,I239613,I353991,I239630,I239661,I239692,I353988,I354003,I239709,I354000,I239726,I239743,I239760,I239791,I354018,I239808,I353997,I239825,I239842,I239901,I353994,I239918,I239935,I239980,I239997,I240075,I240092,I240109,I240126,I240143,I240043,I240174,I240191,I240208,I240046,I240239,I240040,I240270,I240287,I240304,I240321,I240338,I240049,I240369,I240386,I240403,I240420,I240055,I240058,I240037,I240479,I240496,I240513,I240067,I240064,I240558,I240575,I240052,I240061,I240653,I240670,I359038,I359041,I240687,I359047,I240704,I240721,I240752,I359044,I240769,I359023,I240786,I240817,I240848,I359020,I359035,I240865,I359032,I240882,I240899,I240916,I240947,I359050,I240964,I359029,I240981,I240998,I241057,I359026,I241074,I241091,I241136,I241153,I241231,I241248,I241265,I241282,I241299,I241330,I241347,I241364,I241395,I241426,I241443,I241460,I241477,I241494,I241525,I241542,I241559,I241576,I241635,I241652,I241669,I241714,I241731,I241809,I241826,I302879,I302867,I241843,I302861,I241860,I241877,I241908,I302858,I241925,I302852,I241942,I241973,I242004,I302855,I302870,I242021,I302882,I242038,I242055,I242072,I242103,I302873,I242120,I302864,I242137,I242154,I242213,I302876,I242230,I242247,I242292,I242309,I242387,I242404,I242421,I242438,I242455,I242355,I242486,I242503,I242520,I242358,I242551,I242352,I242582,I242599,I242616,I242633,I242650,I242361,I242681,I242698,I242715,I242732,I242367,I242370,I242349,I242791,I242808,I242825,I242379,I242376,I242870,I242887,I242364,I242373,I242965,I242982,I242999,I243016,I243033,I243064,I243081,I243098,I243129,I243160,I243177,I243194,I243211,I243228,I243259,I243276,I243293,I243310,I243369,I243386,I243403,I243448,I243465,I243543,I243560,I327256,I327253,I243577,I327247,I243594,I243611,I243511,I243642,I327268,I243659,I327271,I243676,I243514,I243707,I243508,I243738,I327274,I327265,I243755,I327277,I243772,I243789,I243806,I243517,I243837,I327250,I243854,I327259,I243871,I243888,I243523,I243526,I243505,I243947,I327262,I243964,I243981,I243535,I243532,I244026,I244043,I243520,I243529,I244121,I244138,I244155,I244172,I244189,I244220,I244237,I244254,I244285,I244316,I244333,I244350,I244367,I244384,I244415,I244432,I244449,I244466,I244525,I244542,I244559,I244604,I244621,I244699,I244716,I280864,I280852,I244733,I280846,I244750,I244767,I244798,I280843,I244815,I280837,I244832,I244863,I244894,I280840,I280855,I244911,I280867,I244928,I244945,I244962,I244993,I280858,I245010,I280849,I245027,I245044,I245103,I280861,I245120,I245137,I245182,I245199,I245277,I245294,I245311,I245328,I245345,I245376,I245393,I245410,I245441,I245472,I245489,I245506,I245523,I245540,I245571,I245588,I245605,I245622,I245681,I245698,I245715,I245760,I245777,I245855,I245872,I245889,I245906,I245923,I245954,I245971,I245988,I246019,I246050,I246067,I246084,I246101,I246118,I246149,I246166,I246183,I246200,I246259,I246276,I246293,I246338,I246355,I246433,I246450,I246467,I246484,I246501,I246401,I246532,I246549,I246566,I246404,I246597,I246398,I246628,I246645,I246662,I246679,I246696,I246407,I246727,I246744,I246761,I246778,I246413,I246416,I246395,I246837,I246854,I246871,I246425,I246422,I246916,I246933,I246410,I246419,I247011,I247028,I325471,I325468,I247045,I325462,I247062,I247079,I247110,I325483,I247127,I325486,I247144,I247175,I247206,I325489,I325480,I247223,I325492,I247240,I247257,I247274,I247305,I325465,I247322,I325474,I247339,I247356,I247415,I325477,I247432,I247449,I247494,I247511,I247589,I247606,I247623,I247640,I247657,I247688,I247705,I247722,I247753,I247784,I247801,I247818,I247835,I247852,I247883,I247900,I247917,I247934,I247993,I248010,I248027,I248072,I248089,I248167,I248184,I248201,I248218,I248235,I248266,I248283,I248300,I248331,I248362,I248379,I248396,I248413,I248430,I248461,I248478,I248495,I248512,I248571,I248588,I248605,I248650,I248667,I248745,I248762,I394922,I394934,I248779,I394907,I248796,I248813,I248844,I394925,I248861,I394916,I248878,I248909,I248940,I394913,I394919,I248957,I394931,I248974,I248991,I249008,I249039,I394937,I249056,I394928,I249073,I249090,I249149,I394910,I249166,I249183,I249228,I249245,I249323,I249340,I249357,I249374,I249391,I249422,I249439,I249456,I249487,I249518,I249535,I249552,I249569,I249586,I249617,I249634,I249651,I249668,I249727,I249744,I249761,I249806,I249823,I249901,I249918,I249935,I249952,I249969,I250000,I250017,I250034,I250065,I250096,I250113,I250130,I250147,I250164,I250195,I250212,I250229,I250246,I250305,I250322,I250339,I250384,I250401,I250479,I250496,I250513,I250530,I250547,I250447,I250578,I250595,I250612,I250450,I250643,I250444,I250674,I250691,I250708,I250725,I250742,I250453,I250773,I250790,I250807,I250824,I250459,I250462,I250441,I250883,I250900,I250917,I250471,I250468,I250962,I250979,I250456,I250465,I251057,I251074,I340797,I340800,I251091,I340806,I251108,I251125,I251156,I340803,I251173,I340782,I251190,I251221,I251252,I340779,I340794,I251269,I340791,I251286,I251303,I251320,I251351,I340809,I251368,I340788,I251385,I251402,I251461,I340785,I251478,I251495,I251540,I251557,I251635,I251652,I329636,I329633,I251669,I329627,I251686,I251703,I251734,I329648,I251751,I329651,I251768,I251799,I251830,I329654,I329645,I251847,I329657,I251864,I251881,I251898,I251929,I329630,I251946,I329639,I251963,I251980,I252039,I329642,I252056,I252073,I252118,I252135,I252213,I252230,I252247,I252264,I252281,I252312,I252329,I252346,I252377,I252408,I252425,I252442,I252459,I252476,I252507,I252524,I252541,I252558,I252617,I252634,I252651,I252696,I252713,I252791,I252808,I252825,I252842,I252859,I252890,I252907,I252924,I252955,I252986,I253003,I253020,I253037,I253054,I253085,I253102,I253119,I253136,I253195,I253212,I253229,I253274,I253291,I253369,I253386,I253403,I253420,I253437,I253468,I253485,I253502,I253533,I253564,I253581,I253598,I253615,I253632,I253663,I253680,I253697,I253714,I253773,I253790,I253807,I253852,I253869,I253947,I253964,I253981,I253998,I254015,I254046,I254063,I254080,I254111,I254142,I254159,I254176,I254193,I254210,I254241,I254258,I254275,I254292,I254351,I254368,I254385,I254430,I254447,I254525,I254542,I254559,I254576,I254593,I254624,I254641,I254658,I254689,I254720,I254737,I254754,I254771,I254788,I254819,I254836,I254853,I254870,I254929,I254946,I254963,I255008,I255025,I255103,I255120,I255137,I255154,I255171,I255202,I255219,I255236,I255267,I255298,I255315,I255332,I255349,I255366,I255397,I255414,I255431,I255448,I255507,I255524,I255541,I255586,I255603,I255681,I255698,I255715,I255732,I255749,I255780,I255797,I255814,I255845,I255876,I255893,I255910,I255927,I255944,I255975,I255992,I256009,I256026,I256085,I256102,I256119,I256164,I256181,I256259,I256276,I256293,I256310,I256327,I256358,I256375,I256392,I256423,I256454,I256471,I256488,I256505,I256522,I256553,I256570,I256587,I256604,I256663,I256680,I256697,I256742,I256759,I256837,I256854,I311209,I311197,I256871,I311191,I256888,I256905,I256936,I311188,I256953,I311182,I256970,I257001,I257032,I311185,I311200,I257049,I311212,I257066,I257083,I257100,I257131,I311203,I257148,I311194,I257165,I257182,I257241,I311206,I257258,I257275,I257320,I257337,I257415,I257432,I257449,I257466,I257483,I257514,I257531,I257548,I257579,I257610,I257627,I257644,I257661,I257678,I257709,I257726,I257743,I257760,I257819,I257836,I257853,I257898,I257915,I257993,I258010,I258027,I258044,I258061,I257961,I258092,I258109,I258126,I257964,I258157,I257958,I258188,I258205,I258222,I258239,I258256,I257967,I258287,I258304,I258321,I258338,I257973,I257976,I257955,I258397,I258414,I258431,I257985,I257982,I258476,I258493,I257970,I257979,I258571,I258588,I258605,I258622,I258639,I258670,I258687,I258704,I258735,I258766,I258783,I258800,I258817,I258834,I258865,I258882,I258899,I258916,I258975,I258992,I259009,I259054,I259071,I259149,I259166,I283244,I283232,I259183,I283226,I259200,I259217,I259248,I283223,I259265,I283217,I259282,I259313,I259344,I283220,I283235,I259361,I283247,I259378,I259395,I259412,I259443,I283238,I259460,I283229,I259477,I259494,I259553,I283241,I259570,I259587,I259632,I259649,I259727,I259744,I293359,I293347,I259761,I293341,I259778,I259795,I259695,I259826,I293338,I259843,I293332,I259860,I259698,I259891,I259692,I259922,I293335,I293350,I259939,I293362,I259956,I259973,I259990,I259701,I260021,I293353,I260038,I293344,I260055,I260072,I259707,I259710,I259689,I260131,I293356,I260148,I260165,I259719,I259716,I260210,I260227,I259704,I259713,I260305,I260322,I260339,I260356,I260373,I260273,I260404,I260421,I260438,I260276,I260469,I260270,I260500,I260517,I260534,I260551,I260568,I260279,I260599,I260616,I260633,I260650,I260285,I260288,I260267,I260709,I260726,I260743,I260297,I260294,I260788,I260805,I260282,I260291,I260883,I260900,I260917,I260934,I260951,I260851,I260982,I260999,I261016,I260854,I261047,I260848,I261078,I261095,I261112,I261129,I261146,I260857,I261177,I261194,I261211,I261228,I260863,I260866,I260845,I261287,I261304,I261321,I260875,I260872,I261366,I261383,I260860,I260869,I261461,I261478,I261495,I261512,I261529,I261560,I261577,I261594,I261625,I261656,I261673,I261690,I261707,I261724,I261755,I261772,I261789,I261806,I261865,I261882,I261899,I261944,I261961,I262039,I262056,I262073,I262090,I262107,I262007,I262138,I262155,I262172,I262010,I262203,I262004,I262234,I262251,I262268,I262285,I262302,I262013,I262333,I262350,I262367,I262384,I262019,I262022,I262001,I262443,I262460,I262477,I262031,I262028,I262522,I262539,I262016,I262025,I262617,I262634,I262651,I262668,I262685,I262716,I262733,I262750,I262781,I262812,I262829,I262846,I262863,I262880,I262911,I262928,I262945,I262962,I263021,I263038,I263055,I263100,I263117,I263195,I263212,I263229,I263246,I263263,I263294,I263311,I263328,I263359,I263390,I263407,I263424,I263441,I263458,I263489,I263506,I263523,I263540,I263599,I263616,I263633,I263678,I263695,I263773,I263790,I263807,I263824,I263841,I263741,I263872,I263889,I263906,I263744,I263937,I263738,I263968,I263985,I264002,I264019,I264036,I263747,I264067,I264084,I264101,I264118,I263753,I263756,I263735,I264177,I264194,I264211,I263765,I263762,I264256,I264273,I263750,I263759,I264351,I264368,I264385,I264402,I264419,I264450,I264467,I264484,I264515,I264546,I264563,I264580,I264597,I264614,I264645,I264662,I264679,I264696,I264755,I264772,I264789,I264834,I264851,I264929,I264946,I264963,I264980,I264997,I265028,I265045,I265062,I265093,I265124,I265141,I265158,I265175,I265192,I265223,I265240,I265257,I265274,I265333,I265350,I265367,I265412,I265429,I265507,I265524,I387408,I387420,I265541,I387393,I265558,I265575,I265475,I265606,I387411,I265623,I387402,I265640,I265478,I265671,I265472,I265702,I387399,I387405,I265719,I387417,I265736,I265753,I265770,I265481,I265801,I387423,I265818,I387414,I265835,I265852,I265487,I265490,I265469,I265911,I387396,I265928,I265945,I265499,I265496,I265990,I266007,I265484,I265493,I266085,I266102,I266119,I266136,I266153,I266184,I266201,I266218,I266249,I266280,I266297,I266314,I266331,I266348,I266379,I266396,I266413,I266430,I266489,I266506,I266523,I266568,I266585,I266663,I266680,I266697,I266714,I266731,I266762,I266779,I266796,I266813,I266830,I266847,I266864,I266881,I266926,I266943,I266974,I266991,I267022,I267039,I267070,I267101,I267132,I267149,I267180,I267211,I267275,I267292,I267309,I267326,I267343,I267374,I267391,I267408,I267425,I267442,I267459,I267476,I267493,I267538,I267555,I267586,I267603,I267634,I267651,I267682,I267713,I267744,I267761,I267792,I267823,I267887,I267904,I337032,I337026,I267921,I337035,I267938,I337029,I337011,I267955,I267855,I267986,I268003,I268020,I337008,I268037,I268054,I337023,I337005,I268071,I268088,I268105,I267861,I267852,I268150,I268167,I267876,I268198,I268215,I267864,I268246,I337017,I268263,I337020,I267870,I268294,I267858,I268325,I267849,I268356,I337014,I268373,I267879,I268404,I267873,I268435,I267867,I268499,I268516,I297521,I297527,I268533,I297524,I268550,I297497,I297515,I268567,I268467,I268598,I268615,I268632,I297509,I268649,I268666,I297512,I297500,I268683,I268700,I268717,I268473,I268464,I268762,I268779,I268488,I268810,I268827,I268476,I268858,I297503,I268875,I297518,I268482,I268906,I268470,I268937,I268461,I268968,I297506,I268985,I268491,I269016,I268485,I269047,I268479,I269111,I269128,I388549,I388564,I269145,I388558,I269162,I388555,I388552,I269179,I269079,I269210,I269227,I269244,I388570,I269261,I269278,I388561,I388567,I269295,I269312,I269329,I269085,I269076,I269374,I269391,I269100,I269422,I269439,I269088,I269470,I388579,I269487,I388576,I269094,I269518,I269082,I269549,I269073,I269580,I388573,I269597,I269103,I269628,I269097,I269659,I269091,I269723,I269740,I300496,I300502,I269757,I300499,I269774,I300472,I300490,I269791,I269822,I269839,I269856,I300484,I269873,I269890,I300487,I300475,I269907,I269924,I269941,I269986,I270003,I270034,I270051,I270082,I300478,I270099,I300493,I270130,I270161,I270192,I300481,I270209,I270240,I270271,I270335,I270352,I270369,I270386,I270403,I270303,I270434,I270451,I270468,I270485,I270502,I270519,I270536,I270553,I270309,I270300,I270598,I270615,I270324,I270646,I270663,I270312,I270694,I270711,I270318,I270742,I270306,I270773,I270297,I270804,I270821,I270327,I270852,I270321,I270883,I270315,I270947,I270964,I270981,I270998,I271015,I271046,I271063,I271080,I271097,I271114,I271131,I271148,I271165,I271210,I271227,I271258,I271275,I271306,I271323,I271354,I271385,I271416,I271433,I271464,I271495,I271559,I271576,I287998,I287992,I271593,I287986,I271610,I288007,I287995,I271641,I271658,I287980,I271675,I271692,I271709,I287983,I287977,I271726,I271743,I271774,I271805,I271836,I288004,I271853,I288001,I271870,I271915,I271932,I271963,I287989,I271994,I272011,I272042,I272059,I272137,I272154,I272171,I272188,I272126,I272219,I272236,I272253,I272270,I272287,I272304,I272321,I272111,I272352,I272108,I272383,I272120,I272414,I272431,I272448,I272114,I272129,I272493,I272510,I272099,I272541,I272117,I272572,I272589,I272123,I272620,I272637,I272102,I272105,I272715,I272732,I272749,I272766,I272797,I272814,I272831,I272848,I272865,I272882,I272899,I272930,I272961,I272992,I273009,I273026,I273071,I273088,I273119,I273150,I273167,I273198,I273215,I273293,I273310,I337637,I337640,I273327,I337658,I273344,I337652,I337661,I273375,I273392,I337664,I273409,I273426,I273443,I337649,I337634,I273460,I273477,I273508,I273539,I273570,I337646,I273587,I337655,I273604,I273649,I273666,I273697,I337643,I273728,I273745,I273776,I273793,I273871,I273888,I273905,I273922,I273953,I273970,I273987,I274004,I274021,I274038,I274055,I274086,I274117,I274148,I274165,I274182,I274227,I274244,I274275,I274306,I274323,I274354,I274371,I274449,I274466,I274483,I274500,I274438,I274531,I274548,I274565,I274582,I274599,I274616,I274633,I274423,I274664,I274420,I274695,I274432,I274726,I274743,I274760,I274426,I274441,I274805,I274822,I274411,I274853,I274429,I274884,I274901,I274435,I274932,I274949,I274414,I274417,I275027,I275044,I357136,I357139,I275061,I357157,I275078,I357151,I357160,I275109,I275126,I357163,I275143,I275160,I275177,I357148,I357133,I275194,I275211,I275242,I275273,I275304,I357145,I275321,I357154,I275338,I275383,I275400,I275431,I357142,I275462,I275479,I275510,I275527,I275605,I275622,I275639,I275656,I275594,I275687,I275704,I275721,I275738,I275755,I275772,I275789,I275579,I275820,I275576,I275851,I275588,I275882,I275899,I275916,I275582,I275597,I275961,I275978,I275567,I276009,I275585,I276040,I276057,I275591,I276088,I276105,I275570,I275573,I276183,I276200,I386249,I386240,I276217,I386255,I276234,I386246,I386243,I276172,I276265,I276282,I386237,I276299,I276316,I276333,I386258,I386264,I276350,I276367,I276157,I276398,I276154,I276429,I276166,I276460,I386252,I276477,I386261,I276494,I276160,I276175,I276539,I276556,I276145,I276587,I386267,I276163,I276618,I276635,I276169,I276666,I276683,I276148,I276151,I276761,I276778,I350217,I350220,I276795,I350238,I276812,I350232,I350241,I276843,I276860,I350244,I276877,I276894,I276911,I350229,I350214,I276928,I276945,I276976,I277007,I277038,I350226,I277055,I350235,I277072,I277117,I277134,I277165,I350223,I277196,I277213,I277244,I277261,I277339,I277356,I347072,I347075,I277373,I347093,I277390,I347087,I347096,I277421,I277438,I347099,I277455,I277472,I277489,I347084,I347069,I277506,I277523,I277554,I277585,I277616,I347081,I277633,I347090,I277650,I277695,I277712,I277743,I347078,I277774,I277791,I277822,I277839,I277917,I277934,I277951,I277968,I277999,I278016,I278033,I278050,I278067,I278084,I278101,I278132,I278163,I278194,I278211,I278228,I278273,I278290,I278321,I278352,I278369,I278400,I278417,I278495,I278512,I278529,I278546,I278563,I278580,I278611,I278628,I278645,I278690,I278707,I278724,I278769,I278786,I278803,I278834,I278851,I278882,I278899,I278916,I278947,I278964,I278981,I278998,I279090,I279107,I375392,I375383,I279124,I375401,I279141,I279158,I375398,I279175,I279073,I279206,I375380,I279223,I279240,I279076,I279058,I279285,I375389,I375404,I279302,I375395,I279319,I279079,I279070,I279364,I375377,I279381,I375386,I279398,I279061,I279429,I279446,I279052,I279477,I375374,I279494,I279511,I279082,I279542,I279559,I279576,I279593,I279067,I279064,I279055,I279685,I279702,I279719,I279736,I279753,I279770,I279801,I279818,I279835,I279880,I279897,I279914,I279959,I279976,I279993,I280024,I280041,I280072,I280089,I280106,I280137,I280154,I280171,I280188,I280280,I280297,I280314,I280331,I280348,I280365,I280396,I280413,I280430,I280475,I280492,I280509,I280554,I280571,I280588,I280619,I280636,I280667,I280684,I280701,I280732,I280749,I280766,I280783,I280875,I280892,I280909,I280926,I280943,I280960,I280991,I281008,I281025,I281070,I281087,I281104,I281149,I281166,I281183,I281214,I281231,I281262,I281279,I281296,I281327,I281344,I281361,I281378,I281470,I281487,I281504,I281521,I281538,I281555,I281453,I281586,I281603,I281620,I281456,I281438,I281665,I281682,I281699,I281459,I281450,I281744,I281761,I281778,I281441,I281809,I281826,I281432,I281857,I281874,I281891,I281462,I281922,I281939,I281956,I281973,I281447,I281444,I281435,I282065,I282082,I282099,I282116,I282133,I282150,I282048,I282181,I282198,I282215,I282051,I282033,I282260,I282277,I282294,I282054,I282045,I282339,I282356,I282373,I282036,I282404,I282421,I282027,I282452,I282469,I282486,I282057,I282517,I282534,I282551,I282568,I282042,I282039,I282030,I282660,I282677,I282694,I282711,I282728,I282745,I282643,I282776,I282793,I282810,I282646,I282628,I282855,I282872,I282889,I282649,I282640,I282934,I282951,I282968,I282631,I282999,I283016,I282622,I283047,I283064,I283081,I282652,I283112,I283129,I283146,I283163,I282637,I282634,I282625,I283255,I283272,I283289,I283306,I283323,I283340,I283371,I283388,I283405,I283450,I283467,I283484,I283529,I283546,I283563,I283594,I283611,I283642,I283659,I283676,I283707,I283724,I283741,I283758,I283850,I283867,I394341,I394347,I283884,I394338,I283901,I283918,I394350,I283935,I283966,I394329,I283983,I284000,I284045,I394353,I394335,I284062,I394344,I284079,I284124,I394359,I284141,I394332,I284158,I284189,I284206,I284237,I394356,I284254,I284271,I284302,I284319,I284336,I284353,I284445,I284462,I284479,I284496,I284513,I284530,I284428,I284561,I284578,I284595,I284431,I284413,I284640,I284657,I284674,I284434,I284425,I284719,I284736,I284753,I284416,I284784,I284801,I284407,I284832,I284849,I284866,I284437,I284897,I284914,I284931,I284948,I284422,I284419,I284410,I285040,I285057,I285074,I285091,I285108,I285125,I285023,I285156,I285173,I285190,I285026,I285008,I285235,I285252,I285269,I285029,I285020,I285314,I285331,I285348,I285011,I285379,I285396,I285002,I285427,I285444,I285461,I285032,I285492,I285509,I285526,I285543,I285017,I285014,I285005,I285635,I285652,I285669,I285686,I285703,I285720,I285751,I285768,I285785,I285830,I285847,I285864,I285909,I285926,I285943,I285974,I285991,I286022,I286039,I286056,I286087,I286104,I286121,I286138,I286230,I286247,I286264,I286281,I286298,I286315,I286346,I286363,I286380,I286425,I286442,I286459,I286504,I286521,I286538,I286569,I286586,I286617,I286634,I286651,I286682,I286699,I286716,I286733,I286825,I286842,I286859,I286876,I286893,I286910,I286808,I286941,I286958,I286975,I286811,I286793,I287020,I287037,I287054,I286814,I286805,I287099,I287116,I287133,I286796,I287164,I287181,I286787,I287212,I287229,I287246,I286817,I287277,I287294,I287311,I287328,I286802,I286799,I286790,I287420,I287437,I341426,I341417,I287454,I341435,I287471,I287488,I341432,I287505,I287536,I341414,I287553,I287570,I287615,I341423,I341438,I287632,I341429,I287649,I287694,I341411,I287711,I341420,I287728,I287759,I287776,I287807,I341408,I287824,I287841,I287872,I287889,I287906,I287923,I288015,I288032,I288049,I288066,I288083,I288100,I288131,I288148,I288165,I288210,I288227,I288244,I288289,I288306,I288323,I288354,I288371,I288402,I288419,I288436,I288467,I288484,I288501,I288518,I288610,I288627,I288644,I288661,I288678,I288695,I288726,I288743,I288760,I288805,I288822,I288839,I288884,I288901,I288918,I288949,I288966,I288997,I289014,I289031,I289062,I289079,I289096,I289113,I289205,I289222,I318932,I318923,I289239,I318941,I289256,I289273,I318920,I289290,I289188,I289321,I318929,I289338,I289355,I289191,I289173,I289400,I318944,I318926,I289417,I318947,I289434,I289194,I289185,I289479,I318935,I289496,I318917,I289513,I289176,I289544,I289561,I289167,I289592,I318938,I289609,I289626,I289197,I289657,I289674,I289691,I289708,I289182,I289179,I289170,I289800,I289817,I322502,I322493,I289834,I322511,I289851,I289868,I322490,I289885,I289916,I322499,I289933,I289950,I289995,I322514,I322496,I290012,I322517,I290029,I290074,I322505,I290091,I322487,I290108,I290139,I290156,I290187,I322508,I290204,I290221,I290252,I290269,I290286,I290303,I290395,I290412,I290429,I290446,I290463,I290480,I290511,I290528,I290545,I290590,I290607,I290624,I290669,I290686,I290703,I290734,I290751,I290782,I290799,I290816,I290847,I290864,I290881,I290898,I290990,I291007,I291024,I291041,I291058,I291075,I291106,I291123,I291140,I291185,I291202,I291219,I291264,I291281,I291298,I291329,I291346,I291377,I291394,I291411,I291442,I291459,I291476,I291493,I291585,I291602,I372876,I372867,I291619,I372885,I291636,I291653,I372882,I291670,I291701,I372864,I291718,I291735,I291780,I372873,I372888,I291797,I372879,I291814,I291859,I372861,I291876,I372870,I291893,I291924,I291941,I291972,I372858,I291989,I292006,I292037,I292054,I292071,I292088,I292180,I292197,I292214,I292231,I292248,I292265,I292296,I292313,I292330,I292375,I292392,I292409,I292454,I292471,I292488,I292519,I292536,I292567,I292584,I292601,I292632,I292649,I292666,I292683,I292775,I292792,I292809,I292826,I292843,I292860,I292891,I292908,I292925,I292970,I292987,I293004,I293049,I293066,I293083,I293114,I293131,I293162,I293179,I293196,I293227,I293244,I293261,I293278,I293370,I293387,I374763,I374754,I293404,I374772,I293421,I293438,I374769,I293455,I293486,I374751,I293503,I293520,I293565,I374760,I374775,I293582,I374766,I293599,I293644,I374748,I293661,I374757,I293678,I293709,I293726,I293757,I374745,I293774,I293791,I293822,I293839,I293856,I293873,I293965,I293982,I391451,I391457,I293999,I391448,I294016,I294033,I391460,I294050,I293948,I294081,I391439,I294098,I294115,I293951,I293933,I294160,I391463,I391445,I294177,I391454,I294194,I293954,I293945,I294239,I391469,I294256,I391442,I294273,I293936,I294304,I294321,I293927,I294352,I391466,I294369,I294386,I293957,I294417,I294434,I294451,I294468,I293942,I293939,I293930,I294560,I294577,I335765,I335756,I294594,I335774,I294611,I294628,I335771,I294645,I294676,I335753,I294693,I294710,I294755,I335762,I335777,I294772,I335768,I294789,I294834,I335750,I294851,I335759,I294868,I294899,I294916,I294947,I335747,I294964,I294981,I295012,I295029,I295046,I295063,I295155,I295172,I331427,I331418,I295189,I331436,I295206,I295223,I331415,I295240,I295271,I331424,I295288,I295305,I295350,I331439,I331421,I295367,I331442,I295384,I295429,I331430,I295446,I331412,I295463,I295494,I295511,I295542,I331433,I295559,I295576,I295607,I295624,I295641,I295658,I295750,I295767,I295784,I295801,I295818,I295835,I295866,I295883,I295900,I295945,I295962,I295979,I296024,I296041,I296058,I296089,I296106,I296137,I296154,I296171,I296202,I296219,I296236,I296253,I296345,I296362,I296379,I296396,I296413,I296430,I296328,I296461,I296478,I296495,I296331,I296313,I296540,I296557,I296574,I296334,I296325,I296619,I296636,I296653,I296316,I296684,I296701,I296307,I296732,I296749,I296766,I296337,I296797,I296814,I296831,I296848,I296322,I296319,I296310,I296940,I296957,I296974,I296991,I297008,I297025,I297056,I297073,I297090,I297135,I297152,I297169,I297214,I297231,I297248,I297279,I297296,I297327,I297344,I297361,I297392,I297409,I297426,I297443,I297535,I297552,I297569,I297586,I297603,I297620,I297651,I297668,I297685,I297730,I297747,I297764,I297809,I297826,I297843,I297874,I297891,I297922,I297939,I297956,I297987,I298004,I298021,I298038,I298130,I298147,I298164,I298181,I298198,I298215,I298113,I298246,I298263,I298280,I298116,I298098,I298325,I298342,I298359,I298119,I298110,I298404,I298421,I298438,I298101,I298469,I298486,I298092,I298517,I298534,I298551,I298122,I298582,I298599,I298616,I298633,I298107,I298104,I298095,I298725,I298742,I298759,I298776,I298793,I298810,I298841,I298858,I298875,I298920,I298937,I298954,I298999,I299016,I299033,I299064,I299081,I299112,I299129,I299146,I299177,I299194,I299211,I299228,I299320,I299337,I299354,I299371,I299388,I299405,I299436,I299453,I299470,I299515,I299532,I299549,I299594,I299611,I299628,I299659,I299676,I299707,I299724,I299741,I299772,I299789,I299806,I299823,I299915,I299932,I299949,I299966,I299983,I300000,I299898,I300031,I300048,I300065,I299901,I299883,I300110,I300127,I300144,I299904,I299895,I300189,I300206,I300223,I299886,I300254,I300271,I299877,I300302,I300319,I300336,I299907,I300367,I300384,I300401,I300418,I299892,I299889,I299880,I300510,I300527,I370360,I370351,I300544,I370369,I300561,I300578,I370366,I300595,I300626,I370348,I300643,I300660,I300705,I370357,I370372,I300722,I370363,I300739,I300784,I370345,I300801,I370354,I300818,I300849,I300866,I300897,I370342,I300914,I300931,I300962,I300979,I300996,I301013,I301105,I301122,I378537,I378528,I301139,I378546,I301156,I301173,I378543,I301190,I301221,I378525,I301238,I301255,I301300,I378534,I378549,I301317,I378540,I301334,I301379,I378522,I301396,I378531,I301413,I301444,I301461,I301492,I378519,I301509,I301526,I301557,I301574,I301591,I301608,I301700,I301717,I301734,I301751,I301768,I301785,I301816,I301833,I301850,I301895,I301912,I301929,I301974,I301991,I302008,I302039,I302056,I302087,I302104,I302121,I302152,I302169,I302186,I302203,I302295,I302312,I302329,I302346,I302363,I302380,I302411,I302428,I302445,I302490,I302507,I302524,I302569,I302586,I302603,I302634,I302651,I302682,I302699,I302716,I302747,I302764,I302781,I302798,I302890,I302907,I302924,I302941,I302958,I302975,I303006,I303023,I303040,I303085,I303102,I303119,I303164,I303181,I303198,I303229,I303246,I303277,I303294,I303311,I303342,I303359,I303376,I303393,I303485,I303502,I303519,I303536,I303553,I303570,I303468,I303601,I303618,I303635,I303471,I303453,I303680,I303697,I303714,I303474,I303465,I303759,I303776,I303793,I303456,I303824,I303841,I303447,I303872,I303889,I303906,I303477,I303937,I303954,I303971,I303988,I303462,I303459,I303450,I304080,I304097,I304114,I304131,I304148,I304165,I304063,I304196,I304213,I304230,I304066,I304048,I304275,I304292,I304309,I304069,I304060,I304354,I304371,I304388,I304051,I304419,I304436,I304042,I304467,I304484,I304501,I304072,I304532,I304549,I304566,I304583,I304057,I304054,I304045,I304675,I304692,I369731,I369722,I304709,I369740,I304726,I304743,I369737,I304760,I304791,I369719,I304808,I304825,I304870,I369728,I369743,I304887,I369734,I304904,I304949,I369716,I304966,I369725,I304983,I305014,I305031,I305062,I369713,I305079,I305096,I305127,I305144,I305161,I305178,I305270,I305287,I305304,I305321,I305338,I305355,I305386,I305403,I305420,I305465,I305482,I305499,I305544,I305561,I305578,I305609,I305626,I305657,I305674,I305691,I305722,I305739,I305756,I305773,I305865,I305882,I305899,I305916,I305933,I305950,I305981,I305998,I306015,I306060,I306077,I306094,I306139,I306156,I306173,I306204,I306221,I306252,I306269,I306286,I306317,I306334,I306351,I306368,I306460,I306477,I306494,I306511,I306528,I306545,I306576,I306593,I306610,I306655,I306672,I306689,I306734,I306751,I306768,I306799,I306816,I306847,I306864,I306881,I306912,I306929,I306946,I306963,I307055,I307072,I339539,I339530,I307089,I339548,I307106,I307123,I339545,I307140,I307038,I307171,I339527,I307188,I307205,I307041,I307023,I307250,I339536,I339551,I307267,I339542,I307284,I307044,I307035,I307329,I339524,I307346,I339533,I307363,I307026,I307394,I307411,I307017,I307442,I339521,I307459,I307476,I307047,I307507,I307524,I307541,I307558,I307032,I307029,I307020,I307650,I307667,I307684,I307701,I307718,I307735,I307633,I307766,I307783,I307800,I307636,I307618,I307845,I307862,I307879,I307639,I307630,I307924,I307941,I307958,I307621,I307989,I308006,I307612,I308037,I308054,I308071,I307642,I308102,I308119,I308136,I308153,I307627,I307624,I307615,I308245,I308262,I308279,I308296,I308313,I308330,I308361,I308378,I308395,I308440,I308457,I308474,I308519,I308536,I308553,I308584,I308601,I308632,I308649,I308666,I308697,I308714,I308731,I308748,I308840,I308857,I308874,I308891,I308908,I308925,I308956,I308973,I308990,I309035,I309052,I309069,I309114,I309131,I309148,I309179,I309196,I309227,I309244,I309261,I309292,I309309,I309326,I309343,I309435,I309452,I309469,I309486,I309503,I309520,I309418,I309551,I309568,I309585,I309421,I309403,I309630,I309647,I309664,I309424,I309415,I309709,I309726,I309743,I309406,I309774,I309791,I309397,I309822,I309839,I309856,I309427,I309887,I309904,I309921,I309938,I309412,I309409,I309400,I310030,I310047,I310064,I310081,I310098,I310115,I310146,I310163,I310180,I310225,I310242,I310259,I310304,I310321,I310338,I310369,I310386,I310417,I310434,I310451,I310482,I310499,I310516,I310533,I310625,I310642,I310659,I310676,I310693,I310710,I310741,I310758,I310775,I310820,I310837,I310854,I310899,I310916,I310933,I310964,I310981,I311012,I311029,I311046,I311077,I311094,I311111,I311128,I311220,I311237,I311254,I311271,I311288,I311305,I311336,I311353,I311370,I311415,I311432,I311449,I311494,I311511,I311528,I311559,I311576,I311607,I311624,I311641,I311672,I311689,I311706,I311723,I311815,I311832,I330832,I330823,I311849,I330841,I311866,I311883,I330820,I311900,I311931,I330829,I311948,I311965,I312010,I330844,I330826,I312027,I330847,I312044,I312089,I330835,I312106,I330817,I312123,I312154,I312171,I312202,I330838,I312219,I312236,I312267,I312284,I312301,I312318,I312410,I312427,I312444,I312461,I312478,I312495,I312526,I312543,I312560,I312605,I312622,I312639,I312684,I312701,I312718,I312749,I312766,I312797,I312814,I312831,I312862,I312879,I312896,I312913,I313005,I313022,I313039,I313056,I313073,I313090,I313121,I313138,I313155,I313200,I313217,I313234,I313279,I313296,I313313,I313344,I313361,I313392,I313409,I313426,I313457,I313474,I313491,I313508,I313600,I313617,I313634,I313651,I313668,I313685,I313702,I313733,I313750,I313767,I313784,I313801,I313818,I313835,I313880,I313897,I313914,I313945,I313962,I314007,I314038,I314055,I314086,I314131,I314195,I314212,I314229,I314246,I314263,I314280,I314297,I314328,I314345,I314362,I314379,I314396,I314413,I314430,I314475,I314492,I314509,I314540,I314557,I314602,I314633,I314650,I314681,I314726,I314790,I314807,I314824,I314841,I314858,I314875,I314892,I314761,I314923,I314940,I314957,I314974,I314991,I315008,I315025,I314758,I314752,I315070,I315087,I315104,I314779,I315135,I315152,I314770,I314764,I315197,I314767,I315228,I315245,I314782,I315276,I314776,I314773,I315321,I314755,I315385,I315402,I315419,I315436,I315453,I315470,I315487,I315518,I315535,I315552,I315569,I315586,I315603,I315620,I315665,I315682,I315699,I315730,I315747,I315792,I315823,I315840,I315871,I315916,I315980,I315997,I367856,I367844,I316014,I367829,I316031,I316048,I367841,I316065,I367853,I316082,I315951,I316113,I367826,I367850,I316130,I367835,I316147,I316164,I316181,I316198,I316215,I315948,I315942,I316260,I367838,I316277,I367847,I316294,I315969,I316325,I316342,I315960,I315954,I316387,I315957,I316418,I367832,I316435,I315972,I316466,I315966,I315963,I316511,I315945,I316575,I316592,I316609,I316626,I316643,I316660,I316677,I316708,I316725,I316742,I316759,I316776,I316793,I316810,I316855,I316872,I316889,I316920,I316937,I316982,I317013,I317030,I317061,I317106,I317170,I317187,I317204,I317221,I317238,I317255,I317272,I317303,I317320,I317337,I317354,I317371,I317388,I317405,I317450,I317467,I317484,I317515,I317532,I317577,I317608,I317625,I317656,I317701,I317765,I317782,I317799,I317816,I317833,I317850,I317867,I317898,I317915,I317932,I317949,I317966,I317983,I318000,I318045,I318062,I318079,I318110,I318127,I318172,I318203,I318220,I318251,I318296,I318360,I318377,I318394,I318411,I318428,I318445,I318462,I318493,I318510,I318527,I318544,I318561,I318578,I318595,I318640,I318657,I318674,I318705,I318722,I318767,I318798,I318815,I318846,I318891,I318955,I318972,I397219,I397222,I318989,I397231,I319006,I319023,I397225,I319040,I397246,I319057,I319088,I397243,I397249,I319105,I397234,I319122,I319139,I319156,I319173,I319190,I319235,I397237,I319252,I397240,I319269,I319300,I319317,I319362,I319393,I397228,I319410,I319441,I319486,I319550,I319567,I319584,I319601,I319618,I319635,I319652,I319683,I319700,I319717,I319734,I319751,I319768,I319785,I319830,I319847,I319864,I319895,I319912,I319957,I319988,I320005,I320036,I320081,I320145,I320162,I320179,I320196,I320213,I320230,I320247,I320278,I320295,I320312,I320329,I320346,I320363,I320380,I320425,I320442,I320459,I320490,I320507,I320552,I320583,I320600,I320631,I320676,I320740,I320757,I320774,I320791,I320808,I320825,I320842,I320873,I320890,I320907,I320924,I320941,I320958,I320975,I321020,I321037,I321054,I321085,I321102,I321147,I321178,I321195,I321226,I321271,I321335,I321352,I321369,I321386,I321403,I321420,I321437,I321468,I321485,I321502,I321519,I321536,I321553,I321570,I321615,I321632,I321649,I321680,I321697,I321742,I321773,I321790,I321821,I321866,I321930,I321947,I321964,I321981,I321998,I322015,I322032,I322063,I322080,I322097,I322114,I322131,I322148,I322165,I322210,I322227,I322244,I322275,I322292,I322337,I322368,I322385,I322416,I322461,I322525,I322542,I386815,I386818,I322559,I386827,I322576,I322593,I386821,I322610,I386842,I322627,I322658,I386839,I386845,I322675,I386830,I322692,I322709,I322726,I322743,I322760,I322805,I386833,I322822,I386836,I322839,I322870,I322887,I322932,I322963,I386824,I322980,I323011,I323056,I323120,I323137,I323154,I323171,I323188,I323205,I323222,I323253,I323270,I323287,I323304,I323321,I323338,I323355,I323400,I323417,I323434,I323465,I323482,I323527,I323558,I323575,I323606,I323651,I323715,I323732,I334519,I334507,I323749,I334492,I323766,I323783,I334504,I323800,I334516,I323817,I323848,I334489,I334513,I323865,I334498,I323882,I323899,I323916,I323933,I323950,I323995,I334501,I324012,I334510,I324029,I324060,I324077,I324122,I324153,I334495,I324170,I324201,I324246,I324310,I324327,I324344,I324361,I324378,I324395,I324412,I324443,I324460,I324477,I324494,I324511,I324528,I324545,I324590,I324607,I324624,I324655,I324672,I324717,I324748,I324765,I324796,I324841,I324905,I324922,I324939,I324956,I324973,I324990,I325007,I325038,I325055,I325072,I325089,I325106,I325123,I325140,I325185,I325202,I325219,I325250,I325267,I325312,I325343,I325360,I325391,I325436,I325500,I325517,I325534,I325551,I325568,I325585,I325602,I325633,I325650,I325667,I325684,I325701,I325718,I325735,I325780,I325797,I325814,I325845,I325862,I325907,I325938,I325955,I325986,I326031,I326095,I326112,I349615,I349603,I326129,I349588,I326146,I326163,I349600,I326180,I349612,I326197,I326228,I349585,I349609,I326245,I349594,I326262,I326279,I326296,I326313,I326330,I326375,I349597,I326392,I349606,I326409,I326440,I326457,I326502,I326533,I349591,I326550,I326581,I326626,I326690,I326707,I326724,I326741,I326758,I326775,I326792,I326823,I326840,I326857,I326874,I326891,I326908,I326925,I326970,I326987,I327004,I327035,I327052,I327097,I327128,I327145,I327176,I327221,I327285,I327302,I327319,I327336,I327353,I327370,I327387,I327418,I327435,I327452,I327469,I327486,I327503,I327520,I327565,I327582,I327599,I327630,I327647,I327692,I327723,I327740,I327771,I327816,I327880,I327897,I327914,I327931,I327948,I327965,I327982,I328013,I328030,I328047,I328064,I328081,I328098,I328115,I328160,I328177,I328194,I328225,I328242,I328287,I328318,I328335,I328366,I328411,I328475,I328492,I328509,I328526,I328543,I328560,I328577,I328608,I328625,I328642,I328659,I328676,I328693,I328710,I328755,I328772,I328789,I328820,I328837,I328882,I328913,I328930,I328961,I329006,I329070,I329087,I329104,I329121,I329138,I329155,I329172,I329203,I329220,I329237,I329254,I329271,I329288,I329305,I329350,I329367,I329384,I329415,I329432,I329477,I329508,I329525,I329556,I329601,I329665,I329682,I350873,I350861,I329699,I350846,I329716,I329733,I350858,I329750,I350870,I329767,I329798,I350843,I350867,I329815,I350852,I329832,I329849,I329866,I329883,I329900,I329945,I350855,I329962,I350864,I329979,I330010,I330027,I330072,I330103,I350849,I330120,I330151,I330196,I330260,I330277,I389705,I389708,I330294,I389717,I330311,I330328,I389711,I330345,I389732,I330362,I330393,I389729,I389735,I330410,I389720,I330427,I330444,I330461,I330478,I330495,I330540,I389723,I330557,I389726,I330574,I330605,I330622,I330667,I330698,I389714,I330715,I330746,I330791,I330855,I330872,I330889,I330906,I330923,I330940,I330957,I330988,I331005,I331022,I331039,I331056,I331073,I331090,I331135,I331152,I331169,I331200,I331217,I331262,I331293,I331310,I331341,I331386,I331450,I331467,I331484,I331501,I331518,I331535,I331552,I331583,I331600,I331617,I331634,I331651,I331668,I331685,I331730,I331747,I331764,I331795,I331812,I331857,I331888,I331905,I331936,I331981,I332045,I332062,I332079,I332096,I332113,I332130,I332147,I332016,I332178,I332195,I332212,I332229,I332246,I332263,I332280,I332013,I332007,I332325,I332342,I332359,I332034,I332390,I332407,I332025,I332019,I332452,I332022,I332483,I332500,I332037,I332531,I332031,I332028,I332576,I332010,I332640,I332657,I332674,I332691,I332708,I332725,I332742,I332759,I332776,I332793,I332810,I332827,I332844,I332861,I332892,I332909,I332926,I332957,I332988,I333005,I333036,I333081,I333098,I333115,I333174,I333191,I333269,I333286,I333303,I333320,I333337,I333354,I333371,I333388,I333405,I333422,I333439,I333456,I333473,I333490,I333521,I333538,I333555,I333586,I333617,I333634,I333665,I333710,I333727,I333744,I333803,I333820,I333898,I333915,I333932,I333949,I333966,I333983,I334000,I334017,I334034,I334051,I334068,I334085,I334102,I334119,I334150,I334167,I334184,I334215,I334246,I334263,I334294,I334339,I334356,I334373,I334432,I334449,I334527,I334544,I334561,I334578,I334595,I334612,I334629,I334646,I334663,I334680,I334697,I334714,I334731,I334748,I334779,I334796,I334813,I334844,I334875,I334892,I334923,I334968,I334985,I335002,I335061,I335078,I335156,I335173,I335190,I335207,I335224,I335241,I335258,I335275,I335292,I335309,I335326,I335343,I335360,I335377,I335408,I335425,I335442,I335473,I335504,I335521,I335552,I335597,I335614,I335631,I335690,I335707,I335785,I335802,I335819,I335836,I335853,I335870,I335887,I335904,I335921,I335938,I335955,I335972,I335989,I336006,I336037,I336054,I336071,I336102,I336133,I336150,I336181,I336226,I336243,I336260,I336319,I336336,I336414,I336431,I336448,I336465,I336482,I336499,I336516,I336533,I336550,I336567,I336584,I336601,I336618,I336635,I336666,I336683,I336700,I336731,I336762,I336779,I336810,I336855,I336872,I336889,I336948,I336965,I337043,I337060,I337077,I337094,I337111,I337128,I337145,I337162,I337179,I337196,I337213,I337230,I337247,I337264,I337295,I337312,I337329,I337360,I337391,I337408,I337439,I337484,I337501,I337518,I337577,I337594,I337672,I337689,I384509,I337706,I384533,I384518,I337723,I384503,I337740,I337757,I384530,I337774,I337791,I337808,I384512,I337825,I384506,I337842,I384527,I337859,I384515,I337876,I337893,I337924,I337941,I337958,I337989,I384524,I338020,I338037,I338068,I338113,I384521,I338130,I338147,I338206,I338223,I338301,I338318,I338335,I338352,I338369,I338386,I338403,I338420,I338437,I338454,I338471,I338488,I338505,I338522,I338553,I338570,I338587,I338618,I338649,I338666,I338697,I338742,I338759,I338776,I338835,I338852,I338930,I338947,I396647,I338964,I396671,I396656,I338981,I396641,I338998,I339015,I396668,I339032,I339049,I339066,I396650,I339083,I396644,I339100,I396665,I339117,I396653,I339134,I339151,I339182,I339199,I339216,I339247,I396662,I339278,I339295,I339326,I339371,I396659,I339388,I339405,I339464,I339481,I339559,I339576,I339593,I339610,I339627,I339644,I339661,I339678,I339695,I339712,I339729,I339746,I339763,I339780,I339811,I339828,I339845,I339876,I339907,I339924,I339955,I340000,I340017,I340034,I340093,I340110,I340188,I340205,I340222,I340239,I340256,I340273,I340290,I340307,I340324,I340341,I340358,I340375,I340392,I340409,I340440,I340457,I340474,I340505,I340536,I340553,I340584,I340629,I340646,I340663,I340722,I340739,I340817,I340834,I340851,I340868,I340885,I340902,I340919,I340936,I340953,I340970,I340987,I341004,I341021,I341038,I341069,I341086,I341103,I341134,I341165,I341182,I341213,I341258,I341275,I341292,I341351,I341368,I341446,I341463,I341480,I341497,I341514,I341531,I341548,I341565,I341582,I341599,I341616,I341633,I341650,I341667,I341698,I341715,I341732,I341763,I341794,I341811,I341842,I341887,I341904,I341921,I341980,I341997,I342075,I342092,I342109,I342126,I342143,I342160,I342177,I342194,I342211,I342228,I342245,I342262,I342279,I342296,I342327,I342344,I342361,I342392,I342423,I342440,I342471,I342516,I342533,I342550,I342609,I342626,I342704,I342721,I342738,I342755,I342772,I342789,I342806,I342823,I342840,I342857,I342874,I342891,I342908,I342925,I342956,I342973,I342990,I343021,I343052,I343069,I343100,I343145,I343162,I343179,I343238,I343255,I343333,I343350,I343367,I343384,I343401,I343418,I343435,I343452,I343469,I343486,I343503,I343520,I343537,I343554,I343585,I343602,I343619,I343650,I343681,I343698,I343729,I343774,I343791,I343808,I343867,I343884,I343962,I343979,I343996,I344013,I344030,I344047,I344064,I344081,I344098,I344115,I344132,I344149,I344166,I344183,I344214,I344231,I344248,I344279,I344310,I344327,I344358,I344403,I344420,I344437,I344496,I344513,I344591,I344608,I344625,I344642,I344659,I344676,I344693,I344710,I344727,I344744,I344761,I344778,I344795,I344812,I344843,I344860,I344877,I344908,I344939,I344956,I344987,I345032,I345049,I345066,I345125,I345142,I345220,I345237,I381619,I345254,I381643,I381628,I345271,I381613,I345288,I345305,I381640,I345322,I345339,I345356,I381622,I345373,I381616,I345390,I381637,I345407,I381625,I345424,I345441,I345472,I345489,I345506,I345537,I381634,I345568,I345585,I345616,I345661,I381631,I345678,I345695,I345754,I345771,I345849,I345866,I345883,I345900,I345917,I345934,I345951,I345968,I345985,I346002,I346019,I346036,I346053,I346070,I346101,I346118,I346135,I346166,I346197,I346214,I346245,I346290,I346307,I346324,I346383,I346400,I346478,I346495,I346512,I346529,I346546,I346563,I346580,I346597,I346614,I346631,I346648,I346665,I346682,I346699,I346730,I346747,I346764,I346795,I346826,I346843,I346874,I346919,I346936,I346953,I347012,I347029,I347107,I347124,I347141,I347158,I347175,I347192,I347209,I347226,I347243,I347260,I347277,I347294,I347311,I347328,I347359,I347376,I347393,I347424,I347455,I347472,I347503,I347548,I347565,I347582,I347641,I347658,I347736,I347753,I347770,I347787,I347804,I347821,I347838,I347855,I347872,I347889,I347906,I347923,I347940,I347957,I347988,I348005,I348022,I348053,I348084,I348101,I348132,I348177,I348194,I348211,I348270,I348287,I348365,I348382,I348399,I348416,I348433,I348450,I348467,I348484,I348501,I348518,I348535,I348552,I348569,I348586,I348617,I348634,I348651,I348682,I348713,I348730,I348761,I348806,I348823,I348840,I348899,I348916,I348994,I349011,I349028,I349045,I349062,I349079,I349096,I349113,I349130,I349147,I349164,I349181,I349198,I349215,I349246,I349263,I349280,I349311,I349342,I349359,I349390,I349435,I349452,I349469,I349528,I349545,I349623,I349640,I349657,I349674,I349691,I349708,I349725,I349742,I349759,I349776,I349793,I349810,I349827,I349844,I349875,I349892,I349909,I349940,I349971,I349988,I350019,I350064,I350081,I350098,I350157,I350174,I350252,I350269,I350286,I350303,I350320,I350337,I350354,I350371,I350388,I350405,I350422,I350439,I350456,I350473,I350504,I350521,I350538,I350569,I350600,I350617,I350648,I350693,I350710,I350727,I350786,I350803,I350881,I350898,I350915,I350932,I350949,I350966,I350983,I351000,I351017,I351034,I351051,I351068,I351085,I351102,I351133,I351150,I351167,I351198,I351229,I351246,I351277,I351322,I351339,I351356,I351415,I351432,I351510,I351527,I351544,I351561,I351578,I351595,I351612,I351629,I351646,I351663,I351680,I351697,I351714,I351731,I351762,I351779,I351796,I351827,I351858,I351875,I351906,I351951,I351968,I351985,I352044,I352061,I352139,I352156,I352173,I352190,I352207,I352224,I352241,I352258,I352275,I352292,I352309,I352326,I352343,I352360,I352391,I352408,I352425,I352456,I352487,I352504,I352535,I352580,I352597,I352614,I352673,I352690,I352768,I352785,I352802,I352819,I352836,I352853,I352870,I352887,I352904,I352921,I352938,I352955,I352972,I352989,I353020,I353037,I353054,I353085,I353116,I353133,I353164,I353209,I353226,I353243,I353302,I353319,I353397,I353414,I353431,I353448,I353465,I353482,I353499,I353516,I353533,I353550,I353567,I353584,I353601,I353618,I353649,I353666,I353683,I353714,I353745,I353762,I353793,I353838,I353855,I353872,I353931,I353948,I354026,I354043,I354060,I354077,I354094,I354111,I354128,I354145,I354162,I354179,I354196,I354213,I354230,I354247,I354278,I354295,I354312,I354343,I354374,I354391,I354422,I354467,I354484,I354501,I354560,I354577,I354655,I354672,I354689,I354706,I354723,I354740,I354757,I354774,I354791,I354808,I354825,I354842,I354859,I354876,I354907,I354924,I354941,I354972,I355003,I355020,I355051,I355096,I355113,I355130,I355189,I355206,I355284,I355301,I355318,I355335,I355352,I355369,I355386,I355403,I355420,I355437,I355454,I355471,I355488,I355505,I355536,I355553,I355570,I355601,I355632,I355649,I355680,I355725,I355742,I355759,I355818,I355835,I355913,I355930,I355947,I355964,I355981,I355998,I356015,I356032,I356049,I356066,I356083,I356100,I356117,I356134,I356165,I356182,I356199,I356230,I356261,I356278,I356309,I356354,I356371,I356388,I356447,I356464,I356542,I356559,I356576,I356593,I356610,I356627,I356644,I356661,I356678,I356695,I356712,I356729,I356746,I356763,I356794,I356811,I356828,I356859,I356890,I356907,I356938,I356983,I357000,I357017,I357076,I357093,I357171,I357188,I357205,I357222,I357239,I357256,I357273,I357290,I357307,I357324,I357341,I357358,I357375,I357392,I357423,I357440,I357457,I357488,I357519,I357536,I357567,I357612,I357629,I357646,I357705,I357722,I357800,I357817,I357834,I357851,I357868,I357885,I357902,I357919,I357936,I357953,I357970,I357987,I358004,I358021,I358052,I358069,I358086,I358117,I358148,I358165,I358196,I358241,I358258,I358275,I358334,I358351,I358429,I358446,I358463,I358480,I358497,I358514,I358531,I358548,I358565,I358582,I358599,I358616,I358633,I358650,I358681,I358698,I358715,I358746,I358777,I358794,I358825,I358870,I358887,I358904,I358963,I358980,I359058,I359075,I359092,I359109,I359126,I359143,I359160,I359177,I359194,I359211,I359228,I359245,I359262,I359279,I359310,I359327,I359344,I359375,I359406,I359423,I359454,I359499,I359516,I359533,I359592,I359609,I359687,I359704,I359721,I359738,I359755,I359772,I359789,I359806,I359823,I359840,I359857,I359874,I359891,I359908,I359939,I359956,I359973,I360004,I360035,I360052,I360083,I360128,I360145,I360162,I360221,I360238,I360316,I360333,I360350,I360367,I360384,I360401,I360418,I360435,I360452,I360469,I360486,I360503,I360520,I360537,I360568,I360585,I360602,I360633,I360664,I360681,I360712,I360757,I360774,I360791,I360850,I360867,I360945,I360962,I360979,I360996,I361013,I361030,I361047,I361064,I361081,I361098,I361115,I361132,I361149,I361166,I361197,I361214,I361231,I361262,I361293,I361310,I361341,I361386,I361403,I361420,I361479,I361496,I361574,I361591,I361608,I361625,I361642,I361659,I361676,I361693,I361710,I361727,I361744,I361761,I361778,I361795,I361826,I361843,I361860,I361891,I361922,I361939,I361970,I362015,I362032,I362049,I362108,I362125,I362203,I362220,I362237,I362254,I362271,I362288,I362305,I362322,I362339,I362356,I362373,I362390,I362407,I362424,I362455,I362472,I362489,I362520,I362551,I362568,I362599,I362644,I362661,I362678,I362737,I362754,I362832,I362849,I362866,I362883,I362900,I362917,I362934,I362951,I362968,I362985,I363002,I363019,I363036,I363053,I363084,I363101,I363118,I363149,I363180,I363197,I363228,I363273,I363290,I363307,I363366,I363383,I363461,I363478,I363495,I363512,I363529,I363546,I363563,I363580,I363597,I363614,I363631,I363648,I363665,I363682,I363713,I363730,I363747,I363778,I363809,I363826,I363857,I363902,I363919,I363936,I363995,I364012,I364090,I364107,I395491,I364124,I395515,I395500,I364141,I395485,I364158,I364175,I395512,I364192,I364209,I364226,I395494,I364243,I395488,I364260,I395509,I364277,I395497,I364294,I364311,I364342,I364359,I364376,I364407,I395506,I364438,I364455,I364486,I364531,I395503,I364548,I364565,I364624,I364641,I364719,I364736,I364753,I364770,I364787,I364804,I364821,I364838,I364855,I364872,I364889,I364906,I364923,I364940,I364971,I364988,I365005,I365036,I365067,I365084,I365115,I365160,I365177,I365194,I365253,I365270,I365348,I365365,I365382,I365399,I365416,I365433,I365450,I365467,I365484,I365501,I365518,I365535,I365552,I365569,I365600,I365617,I365634,I365665,I365696,I365713,I365744,I365789,I365806,I365823,I365882,I365899,I365977,I365994,I366011,I366028,I366045,I366062,I366079,I366096,I366113,I366130,I366147,I366164,I366181,I366198,I366229,I366246,I366263,I366294,I366325,I366342,I366373,I366418,I366435,I366452,I366511,I366528,I366606,I366623,I366640,I366657,I366674,I366691,I366708,I366725,I366742,I366759,I366776,I366793,I366810,I366827,I366858,I366875,I366892,I366923,I366954,I366971,I367002,I367047,I367064,I367081,I367140,I367157,I367235,I367252,I367269,I367286,I367303,I367320,I367337,I367354,I367371,I367388,I367405,I367422,I367439,I367456,I367487,I367504,I367521,I367552,I367583,I367600,I367631,I367676,I367693,I367710,I367769,I367786,I367864,I367881,I367898,I367915,I367932,I367949,I367966,I367983,I368000,I368017,I368034,I368051,I368068,I368085,I368116,I368133,I368150,I368181,I368212,I368229,I368260,I368305,I368322,I368339,I368398,I368415,I368493,I368510,I368527,I368544,I368561,I368578,I368595,I368612,I368629,I368646,I368663,I368680,I368697,I368714,I368745,I368762,I368779,I368810,I368841,I368858,I368889,I368934,I368951,I368968,I369027,I369044,I369122,I369139,I369156,I369173,I369190,I369207,I369224,I369241,I369258,I369275,I369292,I369309,I369326,I369343,I369374,I369391,I369408,I369439,I369470,I369487,I369518,I369563,I369580,I369597,I369656,I369673,I369751,I369768,I369785,I369802,I369819,I369836,I369853,I369870,I369887,I369904,I369921,I369938,I369955,I369972,I370003,I370020,I370037,I370068,I370099,I370116,I370147,I370192,I370209,I370226,I370285,I370302,I370380,I370397,I370414,I370431,I370448,I370465,I370482,I370499,I370516,I370533,I370550,I370567,I370584,I370601,I370632,I370649,I370666,I370697,I370728,I370745,I370776,I370821,I370838,I370855,I370914,I370931,I371009,I371026,I371043,I371060,I371077,I371094,I371111,I371128,I371145,I371162,I371179,I371196,I371213,I371230,I371261,I371278,I371295,I371326,I371357,I371374,I371405,I371450,I371467,I371484,I371543,I371560,I371638,I371655,I371672,I371689,I371706,I371723,I371740,I371757,I371774,I371791,I371808,I371825,I371842,I371859,I371890,I371907,I371924,I371955,I371986,I372003,I372034,I372079,I372096,I372113,I372172,I372189,I372267,I372284,I372301,I372318,I372335,I372352,I372369,I372386,I372403,I372420,I372437,I372454,I372471,I372488,I372519,I372536,I372553,I372584,I372615,I372632,I372663,I372708,I372725,I372742,I372801,I372818,I372896,I372913,I372930,I372947,I372964,I372981,I372998,I373015,I373032,I373049,I373066,I373083,I373100,I373117,I373148,I373165,I373182,I373213,I373244,I373261,I373292,I373337,I373354,I373371,I373430,I373447,I373525,I373542,I373559,I373576,I373593,I373610,I373627,I373644,I373661,I373678,I373695,I373712,I373729,I373746,I373777,I373794,I373811,I373842,I373873,I373890,I373921,I373966,I373983,I374000,I374059,I374076,I374154,I374171,I374188,I374205,I374222,I374239,I374256,I374273,I374290,I374307,I374324,I374341,I374358,I374375,I374406,I374423,I374440,I374471,I374502,I374519,I374550,I374595,I374612,I374629,I374688,I374705,I374783,I374800,I374817,I374834,I374851,I374868,I374885,I374902,I374919,I374936,I374953,I374970,I374987,I375004,I375035,I375052,I375069,I375100,I375131,I375148,I375179,I375224,I375241,I375258,I375317,I375334,I375412,I375429,I375446,I375463,I375480,I375497,I375514,I375531,I375548,I375565,I375582,I375599,I375616,I375633,I375664,I375681,I375698,I375729,I375760,I375777,I375808,I375853,I375870,I375887,I375946,I375963,I376041,I376058,I376075,I376092,I376109,I376126,I376143,I376160,I376177,I376194,I376211,I376228,I376245,I376262,I376293,I376310,I376327,I376358,I376389,I376406,I376437,I376482,I376499,I376516,I376575,I376592,I376670,I376687,I376704,I376721,I376738,I376755,I376772,I376789,I376806,I376823,I376840,I376857,I376874,I376891,I376922,I376939,I376956,I376987,I377018,I377035,I377066,I377111,I377128,I377145,I377204,I377221,I377299,I377316,I377333,I377350,I377367,I377384,I377401,I377418,I377435,I377452,I377469,I377486,I377503,I377520,I377551,I377568,I377585,I377616,I377647,I377664,I377695,I377740,I377757,I377774,I377833,I377850,I377928,I377945,I377962,I377979,I377996,I378013,I378030,I378047,I378064,I378081,I378098,I378115,I378132,I378149,I378180,I378197,I378214,I378245,I378276,I378293,I378324,I378369,I378386,I378403,I378462,I378479,I378557,I378574,I378591,I378608,I378625,I378642,I378659,I378676,I378693,I378710,I378727,I378744,I378761,I378778,I378809,I378826,I378843,I378874,I378905,I378922,I378953,I378998,I379015,I379032,I379091,I379108,I379186,I379203,I379220,I379237,I379254,I379271,I379288,I379305,I379322,I379339,I379356,I379373,I379390,I379407,I379438,I379455,I379472,I379503,I379534,I379551,I379582,I379627,I379644,I379661,I379720,I379737,I379815,I379832,I379849,I379866,I379883,I379900,I379917,I379934,I379951,I379968,I379985,I380002,I380019,I380036,I380067,I380084,I380101,I380132,I380163,I380180,I380211,I380256,I380273,I380290,I380349,I380366,I380444,I380461,I380478,I380495,I380512,I380529,I380546,I380563,I380580,I380597,I380614,I380631,I380648,I380665,I380696,I380713,I380730,I380761,I380792,I380809,I380840,I380885,I380902,I380919,I380978,I380995,I381073,I381090,I381107,I381124,I381155,I381186,I381203,I381220,I381237,I381254,I381285,I381316,I381333,I381350,I381367,I381384,I381401,I381432,I381449,I381466,I381525,I381570,I381587,I381651,I381668,I381685,I381702,I381733,I381764,I381781,I381798,I381815,I381832,I381863,I381894,I381911,I381928,I381945,I381962,I381979,I382010,I382027,I382044,I382103,I382148,I382165,I382229,I382246,I382263,I382280,I382311,I382342,I382359,I382376,I382393,I382410,I382441,I382472,I382489,I382506,I382523,I382540,I382557,I382588,I382605,I382622,I382681,I382726,I382743,I382807,I382824,I382841,I382858,I382889,I382920,I382937,I382954,I382971,I382988,I383019,I383050,I383067,I383084,I383101,I383118,I383135,I383166,I383183,I383200,I383259,I383304,I383321,I383385,I383402,I383419,I383436,I383467,I383498,I383515,I383532,I383549,I383566,I383597,I383628,I383645,I383662,I383679,I383696,I383713,I383744,I383761,I383778,I383837,I383882,I383899,I383963,I383980,I383997,I384014,I384045,I384076,I384093,I384110,I384127,I384144,I384175,I384206,I384223,I384240,I384257,I384274,I384291,I384322,I384339,I384356,I384415,I384460,I384477,I384541,I384558,I384575,I384592,I384623,I384654,I384671,I384688,I384705,I384722,I384753,I384784,I384801,I384818,I384835,I384852,I384869,I384900,I384917,I384934,I384993,I385038,I385055,I385119,I385136,I385153,I385170,I385201,I385232,I385249,I385266,I385283,I385300,I385331,I385362,I385379,I385396,I385413,I385430,I385447,I385478,I385495,I385512,I385571,I385616,I385633,I385697,I385714,I385731,I385748,I385779,I385810,I385827,I385844,I385861,I385878,I385909,I385940,I385957,I385974,I385991,I386008,I386025,I386056,I386073,I386090,I386149,I386194,I386211,I386275,I386292,I386309,I386326,I386357,I386388,I386405,I386422,I386439,I386456,I386487,I386518,I386535,I386552,I386569,I386586,I386603,I386634,I386651,I386668,I386727,I386772,I386789,I386853,I386870,I386887,I386904,I386935,I386966,I386983,I387000,I387017,I387034,I387065,I387096,I387113,I387130,I387147,I387164,I387181,I387212,I387229,I387246,I387305,I387350,I387367,I387431,I387448,I387465,I387482,I387513,I387544,I387561,I387578,I387595,I387612,I387643,I387674,I387691,I387708,I387725,I387742,I387759,I387790,I387807,I387824,I387883,I387928,I387945,I388009,I388026,I388043,I388060,I388091,I388122,I388139,I388156,I388173,I388190,I388221,I388252,I388269,I388286,I388303,I388320,I388337,I388368,I388385,I388402,I388461,I388506,I388523,I388587,I388604,I388621,I388638,I388669,I388700,I388717,I388734,I388751,I388768,I388799,I388830,I388847,I388864,I388881,I388898,I388915,I388946,I388963,I388980,I389039,I389084,I389101,I389165,I389182,I389199,I389216,I389247,I389278,I389295,I389312,I389329,I389346,I389377,I389408,I389425,I389442,I389459,I389476,I389493,I389524,I389541,I389558,I389617,I389662,I389679,I389743,I389760,I389777,I389794,I389825,I389856,I389873,I389890,I389907,I389924,I389955,I389986,I390003,I390020,I390037,I390054,I390071,I390102,I390119,I390136,I390195,I390240,I390257,I390321,I390338,I390355,I390372,I390403,I390434,I390451,I390468,I390485,I390502,I390533,I390564,I390581,I390598,I390615,I390632,I390649,I390680,I390697,I390714,I390773,I390818,I390835,I390899,I390916,I390933,I390950,I390981,I391012,I391029,I391046,I391063,I391080,I391111,I391142,I391159,I391176,I391193,I391210,I391227,I391258,I391275,I391292,I391351,I391396,I391413,I391477,I391494,I391511,I391528,I391559,I391590,I391607,I391624,I391641,I391658,I391689,I391720,I391737,I391754,I391771,I391788,I391805,I391836,I391853,I391870,I391929,I391974,I391991,I392055,I392072,I392089,I392106,I392137,I392168,I392185,I392202,I392219,I392236,I392267,I392298,I392315,I392332,I392349,I392366,I392383,I392414,I392431,I392448,I392507,I392552,I392569,I392633,I392650,I392667,I392684,I392715,I392746,I392763,I392780,I392797,I392814,I392845,I392876,I392893,I392910,I392927,I392944,I392961,I392992,I393009,I393026,I393085,I393130,I393147,I393211,I393228,I393245,I393262,I393293,I393324,I393341,I393358,I393375,I393392,I393423,I393454,I393471,I393488,I393505,I393522,I393539,I393570,I393587,I393604,I393663,I393708,I393725,I393789,I393806,I393823,I393840,I393871,I393902,I393919,I393936,I393953,I393970,I394001,I394032,I394049,I394066,I394083,I394100,I394117,I394148,I394165,I394182,I394241,I394286,I394303,I394367,I394384,I394401,I394418,I394449,I394480,I394497,I394514,I394531,I394548,I394579,I394610,I394627,I394644,I394661,I394678,I394695,I394726,I394743,I394760,I394819,I394864,I394881,I394945,I394962,I394979,I394996,I395027,I395058,I395075,I395092,I395109,I395126,I395157,I395188,I395205,I395222,I395239,I395256,I395273,I395304,I395321,I395338,I395397,I395442,I395459,I395523,I395540,I395557,I395574,I395605,I395636,I395653,I395670,I395687,I395704,I395735,I395766,I395783,I395800,I395817,I395834,I395851,I395882,I395899,I395916,I395975,I396020,I396037,I396101,I396118,I396135,I396152,I396183,I396214,I396231,I396248,I396265,I396282,I396313,I396344,I396361,I396378,I396395,I396412,I396429,I396460,I396477,I396494,I396553,I396598,I396615,I396679,I396696,I396713,I396730,I396761,I396792,I396809,I396826,I396843,I396860,I396891,I396922,I396939,I396956,I396973,I396990,I397007,I397038,I397055,I397072,I397131,I397176,I397193,I397257,I397274,I397291,I397308,I397339,I397370,I397387,I397404,I397421,I397438,I397469,I397500,I397517,I397534,I397551,I397568,I397585,I397616,I397633,I397650,I397709,I397754,I397771;
not I_0 (I2398,I2357);
nand I_1 (I2415,I363423,I363426);
and I_2 (I2432,I2415,I363432);
DFFARX1 I_3  ( .D(I2432), .CLK(I2350), .RSTB(I2398), .Q(I2449) );
not I_4 (I2466,I2449);
nor I_5 (I2483,I363444,I363426);
or I_6 (I2381,I2483,I2449);
not I_7 (I2369,I2483);
DFFARX1 I_8  ( .D(I363453), .CLK(I2350), .RSTB(I2398), .Q(I2528) );
nor I_9 (I2545,I2528,I2483);
nand I_10 (I2562,I363441,I363438);
and I_11 (I2579,I2562,I363450);
DFFARX1 I_12  ( .D(I2579), .CLK(I2350), .RSTB(I2398), .Q(I2596) );
nor I_13 (I2378,I2596,I2449);
not I_14 (I2627,I2596);
nor I_15 (I2644,I2528,I2627);
DFFARX1 I_16  ( .D(I363447), .CLK(I2350), .RSTB(I2398), .Q(I2661) );
and I_17 (I2678,I2661,I363435);
or I_18 (I2387,I2678,I2483);
nand I_19 (I2366,I2678,I2644);
DFFARX1 I_20  ( .D(I363429), .CLK(I2350), .RSTB(I2398), .Q(I2723) );
and I_21 (I2740,I2723,I2466);
nor I_22 (I2384,I2678,I2740);
nor I_23 (I2771,I2723,I2528);
DFFARX1 I_24  ( .D(I2771), .CLK(I2350), .RSTB(I2398), .Q(I2375) );
nor I_25 (I2390,I2723,I2449);
not I_26 (I2816,I2723);
nor I_27 (I2833,I2596,I2816);
and I_28 (I2850,I2483,I2833);
or I_29 (I2867,I2678,I2850);
DFFARX1 I_30  ( .D(I2867), .CLK(I2350), .RSTB(I2398), .Q(I2363) );
nand I_31 (I2372,I2723,I2545);
nand I_32 (I2360,I2723,I2627);
not I_33 (I2959,I2357);
nand I_34 (I2976,I226977,I226968);
and I_35 (I2993,I2976,I226971);
DFFARX1 I_36  ( .D(I2993), .CLK(I2350), .RSTB(I2959), .Q(I3010) );
not I_37 (I3027,I3010);
nor I_38 (I3044,I226947,I226968);
or I_39 (I2942,I3044,I3010);
not I_40 (I2930,I3044);
DFFARX1 I_41  ( .D(I226962), .CLK(I2350), .RSTB(I2959), .Q(I3089) );
nor I_42 (I3106,I3089,I3044);
nand I_43 (I3123,I226950,I226965);
and I_44 (I3140,I3123,I226959);
DFFARX1 I_45  ( .D(I3140), .CLK(I2350), .RSTB(I2959), .Q(I3157) );
nor I_46 (I2939,I3157,I3010);
not I_47 (I3188,I3157);
nor I_48 (I3205,I3089,I3188);
DFFARX1 I_49  ( .D(I226974), .CLK(I2350), .RSTB(I2959), .Q(I3222) );
and I_50 (I3239,I3222,I226953);
or I_51 (I2948,I3239,I3044);
nand I_52 (I2927,I3239,I3205);
DFFARX1 I_53  ( .D(I226956), .CLK(I2350), .RSTB(I2959), .Q(I3284) );
and I_54 (I3301,I3284,I3027);
nor I_55 (I2945,I3239,I3301);
nor I_56 (I3332,I3284,I3089);
DFFARX1 I_57  ( .D(I3332), .CLK(I2350), .RSTB(I2959), .Q(I2936) );
nor I_58 (I2951,I3284,I3010);
not I_59 (I3377,I3284);
nor I_60 (I3394,I3157,I3377);
and I_61 (I3411,I3044,I3394);
or I_62 (I3428,I3239,I3411);
DFFARX1 I_63  ( .D(I3428), .CLK(I2350), .RSTB(I2959), .Q(I2924) );
nand I_64 (I2933,I3284,I3106);
nand I_65 (I2921,I3284,I3188);
not I_66 (I3520,I2357);
nand I_67 (I3537,I362794,I362797);
and I_68 (I3554,I3537,I362803);
DFFARX1 I_69  ( .D(I3554), .CLK(I2350), .RSTB(I3520), .Q(I3571) );
not I_70 (I3588,I3571);
nor I_71 (I3605,I362815,I362797);
or I_72 (I3503,I3605,I3571);
not I_73 (I3491,I3605);
DFFARX1 I_74  ( .D(I362824), .CLK(I2350), .RSTB(I3520), .Q(I3650) );
nor I_75 (I3667,I3650,I3605);
nand I_76 (I3684,I362812,I362809);
and I_77 (I3701,I3684,I362821);
DFFARX1 I_78  ( .D(I3701), .CLK(I2350), .RSTB(I3520), .Q(I3718) );
nor I_79 (I3500,I3718,I3571);
not I_80 (I3749,I3718);
nor I_81 (I3766,I3650,I3749);
DFFARX1 I_82  ( .D(I362818), .CLK(I2350), .RSTB(I3520), .Q(I3783) );
and I_83 (I3800,I3783,I362806);
or I_84 (I3509,I3800,I3605);
nand I_85 (I3488,I3800,I3766);
DFFARX1 I_86  ( .D(I362800), .CLK(I2350), .RSTB(I3520), .Q(I3845) );
and I_87 (I3862,I3845,I3588);
nor I_88 (I3506,I3800,I3862);
nor I_89 (I3893,I3845,I3650);
DFFARX1 I_90  ( .D(I3893), .CLK(I2350), .RSTB(I3520), .Q(I3497) );
nor I_91 (I3512,I3845,I3571);
not I_92 (I3938,I3845);
nor I_93 (I3955,I3718,I3938);
and I_94 (I3972,I3605,I3955);
or I_95 (I3989,I3800,I3972);
DFFARX1 I_96  ( .D(I3989), .CLK(I2350), .RSTB(I3520), .Q(I3485) );
nand I_97 (I3494,I3845,I3667);
nand I_98 (I3482,I3845,I3749);
not I_99 (I4081,I2357);
nand I_100 (I4098,I333860,I333863);
and I_101 (I4115,I4098,I333869);
DFFARX1 I_102  ( .D(I4115), .CLK(I2350), .RSTB(I4081), .Q(I4132) );
not I_103 (I4149,I4132);
nor I_104 (I4166,I333881,I333863);
or I_105 (I4064,I4166,I4132);
not I_106 (I4052,I4166);
DFFARX1 I_107  ( .D(I333890), .CLK(I2350), .RSTB(I4081), .Q(I4211) );
nor I_108 (I4228,I4211,I4166);
nand I_109 (I4245,I333878,I333875);
and I_110 (I4262,I4245,I333887);
DFFARX1 I_111  ( .D(I4262), .CLK(I2350), .RSTB(I4081), .Q(I4279) );
nor I_112 (I4061,I4279,I4132);
not I_113 (I4310,I4279);
nor I_114 (I4327,I4211,I4310);
DFFARX1 I_115  ( .D(I333884), .CLK(I2350), .RSTB(I4081), .Q(I4344) );
and I_116 (I4361,I4344,I333872);
or I_117 (I4070,I4361,I4166);
nand I_118 (I4049,I4361,I4327);
DFFARX1 I_119  ( .D(I333866), .CLK(I2350), .RSTB(I4081), .Q(I4406) );
and I_120 (I4423,I4406,I4149);
nor I_121 (I4067,I4361,I4423);
nor I_122 (I4454,I4406,I4211);
DFFARX1 I_123  ( .D(I4454), .CLK(I2350), .RSTB(I4081), .Q(I4058) );
nor I_124 (I4073,I4406,I4132);
not I_125 (I4499,I4406);
nor I_126 (I4516,I4279,I4499);
and I_127 (I4533,I4166,I4516);
or I_128 (I4550,I4361,I4533);
DFFARX1 I_129  ( .D(I4550), .CLK(I2350), .RSTB(I4081), .Q(I4046) );
nand I_130 (I4055,I4406,I4228);
nand I_131 (I4043,I4406,I4310);
not I_132 (I4642,I2357);
nand I_133 (I4659,I125804,I125807);
and I_134 (I4676,I4659,I125801);
DFFARX1 I_135  ( .D(I4676), .CLK(I2350), .RSTB(I4642), .Q(I4693) );
not I_136 (I4710,I4693);
nor I_137 (I4727,I125792,I125807);
or I_138 (I4625,I4727,I4693);
not I_139 (I4613,I4727);
DFFARX1 I_140  ( .D(I125780), .CLK(I2350), .RSTB(I4642), .Q(I4772) );
nor I_141 (I4789,I4772,I4727);
nand I_142 (I4806,I125789,I125783);
and I_143 (I4823,I4806,I125795);
DFFARX1 I_144  ( .D(I4823), .CLK(I2350), .RSTB(I4642), .Q(I4840) );
nor I_145 (I4622,I4840,I4693);
not I_146 (I4871,I4840);
nor I_147 (I4888,I4772,I4871);
DFFARX1 I_148  ( .D(I125810), .CLK(I2350), .RSTB(I4642), .Q(I4905) );
and I_149 (I4922,I4905,I125798);
or I_150 (I4631,I4922,I4727);
nand I_151 (I4610,I4922,I4888);
DFFARX1 I_152  ( .D(I125786), .CLK(I2350), .RSTB(I4642), .Q(I4967) );
and I_153 (I4984,I4967,I4710);
nor I_154 (I4628,I4922,I4984);
nor I_155 (I5015,I4967,I4772);
DFFARX1 I_156  ( .D(I5015), .CLK(I2350), .RSTB(I4642), .Q(I4619) );
nor I_157 (I4634,I4967,I4693);
not I_158 (I5060,I4967);
nor I_159 (I5077,I4840,I5060);
and I_160 (I5094,I4727,I5077);
or I_161 (I5111,I4922,I5094);
DFFARX1 I_162  ( .D(I5111), .CLK(I2350), .RSTB(I4642), .Q(I4607) );
nand I_163 (I4616,I4967,I4789);
nand I_164 (I4604,I4967,I4871);
not I_165 (I5203,I2357);
nand I_166 (I5220,I169528,I169519);
and I_167 (I5237,I5220,I169534);
DFFARX1 I_168  ( .D(I5237), .CLK(I2350), .RSTB(I5203), .Q(I5254) );
not I_169 (I5271,I5254);
nor I_170 (I5288,I169504,I169519);
or I_171 (I5186,I5288,I5254);
not I_172 (I5174,I5288);
DFFARX1 I_173  ( .D(I169507), .CLK(I2350), .RSTB(I5203), .Q(I5333) );
nor I_174 (I5350,I5333,I5288);
nand I_175 (I5367,I169525,I169522);
and I_176 (I5384,I5367,I169510);
DFFARX1 I_177  ( .D(I5384), .CLK(I2350), .RSTB(I5203), .Q(I5401) );
nor I_178 (I5183,I5401,I5254);
not I_179 (I5432,I5401);
nor I_180 (I5449,I5333,I5432);
DFFARX1 I_181  ( .D(I169531), .CLK(I2350), .RSTB(I5203), .Q(I5466) );
and I_182 (I5483,I5466,I169516);
or I_183 (I5192,I5483,I5288);
nand I_184 (I5171,I5483,I5449);
DFFARX1 I_185  ( .D(I169513), .CLK(I2350), .RSTB(I5203), .Q(I5528) );
and I_186 (I5545,I5528,I5271);
nor I_187 (I5189,I5483,I5545);
nor I_188 (I5576,I5528,I5333);
DFFARX1 I_189  ( .D(I5576), .CLK(I2350), .RSTB(I5203), .Q(I5180) );
nor I_190 (I5195,I5528,I5254);
not I_191 (I5621,I5528);
nor I_192 (I5638,I5401,I5621);
and I_193 (I5655,I5288,I5638);
or I_194 (I5672,I5483,I5655);
DFFARX1 I_195  ( .D(I5672), .CLK(I2350), .RSTB(I5203), .Q(I5168) );
nand I_196 (I5177,I5528,I5350);
nand I_197 (I5165,I5528,I5432);
not I_198 (I5764,I2357);
nand I_199 (I5781,I221809,I221800);
and I_200 (I5798,I5781,I221803);
DFFARX1 I_201  ( .D(I5798), .CLK(I2350), .RSTB(I5764), .Q(I5815) );
not I_202 (I5832,I5815);
nor I_203 (I5849,I221779,I221800);
or I_204 (I5747,I5849,I5815);
not I_205 (I5735,I5849);
DFFARX1 I_206  ( .D(I221794), .CLK(I2350), .RSTB(I5764), .Q(I5894) );
nor I_207 (I5911,I5894,I5849);
nand I_208 (I5928,I221782,I221797);
and I_209 (I5945,I5928,I221791);
DFFARX1 I_210  ( .D(I5945), .CLK(I2350), .RSTB(I5764), .Q(I5962) );
nor I_211 (I5744,I5962,I5815);
not I_212 (I5993,I5962);
nor I_213 (I6010,I5894,I5993);
DFFARX1 I_214  ( .D(I221806), .CLK(I2350), .RSTB(I5764), .Q(I6027) );
and I_215 (I6044,I6027,I221785);
or I_216 (I5753,I6044,I5849);
nand I_217 (I5732,I6044,I6010);
DFFARX1 I_218  ( .D(I221788), .CLK(I2350), .RSTB(I5764), .Q(I6089) );
and I_219 (I6106,I6089,I5832);
nor I_220 (I5750,I6044,I6106);
nor I_221 (I6137,I6089,I5894);
DFFARX1 I_222  ( .D(I6137), .CLK(I2350), .RSTB(I5764), .Q(I5741) );
nor I_223 (I5756,I6089,I5815);
not I_224 (I6182,I6089);
nor I_225 (I6199,I5962,I6182);
and I_226 (I6216,I5849,I6199);
or I_227 (I6233,I6044,I6216);
DFFARX1 I_228  ( .D(I6233), .CLK(I2350), .RSTB(I5764), .Q(I5729) );
nand I_229 (I5738,I6089,I5911);
nand I_230 (I5726,I6089,I5993);
not I_231 (I6325,I2357);
nand I_232 (I6342,I319533,I319521);
and I_233 (I6359,I6342,I319518);
DFFARX1 I_234  ( .D(I6359), .CLK(I2350), .RSTB(I6325), .Q(I6376) );
not I_235 (I6393,I6376);
nor I_236 (I6410,I319539,I319521);
or I_237 (I6308,I6410,I6376);
not I_238 (I6296,I6410);
DFFARX1 I_239  ( .D(I319542), .CLK(I2350), .RSTB(I6325), .Q(I6455) );
nor I_240 (I6472,I6455,I6410);
nand I_241 (I6489,I319512,I319530);
and I_242 (I6506,I6489,I319527);
DFFARX1 I_243  ( .D(I6506), .CLK(I2350), .RSTB(I6325), .Q(I6523) );
nor I_244 (I6305,I6523,I6376);
not I_245 (I6554,I6523);
nor I_246 (I6571,I6455,I6554);
DFFARX1 I_247  ( .D(I319536), .CLK(I2350), .RSTB(I6325), .Q(I6588) );
and I_248 (I6605,I6588,I319524);
or I_249 (I6314,I6605,I6410);
nand I_250 (I6293,I6605,I6571);
DFFARX1 I_251  ( .D(I319515), .CLK(I2350), .RSTB(I6325), .Q(I6650) );
and I_252 (I6667,I6650,I6393);
nor I_253 (I6311,I6605,I6667);
nor I_254 (I6698,I6650,I6455);
DFFARX1 I_255  ( .D(I6698), .CLK(I2350), .RSTB(I6325), .Q(I6302) );
nor I_256 (I6317,I6650,I6376);
not I_257 (I6743,I6650);
nor I_258 (I6760,I6523,I6743);
and I_259 (I6777,I6410,I6760);
or I_260 (I6794,I6605,I6777);
DFFARX1 I_261  ( .D(I6794), .CLK(I2350), .RSTB(I6325), .Q(I6290) );
nand I_262 (I6299,I6650,I6472);
nand I_263 (I6287,I6650,I6554);
not I_264 (I6886,I2357);
nand I_265 (I6903,I215349,I215340);
and I_266 (I6920,I6903,I215343);
DFFARX1 I_267  ( .D(I6920), .CLK(I2350), .RSTB(I6886), .Q(I6937) );
not I_268 (I6954,I6937);
nor I_269 (I6971,I215319,I215340);
or I_270 (I6869,I6971,I6937);
not I_271 (I6857,I6971);
DFFARX1 I_272  ( .D(I215334), .CLK(I2350), .RSTB(I6886), .Q(I7016) );
nor I_273 (I7033,I7016,I6971);
nand I_274 (I7050,I215322,I215337);
and I_275 (I7067,I7050,I215331);
DFFARX1 I_276  ( .D(I7067), .CLK(I2350), .RSTB(I6886), .Q(I7084) );
nor I_277 (I6866,I7084,I6937);
not I_278 (I7115,I7084);
nor I_279 (I7132,I7016,I7115);
DFFARX1 I_280  ( .D(I215346), .CLK(I2350), .RSTB(I6886), .Q(I7149) );
and I_281 (I7166,I7149,I215325);
or I_282 (I6875,I7166,I6971);
nand I_283 (I6854,I7166,I7132);
DFFARX1 I_284  ( .D(I215328), .CLK(I2350), .RSTB(I6886), .Q(I7211) );
and I_285 (I7228,I7211,I6954);
nor I_286 (I6872,I7166,I7228);
nor I_287 (I7259,I7211,I7016);
DFFARX1 I_288  ( .D(I7259), .CLK(I2350), .RSTB(I6886), .Q(I6863) );
nor I_289 (I6878,I7211,I6937);
not I_290 (I7304,I7211);
nor I_291 (I7321,I7084,I7304);
and I_292 (I7338,I6971,I7321);
or I_293 (I7355,I7166,I7338);
DFFARX1 I_294  ( .D(I7355), .CLK(I2350), .RSTB(I6886), .Q(I6851) );
nand I_295 (I6860,I7211,I7033);
nand I_296 (I6848,I7211,I7115);
not I_297 (I7447,I2357);
nand I_298 (I7464,I36925,I36928);
and I_299 (I7481,I7464,I36910);
DFFARX1 I_300  ( .D(I7481), .CLK(I2350), .RSTB(I7447), .Q(I7498) );
not I_301 (I7515,I7498);
nor I_302 (I7532,I36907,I36928);
or I_303 (I7430,I7532,I7498);
not I_304 (I7418,I7532);
DFFARX1 I_305  ( .D(I36931), .CLK(I2350), .RSTB(I7447), .Q(I7577) );
nor I_306 (I7594,I7577,I7532);
nand I_307 (I7611,I36916,I36922);
and I_308 (I7628,I7611,I36934);
DFFARX1 I_309  ( .D(I7628), .CLK(I2350), .RSTB(I7447), .Q(I7645) );
nor I_310 (I7427,I7645,I7498);
not I_311 (I7676,I7645);
nor I_312 (I7693,I7577,I7676);
DFFARX1 I_313  ( .D(I36913), .CLK(I2350), .RSTB(I7447), .Q(I7710) );
and I_314 (I7727,I7710,I36904);
or I_315 (I7436,I7727,I7532);
nand I_316 (I7415,I7727,I7693);
DFFARX1 I_317  ( .D(I36919), .CLK(I2350), .RSTB(I7447), .Q(I7772) );
and I_318 (I7789,I7772,I7515);
nor I_319 (I7433,I7727,I7789);
nor I_320 (I7820,I7772,I7577);
DFFARX1 I_321  ( .D(I7820), .CLK(I2350), .RSTB(I7447), .Q(I7424) );
nor I_322 (I7439,I7772,I7498);
not I_323 (I7865,I7772);
nor I_324 (I7882,I7645,I7865);
and I_325 (I7899,I7532,I7882);
or I_326 (I7916,I7727,I7899);
DFFARX1 I_327  ( .D(I7916), .CLK(I2350), .RSTB(I7447), .Q(I7412) );
nand I_328 (I7421,I7772,I7594);
nand I_329 (I7409,I7772,I7676);
not I_330 (I8008,I2357);
nand I_331 (I8025,I45323,I45326);
and I_332 (I8042,I8025,I45308);
DFFARX1 I_333  ( .D(I8042), .CLK(I2350), .RSTB(I8008), .Q(I8059) );
not I_334 (I8076,I8059);
nor I_335 (I8093,I45305,I45326);
or I_336 (I7991,I8093,I8059);
not I_337 (I7979,I8093);
DFFARX1 I_338  ( .D(I45329), .CLK(I2350), .RSTB(I8008), .Q(I8138) );
nor I_339 (I8155,I8138,I8093);
nand I_340 (I8172,I45314,I45320);
and I_341 (I8189,I8172,I45332);
DFFARX1 I_342  ( .D(I8189), .CLK(I2350), .RSTB(I8008), .Q(I8206) );
nor I_343 (I7988,I8206,I8059);
not I_344 (I8237,I8206);
nor I_345 (I8254,I8138,I8237);
DFFARX1 I_346  ( .D(I45311), .CLK(I2350), .RSTB(I8008), .Q(I8271) );
and I_347 (I8288,I8271,I45302);
or I_348 (I7997,I8288,I8093);
nand I_349 (I7976,I8288,I8254);
DFFARX1 I_350  ( .D(I45317), .CLK(I2350), .RSTB(I8008), .Q(I8333) );
and I_351 (I8350,I8333,I8076);
nor I_352 (I7994,I8288,I8350);
nor I_353 (I8381,I8333,I8138);
DFFARX1 I_354  ( .D(I8381), .CLK(I2350), .RSTB(I8008), .Q(I7985) );
nor I_355 (I8000,I8333,I8059);
not I_356 (I8426,I8333);
nor I_357 (I8443,I8206,I8426);
and I_358 (I8460,I8093,I8443);
or I_359 (I8477,I8288,I8460);
DFFARX1 I_360  ( .D(I8477), .CLK(I2350), .RSTB(I8008), .Q(I7973) );
nand I_361 (I7982,I8333,I8155);
nand I_362 (I7970,I8333,I8237);
not I_363 (I8569,I2357);
nand I_364 (I8586,I111900,I111897);
and I_365 (I8603,I8586,I111894);
DFFARX1 I_366  ( .D(I8603), .CLK(I2350), .RSTB(I8569), .Q(I8620) );
not I_367 (I8637,I8620);
nor I_368 (I8654,I111918,I111897);
or I_369 (I8552,I8654,I8620);
not I_370 (I8540,I8654);
DFFARX1 I_371  ( .D(I111912), .CLK(I2350), .RSTB(I8569), .Q(I8699) );
nor I_372 (I8716,I8699,I8654);
nand I_373 (I8733,I111891,I111903);
and I_374 (I8750,I8733,I111906);
DFFARX1 I_375  ( .D(I8750), .CLK(I2350), .RSTB(I8569), .Q(I8767) );
nor I_376 (I8549,I8767,I8620);
not I_377 (I8798,I8767);
nor I_378 (I8815,I8699,I8798);
DFFARX1 I_379  ( .D(I111915), .CLK(I2350), .RSTB(I8569), .Q(I8832) );
and I_380 (I8849,I8832,I111921);
or I_381 (I8558,I8849,I8654);
nand I_382 (I8537,I8849,I8815);
DFFARX1 I_383  ( .D(I111909), .CLK(I2350), .RSTB(I8569), .Q(I8894) );
and I_384 (I8911,I8894,I8637);
nor I_385 (I8555,I8849,I8911);
nor I_386 (I8942,I8894,I8699);
DFFARX1 I_387  ( .D(I8942), .CLK(I2350), .RSTB(I8569), .Q(I8546) );
nor I_388 (I8561,I8894,I8620);
not I_389 (I8987,I8894);
nor I_390 (I9004,I8767,I8987);
and I_391 (I9021,I8654,I9004);
or I_392 (I9038,I8849,I9021);
DFFARX1 I_393  ( .D(I9038), .CLK(I2350), .RSTB(I8569), .Q(I8534) );
nand I_394 (I8543,I8894,I8716);
nand I_395 (I8531,I8894,I8798);
not I_396 (I9130,I2357);
nand I_397 (I9147,I345182,I345185);
and I_398 (I9164,I9147,I345191);
DFFARX1 I_399  ( .D(I9164), .CLK(I2350), .RSTB(I9130), .Q(I9181) );
not I_400 (I9198,I9181);
nor I_401 (I9215,I345203,I345185);
or I_402 (I9113,I9215,I9181);
not I_403 (I9101,I9215);
DFFARX1 I_404  ( .D(I345212), .CLK(I2350), .RSTB(I9130), .Q(I9260) );
nor I_405 (I9277,I9260,I9215);
nand I_406 (I9294,I345200,I345197);
and I_407 (I9311,I9294,I345209);
DFFARX1 I_408  ( .D(I9311), .CLK(I2350), .RSTB(I9130), .Q(I9328) );
nor I_409 (I9110,I9328,I9181);
not I_410 (I9359,I9328);
nor I_411 (I9376,I9260,I9359);
DFFARX1 I_412  ( .D(I345206), .CLK(I2350), .RSTB(I9130), .Q(I9393) );
and I_413 (I9410,I9393,I345194);
or I_414 (I9119,I9410,I9215);
nand I_415 (I9098,I9410,I9376);
DFFARX1 I_416  ( .D(I345188), .CLK(I2350), .RSTB(I9130), .Q(I9455) );
and I_417 (I9472,I9455,I9198);
nor I_418 (I9116,I9410,I9472);
nor I_419 (I9503,I9455,I9260);
DFFARX1 I_420  ( .D(I9503), .CLK(I2350), .RSTB(I9130), .Q(I9107) );
nor I_421 (I9122,I9455,I9181);
not I_422 (I9548,I9455);
nor I_423 (I9565,I9328,I9548);
and I_424 (I9582,I9215,I9565);
or I_425 (I9599,I9410,I9582);
DFFARX1 I_426  ( .D(I9599), .CLK(I2350), .RSTB(I9130), .Q(I9095) );
nand I_427 (I9104,I9455,I9277);
nand I_428 (I9092,I9455,I9359);
not I_429 (I9691,I2357);
nand I_430 (I9708,I119259,I119262);
and I_431 (I9725,I9708,I119256);
DFFARX1 I_432  ( .D(I9725), .CLK(I2350), .RSTB(I9691), .Q(I9742) );
not I_433 (I9759,I9742);
nor I_434 (I9776,I119247,I119262);
or I_435 (I9674,I9776,I9742);
not I_436 (I9662,I9776);
DFFARX1 I_437  ( .D(I119235), .CLK(I2350), .RSTB(I9691), .Q(I9821) );
nor I_438 (I9838,I9821,I9776);
nand I_439 (I9855,I119244,I119238);
and I_440 (I9872,I9855,I119250);
DFFARX1 I_441  ( .D(I9872), .CLK(I2350), .RSTB(I9691), .Q(I9889) );
nor I_442 (I9671,I9889,I9742);
not I_443 (I9920,I9889);
nor I_444 (I9937,I9821,I9920);
DFFARX1 I_445  ( .D(I119265), .CLK(I2350), .RSTB(I9691), .Q(I9954) );
and I_446 (I9971,I9954,I119253);
or I_447 (I9680,I9971,I9776);
nand I_448 (I9659,I9971,I9937);
DFFARX1 I_449  ( .D(I119241), .CLK(I2350), .RSTB(I9691), .Q(I10016) );
and I_450 (I10033,I10016,I9759);
nor I_451 (I9677,I9971,I10033);
nor I_452 (I10064,I10016,I9821);
DFFARX1 I_453  ( .D(I10064), .CLK(I2350), .RSTB(I9691), .Q(I9668) );
nor I_454 (I9683,I10016,I9742);
not I_455 (I10109,I10016);
nor I_456 (I10126,I9889,I10109);
and I_457 (I10143,I9776,I10126);
or I_458 (I10160,I9971,I10143);
DFFARX1 I_459  ( .D(I10160), .CLK(I2350), .RSTB(I9691), .Q(I9656) );
nand I_460 (I9665,I10016,I9838);
nand I_461 (I9653,I10016,I9920);
not I_462 (I10252,I2357);
nand I_463 (I10269,I78269,I78272);
and I_464 (I10286,I10269,I78254);
DFFARX1 I_465  ( .D(I10286), .CLK(I2350), .RSTB(I10252), .Q(I10303) );
not I_466 (I10320,I10303);
nor I_467 (I10337,I78251,I78272);
or I_468 (I10235,I10337,I10303);
not I_469 (I10223,I10337);
DFFARX1 I_470  ( .D(I78275), .CLK(I2350), .RSTB(I10252), .Q(I10382) );
nor I_471 (I10399,I10382,I10337);
nand I_472 (I10416,I78260,I78266);
and I_473 (I10433,I10416,I78278);
DFFARX1 I_474  ( .D(I10433), .CLK(I2350), .RSTB(I10252), .Q(I10450) );
nor I_475 (I10232,I10450,I10303);
not I_476 (I10481,I10450);
nor I_477 (I10498,I10382,I10481);
DFFARX1 I_478  ( .D(I78257), .CLK(I2350), .RSTB(I10252), .Q(I10515) );
and I_479 (I10532,I10515,I78248);
or I_480 (I10241,I10532,I10337);
nand I_481 (I10220,I10532,I10498);
DFFARX1 I_482  ( .D(I78263), .CLK(I2350), .RSTB(I10252), .Q(I10577) );
and I_483 (I10594,I10577,I10320);
nor I_484 (I10238,I10532,I10594);
nor I_485 (I10625,I10577,I10382);
DFFARX1 I_486  ( .D(I10625), .CLK(I2350), .RSTB(I10252), .Q(I10229) );
nor I_487 (I10244,I10577,I10303);
not I_488 (I10670,I10577);
nor I_489 (I10687,I10450,I10670);
and I_490 (I10704,I10337,I10687);
or I_491 (I10721,I10532,I10704);
DFFARX1 I_492  ( .D(I10721), .CLK(I2350), .RSTB(I10252), .Q(I10217) );
nand I_493 (I10226,I10577,I10399);
nand I_494 (I10214,I10577,I10481);
not I_495 (I10813,I2357);
nand I_496 (I10830,I242939,I242936);
and I_497 (I10847,I10830,I242930);
DFFARX1 I_498  ( .D(I10847), .CLK(I2350), .RSTB(I10813), .Q(I10864) );
not I_499 (I10881,I10864);
nor I_500 (I10898,I242942,I242936);
or I_501 (I10796,I10898,I10864);
not I_502 (I10784,I10898);
DFFARX1 I_503  ( .D(I242954), .CLK(I2350), .RSTB(I10813), .Q(I10943) );
nor I_504 (I10960,I10943,I10898);
nand I_505 (I10977,I242945,I242927);
and I_506 (I10994,I10977,I242957);
DFFARX1 I_507  ( .D(I10994), .CLK(I2350), .RSTB(I10813), .Q(I11011) );
nor I_508 (I10793,I11011,I10864);
not I_509 (I11042,I11011);
nor I_510 (I11059,I10943,I11042);
DFFARX1 I_511  ( .D(I242933), .CLK(I2350), .RSTB(I10813), .Q(I11076) );
and I_512 (I11093,I11076,I242951);
or I_513 (I10802,I11093,I10898);
nand I_514 (I10781,I11093,I11059);
DFFARX1 I_515  ( .D(I242948), .CLK(I2350), .RSTB(I10813), .Q(I11138) );
and I_516 (I11155,I11138,I10881);
nor I_517 (I10799,I11093,I11155);
nor I_518 (I11186,I11138,I10943);
DFFARX1 I_519  ( .D(I11186), .CLK(I2350), .RSTB(I10813), .Q(I10790) );
nor I_520 (I10805,I11138,I10864);
not I_521 (I11231,I11138);
nor I_522 (I11248,I11011,I11231);
and I_523 (I11265,I10898,I11248);
or I_524 (I11282,I11093,I11265);
DFFARX1 I_525  ( .D(I11282), .CLK(I2350), .RSTB(I10813), .Q(I10778) );
nand I_526 (I10787,I11138,I10960);
nand I_527 (I10775,I11138,I11042);
not I_528 (I11374,I2357);
nand I_529 (I11391,I175495,I175486);
and I_530 (I11408,I11391,I175501);
DFFARX1 I_531  ( .D(I11408), .CLK(I2350), .RSTB(I11374), .Q(I11425) );
not I_532 (I11442,I11425);
nor I_533 (I11459,I175471,I175486);
or I_534 (I11357,I11459,I11425);
not I_535 (I11345,I11459);
DFFARX1 I_536  ( .D(I175474), .CLK(I2350), .RSTB(I11374), .Q(I11504) );
nor I_537 (I11521,I11504,I11459);
nand I_538 (I11538,I175492,I175489);
and I_539 (I11555,I11538,I175477);
DFFARX1 I_540  ( .D(I11555), .CLK(I2350), .RSTB(I11374), .Q(I11572) );
nor I_541 (I11354,I11572,I11425);
not I_542 (I11603,I11572);
nor I_543 (I11620,I11504,I11603);
DFFARX1 I_544  ( .D(I175498), .CLK(I2350), .RSTB(I11374), .Q(I11637) );
and I_545 (I11654,I11637,I175483);
or I_546 (I11363,I11654,I11459);
nand I_547 (I11342,I11654,I11620);
DFFARX1 I_548  ( .D(I175480), .CLK(I2350), .RSTB(I11374), .Q(I11699) );
and I_549 (I11716,I11699,I11442);
nor I_550 (I11360,I11654,I11716);
nor I_551 (I11747,I11699,I11504);
DFFARX1 I_552  ( .D(I11747), .CLK(I2350), .RSTB(I11374), .Q(I11351) );
nor I_553 (I11366,I11699,I11425);
not I_554 (I11792,I11699);
nor I_555 (I11809,I11572,I11792);
and I_556 (I11826,I11459,I11809);
or I_557 (I11843,I11654,I11826);
DFFARX1 I_558  ( .D(I11843), .CLK(I2350), .RSTB(I11374), .Q(I11339) );
nand I_559 (I11348,I11699,I11521);
nand I_560 (I11336,I11699,I11603);
not I_561 (I11935,I2357);
nand I_562 (I11952,I157594,I157585);
and I_563 (I11969,I11952,I157600);
DFFARX1 I_564  ( .D(I11969), .CLK(I2350), .RSTB(I11935), .Q(I11986) );
not I_565 (I12003,I11986);
nor I_566 (I12020,I157570,I157585);
or I_567 (I11918,I12020,I11986);
not I_568 (I11906,I12020);
DFFARX1 I_569  ( .D(I157573), .CLK(I2350), .RSTB(I11935), .Q(I12065) );
nor I_570 (I12082,I12065,I12020);
nand I_571 (I12099,I157591,I157588);
and I_572 (I12116,I12099,I157576);
DFFARX1 I_573  ( .D(I12116), .CLK(I2350), .RSTB(I11935), .Q(I12133) );
nor I_574 (I11915,I12133,I11986);
not I_575 (I12164,I12133);
nor I_576 (I12181,I12065,I12164);
DFFARX1 I_577  ( .D(I157597), .CLK(I2350), .RSTB(I11935), .Q(I12198) );
and I_578 (I12215,I12198,I157582);
or I_579 (I11924,I12215,I12020);
nand I_580 (I11903,I12215,I12181);
DFFARX1 I_581  ( .D(I157579), .CLK(I2350), .RSTB(I11935), .Q(I12260) );
and I_582 (I12277,I12260,I12003);
nor I_583 (I11921,I12215,I12277);
nor I_584 (I12308,I12260,I12065);
DFFARX1 I_585  ( .D(I12308), .CLK(I2350), .RSTB(I11935), .Q(I11912) );
nor I_586 (I11927,I12260,I11986);
not I_587 (I12353,I12260);
nor I_588 (I12370,I12133,I12353);
and I_589 (I12387,I12020,I12370);
or I_590 (I12404,I12215,I12387);
DFFARX1 I_591  ( .D(I12404), .CLK(I2350), .RSTB(I11935), .Q(I11900) );
nand I_592 (I11909,I12260,I12082);
nand I_593 (I11897,I12260,I12164);
not I_594 (I12496,I2357);
nand I_595 (I12513,I311780,I311783);
and I_596 (I12530,I12513,I311795);
DFFARX1 I_597  ( .D(I12530), .CLK(I2350), .RSTB(I12496), .Q(I12547) );
not I_598 (I12564,I12547);
nor I_599 (I12581,I311789,I311783);
or I_600 (I12479,I12581,I12547);
not I_601 (I12467,I12581);
DFFARX1 I_602  ( .D(I311792), .CLK(I2350), .RSTB(I12496), .Q(I12626) );
nor I_603 (I12643,I12626,I12581);
nand I_604 (I12660,I311786,I311804);
and I_605 (I12677,I12660,I311807);
DFFARX1 I_606  ( .D(I12677), .CLK(I2350), .RSTB(I12496), .Q(I12694) );
nor I_607 (I12476,I12694,I12547);
not I_608 (I12725,I12694);
nor I_609 (I12742,I12626,I12725);
DFFARX1 I_610  ( .D(I311777), .CLK(I2350), .RSTB(I12496), .Q(I12759) );
and I_611 (I12776,I12759,I311798);
or I_612 (I12485,I12776,I12581);
nand I_613 (I12464,I12776,I12742);
DFFARX1 I_614  ( .D(I311801), .CLK(I2350), .RSTB(I12496), .Q(I12821) );
and I_615 (I12838,I12821,I12564);
nor I_616 (I12482,I12776,I12838);
nor I_617 (I12869,I12821,I12626);
DFFARX1 I_618  ( .D(I12869), .CLK(I2350), .RSTB(I12496), .Q(I12473) );
nor I_619 (I12488,I12821,I12547);
not I_620 (I12914,I12821);
nor I_621 (I12931,I12694,I12914);
and I_622 (I12948,I12581,I12931);
or I_623 (I12965,I12776,I12948);
DFFARX1 I_624  ( .D(I12965), .CLK(I2350), .RSTB(I12496), .Q(I12461) );
nand I_625 (I12470,I12821,I12643);
nand I_626 (I12458,I12821,I12725);
not I_627 (I13057,I2357);
nand I_628 (I13074,I128779,I128782);
and I_629 (I13091,I13074,I128776);
DFFARX1 I_630  ( .D(I13091), .CLK(I2350), .RSTB(I13057), .Q(I13108) );
not I_631 (I13125,I13108);
nor I_632 (I13142,I128767,I128782);
or I_633 (I13040,I13142,I13108);
not I_634 (I13028,I13142);
DFFARX1 I_635  ( .D(I128755), .CLK(I2350), .RSTB(I13057), .Q(I13187) );
nor I_636 (I13204,I13187,I13142);
nand I_637 (I13221,I128764,I128758);
and I_638 (I13238,I13221,I128770);
DFFARX1 I_639  ( .D(I13238), .CLK(I2350), .RSTB(I13057), .Q(I13255) );
nor I_640 (I13037,I13255,I13108);
not I_641 (I13286,I13255);
nor I_642 (I13303,I13187,I13286);
DFFARX1 I_643  ( .D(I128785), .CLK(I2350), .RSTB(I13057), .Q(I13320) );
and I_644 (I13337,I13320,I128773);
or I_645 (I13046,I13337,I13142);
nand I_646 (I13025,I13337,I13303);
DFFARX1 I_647  ( .D(I128761), .CLK(I2350), .RSTB(I13057), .Q(I13382) );
and I_648 (I13399,I13382,I13125);
nor I_649 (I13043,I13337,I13399);
nor I_650 (I13430,I13382,I13187);
DFFARX1 I_651  ( .D(I13430), .CLK(I2350), .RSTB(I13057), .Q(I13034) );
nor I_652 (I13049,I13382,I13108);
not I_653 (I13475,I13382);
nor I_654 (I13492,I13255,I13475);
and I_655 (I13509,I13142,I13492);
or I_656 (I13526,I13337,I13509);
DFFARX1 I_657  ( .D(I13526), .CLK(I2350), .RSTB(I13057), .Q(I13022) );
nand I_658 (I13031,I13382,I13204);
nand I_659 (I13019,I13382,I13286);
not I_660 (I13618,I2357);
nand I_661 (I13635,I336376,I336379);
and I_662 (I13652,I13635,I336385);
DFFARX1 I_663  ( .D(I13652), .CLK(I2350), .RSTB(I13618), .Q(I13669) );
not I_664 (I13686,I13669);
nor I_665 (I13703,I336397,I336379);
or I_666 (I13601,I13703,I13669);
not I_667 (I13589,I13703);
DFFARX1 I_668  ( .D(I336406), .CLK(I2350), .RSTB(I13618), .Q(I13748) );
nor I_669 (I13765,I13748,I13703);
nand I_670 (I13782,I336394,I336391);
and I_671 (I13799,I13782,I336403);
DFFARX1 I_672  ( .D(I13799), .CLK(I2350), .RSTB(I13618), .Q(I13816) );
nor I_673 (I13598,I13816,I13669);
not I_674 (I13847,I13816);
nor I_675 (I13864,I13748,I13847);
DFFARX1 I_676  ( .D(I336400), .CLK(I2350), .RSTB(I13618), .Q(I13881) );
and I_677 (I13898,I13881,I336388);
or I_678 (I13607,I13898,I13703);
nand I_679 (I13586,I13898,I13864);
DFFARX1 I_680  ( .D(I336382), .CLK(I2350), .RSTB(I13618), .Q(I13943) );
and I_681 (I13960,I13943,I13686);
nor I_682 (I13604,I13898,I13960);
nor I_683 (I13991,I13943,I13748);
DFFARX1 I_684  ( .D(I13991), .CLK(I2350), .RSTB(I13618), .Q(I13595) );
nor I_685 (I13610,I13943,I13669);
not I_686 (I14036,I13943);
nor I_687 (I14053,I13816,I14036);
and I_688 (I14070,I13703,I14053);
or I_689 (I14087,I13898,I14070);
DFFARX1 I_690  ( .D(I14087), .CLK(I2350), .RSTB(I13618), .Q(I13583) );
nand I_691 (I13592,I13943,I13765);
nand I_692 (I13580,I13943,I13847);
not I_693 (I14179,I2357);
nand I_694 (I14196,I195969,I195960);
and I_695 (I14213,I14196,I195963);
DFFARX1 I_696  ( .D(I14213), .CLK(I2350), .RSTB(I14179), .Q(I14230) );
not I_697 (I14247,I14230);
nor I_698 (I14264,I195939,I195960);
or I_699 (I14162,I14264,I14230);
not I_700 (I14150,I14264);
DFFARX1 I_701  ( .D(I195954), .CLK(I2350), .RSTB(I14179), .Q(I14309) );
nor I_702 (I14326,I14309,I14264);
nand I_703 (I14343,I195942,I195957);
and I_704 (I14360,I14343,I195951);
DFFARX1 I_705  ( .D(I14360), .CLK(I2350), .RSTB(I14179), .Q(I14377) );
nor I_706 (I14159,I14377,I14230);
not I_707 (I14408,I14377);
nor I_708 (I14425,I14309,I14408);
DFFARX1 I_709  ( .D(I195966), .CLK(I2350), .RSTB(I14179), .Q(I14442) );
and I_710 (I14459,I14442,I195945);
or I_711 (I14168,I14459,I14264);
nand I_712 (I14147,I14459,I14425);
DFFARX1 I_713  ( .D(I195948), .CLK(I2350), .RSTB(I14179), .Q(I14504) );
and I_714 (I14521,I14504,I14247);
nor I_715 (I14165,I14459,I14521);
nor I_716 (I14552,I14504,I14309);
DFFARX1 I_717  ( .D(I14552), .CLK(I2350), .RSTB(I14179), .Q(I14156) );
nor I_718 (I14171,I14504,I14230);
not I_719 (I14597,I14504);
nor I_720 (I14614,I14377,I14597);
and I_721 (I14631,I14264,I14614);
or I_722 (I14648,I14459,I14631);
DFFARX1 I_723  ( .D(I14648), .CLK(I2350), .RSTB(I14179), .Q(I14144) );
nand I_724 (I14153,I14504,I14326);
nand I_725 (I14141,I14504,I14408);
not I_726 (I14740,I2357);
nand I_727 (I14757,I244673,I244670);
and I_728 (I14774,I14757,I244664);
DFFARX1 I_729  ( .D(I14774), .CLK(I2350), .RSTB(I14740), .Q(I14791) );
not I_730 (I14808,I14791);
nor I_731 (I14825,I244676,I244670);
or I_732 (I14723,I14825,I14791);
not I_733 (I14711,I14825);
DFFARX1 I_734  ( .D(I244688), .CLK(I2350), .RSTB(I14740), .Q(I14870) );
nor I_735 (I14887,I14870,I14825);
nand I_736 (I14904,I244679,I244661);
and I_737 (I14921,I14904,I244691);
DFFARX1 I_738  ( .D(I14921), .CLK(I2350), .RSTB(I14740), .Q(I14938) );
nor I_739 (I14720,I14938,I14791);
not I_740 (I14969,I14938);
nor I_741 (I14986,I14870,I14969);
DFFARX1 I_742  ( .D(I244667), .CLK(I2350), .RSTB(I14740), .Q(I15003) );
and I_743 (I15020,I15003,I244685);
or I_744 (I14729,I15020,I14825);
nand I_745 (I14708,I15020,I14986);
DFFARX1 I_746  ( .D(I244682), .CLK(I2350), .RSTB(I14740), .Q(I15065) );
and I_747 (I15082,I15065,I14808);
nor I_748 (I14726,I15020,I15082);
nor I_749 (I15113,I15065,I14870);
DFFARX1 I_750  ( .D(I15113), .CLK(I2350), .RSTB(I14740), .Q(I14717) );
nor I_751 (I14732,I15065,I14791);
not I_752 (I15158,I15065);
nor I_753 (I15175,I14938,I15158);
and I_754 (I15192,I14825,I15175);
or I_755 (I15209,I15020,I15192);
DFFARX1 I_756  ( .D(I15209), .CLK(I2350), .RSTB(I14740), .Q(I14705) );
nand I_757 (I14714,I15065,I14887);
nand I_758 (I14702,I15065,I14969);
not I_759 (I15301,I2357);
nand I_760 (I15318,I390870,I390891);
and I_761 (I15335,I15318,I390879);
DFFARX1 I_762  ( .D(I15335), .CLK(I2350), .RSTB(I15301), .Q(I15352) );
not I_763 (I15369,I15352);
nor I_764 (I15386,I390885,I390891);
or I_765 (I15284,I15386,I15352);
not I_766 (I15272,I15386);
DFFARX1 I_767  ( .D(I390873), .CLK(I2350), .RSTB(I15301), .Q(I15431) );
nor I_768 (I15448,I15431,I15386);
nand I_769 (I15465,I390864,I390882);
and I_770 (I15482,I15465,I390876);
DFFARX1 I_771  ( .D(I15482), .CLK(I2350), .RSTB(I15301), .Q(I15499) );
nor I_772 (I15281,I15499,I15352);
not I_773 (I15530,I15499);
nor I_774 (I15547,I15431,I15530);
DFFARX1 I_775  ( .D(I390888), .CLK(I2350), .RSTB(I15301), .Q(I15564) );
and I_776 (I15581,I15564,I390861);
or I_777 (I15290,I15581,I15386);
nand I_778 (I15269,I15581,I15547);
DFFARX1 I_779  ( .D(I390867), .CLK(I2350), .RSTB(I15301), .Q(I15626) );
and I_780 (I15643,I15626,I15369);
nor I_781 (I15287,I15581,I15643);
nor I_782 (I15674,I15626,I15431);
DFFARX1 I_783  ( .D(I15674), .CLK(I2350), .RSTB(I15301), .Q(I15278) );
nor I_784 (I15293,I15626,I15352);
not I_785 (I15719,I15626);
nor I_786 (I15736,I15499,I15719);
and I_787 (I15753,I15386,I15736);
or I_788 (I15770,I15581,I15753);
DFFARX1 I_789  ( .D(I15770), .CLK(I2350), .RSTB(I15301), .Q(I15266) );
nand I_790 (I15275,I15626,I15448);
nand I_791 (I15263,I15626,I15530);
not I_792 (I15862,I2357);
nand I_793 (I15879,I326673,I326661);
and I_794 (I15896,I15879,I326658);
DFFARX1 I_795  ( .D(I15896), .CLK(I2350), .RSTB(I15862), .Q(I15913) );
not I_796 (I15930,I15913);
nor I_797 (I15947,I326679,I326661);
or I_798 (I15845,I15947,I15913);
not I_799 (I15833,I15947);
DFFARX1 I_800  ( .D(I326682), .CLK(I2350), .RSTB(I15862), .Q(I15992) );
nor I_801 (I16009,I15992,I15947);
nand I_802 (I16026,I326652,I326670);
and I_803 (I16043,I16026,I326667);
DFFARX1 I_804  ( .D(I16043), .CLK(I2350), .RSTB(I15862), .Q(I16060) );
nor I_805 (I15842,I16060,I15913);
not I_806 (I16091,I16060);
nor I_807 (I16108,I15992,I16091);
DFFARX1 I_808  ( .D(I326676), .CLK(I2350), .RSTB(I15862), .Q(I16125) );
and I_809 (I16142,I16125,I326664);
or I_810 (I15851,I16142,I15947);
nand I_811 (I15830,I16142,I16108);
DFFARX1 I_812  ( .D(I326655), .CLK(I2350), .RSTB(I15862), .Q(I16187) );
and I_813 (I16204,I16187,I15930);
nor I_814 (I15848,I16142,I16204);
nor I_815 (I16235,I16187,I15992);
DFFARX1 I_816  ( .D(I16235), .CLK(I2350), .RSTB(I15862), .Q(I15839) );
nor I_817 (I15854,I16187,I15913);
not I_818 (I16280,I16187);
nor I_819 (I16297,I16060,I16280);
and I_820 (I16314,I15947,I16297);
or I_821 (I16331,I16142,I16314);
DFFARX1 I_822  ( .D(I16331), .CLK(I2350), .RSTB(I15862), .Q(I15827) );
nand I_823 (I15836,I16187,I16009);
nand I_824 (I15824,I16187,I16091);
not I_825 (I16423,I2357);
nand I_826 (I16440,I224393,I224384);
and I_827 (I16457,I16440,I224387);
DFFARX1 I_828  ( .D(I16457), .CLK(I2350), .RSTB(I16423), .Q(I16474) );
not I_829 (I16491,I16474);
nor I_830 (I16508,I224363,I224384);
or I_831 (I16406,I16508,I16474);
not I_832 (I16394,I16508);
DFFARX1 I_833  ( .D(I224378), .CLK(I2350), .RSTB(I16423), .Q(I16553) );
nor I_834 (I16570,I16553,I16508);
nand I_835 (I16587,I224366,I224381);
and I_836 (I16604,I16587,I224375);
DFFARX1 I_837  ( .D(I16604), .CLK(I2350), .RSTB(I16423), .Q(I16621) );
nor I_838 (I16403,I16621,I16474);
not I_839 (I16652,I16621);
nor I_840 (I16669,I16553,I16652);
DFFARX1 I_841  ( .D(I224390), .CLK(I2350), .RSTB(I16423), .Q(I16686) );
and I_842 (I16703,I16686,I224369);
or I_843 (I16412,I16703,I16508);
nand I_844 (I16391,I16703,I16669);
DFFARX1 I_845  ( .D(I224372), .CLK(I2350), .RSTB(I16423), .Q(I16748) );
and I_846 (I16765,I16748,I16491);
nor I_847 (I16409,I16703,I16765);
nor I_848 (I16796,I16748,I16553);
DFFARX1 I_849  ( .D(I16796), .CLK(I2350), .RSTB(I16423), .Q(I16400) );
nor I_850 (I16415,I16748,I16474);
not I_851 (I16841,I16748);
nor I_852 (I16858,I16621,I16841);
and I_853 (I16875,I16508,I16858);
or I_854 (I16892,I16703,I16875);
DFFARX1 I_855  ( .D(I16892), .CLK(I2350), .RSTB(I16423), .Q(I16388) );
nand I_856 (I16397,I16748,I16570);
nand I_857 (I16385,I16748,I16652);
not I_858 (I16984,I2357);
nand I_859 (I17001,I78915,I78918);
and I_860 (I17018,I17001,I78900);
DFFARX1 I_861  ( .D(I17018), .CLK(I2350), .RSTB(I16984), .Q(I17035) );
not I_862 (I17052,I17035);
nor I_863 (I17069,I78897,I78918);
or I_864 (I16967,I17069,I17035);
not I_865 (I16955,I17069);
DFFARX1 I_866  ( .D(I78921), .CLK(I2350), .RSTB(I16984), .Q(I17114) );
nor I_867 (I17131,I17114,I17069);
nand I_868 (I17148,I78906,I78912);
and I_869 (I17165,I17148,I78924);
DFFARX1 I_870  ( .D(I17165), .CLK(I2350), .RSTB(I16984), .Q(I17182) );
nor I_871 (I16964,I17182,I17035);
not I_872 (I17213,I17182);
nor I_873 (I17230,I17114,I17213);
DFFARX1 I_874  ( .D(I78903), .CLK(I2350), .RSTB(I16984), .Q(I17247) );
and I_875 (I17264,I17247,I78894);
or I_876 (I16973,I17264,I17069);
nand I_877 (I16952,I17264,I17230);
DFFARX1 I_878  ( .D(I78909), .CLK(I2350), .RSTB(I16984), .Q(I17309) );
and I_879 (I17326,I17309,I17052);
nor I_880 (I16970,I17264,I17326);
nor I_881 (I17357,I17309,I17114);
DFFARX1 I_882  ( .D(I17357), .CLK(I2350), .RSTB(I16984), .Q(I16961) );
nor I_883 (I16976,I17309,I17035);
not I_884 (I17402,I17309);
nor I_885 (I17419,I17182,I17402);
and I_886 (I17436,I17069,I17419);
or I_887 (I17453,I17264,I17436);
DFFARX1 I_888  ( .D(I17453), .CLK(I2350), .RSTB(I16984), .Q(I16949) );
nand I_889 (I16958,I17309,I17131);
nand I_890 (I16946,I17309,I17213);
not I_891 (I17545,I2357);
nand I_892 (I17562,I197907,I197898);
and I_893 (I17579,I17562,I197901);
DFFARX1 I_894  ( .D(I17579), .CLK(I2350), .RSTB(I17545), .Q(I17596) );
not I_895 (I17613,I17596);
nor I_896 (I17630,I197877,I197898);
or I_897 (I17528,I17630,I17596);
not I_898 (I17516,I17630);
DFFARX1 I_899  ( .D(I197892), .CLK(I2350), .RSTB(I17545), .Q(I17675) );
nor I_900 (I17692,I17675,I17630);
nand I_901 (I17709,I197880,I197895);
and I_902 (I17726,I17709,I197889);
DFFARX1 I_903  ( .D(I17726), .CLK(I2350), .RSTB(I17545), .Q(I17743) );
nor I_904 (I17525,I17743,I17596);
not I_905 (I17774,I17743);
nor I_906 (I17791,I17675,I17774);
DFFARX1 I_907  ( .D(I197904), .CLK(I2350), .RSTB(I17545), .Q(I17808) );
and I_908 (I17825,I17808,I197883);
or I_909 (I17534,I17825,I17630);
nand I_910 (I17513,I17825,I17791);
DFFARX1 I_911  ( .D(I197886), .CLK(I2350), .RSTB(I17545), .Q(I17870) );
and I_912 (I17887,I17870,I17613);
nor I_913 (I17531,I17825,I17887);
nor I_914 (I17918,I17870,I17675);
DFFARX1 I_915  ( .D(I17918), .CLK(I2350), .RSTB(I17545), .Q(I17522) );
nor I_916 (I17537,I17870,I17596);
not I_917 (I17963,I17870);
nor I_918 (I17980,I17743,I17963);
and I_919 (I17997,I17630,I17980);
or I_920 (I18014,I17825,I17997);
DFFARX1 I_921  ( .D(I18014), .CLK(I2350), .RSTB(I17545), .Q(I17510) );
nand I_922 (I17519,I17870,I17692);
nand I_923 (I17507,I17870,I17774);
not I_924 (I18106,I2357);
nand I_925 (I18123,I306425,I306428);
and I_926 (I18140,I18123,I306440);
DFFARX1 I_927  ( .D(I18140), .CLK(I2350), .RSTB(I18106), .Q(I18157) );
not I_928 (I18174,I18157);
nor I_929 (I18191,I306434,I306428);
or I_930 (I18089,I18191,I18157);
not I_931 (I18077,I18191);
DFFARX1 I_932  ( .D(I306437), .CLK(I2350), .RSTB(I18106), .Q(I18236) );
nor I_933 (I18253,I18236,I18191);
nand I_934 (I18270,I306431,I306449);
and I_935 (I18287,I18270,I306452);
DFFARX1 I_936  ( .D(I18287), .CLK(I2350), .RSTB(I18106), .Q(I18304) );
nor I_937 (I18086,I18304,I18157);
not I_938 (I18335,I18304);
nor I_939 (I18352,I18236,I18335);
DFFARX1 I_940  ( .D(I306422), .CLK(I2350), .RSTB(I18106), .Q(I18369) );
and I_941 (I18386,I18369,I306443);
or I_942 (I18095,I18386,I18191);
nand I_943 (I18074,I18386,I18352);
DFFARX1 I_944  ( .D(I306446), .CLK(I2350), .RSTB(I18106), .Q(I18431) );
and I_945 (I18448,I18431,I18174);
nor I_946 (I18092,I18386,I18448);
nor I_947 (I18479,I18431,I18236);
DFFARX1 I_948  ( .D(I18479), .CLK(I2350), .RSTB(I18106), .Q(I18083) );
nor I_949 (I18098,I18431,I18157);
not I_950 (I18524,I18431);
nor I_951 (I18541,I18304,I18524);
and I_952 (I18558,I18191,I18541);
or I_953 (I18575,I18386,I18558);
DFFARX1 I_954  ( .D(I18575), .CLK(I2350), .RSTB(I18106), .Q(I18071) );
nand I_955 (I18080,I18431,I18253);
nand I_956 (I18068,I18431,I18335);
not I_957 (I18667,I2357);
nand I_958 (I18684,I278460,I278463);
and I_959 (I18701,I18684,I278475);
DFFARX1 I_960  ( .D(I18701), .CLK(I2350), .RSTB(I18667), .Q(I18718) );
not I_961 (I18735,I18718);
nor I_962 (I18752,I278469,I278463);
or I_963 (I18650,I18752,I18718);
not I_964 (I18638,I18752);
DFFARX1 I_965  ( .D(I278472), .CLK(I2350), .RSTB(I18667), .Q(I18797) );
nor I_966 (I18814,I18797,I18752);
nand I_967 (I18831,I278466,I278484);
and I_968 (I18848,I18831,I278487);
DFFARX1 I_969  ( .D(I18848), .CLK(I2350), .RSTB(I18667), .Q(I18865) );
nor I_970 (I18647,I18865,I18718);
not I_971 (I18896,I18865);
nor I_972 (I18913,I18797,I18896);
DFFARX1 I_973  ( .D(I278457), .CLK(I2350), .RSTB(I18667), .Q(I18930) );
and I_974 (I18947,I18930,I278478);
or I_975 (I18656,I18947,I18752);
nand I_976 (I18635,I18947,I18913);
DFFARX1 I_977  ( .D(I278481), .CLK(I2350), .RSTB(I18667), .Q(I18992) );
and I_978 (I19009,I18992,I18735);
nor I_979 (I18653,I18947,I19009);
nor I_980 (I19040,I18992,I18797);
DFFARX1 I_981  ( .D(I19040), .CLK(I2350), .RSTB(I18667), .Q(I18644) );
nor I_982 (I18659,I18992,I18718);
not I_983 (I19085,I18992);
nor I_984 (I19102,I18865,I19085);
and I_985 (I19119,I18752,I19102);
or I_986 (I19136,I18947,I19119);
DFFARX1 I_987  ( .D(I19136), .CLK(I2350), .RSTB(I18667), .Q(I18632) );
nand I_988 (I18641,I18992,I18814);
nand I_989 (I18629,I18992,I18896);
not I_990 (I19228,I2357);
nand I_991 (I19245,I382200,I382221);
and I_992 (I19262,I19245,I382209);
DFFARX1 I_993  ( .D(I19262), .CLK(I2350), .RSTB(I19228), .Q(I19279) );
not I_994 (I19296,I19279);
nor I_995 (I19313,I382215,I382221);
or I_996 (I19211,I19313,I19279);
not I_997 (I19199,I19313);
DFFARX1 I_998  ( .D(I382203), .CLK(I2350), .RSTB(I19228), .Q(I19358) );
nor I_999 (I19375,I19358,I19313);
nand I_1000 (I19392,I382194,I382212);
and I_1001 (I19409,I19392,I382206);
DFFARX1 I_1002  ( .D(I19409), .CLK(I2350), .RSTB(I19228), .Q(I19426) );
nor I_1003 (I19208,I19426,I19279);
not I_1004 (I19457,I19426);
nor I_1005 (I19474,I19358,I19457);
DFFARX1 I_1006  ( .D(I382218), .CLK(I2350), .RSTB(I19228), .Q(I19491) );
and I_1007 (I19508,I19491,I382191);
or I_1008 (I19217,I19508,I19313);
nand I_1009 (I19196,I19508,I19474);
DFFARX1 I_1010  ( .D(I382197), .CLK(I2350), .RSTB(I19228), .Q(I19553) );
and I_1011 (I19570,I19553,I19296);
nor I_1012 (I19214,I19508,I19570);
nor I_1013 (I19601,I19553,I19358);
DFFARX1 I_1014  ( .D(I19601), .CLK(I2350), .RSTB(I19228), .Q(I19205) );
nor I_1015 (I19220,I19553,I19279);
not I_1016 (I19646,I19553);
nor I_1017 (I19663,I19426,I19646);
and I_1018 (I19680,I19313,I19663);
or I_1019 (I19697,I19508,I19680);
DFFARX1 I_1020  ( .D(I19697), .CLK(I2350), .RSTB(I19228), .Q(I19193) );
nand I_1021 (I19202,I19553,I19375);
nand I_1022 (I19190,I19553,I19457);
not I_1023 (I19789,I2357);
nand I_1024 (I19806,I109911,I109908);
and I_1025 (I19823,I19806,I109905);
DFFARX1 I_1026  ( .D(I19823), .CLK(I2350), .RSTB(I19789), .Q(I19840) );
not I_1027 (I19857,I19840);
nor I_1028 (I19874,I109929,I109908);
or I_1029 (I19772,I19874,I19840);
not I_1030 (I19760,I19874);
DFFARX1 I_1031  ( .D(I109923), .CLK(I2350), .RSTB(I19789), .Q(I19919) );
nor I_1032 (I19936,I19919,I19874);
nand I_1033 (I19953,I109902,I109914);
and I_1034 (I19970,I19953,I109917);
DFFARX1 I_1035  ( .D(I19970), .CLK(I2350), .RSTB(I19789), .Q(I19987) );
nor I_1036 (I19769,I19987,I19840);
not I_1037 (I20018,I19987);
nor I_1038 (I20035,I19919,I20018);
DFFARX1 I_1039  ( .D(I109926), .CLK(I2350), .RSTB(I19789), .Q(I20052) );
and I_1040 (I20069,I20052,I109932);
or I_1041 (I19778,I20069,I19874);
nand I_1042 (I19757,I20069,I20035);
DFFARX1 I_1043  ( .D(I109920), .CLK(I2350), .RSTB(I19789), .Q(I20114) );
and I_1044 (I20131,I20114,I19857);
nor I_1045 (I19775,I20069,I20131);
nor I_1046 (I20162,I20114,I19919);
DFFARX1 I_1047  ( .D(I20162), .CLK(I2350), .RSTB(I19789), .Q(I19766) );
nor I_1048 (I19781,I20114,I19840);
not I_1049 (I20207,I20114);
nor I_1050 (I20224,I19987,I20207);
and I_1051 (I20241,I19874,I20224);
or I_1052 (I20258,I20069,I20241);
DFFARX1 I_1053  ( .D(I20258), .CLK(I2350), .RSTB(I19789), .Q(I19754) );
nand I_1054 (I19763,I20114,I19936);
nand I_1055 (I19751,I20114,I20018);
not I_1056 (I20350,I2357);
nand I_1057 (I20367,I226331,I226322);
and I_1058 (I20384,I20367,I226325);
DFFARX1 I_1059  ( .D(I20384), .CLK(I2350), .RSTB(I20350), .Q(I20401) );
not I_1060 (I20418,I20401);
nor I_1061 (I20435,I226301,I226322);
or I_1062 (I20333,I20435,I20401);
not I_1063 (I20321,I20435);
DFFARX1 I_1064  ( .D(I226316), .CLK(I2350), .RSTB(I20350), .Q(I20480) );
nor I_1065 (I20497,I20480,I20435);
nand I_1066 (I20514,I226304,I226319);
and I_1067 (I20531,I20514,I226313);
DFFARX1 I_1068  ( .D(I20531), .CLK(I2350), .RSTB(I20350), .Q(I20548) );
nor I_1069 (I20330,I20548,I20401);
not I_1070 (I20579,I20548);
nor I_1071 (I20596,I20480,I20579);
DFFARX1 I_1072  ( .D(I226328), .CLK(I2350), .RSTB(I20350), .Q(I20613) );
and I_1073 (I20630,I20613,I226307);
or I_1074 (I20339,I20630,I20435);
nand I_1075 (I20318,I20630,I20596);
DFFARX1 I_1076  ( .D(I226310), .CLK(I2350), .RSTB(I20350), .Q(I20675) );
and I_1077 (I20692,I20675,I20418);
nor I_1078 (I20336,I20630,I20692);
nor I_1079 (I20723,I20675,I20480);
DFFARX1 I_1080  ( .D(I20723), .CLK(I2350), .RSTB(I20350), .Q(I20327) );
nor I_1081 (I20342,I20675,I20401);
not I_1082 (I20768,I20675);
nor I_1083 (I20785,I20548,I20768);
and I_1084 (I20802,I20435,I20785);
or I_1085 (I20819,I20630,I20802);
DFFARX1 I_1086  ( .D(I20819), .CLK(I2350), .RSTB(I20350), .Q(I20315) );
nand I_1087 (I20324,I20675,I20497);
nand I_1088 (I20312,I20675,I20579);
not I_1089 (I20911,I2357);
nand I_1090 (I20928,I353359,I353362);
and I_1091 (I20945,I20928,I353368);
DFFARX1 I_1092  ( .D(I20945), .CLK(I2350), .RSTB(I20911), .Q(I20962) );
not I_1093 (I20979,I20962);
nor I_1094 (I20996,I353380,I353362);
or I_1095 (I20894,I20996,I20962);
not I_1096 (I20882,I20996);
DFFARX1 I_1097  ( .D(I353389), .CLK(I2350), .RSTB(I20911), .Q(I21041) );
nor I_1098 (I21058,I21041,I20996);
nand I_1099 (I21075,I353377,I353374);
and I_1100 (I21092,I21075,I353386);
DFFARX1 I_1101  ( .D(I21092), .CLK(I2350), .RSTB(I20911), .Q(I21109) );
nor I_1102 (I20891,I21109,I20962);
not I_1103 (I21140,I21109);
nor I_1104 (I21157,I21041,I21140);
DFFARX1 I_1105  ( .D(I353383), .CLK(I2350), .RSTB(I20911), .Q(I21174) );
and I_1106 (I21191,I21174,I353371);
or I_1107 (I20900,I21191,I20996);
nand I_1108 (I20879,I21191,I21157);
DFFARX1 I_1109  ( .D(I353365), .CLK(I2350), .RSTB(I20911), .Q(I21236) );
and I_1110 (I21253,I21236,I20979);
nor I_1111 (I20897,I21191,I21253);
nor I_1112 (I21284,I21236,I21041);
DFFARX1 I_1113  ( .D(I21284), .CLK(I2350), .RSTB(I20911), .Q(I20888) );
nor I_1114 (I20903,I21236,I20962);
not I_1115 (I21329,I21236);
nor I_1116 (I21346,I21109,I21329);
and I_1117 (I21363,I20996,I21346);
or I_1118 (I21380,I21191,I21363);
DFFARX1 I_1119  ( .D(I21380), .CLK(I2350), .RSTB(I20911), .Q(I20876) );
nand I_1120 (I20885,I21236,I21058);
nand I_1121 (I20873,I21236,I21140);
not I_1122 (I21472,I2357);
nand I_1123 (I21489,I280245,I280248);
and I_1124 (I21506,I21489,I280260);
DFFARX1 I_1125  ( .D(I21506), .CLK(I2350), .RSTB(I21472), .Q(I21523) );
not I_1126 (I21540,I21523);
nor I_1127 (I21557,I280254,I280248);
or I_1128 (I21455,I21557,I21523);
not I_1129 (I21443,I21557);
DFFARX1 I_1130  ( .D(I280257), .CLK(I2350), .RSTB(I21472), .Q(I21602) );
nor I_1131 (I21619,I21602,I21557);
nand I_1132 (I21636,I280251,I280269);
and I_1133 (I21653,I21636,I280272);
DFFARX1 I_1134  ( .D(I21653), .CLK(I2350), .RSTB(I21472), .Q(I21670) );
nor I_1135 (I21452,I21670,I21523);
not I_1136 (I21701,I21670);
nor I_1137 (I21718,I21602,I21701);
DFFARX1 I_1138  ( .D(I280242), .CLK(I2350), .RSTB(I21472), .Q(I21735) );
and I_1139 (I21752,I21735,I280263);
or I_1140 (I21461,I21752,I21557);
nand I_1141 (I21440,I21752,I21718);
DFFARX1 I_1142  ( .D(I280266), .CLK(I2350), .RSTB(I21472), .Q(I21797) );
and I_1143 (I21814,I21797,I21540);
nor I_1144 (I21458,I21752,I21814);
nor I_1145 (I21845,I21797,I21602);
DFFARX1 I_1146  ( .D(I21845), .CLK(I2350), .RSTB(I21472), .Q(I21449) );
nor I_1147 (I21464,I21797,I21523);
not I_1148 (I21890,I21797);
nor I_1149 (I21907,I21670,I21890);
and I_1150 (I21924,I21557,I21907);
or I_1151 (I21941,I21752,I21924);
DFFARX1 I_1152  ( .D(I21941), .CLK(I2350), .RSTB(I21472), .Q(I21437) );
nand I_1153 (I21446,I21797,I21619);
nand I_1154 (I21434,I21797,I21701);
not I_1155 (I22033,I2357);
nand I_1156 (I22050,I237066,I237060);
and I_1157 (I22067,I22050,I237072);
DFFARX1 I_1158  ( .D(I22067), .CLK(I2350), .RSTB(I22033), .Q(I22084) );
not I_1159 (I22101,I22084);
nor I_1160 (I22118,I237069,I237060);
or I_1161 (I22016,I22118,I22084);
not I_1162 (I22004,I22118);
DFFARX1 I_1163  ( .D(I237048), .CLK(I2350), .RSTB(I22033), .Q(I22163) );
nor I_1164 (I22180,I22163,I22118);
nand I_1165 (I22197,I237054,I237063);
and I_1166 (I22214,I22197,I237051);
DFFARX1 I_1167  ( .D(I22214), .CLK(I2350), .RSTB(I22033), .Q(I22231) );
nor I_1168 (I22013,I22231,I22084);
not I_1169 (I22262,I22231);
nor I_1170 (I22279,I22163,I22262);
DFFARX1 I_1171  ( .D(I237075), .CLK(I2350), .RSTB(I22033), .Q(I22296) );
and I_1172 (I22313,I22296,I237045);
or I_1173 (I22022,I22313,I22118);
nand I_1174 (I22001,I22313,I22279);
DFFARX1 I_1175  ( .D(I237057), .CLK(I2350), .RSTB(I22033), .Q(I22358) );
and I_1176 (I22375,I22358,I22101);
nor I_1177 (I22019,I22313,I22375);
nor I_1178 (I22406,I22358,I22163);
DFFARX1 I_1179  ( .D(I22406), .CLK(I2350), .RSTB(I22033), .Q(I22010) );
nor I_1180 (I22025,I22358,I22084);
not I_1181 (I22451,I22358);
nor I_1182 (I22468,I22231,I22451);
and I_1183 (I22485,I22118,I22468);
or I_1184 (I22502,I22313,I22485);
DFFARX1 I_1185  ( .D(I22502), .CLK(I2350), .RSTB(I22033), .Q(I21998) );
nand I_1186 (I22007,I22358,I22180);
nand I_1187 (I21995,I22358,I22262);
not I_1188 (I22594,I2357);
nand I_1189 (I22611,I249297,I249294);
and I_1190 (I22628,I22611,I249288);
DFFARX1 I_1191  ( .D(I22628), .CLK(I2350), .RSTB(I22594), .Q(I22645) );
not I_1192 (I22662,I22645);
nor I_1193 (I22679,I249300,I249294);
or I_1194 (I22577,I22679,I22645);
not I_1195 (I22565,I22679);
DFFARX1 I_1196  ( .D(I249312), .CLK(I2350), .RSTB(I22594), .Q(I22724) );
nor I_1197 (I22741,I22724,I22679);
nand I_1198 (I22758,I249303,I249285);
and I_1199 (I22775,I22758,I249315);
DFFARX1 I_1200  ( .D(I22775), .CLK(I2350), .RSTB(I22594), .Q(I22792) );
nor I_1201 (I22574,I22792,I22645);
not I_1202 (I22823,I22792);
nor I_1203 (I22840,I22724,I22823);
DFFARX1 I_1204  ( .D(I249291), .CLK(I2350), .RSTB(I22594), .Q(I22857) );
and I_1205 (I22874,I22857,I249309);
or I_1206 (I22583,I22874,I22679);
nand I_1207 (I22562,I22874,I22840);
DFFARX1 I_1208  ( .D(I249306), .CLK(I2350), .RSTB(I22594), .Q(I22919) );
and I_1209 (I22936,I22919,I22662);
nor I_1210 (I22580,I22874,I22936);
nor I_1211 (I22967,I22919,I22724);
DFFARX1 I_1212  ( .D(I22967), .CLK(I2350), .RSTB(I22594), .Q(I22571) );
nor I_1213 (I22586,I22919,I22645);
not I_1214 (I23012,I22919);
nor I_1215 (I23029,I22792,I23012);
and I_1216 (I23046,I22679,I23029);
or I_1217 (I23063,I22874,I23046);
DFFARX1 I_1218  ( .D(I23063), .CLK(I2350), .RSTB(I22594), .Q(I22559) );
nand I_1219 (I22568,I22919,I22741);
nand I_1220 (I22556,I22919,I22823);
not I_1221 (I23155,I2357);
nand I_1222 (I23172,I231499,I231490);
and I_1223 (I23189,I23172,I231493);
DFFARX1 I_1224  ( .D(I23189), .CLK(I2350), .RSTB(I23155), .Q(I23206) );
not I_1225 (I23223,I23206);
nor I_1226 (I23240,I231469,I231490);
or I_1227 (I23138,I23240,I23206);
not I_1228 (I23126,I23240);
DFFARX1 I_1229  ( .D(I231484), .CLK(I2350), .RSTB(I23155), .Q(I23285) );
nor I_1230 (I23302,I23285,I23240);
nand I_1231 (I23319,I231472,I231487);
and I_1232 (I23336,I23319,I231481);
DFFARX1 I_1233  ( .D(I23336), .CLK(I2350), .RSTB(I23155), .Q(I23353) );
nor I_1234 (I23135,I23353,I23206);
not I_1235 (I23384,I23353);
nor I_1236 (I23401,I23285,I23384);
DFFARX1 I_1237  ( .D(I231496), .CLK(I2350), .RSTB(I23155), .Q(I23418) );
and I_1238 (I23435,I23418,I231475);
or I_1239 (I23144,I23435,I23240);
nand I_1240 (I23123,I23435,I23401);
DFFARX1 I_1241  ( .D(I231478), .CLK(I2350), .RSTB(I23155), .Q(I23480) );
and I_1242 (I23497,I23480,I23223);
nor I_1243 (I23141,I23435,I23497);
nor I_1244 (I23528,I23480,I23285);
DFFARX1 I_1245  ( .D(I23528), .CLK(I2350), .RSTB(I23155), .Q(I23132) );
nor I_1246 (I23147,I23480,I23206);
not I_1247 (I23573,I23480);
nor I_1248 (I23590,I23353,I23573);
and I_1249 (I23607,I23240,I23590);
or I_1250 (I23624,I23435,I23607);
DFFARX1 I_1251  ( .D(I23624), .CLK(I2350), .RSTB(I23155), .Q(I23120) );
nand I_1252 (I23129,I23480,I23302);
nand I_1253 (I23117,I23480,I23384);
not I_1254 (I23716,I2357);
nand I_1255 (I23733,I338892,I338895);
and I_1256 (I23750,I23733,I338901);
DFFARX1 I_1257  ( .D(I23750), .CLK(I2350), .RSTB(I23716), .Q(I23767) );
not I_1258 (I23784,I23767);
nor I_1259 (I23801,I338913,I338895);
or I_1260 (I23699,I23801,I23767);
not I_1261 (I23687,I23801);
DFFARX1 I_1262  ( .D(I338922), .CLK(I2350), .RSTB(I23716), .Q(I23846) );
nor I_1263 (I23863,I23846,I23801);
nand I_1264 (I23880,I338910,I338907);
and I_1265 (I23897,I23880,I338919);
DFFARX1 I_1266  ( .D(I23897), .CLK(I2350), .RSTB(I23716), .Q(I23914) );
nor I_1267 (I23696,I23914,I23767);
not I_1268 (I23945,I23914);
nor I_1269 (I23962,I23846,I23945);
DFFARX1 I_1270  ( .D(I338916), .CLK(I2350), .RSTB(I23716), .Q(I23979) );
and I_1271 (I23996,I23979,I338904);
or I_1272 (I23705,I23996,I23801);
nand I_1273 (I23684,I23996,I23962);
DFFARX1 I_1274  ( .D(I338898), .CLK(I2350), .RSTB(I23716), .Q(I24041) );
and I_1275 (I24058,I24041,I23784);
nor I_1276 (I23702,I23996,I24058);
nor I_1277 (I24089,I24041,I23846);
DFFARX1 I_1278  ( .D(I24089), .CLK(I2350), .RSTB(I23716), .Q(I23693) );
nor I_1279 (I23708,I24041,I23767);
not I_1280 (I24134,I24041);
nor I_1281 (I24151,I23914,I24134);
and I_1282 (I24168,I23801,I24151);
or I_1283 (I24185,I23996,I24168);
DFFARX1 I_1284  ( .D(I24185), .CLK(I2350), .RSTB(I23716), .Q(I23681) );
nand I_1285 (I23690,I24041,I23863);
nand I_1286 (I23678,I24041,I23945);
not I_1287 (I24277,I2357);
nand I_1288 (I24294,I192070,I192061);
and I_1289 (I24311,I24294,I192076);
DFFARX1 I_1290  ( .D(I24311), .CLK(I2350), .RSTB(I24277), .Q(I24328) );
not I_1291 (I24345,I24328);
nor I_1292 (I24362,I192046,I192061);
or I_1293 (I24260,I24362,I24328);
not I_1294 (I24248,I24362);
DFFARX1 I_1295  ( .D(I192049), .CLK(I2350), .RSTB(I24277), .Q(I24407) );
nor I_1296 (I24424,I24407,I24362);
nand I_1297 (I24441,I192067,I192064);
and I_1298 (I24458,I24441,I192052);
DFFARX1 I_1299  ( .D(I24458), .CLK(I2350), .RSTB(I24277), .Q(I24475) );
nor I_1300 (I24257,I24475,I24328);
not I_1301 (I24506,I24475);
nor I_1302 (I24523,I24407,I24506);
DFFARX1 I_1303  ( .D(I192073), .CLK(I2350), .RSTB(I24277), .Q(I24540) );
and I_1304 (I24557,I24540,I192058);
or I_1305 (I24266,I24557,I24362);
nand I_1306 (I24245,I24557,I24523);
DFFARX1 I_1307  ( .D(I192055), .CLK(I2350), .RSTB(I24277), .Q(I24602) );
and I_1308 (I24619,I24602,I24345);
nor I_1309 (I24263,I24557,I24619);
nor I_1310 (I24650,I24602,I24407);
DFFARX1 I_1311  ( .D(I24650), .CLK(I2350), .RSTB(I24277), .Q(I24254) );
nor I_1312 (I24269,I24602,I24328);
not I_1313 (I24695,I24602);
nor I_1314 (I24712,I24475,I24695);
and I_1315 (I24729,I24362,I24712);
or I_1316 (I24746,I24557,I24729);
DFFARX1 I_1317  ( .D(I24746), .CLK(I2350), .RSTB(I24277), .Q(I24242) );
nand I_1318 (I24251,I24602,I24424);
nand I_1319 (I24239,I24602,I24506);
not I_1320 (I24838,I2357);
nand I_1321 (I24855,I113226,I113223);
and I_1322 (I24872,I24855,I113220);
DFFARX1 I_1323  ( .D(I24872), .CLK(I2350), .RSTB(I24838), .Q(I24889) );
not I_1324 (I24906,I24889);
nor I_1325 (I24923,I113244,I113223);
or I_1326 (I24821,I24923,I24889);
not I_1327 (I24809,I24923);
DFFARX1 I_1328  ( .D(I113238), .CLK(I2350), .RSTB(I24838), .Q(I24968) );
nor I_1329 (I24985,I24968,I24923);
nand I_1330 (I25002,I113217,I113229);
and I_1331 (I25019,I25002,I113232);
DFFARX1 I_1332  ( .D(I25019), .CLK(I2350), .RSTB(I24838), .Q(I25036) );
nor I_1333 (I24818,I25036,I24889);
not I_1334 (I25067,I25036);
nor I_1335 (I25084,I24968,I25067);
DFFARX1 I_1336  ( .D(I113241), .CLK(I2350), .RSTB(I24838), .Q(I25101) );
and I_1337 (I25118,I25101,I113247);
or I_1338 (I24827,I25118,I24923);
nand I_1339 (I24806,I25118,I25084);
DFFARX1 I_1340  ( .D(I113235), .CLK(I2350), .RSTB(I24838), .Q(I25163) );
and I_1341 (I25180,I25163,I24906);
nor I_1342 (I24824,I25118,I25180);
nor I_1343 (I25211,I25163,I24968);
DFFARX1 I_1344  ( .D(I25211), .CLK(I2350), .RSTB(I24838), .Q(I24815) );
nor I_1345 (I24830,I25163,I24889);
not I_1346 (I25256,I25163);
nor I_1347 (I25273,I25036,I25256);
and I_1348 (I25290,I24923,I25273);
or I_1349 (I25307,I25118,I25290);
DFFARX1 I_1350  ( .D(I25307), .CLK(I2350), .RSTB(I24838), .Q(I24803) );
nand I_1351 (I24812,I25163,I24985);
nand I_1352 (I24800,I25163,I25067);
not I_1353 (I25399,I2357);
nand I_1354 (I25416,I156931,I156922);
and I_1355 (I25433,I25416,I156937);
DFFARX1 I_1356  ( .D(I25433), .CLK(I2350), .RSTB(I25399), .Q(I25450) );
not I_1357 (I25467,I25450);
nor I_1358 (I25484,I156907,I156922);
or I_1359 (I25382,I25484,I25450);
not I_1360 (I25370,I25484);
DFFARX1 I_1361  ( .D(I156910), .CLK(I2350), .RSTB(I25399), .Q(I25529) );
nor I_1362 (I25546,I25529,I25484);
nand I_1363 (I25563,I156928,I156925);
and I_1364 (I25580,I25563,I156913);
DFFARX1 I_1365  ( .D(I25580), .CLK(I2350), .RSTB(I25399), .Q(I25597) );
nor I_1366 (I25379,I25597,I25450);
not I_1367 (I25628,I25597);
nor I_1368 (I25645,I25529,I25628);
DFFARX1 I_1369  ( .D(I156934), .CLK(I2350), .RSTB(I25399), .Q(I25662) );
and I_1370 (I25679,I25662,I156919);
or I_1371 (I25388,I25679,I25484);
nand I_1372 (I25367,I25679,I25645);
DFFARX1 I_1373  ( .D(I156916), .CLK(I2350), .RSTB(I25399), .Q(I25724) );
and I_1374 (I25741,I25724,I25467);
nor I_1375 (I25385,I25679,I25741);
nor I_1376 (I25772,I25724,I25529);
DFFARX1 I_1377  ( .D(I25772), .CLK(I2350), .RSTB(I25399), .Q(I25376) );
nor I_1378 (I25391,I25724,I25450);
not I_1379 (I25817,I25724);
nor I_1380 (I25834,I25597,I25817);
and I_1381 (I25851,I25484,I25834);
or I_1382 (I25868,I25679,I25851);
DFFARX1 I_1383  ( .D(I25868), .CLK(I2350), .RSTB(I25399), .Q(I25364) );
nand I_1384 (I25373,I25724,I25546);
nand I_1385 (I25361,I25724,I25628);
not I_1386 (I25960,I2357);
not I_1387 (I25977,I241208);
nor I_1388 (I25994,I241196,I241202);
nand I_1389 (I26011,I25994,I241193);
DFFARX1 I_1390  ( .D(I26011), .CLK(I2350), .RSTB(I25960), .Q(I25934) );
nor I_1391 (I26042,I25977,I241196);
nand I_1392 (I26059,I26042,I241199);
not I_1393 (I25949,I26059);
DFFARX1 I_1394  ( .D(I26059), .CLK(I2350), .RSTB(I25960), .Q(I25931) );
not I_1395 (I26104,I241196);
not I_1396 (I26121,I26104);
not I_1397 (I26138,I241211);
nor I_1398 (I26155,I26138,I241223);
and I_1399 (I26172,I26155,I241205);
or I_1400 (I26189,I26172,I241220);
DFFARX1 I_1401  ( .D(I26189), .CLK(I2350), .RSTB(I25960), .Q(I26206) );
nor I_1402 (I26223,I26206,I26059);
nor I_1403 (I26240,I26206,I26121);
nand I_1404 (I25946,I26011,I26240);
nand I_1405 (I26271,I25977,I241211);
nand I_1406 (I26288,I26271,I26206);
and I_1407 (I26305,I26271,I26288);
DFFARX1 I_1408  ( .D(I26305), .CLK(I2350), .RSTB(I25960), .Q(I25928) );
DFFARX1 I_1409  ( .D(I26271), .CLK(I2350), .RSTB(I25960), .Q(I26336) );
and I_1410 (I25925,I26104,I26336);
DFFARX1 I_1411  ( .D(I241214), .CLK(I2350), .RSTB(I25960), .Q(I26367) );
not I_1412 (I26384,I26367);
nor I_1413 (I26401,I26059,I26384);
and I_1414 (I26418,I26367,I26401);
nand I_1415 (I25940,I26367,I26121);
DFFARX1 I_1416  ( .D(I26367), .CLK(I2350), .RSTB(I25960), .Q(I26449) );
not I_1417 (I25937,I26449);
DFFARX1 I_1418  ( .D(I241217), .CLK(I2350), .RSTB(I25960), .Q(I26480) );
not I_1419 (I26497,I26480);
or I_1420 (I26514,I26497,I26418);
DFFARX1 I_1421  ( .D(I26514), .CLK(I2350), .RSTB(I25960), .Q(I25943) );
nand I_1422 (I25952,I26497,I26223);
DFFARX1 I_1423  ( .D(I26497), .CLK(I2350), .RSTB(I25960), .Q(I25922) );
not I_1424 (I26606,I2357);
not I_1425 (I26623,I163555);
nor I_1426 (I26640,I163552,I163540);
nand I_1427 (I26657,I26640,I163543);
DFFARX1 I_1428  ( .D(I26657), .CLK(I2350), .RSTB(I26606), .Q(I26580) );
nor I_1429 (I26688,I26623,I163552);
nand I_1430 (I26705,I26688,I163549);
not I_1431 (I26595,I26705);
DFFARX1 I_1432  ( .D(I26705), .CLK(I2350), .RSTB(I26606), .Q(I26577) );
not I_1433 (I26750,I163552);
not I_1434 (I26767,I26750);
not I_1435 (I26784,I163561);
nor I_1436 (I26801,I26784,I163537);
and I_1437 (I26818,I26801,I163558);
or I_1438 (I26835,I26818,I163546);
DFFARX1 I_1439  ( .D(I26835), .CLK(I2350), .RSTB(I26606), .Q(I26852) );
nor I_1440 (I26869,I26852,I26705);
nor I_1441 (I26886,I26852,I26767);
nand I_1442 (I26592,I26657,I26886);
nand I_1443 (I26917,I26623,I163561);
nand I_1444 (I26934,I26917,I26852);
and I_1445 (I26951,I26917,I26934);
DFFARX1 I_1446  ( .D(I26951), .CLK(I2350), .RSTB(I26606), .Q(I26574) );
DFFARX1 I_1447  ( .D(I26917), .CLK(I2350), .RSTB(I26606), .Q(I26982) );
and I_1448 (I26571,I26750,I26982);
DFFARX1 I_1449  ( .D(I163567), .CLK(I2350), .RSTB(I26606), .Q(I27013) );
not I_1450 (I27030,I27013);
nor I_1451 (I27047,I26705,I27030);
and I_1452 (I27064,I27013,I27047);
nand I_1453 (I26586,I27013,I26767);
DFFARX1 I_1454  ( .D(I27013), .CLK(I2350), .RSTB(I26606), .Q(I27095) );
not I_1455 (I26583,I27095);
DFFARX1 I_1456  ( .D(I163564), .CLK(I2350), .RSTB(I26606), .Q(I27126) );
not I_1457 (I27143,I27126);
or I_1458 (I27160,I27143,I27064);
DFFARX1 I_1459  ( .D(I27160), .CLK(I2350), .RSTB(I26606), .Q(I26589) );
nand I_1460 (I26598,I27143,I26869);
DFFARX1 I_1461  ( .D(I27143), .CLK(I2350), .RSTB(I26606), .Q(I26568) );
not I_1462 (I27252,I2357);
not I_1463 (I27269,I154936);
nor I_1464 (I27286,I154933,I154921);
nand I_1465 (I27303,I27286,I154924);
DFFARX1 I_1466  ( .D(I27303), .CLK(I2350), .RSTB(I27252), .Q(I27226) );
nor I_1467 (I27334,I27269,I154933);
nand I_1468 (I27351,I27334,I154930);
not I_1469 (I27241,I27351);
DFFARX1 I_1470  ( .D(I27351), .CLK(I2350), .RSTB(I27252), .Q(I27223) );
not I_1471 (I27396,I154933);
not I_1472 (I27413,I27396);
not I_1473 (I27430,I154942);
nor I_1474 (I27447,I27430,I154918);
and I_1475 (I27464,I27447,I154939);
or I_1476 (I27481,I27464,I154927);
DFFARX1 I_1477  ( .D(I27481), .CLK(I2350), .RSTB(I27252), .Q(I27498) );
nor I_1478 (I27515,I27498,I27351);
nor I_1479 (I27532,I27498,I27413);
nand I_1480 (I27238,I27303,I27532);
nand I_1481 (I27563,I27269,I154942);
nand I_1482 (I27580,I27563,I27498);
and I_1483 (I27597,I27563,I27580);
DFFARX1 I_1484  ( .D(I27597), .CLK(I2350), .RSTB(I27252), .Q(I27220) );
DFFARX1 I_1485  ( .D(I27563), .CLK(I2350), .RSTB(I27252), .Q(I27628) );
and I_1486 (I27217,I27396,I27628);
DFFARX1 I_1487  ( .D(I154948), .CLK(I2350), .RSTB(I27252), .Q(I27659) );
not I_1488 (I27676,I27659);
nor I_1489 (I27693,I27351,I27676);
and I_1490 (I27710,I27659,I27693);
nand I_1491 (I27232,I27659,I27413);
DFFARX1 I_1492  ( .D(I27659), .CLK(I2350), .RSTB(I27252), .Q(I27741) );
not I_1493 (I27229,I27741);
DFFARX1 I_1494  ( .D(I154945), .CLK(I2350), .RSTB(I27252), .Q(I27772) );
not I_1495 (I27789,I27772);
or I_1496 (I27806,I27789,I27710);
DFFARX1 I_1497  ( .D(I27806), .CLK(I2350), .RSTB(I27252), .Q(I27235) );
nand I_1498 (I27244,I27789,I27515);
DFFARX1 I_1499  ( .D(I27789), .CLK(I2350), .RSTB(I27252), .Q(I27214) );
not I_1500 (I27898,I2357);
not I_1501 (I27915,I312399);
nor I_1502 (I27932,I312375,I312381);
nand I_1503 (I27949,I27932,I312384);
DFFARX1 I_1504  ( .D(I27949), .CLK(I2350), .RSTB(I27898), .Q(I27872) );
nor I_1505 (I27980,I27915,I312375);
nand I_1506 (I27997,I27980,I312393);
not I_1507 (I27887,I27997);
DFFARX1 I_1508  ( .D(I27997), .CLK(I2350), .RSTB(I27898), .Q(I27869) );
not I_1509 (I28042,I312375);
not I_1510 (I28059,I28042);
not I_1511 (I28076,I312372);
nor I_1512 (I28093,I28076,I312387);
and I_1513 (I28110,I28093,I312378);
or I_1514 (I28127,I28110,I312390);
DFFARX1 I_1515  ( .D(I28127), .CLK(I2350), .RSTB(I27898), .Q(I28144) );
nor I_1516 (I28161,I28144,I27997);
nor I_1517 (I28178,I28144,I28059);
nand I_1518 (I27884,I27949,I28178);
nand I_1519 (I28209,I27915,I312372);
nand I_1520 (I28226,I28209,I28144);
and I_1521 (I28243,I28209,I28226);
DFFARX1 I_1522  ( .D(I28243), .CLK(I2350), .RSTB(I27898), .Q(I27866) );
DFFARX1 I_1523  ( .D(I28209), .CLK(I2350), .RSTB(I27898), .Q(I28274) );
and I_1524 (I27863,I28042,I28274);
DFFARX1 I_1525  ( .D(I312402), .CLK(I2350), .RSTB(I27898), .Q(I28305) );
not I_1526 (I28322,I28305);
nor I_1527 (I28339,I27997,I28322);
and I_1528 (I28356,I28305,I28339);
nand I_1529 (I27878,I28305,I28059);
DFFARX1 I_1530  ( .D(I28305), .CLK(I2350), .RSTB(I27898), .Q(I28387) );
not I_1531 (I27875,I28387);
DFFARX1 I_1532  ( .D(I312396), .CLK(I2350), .RSTB(I27898), .Q(I28418) );
not I_1533 (I28435,I28418);
or I_1534 (I28452,I28435,I28356);
DFFARX1 I_1535  ( .D(I28452), .CLK(I2350), .RSTB(I27898), .Q(I27881) );
nand I_1536 (I27890,I28435,I28161);
DFFARX1 I_1537  ( .D(I28435), .CLK(I2350), .RSTB(I27898), .Q(I27860) );
not I_1538 (I28544,I2357);
not I_1539 (I28561,I335118);
nor I_1540 (I28578,I335133,I335148);
nand I_1541 (I28595,I28578,I335136);
DFFARX1 I_1542  ( .D(I28595), .CLK(I2350), .RSTB(I28544), .Q(I28518) );
nor I_1543 (I28626,I28561,I335133);
nand I_1544 (I28643,I28626,I335139);
not I_1545 (I28533,I28643);
DFFARX1 I_1546  ( .D(I28643), .CLK(I2350), .RSTB(I28544), .Q(I28515) );
not I_1547 (I28688,I335133);
not I_1548 (I28705,I28688);
not I_1549 (I28722,I335145);
nor I_1550 (I28739,I28722,I335142);
and I_1551 (I28756,I28739,I335121);
or I_1552 (I28773,I28756,I335130);
DFFARX1 I_1553  ( .D(I28773), .CLK(I2350), .RSTB(I28544), .Q(I28790) );
nor I_1554 (I28807,I28790,I28643);
nor I_1555 (I28824,I28790,I28705);
nand I_1556 (I28530,I28595,I28824);
nand I_1557 (I28855,I28561,I335145);
nand I_1558 (I28872,I28855,I28790);
and I_1559 (I28889,I28855,I28872);
DFFARX1 I_1560  ( .D(I28889), .CLK(I2350), .RSTB(I28544), .Q(I28512) );
DFFARX1 I_1561  ( .D(I28855), .CLK(I2350), .RSTB(I28544), .Q(I28920) );
and I_1562 (I28509,I28688,I28920);
DFFARX1 I_1563  ( .D(I335127), .CLK(I2350), .RSTB(I28544), .Q(I28951) );
not I_1564 (I28968,I28951);
nor I_1565 (I28985,I28643,I28968);
and I_1566 (I29002,I28951,I28985);
nand I_1567 (I28524,I28951,I28705);
DFFARX1 I_1568  ( .D(I28951), .CLK(I2350), .RSTB(I28544), .Q(I29033) );
not I_1569 (I28521,I29033);
DFFARX1 I_1570  ( .D(I335124), .CLK(I2350), .RSTB(I28544), .Q(I29064) );
not I_1571 (I29081,I29064);
or I_1572 (I29098,I29081,I29002);
DFFARX1 I_1573  ( .D(I29098), .CLK(I2350), .RSTB(I28544), .Q(I28527) );
nand I_1574 (I28536,I29081,I28807);
DFFARX1 I_1575  ( .D(I29081), .CLK(I2350), .RSTB(I28544), .Q(I28506) );
not I_1576 (I29190,I2357);
not I_1577 (I29207,I292764);
nor I_1578 (I29224,I292740,I292746);
nand I_1579 (I29241,I29224,I292749);
DFFARX1 I_1580  ( .D(I29241), .CLK(I2350), .RSTB(I29190), .Q(I29164) );
nor I_1581 (I29272,I29207,I292740);
nand I_1582 (I29289,I29272,I292758);
not I_1583 (I29179,I29289);
DFFARX1 I_1584  ( .D(I29289), .CLK(I2350), .RSTB(I29190), .Q(I29161) );
not I_1585 (I29334,I292740);
not I_1586 (I29351,I29334);
not I_1587 (I29368,I292737);
nor I_1588 (I29385,I29368,I292752);
and I_1589 (I29402,I29385,I292743);
or I_1590 (I29419,I29402,I292755);
DFFARX1 I_1591  ( .D(I29419), .CLK(I2350), .RSTB(I29190), .Q(I29436) );
nor I_1592 (I29453,I29436,I29289);
nor I_1593 (I29470,I29436,I29351);
nand I_1594 (I29176,I29241,I29470);
nand I_1595 (I29501,I29207,I292737);
nand I_1596 (I29518,I29501,I29436);
and I_1597 (I29535,I29501,I29518);
DFFARX1 I_1598  ( .D(I29535), .CLK(I2350), .RSTB(I29190), .Q(I29158) );
DFFARX1 I_1599  ( .D(I29501), .CLK(I2350), .RSTB(I29190), .Q(I29566) );
and I_1600 (I29155,I29334,I29566);
DFFARX1 I_1601  ( .D(I292767), .CLK(I2350), .RSTB(I29190), .Q(I29597) );
not I_1602 (I29614,I29597);
nor I_1603 (I29631,I29289,I29614);
and I_1604 (I29648,I29597,I29631);
nand I_1605 (I29170,I29597,I29351);
DFFARX1 I_1606  ( .D(I29597), .CLK(I2350), .RSTB(I29190), .Q(I29679) );
not I_1607 (I29167,I29679);
DFFARX1 I_1608  ( .D(I292761), .CLK(I2350), .RSTB(I29190), .Q(I29710) );
not I_1609 (I29727,I29710);
or I_1610 (I29744,I29727,I29648);
DFFARX1 I_1611  ( .D(I29744), .CLK(I2350), .RSTB(I29190), .Q(I29173) );
nand I_1612 (I29182,I29727,I29453);
DFFARX1 I_1613  ( .D(I29727), .CLK(I2350), .RSTB(I29190), .Q(I29152) );
not I_1614 (I29836,I2357);
not I_1615 (I29853,I287409);
nor I_1616 (I29870,I287385,I287391);
nand I_1617 (I29887,I29870,I287394);
DFFARX1 I_1618  ( .D(I29887), .CLK(I2350), .RSTB(I29836), .Q(I29810) );
nor I_1619 (I29918,I29853,I287385);
nand I_1620 (I29935,I29918,I287403);
not I_1621 (I29825,I29935);
DFFARX1 I_1622  ( .D(I29935), .CLK(I2350), .RSTB(I29836), .Q(I29807) );
not I_1623 (I29980,I287385);
not I_1624 (I29997,I29980);
not I_1625 (I30014,I287382);
nor I_1626 (I30031,I30014,I287397);
and I_1627 (I30048,I30031,I287388);
or I_1628 (I30065,I30048,I287400);
DFFARX1 I_1629  ( .D(I30065), .CLK(I2350), .RSTB(I29836), .Q(I30082) );
nor I_1630 (I30099,I30082,I29935);
nor I_1631 (I30116,I30082,I29997);
nand I_1632 (I29822,I29887,I30116);
nand I_1633 (I30147,I29853,I287382);
nand I_1634 (I30164,I30147,I30082);
and I_1635 (I30181,I30147,I30164);
DFFARX1 I_1636  ( .D(I30181), .CLK(I2350), .RSTB(I29836), .Q(I29804) );
DFFARX1 I_1637  ( .D(I30147), .CLK(I2350), .RSTB(I29836), .Q(I30212) );
and I_1638 (I29801,I29980,I30212);
DFFARX1 I_1639  ( .D(I287412), .CLK(I2350), .RSTB(I29836), .Q(I30243) );
not I_1640 (I30260,I30243);
nor I_1641 (I30277,I29935,I30260);
and I_1642 (I30294,I30243,I30277);
nand I_1643 (I29816,I30243,I29997);
DFFARX1 I_1644  ( .D(I30243), .CLK(I2350), .RSTB(I29836), .Q(I30325) );
not I_1645 (I29813,I30325);
DFFARX1 I_1646  ( .D(I287406), .CLK(I2350), .RSTB(I29836), .Q(I30356) );
not I_1647 (I30373,I30356);
or I_1648 (I30390,I30373,I30294);
DFFARX1 I_1649  ( .D(I30390), .CLK(I2350), .RSTB(I29836), .Q(I29819) );
nand I_1650 (I29828,I30373,I30099);
DFFARX1 I_1651  ( .D(I30373), .CLK(I2350), .RSTB(I29836), .Q(I29798) );
not I_1652 (I30482,I2357);
not I_1653 (I30499,I263172);
nor I_1654 (I30516,I263160,I263166);
nand I_1655 (I30533,I30516,I263157);
DFFARX1 I_1656  ( .D(I30533), .CLK(I2350), .RSTB(I30482), .Q(I30456) );
nor I_1657 (I30564,I30499,I263160);
nand I_1658 (I30581,I30564,I263163);
not I_1659 (I30471,I30581);
DFFARX1 I_1660  ( .D(I30581), .CLK(I2350), .RSTB(I30482), .Q(I30453) );
not I_1661 (I30626,I263160);
not I_1662 (I30643,I30626);
not I_1663 (I30660,I263175);
nor I_1664 (I30677,I30660,I263187);
and I_1665 (I30694,I30677,I263169);
or I_1666 (I30711,I30694,I263184);
DFFARX1 I_1667  ( .D(I30711), .CLK(I2350), .RSTB(I30482), .Q(I30728) );
nor I_1668 (I30745,I30728,I30581);
nor I_1669 (I30762,I30728,I30643);
nand I_1670 (I30468,I30533,I30762);
nand I_1671 (I30793,I30499,I263175);
nand I_1672 (I30810,I30793,I30728);
and I_1673 (I30827,I30793,I30810);
DFFARX1 I_1674  ( .D(I30827), .CLK(I2350), .RSTB(I30482), .Q(I30450) );
DFFARX1 I_1675  ( .D(I30793), .CLK(I2350), .RSTB(I30482), .Q(I30858) );
and I_1676 (I30447,I30626,I30858);
DFFARX1 I_1677  ( .D(I263178), .CLK(I2350), .RSTB(I30482), .Q(I30889) );
not I_1678 (I30906,I30889);
nor I_1679 (I30923,I30581,I30906);
and I_1680 (I30940,I30889,I30923);
nand I_1681 (I30462,I30889,I30643);
DFFARX1 I_1682  ( .D(I30889), .CLK(I2350), .RSTB(I30482), .Q(I30971) );
not I_1683 (I30459,I30971);
DFFARX1 I_1684  ( .D(I263181), .CLK(I2350), .RSTB(I30482), .Q(I31002) );
not I_1685 (I31019,I31002);
or I_1686 (I31036,I31019,I30940);
DFFARX1 I_1687  ( .D(I31036), .CLK(I2350), .RSTB(I30482), .Q(I30465) );
nand I_1688 (I30474,I31019,I30745);
DFFARX1 I_1689  ( .D(I31019), .CLK(I2350), .RSTB(I30482), .Q(I30444) );
not I_1690 (I31128,I2357);
not I_1691 (I31145,I123400);
nor I_1692 (I31162,I123430,I123409);
nand I_1693 (I31179,I31162,I123421);
DFFARX1 I_1694  ( .D(I31179), .CLK(I2350), .RSTB(I31128), .Q(I31102) );
nor I_1695 (I31210,I31145,I123430);
nand I_1696 (I31227,I31210,I123403);
not I_1697 (I31117,I31227);
DFFARX1 I_1698  ( .D(I31227), .CLK(I2350), .RSTB(I31128), .Q(I31099) );
not I_1699 (I31272,I123430);
not I_1700 (I31289,I31272);
not I_1701 (I31306,I123406);
nor I_1702 (I31323,I31306,I123424);
and I_1703 (I31340,I31323,I123415);
or I_1704 (I31357,I31340,I123412);
DFFARX1 I_1705  ( .D(I31357), .CLK(I2350), .RSTB(I31128), .Q(I31374) );
nor I_1706 (I31391,I31374,I31227);
nor I_1707 (I31408,I31374,I31289);
nand I_1708 (I31114,I31179,I31408);
nand I_1709 (I31439,I31145,I123406);
nand I_1710 (I31456,I31439,I31374);
and I_1711 (I31473,I31439,I31456);
DFFARX1 I_1712  ( .D(I31473), .CLK(I2350), .RSTB(I31128), .Q(I31096) );
DFFARX1 I_1713  ( .D(I31439), .CLK(I2350), .RSTB(I31128), .Q(I31504) );
and I_1714 (I31093,I31272,I31504);
DFFARX1 I_1715  ( .D(I123418), .CLK(I2350), .RSTB(I31128), .Q(I31535) );
not I_1716 (I31552,I31535);
nor I_1717 (I31569,I31227,I31552);
and I_1718 (I31586,I31535,I31569);
nand I_1719 (I31108,I31535,I31289);
DFFARX1 I_1720  ( .D(I31535), .CLK(I2350), .RSTB(I31128), .Q(I31617) );
not I_1721 (I31105,I31617);
DFFARX1 I_1722  ( .D(I123427), .CLK(I2350), .RSTB(I31128), .Q(I31648) );
not I_1723 (I31665,I31648);
or I_1724 (I31682,I31665,I31586);
DFFARX1 I_1725  ( .D(I31682), .CLK(I2350), .RSTB(I31128), .Q(I31111) );
nand I_1726 (I31120,I31665,I31391);
DFFARX1 I_1727  ( .D(I31665), .CLK(I2350), .RSTB(I31128), .Q(I31090) );
not I_1728 (I31774,I2357);
not I_1729 (I31791,I356504);
nor I_1730 (I31808,I356519,I356534);
nand I_1731 (I31825,I31808,I356522);
DFFARX1 I_1732  ( .D(I31825), .CLK(I2350), .RSTB(I31774), .Q(I31748) );
nor I_1733 (I31856,I31791,I356519);
nand I_1734 (I31873,I31856,I356525);
not I_1735 (I31763,I31873);
DFFARX1 I_1736  ( .D(I31873), .CLK(I2350), .RSTB(I31774), .Q(I31745) );
not I_1737 (I31918,I356519);
not I_1738 (I31935,I31918);
not I_1739 (I31952,I356531);
nor I_1740 (I31969,I31952,I356528);
and I_1741 (I31986,I31969,I356507);
or I_1742 (I32003,I31986,I356516);
DFFARX1 I_1743  ( .D(I32003), .CLK(I2350), .RSTB(I31774), .Q(I32020) );
nor I_1744 (I32037,I32020,I31873);
nor I_1745 (I32054,I32020,I31935);
nand I_1746 (I31760,I31825,I32054);
nand I_1747 (I32085,I31791,I356531);
nand I_1748 (I32102,I32085,I32020);
and I_1749 (I32119,I32085,I32102);
DFFARX1 I_1750  ( .D(I32119), .CLK(I2350), .RSTB(I31774), .Q(I31742) );
DFFARX1 I_1751  ( .D(I32085), .CLK(I2350), .RSTB(I31774), .Q(I32150) );
and I_1752 (I31739,I31918,I32150);
DFFARX1 I_1753  ( .D(I356513), .CLK(I2350), .RSTB(I31774), .Q(I32181) );
not I_1754 (I32198,I32181);
nor I_1755 (I32215,I31873,I32198);
and I_1756 (I32232,I32181,I32215);
nand I_1757 (I31754,I32181,I31935);
DFFARX1 I_1758  ( .D(I32181), .CLK(I2350), .RSTB(I31774), .Q(I32263) );
not I_1759 (I31751,I32263);
DFFARX1 I_1760  ( .D(I356510), .CLK(I2350), .RSTB(I31774), .Q(I32294) );
not I_1761 (I32311,I32294);
or I_1762 (I32328,I32311,I32232);
DFFARX1 I_1763  ( .D(I32328), .CLK(I2350), .RSTB(I31774), .Q(I31757) );
nand I_1764 (I31766,I32311,I32037);
DFFARX1 I_1765  ( .D(I32311), .CLK(I2350), .RSTB(I31774), .Q(I31736) );
not I_1766 (I32420,I2357);
not I_1767 (I32437,I236451);
nor I_1768 (I32454,I236433,I236448);
nand I_1769 (I32471,I32454,I236457);
DFFARX1 I_1770  ( .D(I32471), .CLK(I2350), .RSTB(I32420), .Q(I32394) );
nor I_1771 (I32502,I32437,I236433);
nand I_1772 (I32519,I32502,I236460);
not I_1773 (I32409,I32519);
DFFARX1 I_1774  ( .D(I32519), .CLK(I2350), .RSTB(I32420), .Q(I32391) );
not I_1775 (I32564,I236433);
not I_1776 (I32581,I32564);
not I_1777 (I32598,I236463);
nor I_1778 (I32615,I32598,I236439);
and I_1779 (I32632,I32615,I236442);
or I_1780 (I32649,I32632,I236436);
DFFARX1 I_1781  ( .D(I32649), .CLK(I2350), .RSTB(I32420), .Q(I32666) );
nor I_1782 (I32683,I32666,I32519);
nor I_1783 (I32700,I32666,I32581);
nand I_1784 (I32406,I32471,I32700);
nand I_1785 (I32731,I32437,I236463);
nand I_1786 (I32748,I32731,I32666);
and I_1787 (I32765,I32731,I32748);
DFFARX1 I_1788  ( .D(I32765), .CLK(I2350), .RSTB(I32420), .Q(I32388) );
DFFARX1 I_1789  ( .D(I32731), .CLK(I2350), .RSTB(I32420), .Q(I32796) );
and I_1790 (I32385,I32564,I32796);
DFFARX1 I_1791  ( .D(I236445), .CLK(I2350), .RSTB(I32420), .Q(I32827) );
not I_1792 (I32844,I32827);
nor I_1793 (I32861,I32519,I32844);
and I_1794 (I32878,I32827,I32861);
nand I_1795 (I32400,I32827,I32581);
DFFARX1 I_1796  ( .D(I32827), .CLK(I2350), .RSTB(I32420), .Q(I32909) );
not I_1797 (I32397,I32909);
DFFARX1 I_1798  ( .D(I236454), .CLK(I2350), .RSTB(I32420), .Q(I32940) );
not I_1799 (I32957,I32940);
or I_1800 (I32974,I32957,I32878);
DFFARX1 I_1801  ( .D(I32974), .CLK(I2350), .RSTB(I32420), .Q(I32403) );
nand I_1802 (I32412,I32957,I32683);
DFFARX1 I_1803  ( .D(I32957), .CLK(I2350), .RSTB(I32420), .Q(I32382) );
not I_1804 (I33066,I2357);
not I_1805 (I33083,I116260);
nor I_1806 (I33100,I116290,I116269);
nand I_1807 (I33117,I33100,I116281);
DFFARX1 I_1808  ( .D(I33117), .CLK(I2350), .RSTB(I33066), .Q(I33040) );
nor I_1809 (I33148,I33083,I116290);
nand I_1810 (I33165,I33148,I116263);
not I_1811 (I33055,I33165);
DFFARX1 I_1812  ( .D(I33165), .CLK(I2350), .RSTB(I33066), .Q(I33037) );
not I_1813 (I33210,I116290);
not I_1814 (I33227,I33210);
not I_1815 (I33244,I116266);
nor I_1816 (I33261,I33244,I116284);
and I_1817 (I33278,I33261,I116275);
or I_1818 (I33295,I33278,I116272);
DFFARX1 I_1819  ( .D(I33295), .CLK(I2350), .RSTB(I33066), .Q(I33312) );
nor I_1820 (I33329,I33312,I33165);
nor I_1821 (I33346,I33312,I33227);
nand I_1822 (I33052,I33117,I33346);
nand I_1823 (I33377,I33083,I116266);
nand I_1824 (I33394,I33377,I33312);
and I_1825 (I33411,I33377,I33394);
DFFARX1 I_1826  ( .D(I33411), .CLK(I2350), .RSTB(I33066), .Q(I33034) );
DFFARX1 I_1827  ( .D(I33377), .CLK(I2350), .RSTB(I33066), .Q(I33442) );
and I_1828 (I33031,I33210,I33442);
DFFARX1 I_1829  ( .D(I116278), .CLK(I2350), .RSTB(I33066), .Q(I33473) );
not I_1830 (I33490,I33473);
nor I_1831 (I33507,I33165,I33490);
and I_1832 (I33524,I33473,I33507);
nand I_1833 (I33046,I33473,I33227);
DFFARX1 I_1834  ( .D(I33473), .CLK(I2350), .RSTB(I33066), .Q(I33555) );
not I_1835 (I33043,I33555);
DFFARX1 I_1836  ( .D(I116287), .CLK(I2350), .RSTB(I33066), .Q(I33586) );
not I_1837 (I33603,I33586);
or I_1838 (I33620,I33603,I33524);
DFFARX1 I_1839  ( .D(I33620), .CLK(I2350), .RSTB(I33066), .Q(I33049) );
nand I_1840 (I33058,I33603,I33329);
DFFARX1 I_1841  ( .D(I33603), .CLK(I2350), .RSTB(I33066), .Q(I33028) );
not I_1842 (I33712,I2357);
not I_1843 (I33729,I323692);
nor I_1844 (I33746,I323677,I323704);
nand I_1845 (I33763,I33746,I323680);
DFFARX1 I_1846  ( .D(I33763), .CLK(I2350), .RSTB(I33712), .Q(I33686) );
nor I_1847 (I33794,I33729,I323677);
nand I_1848 (I33811,I33794,I323695);
not I_1849 (I33701,I33811);
DFFARX1 I_1850  ( .D(I33811), .CLK(I2350), .RSTB(I33712), .Q(I33683) );
not I_1851 (I33856,I323677);
not I_1852 (I33873,I33856);
not I_1853 (I33890,I323707);
nor I_1854 (I33907,I33890,I323689);
and I_1855 (I33924,I33907,I323698);
or I_1856 (I33941,I33924,I323683);
DFFARX1 I_1857  ( .D(I33941), .CLK(I2350), .RSTB(I33712), .Q(I33958) );
nor I_1858 (I33975,I33958,I33811);
nor I_1859 (I33992,I33958,I33873);
nand I_1860 (I33698,I33763,I33992);
nand I_1861 (I34023,I33729,I323707);
nand I_1862 (I34040,I34023,I33958);
and I_1863 (I34057,I34023,I34040);
DFFARX1 I_1864  ( .D(I34057), .CLK(I2350), .RSTB(I33712), .Q(I33680) );
DFFARX1 I_1865  ( .D(I34023), .CLK(I2350), .RSTB(I33712), .Q(I34088) );
and I_1866 (I33677,I33856,I34088);
DFFARX1 I_1867  ( .D(I323686), .CLK(I2350), .RSTB(I33712), .Q(I34119) );
not I_1868 (I34136,I34119);
nor I_1869 (I34153,I33811,I34136);
and I_1870 (I34170,I34119,I34153);
nand I_1871 (I33692,I34119,I33873);
DFFARX1 I_1872  ( .D(I34119), .CLK(I2350), .RSTB(I33712), .Q(I34201) );
not I_1873 (I33689,I34201);
DFFARX1 I_1874  ( .D(I323701), .CLK(I2350), .RSTB(I33712), .Q(I34232) );
not I_1875 (I34249,I34232);
or I_1876 (I34266,I34249,I34170);
DFFARX1 I_1877  ( .D(I34266), .CLK(I2350), .RSTB(I33712), .Q(I33695) );
nand I_1878 (I33704,I34249,I33975);
DFFARX1 I_1879  ( .D(I34249), .CLK(I2350), .RSTB(I33712), .Q(I33674) );
not I_1880 (I34358,I2357);
not I_1881 (I34375,I10217);
nor I_1882 (I34392,I10229,I10214);
nand I_1883 (I34409,I34392,I10226);
DFFARX1 I_1884  ( .D(I34409), .CLK(I2350), .RSTB(I34358), .Q(I34332) );
nor I_1885 (I34440,I34375,I10229);
nand I_1886 (I34457,I34440,I10244);
not I_1887 (I34347,I34457);
DFFARX1 I_1888  ( .D(I34457), .CLK(I2350), .RSTB(I34358), .Q(I34329) );
not I_1889 (I34502,I10229);
not I_1890 (I34519,I34502);
not I_1891 (I34536,I10220);
nor I_1892 (I34553,I34536,I10232);
and I_1893 (I34570,I34553,I10223);
or I_1894 (I34587,I34570,I10238);
DFFARX1 I_1895  ( .D(I34587), .CLK(I2350), .RSTB(I34358), .Q(I34604) );
nor I_1896 (I34621,I34604,I34457);
nor I_1897 (I34638,I34604,I34519);
nand I_1898 (I34344,I34409,I34638);
nand I_1899 (I34669,I34375,I10220);
nand I_1900 (I34686,I34669,I34604);
and I_1901 (I34703,I34669,I34686);
DFFARX1 I_1902  ( .D(I34703), .CLK(I2350), .RSTB(I34358), .Q(I34326) );
DFFARX1 I_1903  ( .D(I34669), .CLK(I2350), .RSTB(I34358), .Q(I34734) );
and I_1904 (I34323,I34502,I34734);
DFFARX1 I_1905  ( .D(I10241), .CLK(I2350), .RSTB(I34358), .Q(I34765) );
not I_1906 (I34782,I34765);
nor I_1907 (I34799,I34457,I34782);
and I_1908 (I34816,I34765,I34799);
nand I_1909 (I34338,I34765,I34519);
DFFARX1 I_1910  ( .D(I34765), .CLK(I2350), .RSTB(I34358), .Q(I34847) );
not I_1911 (I34335,I34847);
DFFARX1 I_1912  ( .D(I10235), .CLK(I2350), .RSTB(I34358), .Q(I34878) );
not I_1913 (I34895,I34878);
or I_1914 (I34912,I34895,I34816);
DFFARX1 I_1915  ( .D(I34912), .CLK(I2350), .RSTB(I34358), .Q(I34341) );
nand I_1916 (I34350,I34895,I34621);
DFFARX1 I_1917  ( .D(I34895), .CLK(I2350), .RSTB(I34358), .Q(I34320) );
not I_1918 (I35004,I2357);
not I_1919 (I35021,I251034);
nor I_1920 (I35038,I251022,I251028);
nand I_1921 (I35055,I35038,I251019);
DFFARX1 I_1922  ( .D(I35055), .CLK(I2350), .RSTB(I35004), .Q(I34978) );
nor I_1923 (I35086,I35021,I251022);
nand I_1924 (I35103,I35086,I251025);
not I_1925 (I34993,I35103);
DFFARX1 I_1926  ( .D(I35103), .CLK(I2350), .RSTB(I35004), .Q(I34975) );
not I_1927 (I35148,I251022);
not I_1928 (I35165,I35148);
not I_1929 (I35182,I251037);
nor I_1930 (I35199,I35182,I251049);
and I_1931 (I35216,I35199,I251031);
or I_1932 (I35233,I35216,I251046);
DFFARX1 I_1933  ( .D(I35233), .CLK(I2350), .RSTB(I35004), .Q(I35250) );
nor I_1934 (I35267,I35250,I35103);
nor I_1935 (I35284,I35250,I35165);
nand I_1936 (I34990,I35055,I35284);
nand I_1937 (I35315,I35021,I251037);
nand I_1938 (I35332,I35315,I35250);
and I_1939 (I35349,I35315,I35332);
DFFARX1 I_1940  ( .D(I35349), .CLK(I2350), .RSTB(I35004), .Q(I34972) );
DFFARX1 I_1941  ( .D(I35315), .CLK(I2350), .RSTB(I35004), .Q(I35380) );
and I_1942 (I34969,I35148,I35380);
DFFARX1 I_1943  ( .D(I251040), .CLK(I2350), .RSTB(I35004), .Q(I35411) );
not I_1944 (I35428,I35411);
nor I_1945 (I35445,I35103,I35428);
and I_1946 (I35462,I35411,I35445);
nand I_1947 (I34984,I35411,I35165);
DFFARX1 I_1948  ( .D(I35411), .CLK(I2350), .RSTB(I35004), .Q(I35493) );
not I_1949 (I34981,I35493);
DFFARX1 I_1950  ( .D(I251043), .CLK(I2350), .RSTB(I35004), .Q(I35524) );
not I_1951 (I35541,I35524);
or I_1952 (I35558,I35541,I35462);
DFFARX1 I_1953  ( .D(I35558), .CLK(I2350), .RSTB(I35004), .Q(I34987) );
nand I_1954 (I34996,I35541,I35267);
DFFARX1 I_1955  ( .D(I35541), .CLK(I2350), .RSTB(I35004), .Q(I34966) );
not I_1956 (I35650,I2357);
not I_1957 (I35667,I1223);
nor I_1958 (I35684,I2311,I1367);
nand I_1959 (I35701,I35684,I2255);
DFFARX1 I_1960  ( .D(I35701), .CLK(I2350), .RSTB(I35650), .Q(I35624) );
nor I_1961 (I35732,I35667,I2311);
nand I_1962 (I35749,I35732,I2127);
not I_1963 (I35639,I35749);
DFFARX1 I_1964  ( .D(I35749), .CLK(I2350), .RSTB(I35650), .Q(I35621) );
not I_1965 (I35794,I2311);
not I_1966 (I35811,I35794);
not I_1967 (I35828,I1335);
nor I_1968 (I35845,I35828,I2239);
and I_1969 (I35862,I35845,I1623);
or I_1970 (I35879,I35862,I1495);
DFFARX1 I_1971  ( .D(I35879), .CLK(I2350), .RSTB(I35650), .Q(I35896) );
nor I_1972 (I35913,I35896,I35749);
nor I_1973 (I35930,I35896,I35811);
nand I_1974 (I35636,I35701,I35930);
nand I_1975 (I35961,I35667,I1335);
nand I_1976 (I35978,I35961,I35896);
and I_1977 (I35995,I35961,I35978);
DFFARX1 I_1978  ( .D(I35995), .CLK(I2350), .RSTB(I35650), .Q(I35618) );
DFFARX1 I_1979  ( .D(I35961), .CLK(I2350), .RSTB(I35650), .Q(I36026) );
and I_1980 (I35615,I35794,I36026);
DFFARX1 I_1981  ( .D(I1991), .CLK(I2350), .RSTB(I35650), .Q(I36057) );
not I_1982 (I36074,I36057);
nor I_1983 (I36091,I35749,I36074);
and I_1984 (I36108,I36057,I36091);
nand I_1985 (I35630,I36057,I35811);
DFFARX1 I_1986  ( .D(I36057), .CLK(I2350), .RSTB(I35650), .Q(I36139) );
not I_1987 (I35627,I36139);
DFFARX1 I_1988  ( .D(I2039), .CLK(I2350), .RSTB(I35650), .Q(I36170) );
not I_1989 (I36187,I36170);
or I_1990 (I36204,I36187,I36108);
DFFARX1 I_1991  ( .D(I36204), .CLK(I2350), .RSTB(I35650), .Q(I35633) );
nand I_1992 (I35642,I36187,I35913);
DFFARX1 I_1993  ( .D(I36187), .CLK(I2350), .RSTB(I35650), .Q(I35612) );
not I_1994 (I36296,I2357);
not I_1995 (I36313,I93345);
nor I_1996 (I36330,I93333,I93339);
nand I_1997 (I36347,I36330,I93348);
DFFARX1 I_1998  ( .D(I36347), .CLK(I2350), .RSTB(I36296), .Q(I36270) );
nor I_1999 (I36378,I36313,I93333);
nand I_2000 (I36395,I36378,I93336);
not I_2001 (I36285,I36395);
DFFARX1 I_2002  ( .D(I36395), .CLK(I2350), .RSTB(I36296), .Q(I36267) );
not I_2003 (I36440,I93333);
not I_2004 (I36457,I36440);
not I_2005 (I36474,I93357);
nor I_2006 (I36491,I36474,I93330);
and I_2007 (I36508,I36491,I93351);
or I_2008 (I36525,I36508,I93342);
DFFARX1 I_2009  ( .D(I36525), .CLK(I2350), .RSTB(I36296), .Q(I36542) );
nor I_2010 (I36559,I36542,I36395);
nor I_2011 (I36576,I36542,I36457);
nand I_2012 (I36282,I36347,I36576);
nand I_2013 (I36607,I36313,I93357);
nand I_2014 (I36624,I36607,I36542);
and I_2015 (I36641,I36607,I36624);
DFFARX1 I_2016  ( .D(I36641), .CLK(I2350), .RSTB(I36296), .Q(I36264) );
DFFARX1 I_2017  ( .D(I36607), .CLK(I2350), .RSTB(I36296), .Q(I36672) );
and I_2018 (I36261,I36440,I36672);
DFFARX1 I_2019  ( .D(I93327), .CLK(I2350), .RSTB(I36296), .Q(I36703) );
not I_2020 (I36720,I36703);
nor I_2021 (I36737,I36395,I36720);
and I_2022 (I36754,I36703,I36737);
nand I_2023 (I36276,I36703,I36457);
DFFARX1 I_2024  ( .D(I36703), .CLK(I2350), .RSTB(I36296), .Q(I36785) );
not I_2025 (I36273,I36785);
DFFARX1 I_2026  ( .D(I93354), .CLK(I2350), .RSTB(I36296), .Q(I36816) );
not I_2027 (I36833,I36816);
or I_2028 (I36850,I36833,I36754);
DFFARX1 I_2029  ( .D(I36850), .CLK(I2350), .RSTB(I36296), .Q(I36279) );
nand I_2030 (I36288,I36833,I36559);
DFFARX1 I_2031  ( .D(I36833), .CLK(I2350), .RSTB(I36296), .Q(I36258) );
not I_2032 (I36942,I2357);
not I_2033 (I36959,I166207);
nor I_2034 (I36976,I166204,I166192);
nand I_2035 (I36993,I36976,I166195);
DFFARX1 I_2036  ( .D(I36993), .CLK(I2350), .RSTB(I36942), .Q(I36916) );
nor I_2037 (I37024,I36959,I166204);
nand I_2038 (I37041,I37024,I166201);
not I_2039 (I36931,I37041);
DFFARX1 I_2040  ( .D(I37041), .CLK(I2350), .RSTB(I36942), .Q(I36913) );
not I_2041 (I37086,I166204);
not I_2042 (I37103,I37086);
not I_2043 (I37120,I166213);
nor I_2044 (I37137,I37120,I166189);
and I_2045 (I37154,I37137,I166210);
or I_2046 (I37171,I37154,I166198);
DFFARX1 I_2047  ( .D(I37171), .CLK(I2350), .RSTB(I36942), .Q(I37188) );
nor I_2048 (I37205,I37188,I37041);
nor I_2049 (I37222,I37188,I37103);
nand I_2050 (I36928,I36993,I37222);
nand I_2051 (I37253,I36959,I166213);
nand I_2052 (I37270,I37253,I37188);
and I_2053 (I37287,I37253,I37270);
DFFARX1 I_2054  ( .D(I37287), .CLK(I2350), .RSTB(I36942), .Q(I36910) );
DFFARX1 I_2055  ( .D(I37253), .CLK(I2350), .RSTB(I36942), .Q(I37318) );
and I_2056 (I36907,I37086,I37318);
DFFARX1 I_2057  ( .D(I166219), .CLK(I2350), .RSTB(I36942), .Q(I37349) );
not I_2058 (I37366,I37349);
nor I_2059 (I37383,I37041,I37366);
and I_2060 (I37400,I37349,I37383);
nand I_2061 (I36922,I37349,I37103);
DFFARX1 I_2062  ( .D(I37349), .CLK(I2350), .RSTB(I36942), .Q(I37431) );
not I_2063 (I36919,I37431);
DFFARX1 I_2064  ( .D(I166216), .CLK(I2350), .RSTB(I36942), .Q(I37462) );
not I_2065 (I37479,I37462);
or I_2066 (I37496,I37479,I37400);
DFFARX1 I_2067  ( .D(I37496), .CLK(I2350), .RSTB(I36942), .Q(I36925) );
nand I_2068 (I36934,I37479,I37205);
DFFARX1 I_2069  ( .D(I37479), .CLK(I2350), .RSTB(I36942), .Q(I36904) );
not I_2070 (I37588,I2357);
not I_2071 (I37605,I202417);
nor I_2072 (I37622,I202429,I202411);
nand I_2073 (I37639,I37622,I202426);
DFFARX1 I_2074  ( .D(I37639), .CLK(I2350), .RSTB(I37588), .Q(I37562) );
nor I_2075 (I37670,I37605,I202429);
nand I_2076 (I37687,I37670,I202414);
not I_2077 (I37577,I37687);
DFFARX1 I_2078  ( .D(I37687), .CLK(I2350), .RSTB(I37588), .Q(I37559) );
not I_2079 (I37732,I202429);
not I_2080 (I37749,I37732);
not I_2081 (I37766,I202423);
nor I_2082 (I37783,I37766,I202402);
and I_2083 (I37800,I37783,I202405);
or I_2084 (I37817,I37800,I202408);
DFFARX1 I_2085  ( .D(I37817), .CLK(I2350), .RSTB(I37588), .Q(I37834) );
nor I_2086 (I37851,I37834,I37687);
nor I_2087 (I37868,I37834,I37749);
nand I_2088 (I37574,I37639,I37868);
nand I_2089 (I37899,I37605,I202423);
nand I_2090 (I37916,I37899,I37834);
and I_2091 (I37933,I37899,I37916);
DFFARX1 I_2092  ( .D(I37933), .CLK(I2350), .RSTB(I37588), .Q(I37556) );
DFFARX1 I_2093  ( .D(I37899), .CLK(I2350), .RSTB(I37588), .Q(I37964) );
and I_2094 (I37553,I37732,I37964);
DFFARX1 I_2095  ( .D(I202399), .CLK(I2350), .RSTB(I37588), .Q(I37995) );
not I_2096 (I38012,I37995);
nor I_2097 (I38029,I37687,I38012);
and I_2098 (I38046,I37995,I38029);
nand I_2099 (I37568,I37995,I37749);
DFFARX1 I_2100  ( .D(I37995), .CLK(I2350), .RSTB(I37588), .Q(I38077) );
not I_2101 (I37565,I38077);
DFFARX1 I_2102  ( .D(I202420), .CLK(I2350), .RSTB(I37588), .Q(I38108) );
not I_2103 (I38125,I38108);
or I_2104 (I38142,I38125,I38046);
DFFARX1 I_2105  ( .D(I38142), .CLK(I2350), .RSTB(I37588), .Q(I37571) );
nand I_2106 (I37580,I38125,I37851);
DFFARX1 I_2107  ( .D(I38125), .CLK(I2350), .RSTB(I37588), .Q(I37550) );
not I_2108 (I38234,I2357);
not I_2109 (I38251,I216629);
nor I_2110 (I38268,I216641,I216623);
nand I_2111 (I38285,I38268,I216638);
DFFARX1 I_2112  ( .D(I38285), .CLK(I2350), .RSTB(I38234), .Q(I38208) );
nor I_2113 (I38316,I38251,I216641);
nand I_2114 (I38333,I38316,I216626);
not I_2115 (I38223,I38333);
DFFARX1 I_2116  ( .D(I38333), .CLK(I2350), .RSTB(I38234), .Q(I38205) );
not I_2117 (I38378,I216641);
not I_2118 (I38395,I38378);
not I_2119 (I38412,I216635);
nor I_2120 (I38429,I38412,I216614);
and I_2121 (I38446,I38429,I216617);
or I_2122 (I38463,I38446,I216620);
DFFARX1 I_2123  ( .D(I38463), .CLK(I2350), .RSTB(I38234), .Q(I38480) );
nor I_2124 (I38497,I38480,I38333);
nor I_2125 (I38514,I38480,I38395);
nand I_2126 (I38220,I38285,I38514);
nand I_2127 (I38545,I38251,I216635);
nand I_2128 (I38562,I38545,I38480);
and I_2129 (I38579,I38545,I38562);
DFFARX1 I_2130  ( .D(I38579), .CLK(I2350), .RSTB(I38234), .Q(I38202) );
DFFARX1 I_2131  ( .D(I38545), .CLK(I2350), .RSTB(I38234), .Q(I38610) );
and I_2132 (I38199,I38378,I38610);
DFFARX1 I_2133  ( .D(I216611), .CLK(I2350), .RSTB(I38234), .Q(I38641) );
not I_2134 (I38658,I38641);
nor I_2135 (I38675,I38333,I38658);
and I_2136 (I38692,I38641,I38675);
nand I_2137 (I38214,I38641,I38395);
DFFARX1 I_2138  ( .D(I38641), .CLK(I2350), .RSTB(I38234), .Q(I38723) );
not I_2139 (I38211,I38723);
DFFARX1 I_2140  ( .D(I216632), .CLK(I2350), .RSTB(I38234), .Q(I38754) );
not I_2141 (I38771,I38754);
or I_2142 (I38788,I38771,I38692);
DFFARX1 I_2143  ( .D(I38788), .CLK(I2350), .RSTB(I38234), .Q(I38217) );
nand I_2144 (I38226,I38771,I38497);
DFFARX1 I_2145  ( .D(I38771), .CLK(I2350), .RSTB(I38234), .Q(I38196) );
not I_2146 (I38880,I2357);
not I_2147 (I38897,I381044);
nor I_2148 (I38914,I381041,I381038);
nand I_2149 (I38931,I38914,I381059);
DFFARX1 I_2150  ( .D(I38931), .CLK(I2350), .RSTB(I38880), .Q(I38854) );
nor I_2151 (I38962,I38897,I381041);
nand I_2152 (I38979,I38962,I381062);
not I_2153 (I38869,I38979);
DFFARX1 I_2154  ( .D(I38979), .CLK(I2350), .RSTB(I38880), .Q(I38851) );
not I_2155 (I39024,I381041);
not I_2156 (I39041,I39024);
not I_2157 (I39058,I381035);
nor I_2158 (I39075,I39058,I381047);
and I_2159 (I39092,I39075,I381056);
or I_2160 (I39109,I39092,I381050);
DFFARX1 I_2161  ( .D(I39109), .CLK(I2350), .RSTB(I38880), .Q(I39126) );
nor I_2162 (I39143,I39126,I38979);
nor I_2163 (I39160,I39126,I39041);
nand I_2164 (I38866,I38931,I39160);
nand I_2165 (I39191,I38897,I381035);
nand I_2166 (I39208,I39191,I39126);
and I_2167 (I39225,I39191,I39208);
DFFARX1 I_2168  ( .D(I39225), .CLK(I2350), .RSTB(I38880), .Q(I38848) );
DFFARX1 I_2169  ( .D(I39191), .CLK(I2350), .RSTB(I38880), .Q(I39256) );
and I_2170 (I38845,I39024,I39256);
DFFARX1 I_2171  ( .D(I381065), .CLK(I2350), .RSTB(I38880), .Q(I39287) );
not I_2172 (I39304,I39287);
nor I_2173 (I39321,I38979,I39304);
and I_2174 (I39338,I39287,I39321);
nand I_2175 (I38860,I39287,I39041);
DFFARX1 I_2176  ( .D(I39287), .CLK(I2350), .RSTB(I38880), .Q(I39369) );
not I_2177 (I38857,I39369);
DFFARX1 I_2178  ( .D(I381053), .CLK(I2350), .RSTB(I38880), .Q(I39400) );
not I_2179 (I39417,I39400);
or I_2180 (I39434,I39417,I39338);
DFFARX1 I_2181  ( .D(I39434), .CLK(I2350), .RSTB(I38880), .Q(I38863) );
nand I_2182 (I38872,I39417,I39143);
DFFARX1 I_2183  ( .D(I39417), .CLK(I2350), .RSTB(I38880), .Q(I38842) );
not I_2184 (I39526,I2357);
not I_2185 (I39543,I310614);
nor I_2186 (I39560,I310590,I310596);
nand I_2187 (I39577,I39560,I310599);
DFFARX1 I_2188  ( .D(I39577), .CLK(I2350), .RSTB(I39526), .Q(I39500) );
nor I_2189 (I39608,I39543,I310590);
nand I_2190 (I39625,I39608,I310608);
not I_2191 (I39515,I39625);
DFFARX1 I_2192  ( .D(I39625), .CLK(I2350), .RSTB(I39526), .Q(I39497) );
not I_2193 (I39670,I310590);
not I_2194 (I39687,I39670);
not I_2195 (I39704,I310587);
nor I_2196 (I39721,I39704,I310602);
and I_2197 (I39738,I39721,I310593);
or I_2198 (I39755,I39738,I310605);
DFFARX1 I_2199  ( .D(I39755), .CLK(I2350), .RSTB(I39526), .Q(I39772) );
nor I_2200 (I39789,I39772,I39625);
nor I_2201 (I39806,I39772,I39687);
nand I_2202 (I39512,I39577,I39806);
nand I_2203 (I39837,I39543,I310587);
nand I_2204 (I39854,I39837,I39772);
and I_2205 (I39871,I39837,I39854);
DFFARX1 I_2206  ( .D(I39871), .CLK(I2350), .RSTB(I39526), .Q(I39494) );
DFFARX1 I_2207  ( .D(I39837), .CLK(I2350), .RSTB(I39526), .Q(I39902) );
and I_2208 (I39491,I39670,I39902);
DFFARX1 I_2209  ( .D(I310617), .CLK(I2350), .RSTB(I39526), .Q(I39933) );
not I_2210 (I39950,I39933);
nor I_2211 (I39967,I39625,I39950);
and I_2212 (I39984,I39933,I39967);
nand I_2213 (I39506,I39933,I39687);
DFFARX1 I_2214  ( .D(I39933), .CLK(I2350), .RSTB(I39526), .Q(I40015) );
not I_2215 (I39503,I40015);
DFFARX1 I_2216  ( .D(I310611), .CLK(I2350), .RSTB(I39526), .Q(I40046) );
not I_2217 (I40063,I40046);
or I_2218 (I40080,I40063,I39984);
DFFARX1 I_2219  ( .D(I40080), .CLK(I2350), .RSTB(I39526), .Q(I39509) );
nand I_2220 (I39518,I40063,I39789);
DFFARX1 I_2221  ( .D(I40063), .CLK(I2350), .RSTB(I39526), .Q(I39488) );
not I_2222 (I40172,I2357);
not I_2223 (I40189,I256236);
nor I_2224 (I40206,I256224,I256230);
nand I_2225 (I40223,I40206,I256221);
DFFARX1 I_2226  ( .D(I40223), .CLK(I2350), .RSTB(I40172), .Q(I40146) );
nor I_2227 (I40254,I40189,I256224);
nand I_2228 (I40271,I40254,I256227);
not I_2229 (I40161,I40271);
DFFARX1 I_2230  ( .D(I40271), .CLK(I2350), .RSTB(I40172), .Q(I40143) );
not I_2231 (I40316,I256224);
not I_2232 (I40333,I40316);
not I_2233 (I40350,I256239);
nor I_2234 (I40367,I40350,I256251);
and I_2235 (I40384,I40367,I256233);
or I_2236 (I40401,I40384,I256248);
DFFARX1 I_2237  ( .D(I40401), .CLK(I2350), .RSTB(I40172), .Q(I40418) );
nor I_2238 (I40435,I40418,I40271);
nor I_2239 (I40452,I40418,I40333);
nand I_2240 (I40158,I40223,I40452);
nand I_2241 (I40483,I40189,I256239);
nand I_2242 (I40500,I40483,I40418);
and I_2243 (I40517,I40483,I40500);
DFFARX1 I_2244  ( .D(I40517), .CLK(I2350), .RSTB(I40172), .Q(I40140) );
DFFARX1 I_2245  ( .D(I40483), .CLK(I2350), .RSTB(I40172), .Q(I40548) );
and I_2246 (I40137,I40316,I40548);
DFFARX1 I_2247  ( .D(I256242), .CLK(I2350), .RSTB(I40172), .Q(I40579) );
not I_2248 (I40596,I40579);
nor I_2249 (I40613,I40271,I40596);
and I_2250 (I40630,I40579,I40613);
nand I_2251 (I40152,I40579,I40333);
DFFARX1 I_2252  ( .D(I40579), .CLK(I2350), .RSTB(I40172), .Q(I40661) );
not I_2253 (I40149,I40661);
DFFARX1 I_2254  ( .D(I256245), .CLK(I2350), .RSTB(I40172), .Q(I40692) );
not I_2255 (I40709,I40692);
or I_2256 (I40726,I40709,I40630);
DFFARX1 I_2257  ( .D(I40726), .CLK(I2350), .RSTB(I40172), .Q(I40155) );
nand I_2258 (I40164,I40709,I40435);
DFFARX1 I_2259  ( .D(I40709), .CLK(I2350), .RSTB(I40172), .Q(I40134) );
not I_2260 (I40818,I2357);
not I_2261 (I40835,I383356);
nor I_2262 (I40852,I383353,I383350);
nand I_2263 (I40869,I40852,I383371);
DFFARX1 I_2264  ( .D(I40869), .CLK(I2350), .RSTB(I40818), .Q(I40792) );
nor I_2265 (I40900,I40835,I383353);
nand I_2266 (I40917,I40900,I383374);
not I_2267 (I40807,I40917);
DFFARX1 I_2268  ( .D(I40917), .CLK(I2350), .RSTB(I40818), .Q(I40789) );
not I_2269 (I40962,I383353);
not I_2270 (I40979,I40962);
not I_2271 (I40996,I383347);
nor I_2272 (I41013,I40996,I383359);
and I_2273 (I41030,I41013,I383368);
or I_2274 (I41047,I41030,I383362);
DFFARX1 I_2275  ( .D(I41047), .CLK(I2350), .RSTB(I40818), .Q(I41064) );
nor I_2276 (I41081,I41064,I40917);
nor I_2277 (I41098,I41064,I40979);
nand I_2278 (I40804,I40869,I41098);
nand I_2279 (I41129,I40835,I383347);
nand I_2280 (I41146,I41129,I41064);
and I_2281 (I41163,I41129,I41146);
DFFARX1 I_2282  ( .D(I41163), .CLK(I2350), .RSTB(I40818), .Q(I40786) );
DFFARX1 I_2283  ( .D(I41129), .CLK(I2350), .RSTB(I40818), .Q(I41194) );
and I_2284 (I40783,I40962,I41194);
DFFARX1 I_2285  ( .D(I383377), .CLK(I2350), .RSTB(I40818), .Q(I41225) );
not I_2286 (I41242,I41225);
nor I_2287 (I41259,I40917,I41242);
and I_2288 (I41276,I41225,I41259);
nand I_2289 (I40798,I41225,I40979);
DFFARX1 I_2290  ( .D(I41225), .CLK(I2350), .RSTB(I40818), .Q(I41307) );
not I_2291 (I40795,I41307);
DFFARX1 I_2292  ( .D(I383365), .CLK(I2350), .RSTB(I40818), .Q(I41338) );
not I_2293 (I41355,I41338);
or I_2294 (I41372,I41355,I41276);
DFFARX1 I_2295  ( .D(I41372), .CLK(I2350), .RSTB(I40818), .Q(I40801) );
nand I_2296 (I40810,I41355,I41081);
DFFARX1 I_2297  ( .D(I41355), .CLK(I2350), .RSTB(I40818), .Q(I40780) );
not I_2298 (I41464,I2357);
not I_2299 (I41481,I308829);
nor I_2300 (I41498,I308805,I308811);
nand I_2301 (I41515,I41498,I308814);
DFFARX1 I_2302  ( .D(I41515), .CLK(I2350), .RSTB(I41464), .Q(I41438) );
nor I_2303 (I41546,I41481,I308805);
nand I_2304 (I41563,I41546,I308823);
not I_2305 (I41453,I41563);
DFFARX1 I_2306  ( .D(I41563), .CLK(I2350), .RSTB(I41464), .Q(I41435) );
not I_2307 (I41608,I308805);
not I_2308 (I41625,I41608);
not I_2309 (I41642,I308802);
nor I_2310 (I41659,I41642,I308817);
and I_2311 (I41676,I41659,I308808);
or I_2312 (I41693,I41676,I308820);
DFFARX1 I_2313  ( .D(I41693), .CLK(I2350), .RSTB(I41464), .Q(I41710) );
nor I_2314 (I41727,I41710,I41563);
nor I_2315 (I41744,I41710,I41625);
nand I_2316 (I41450,I41515,I41744);
nand I_2317 (I41775,I41481,I308802);
nand I_2318 (I41792,I41775,I41710);
and I_2319 (I41809,I41775,I41792);
DFFARX1 I_2320  ( .D(I41809), .CLK(I2350), .RSTB(I41464), .Q(I41432) );
DFFARX1 I_2321  ( .D(I41775), .CLK(I2350), .RSTB(I41464), .Q(I41840) );
and I_2322 (I41429,I41608,I41840);
DFFARX1 I_2323  ( .D(I308832), .CLK(I2350), .RSTB(I41464), .Q(I41871) );
not I_2324 (I41888,I41871);
nor I_2325 (I41905,I41563,I41888);
and I_2326 (I41922,I41871,I41905);
nand I_2327 (I41444,I41871,I41625);
DFFARX1 I_2328  ( .D(I41871), .CLK(I2350), .RSTB(I41464), .Q(I41953) );
not I_2329 (I41441,I41953);
DFFARX1 I_2330  ( .D(I308826), .CLK(I2350), .RSTB(I41464), .Q(I41984) );
not I_2331 (I42001,I41984);
or I_2332 (I42018,I42001,I41922);
DFFARX1 I_2333  ( .D(I42018), .CLK(I2350), .RSTB(I41464), .Q(I41447) );
nand I_2334 (I41456,I42001,I41727);
DFFARX1 I_2335  ( .D(I42001), .CLK(I2350), .RSTB(I41464), .Q(I41426) );
not I_2336 (I42110,I2357);
not I_2337 (I42127,I288599);
nor I_2338 (I42144,I288575,I288581);
nand I_2339 (I42161,I42144,I288584);
DFFARX1 I_2340  ( .D(I42161), .CLK(I2350), .RSTB(I42110), .Q(I42084) );
nor I_2341 (I42192,I42127,I288575);
nand I_2342 (I42209,I42192,I288593);
not I_2343 (I42099,I42209);
DFFARX1 I_2344  ( .D(I42209), .CLK(I2350), .RSTB(I42110), .Q(I42081) );
not I_2345 (I42254,I288575);
not I_2346 (I42271,I42254);
not I_2347 (I42288,I288572);
nor I_2348 (I42305,I42288,I288587);
and I_2349 (I42322,I42305,I288578);
or I_2350 (I42339,I42322,I288590);
DFFARX1 I_2351  ( .D(I42339), .CLK(I2350), .RSTB(I42110), .Q(I42356) );
nor I_2352 (I42373,I42356,I42209);
nor I_2353 (I42390,I42356,I42271);
nand I_2354 (I42096,I42161,I42390);
nand I_2355 (I42421,I42127,I288572);
nand I_2356 (I42438,I42421,I42356);
and I_2357 (I42455,I42421,I42438);
DFFARX1 I_2358  ( .D(I42455), .CLK(I2350), .RSTB(I42110), .Q(I42078) );
DFFARX1 I_2359  ( .D(I42421), .CLK(I2350), .RSTB(I42110), .Q(I42486) );
and I_2360 (I42075,I42254,I42486);
DFFARX1 I_2361  ( .D(I288602), .CLK(I2350), .RSTB(I42110), .Q(I42517) );
not I_2362 (I42534,I42517);
nor I_2363 (I42551,I42209,I42534);
and I_2364 (I42568,I42517,I42551);
nand I_2365 (I42090,I42517,I42271);
DFFARX1 I_2366  ( .D(I42517), .CLK(I2350), .RSTB(I42110), .Q(I42599) );
not I_2367 (I42087,I42599);
DFFARX1 I_2368  ( .D(I288596), .CLK(I2350), .RSTB(I42110), .Q(I42630) );
not I_2369 (I42647,I42630);
or I_2370 (I42664,I42647,I42568);
DFFARX1 I_2371  ( .D(I42664), .CLK(I2350), .RSTB(I42110), .Q(I42093) );
nand I_2372 (I42102,I42647,I42373);
DFFARX1 I_2373  ( .D(I42647), .CLK(I2350), .RSTB(I42110), .Q(I42072) );
not I_2374 (I42756,I2357);
not I_2375 (I42773,I19754);
nor I_2376 (I42790,I19766,I19751);
nand I_2377 (I42807,I42790,I19763);
DFFARX1 I_2378  ( .D(I42807), .CLK(I2350), .RSTB(I42756), .Q(I42730) );
nor I_2379 (I42838,I42773,I19766);
nand I_2380 (I42855,I42838,I19781);
not I_2381 (I42745,I42855);
DFFARX1 I_2382  ( .D(I42855), .CLK(I2350), .RSTB(I42756), .Q(I42727) );
not I_2383 (I42900,I19766);
not I_2384 (I42917,I42900);
not I_2385 (I42934,I19757);
nor I_2386 (I42951,I42934,I19769);
and I_2387 (I42968,I42951,I19760);
or I_2388 (I42985,I42968,I19775);
DFFARX1 I_2389  ( .D(I42985), .CLK(I2350), .RSTB(I42756), .Q(I43002) );
nor I_2390 (I43019,I43002,I42855);
nor I_2391 (I43036,I43002,I42917);
nand I_2392 (I42742,I42807,I43036);
nand I_2393 (I43067,I42773,I19757);
nand I_2394 (I43084,I43067,I43002);
and I_2395 (I43101,I43067,I43084);
DFFARX1 I_2396  ( .D(I43101), .CLK(I2350), .RSTB(I42756), .Q(I42724) );
DFFARX1 I_2397  ( .D(I43067), .CLK(I2350), .RSTB(I42756), .Q(I43132) );
and I_2398 (I42721,I42900,I43132);
DFFARX1 I_2399  ( .D(I19778), .CLK(I2350), .RSTB(I42756), .Q(I43163) );
not I_2400 (I43180,I43163);
nor I_2401 (I43197,I42855,I43180);
and I_2402 (I43214,I43163,I43197);
nand I_2403 (I42736,I43163,I42917);
DFFARX1 I_2404  ( .D(I43163), .CLK(I2350), .RSTB(I42756), .Q(I43245) );
not I_2405 (I42733,I43245);
DFFARX1 I_2406  ( .D(I19772), .CLK(I2350), .RSTB(I42756), .Q(I43276) );
not I_2407 (I43293,I43276);
or I_2408 (I43310,I43293,I43214);
DFFARX1 I_2409  ( .D(I43310), .CLK(I2350), .RSTB(I42756), .Q(I42739) );
nand I_2410 (I42748,I43293,I43019);
DFFARX1 I_2411  ( .D(I43293), .CLK(I2350), .RSTB(I42756), .Q(I42718) );
not I_2412 (I43402,I2357);
not I_2413 (I43419,I364052);
nor I_2414 (I43436,I364067,I364082);
nand I_2415 (I43453,I43436,I364070);
DFFARX1 I_2416  ( .D(I43453), .CLK(I2350), .RSTB(I43402), .Q(I43376) );
nor I_2417 (I43484,I43419,I364067);
nand I_2418 (I43501,I43484,I364073);
not I_2419 (I43391,I43501);
DFFARX1 I_2420  ( .D(I43501), .CLK(I2350), .RSTB(I43402), .Q(I43373) );
not I_2421 (I43546,I364067);
not I_2422 (I43563,I43546);
not I_2423 (I43580,I364079);
nor I_2424 (I43597,I43580,I364076);
and I_2425 (I43614,I43597,I364055);
or I_2426 (I43631,I43614,I364064);
DFFARX1 I_2427  ( .D(I43631), .CLK(I2350), .RSTB(I43402), .Q(I43648) );
nor I_2428 (I43665,I43648,I43501);
nor I_2429 (I43682,I43648,I43563);
nand I_2430 (I43388,I43453,I43682);
nand I_2431 (I43713,I43419,I364079);
nand I_2432 (I43730,I43713,I43648);
and I_2433 (I43747,I43713,I43730);
DFFARX1 I_2434  ( .D(I43747), .CLK(I2350), .RSTB(I43402), .Q(I43370) );
DFFARX1 I_2435  ( .D(I43713), .CLK(I2350), .RSTB(I43402), .Q(I43778) );
and I_2436 (I43367,I43546,I43778);
DFFARX1 I_2437  ( .D(I364061), .CLK(I2350), .RSTB(I43402), .Q(I43809) );
not I_2438 (I43826,I43809);
nor I_2439 (I43843,I43501,I43826);
and I_2440 (I43860,I43809,I43843);
nand I_2441 (I43382,I43809,I43563);
DFFARX1 I_2442  ( .D(I43809), .CLK(I2350), .RSTB(I43402), .Q(I43891) );
not I_2443 (I43379,I43891);
DFFARX1 I_2444  ( .D(I364058), .CLK(I2350), .RSTB(I43402), .Q(I43922) );
not I_2445 (I43939,I43922);
or I_2446 (I43956,I43939,I43860);
DFFARX1 I_2447  ( .D(I43956), .CLK(I2350), .RSTB(I43402), .Q(I43385) );
nand I_2448 (I43394,I43939,I43665);
DFFARX1 I_2449  ( .D(I43939), .CLK(I2350), .RSTB(I43402), .Q(I43364) );
not I_2450 (I44048,I2357);
not I_2451 (I44065,I203063);
nor I_2452 (I44082,I203075,I203057);
nand I_2453 (I44099,I44082,I203072);
DFFARX1 I_2454  ( .D(I44099), .CLK(I2350), .RSTB(I44048), .Q(I44022) );
nor I_2455 (I44130,I44065,I203075);
nand I_2456 (I44147,I44130,I203060);
not I_2457 (I44037,I44147);
DFFARX1 I_2458  ( .D(I44147), .CLK(I2350), .RSTB(I44048), .Q(I44019) );
not I_2459 (I44192,I203075);
not I_2460 (I44209,I44192);
not I_2461 (I44226,I203069);
nor I_2462 (I44243,I44226,I203048);
and I_2463 (I44260,I44243,I203051);
or I_2464 (I44277,I44260,I203054);
DFFARX1 I_2465  ( .D(I44277), .CLK(I2350), .RSTB(I44048), .Q(I44294) );
nor I_2466 (I44311,I44294,I44147);
nor I_2467 (I44328,I44294,I44209);
nand I_2468 (I44034,I44099,I44328);
nand I_2469 (I44359,I44065,I203069);
nand I_2470 (I44376,I44359,I44294);
and I_2471 (I44393,I44359,I44376);
DFFARX1 I_2472  ( .D(I44393), .CLK(I2350), .RSTB(I44048), .Q(I44016) );
DFFARX1 I_2473  ( .D(I44359), .CLK(I2350), .RSTB(I44048), .Q(I44424) );
and I_2474 (I44013,I44192,I44424);
DFFARX1 I_2475  ( .D(I203045), .CLK(I2350), .RSTB(I44048), .Q(I44455) );
not I_2476 (I44472,I44455);
nor I_2477 (I44489,I44147,I44472);
and I_2478 (I44506,I44455,I44489);
nand I_2479 (I44028,I44455,I44209);
DFFARX1 I_2480  ( .D(I44455), .CLK(I2350), .RSTB(I44048), .Q(I44537) );
not I_2481 (I44025,I44537);
DFFARX1 I_2482  ( .D(I203066), .CLK(I2350), .RSTB(I44048), .Q(I44568) );
not I_2483 (I44585,I44568);
or I_2484 (I44602,I44585,I44506);
DFFARX1 I_2485  ( .D(I44602), .CLK(I2350), .RSTB(I44048), .Q(I44031) );
nand I_2486 (I44040,I44585,I44311);
DFFARX1 I_2487  ( .D(I44585), .CLK(I2350), .RSTB(I44048), .Q(I44010) );
not I_2488 (I44694,I2357);
not I_2489 (I44711,I135306);
nor I_2490 (I44728,I135327,I135300);
nand I_2491 (I44745,I44728,I135315);
DFFARX1 I_2492  ( .D(I44745), .CLK(I2350), .RSTB(I44694), .Q(I44668) );
nor I_2493 (I44776,I44711,I135327);
nand I_2494 (I44793,I44776,I135330);
not I_2495 (I44683,I44793);
DFFARX1 I_2496  ( .D(I44793), .CLK(I2350), .RSTB(I44694), .Q(I44665) );
not I_2497 (I44838,I135327);
not I_2498 (I44855,I44838);
not I_2499 (I44872,I135303);
nor I_2500 (I44889,I44872,I135321);
and I_2501 (I44906,I44889,I135309);
or I_2502 (I44923,I44906,I135312);
DFFARX1 I_2503  ( .D(I44923), .CLK(I2350), .RSTB(I44694), .Q(I44940) );
nor I_2504 (I44957,I44940,I44793);
nor I_2505 (I44974,I44940,I44855);
nand I_2506 (I44680,I44745,I44974);
nand I_2507 (I45005,I44711,I135303);
nand I_2508 (I45022,I45005,I44940);
and I_2509 (I45039,I45005,I45022);
DFFARX1 I_2510  ( .D(I45039), .CLK(I2350), .RSTB(I44694), .Q(I44662) );
DFFARX1 I_2511  ( .D(I45005), .CLK(I2350), .RSTB(I44694), .Q(I45070) );
and I_2512 (I44659,I44838,I45070);
DFFARX1 I_2513  ( .D(I135324), .CLK(I2350), .RSTB(I44694), .Q(I45101) );
not I_2514 (I45118,I45101);
nor I_2515 (I45135,I44793,I45118);
and I_2516 (I45152,I45101,I45135);
nand I_2517 (I44674,I45101,I44855);
DFFARX1 I_2518  ( .D(I45101), .CLK(I2350), .RSTB(I44694), .Q(I45183) );
not I_2519 (I44671,I45183);
DFFARX1 I_2520  ( .D(I135318), .CLK(I2350), .RSTB(I44694), .Q(I45214) );
not I_2521 (I45231,I45214);
or I_2522 (I45248,I45231,I45152);
DFFARX1 I_2523  ( .D(I45248), .CLK(I2350), .RSTB(I44694), .Q(I44677) );
nand I_2524 (I44686,I45231,I44957);
DFFARX1 I_2525  ( .D(I45231), .CLK(I2350), .RSTB(I44694), .Q(I44656) );
not I_2526 (I45340,I2357);
not I_2527 (I45357,I256814);
nor I_2528 (I45374,I256802,I256808);
nand I_2529 (I45391,I45374,I256799);
DFFARX1 I_2530  ( .D(I45391), .CLK(I2350), .RSTB(I45340), .Q(I45314) );
nor I_2531 (I45422,I45357,I256802);
nand I_2532 (I45439,I45422,I256805);
not I_2533 (I45329,I45439);
DFFARX1 I_2534  ( .D(I45439), .CLK(I2350), .RSTB(I45340), .Q(I45311) );
not I_2535 (I45484,I256802);
not I_2536 (I45501,I45484);
not I_2537 (I45518,I256817);
nor I_2538 (I45535,I45518,I256829);
and I_2539 (I45552,I45535,I256811);
or I_2540 (I45569,I45552,I256826);
DFFARX1 I_2541  ( .D(I45569), .CLK(I2350), .RSTB(I45340), .Q(I45586) );
nor I_2542 (I45603,I45586,I45439);
nor I_2543 (I45620,I45586,I45501);
nand I_2544 (I45326,I45391,I45620);
nand I_2545 (I45651,I45357,I256817);
nand I_2546 (I45668,I45651,I45586);
and I_2547 (I45685,I45651,I45668);
DFFARX1 I_2548  ( .D(I45685), .CLK(I2350), .RSTB(I45340), .Q(I45308) );
DFFARX1 I_2549  ( .D(I45651), .CLK(I2350), .RSTB(I45340), .Q(I45716) );
and I_2550 (I45305,I45484,I45716);
DFFARX1 I_2551  ( .D(I256820), .CLK(I2350), .RSTB(I45340), .Q(I45747) );
not I_2552 (I45764,I45747);
nor I_2553 (I45781,I45439,I45764);
and I_2554 (I45798,I45747,I45781);
nand I_2555 (I45320,I45747,I45501);
DFFARX1 I_2556  ( .D(I45747), .CLK(I2350), .RSTB(I45340), .Q(I45829) );
not I_2557 (I45317,I45829);
DFFARX1 I_2558  ( .D(I256823), .CLK(I2350), .RSTB(I45340), .Q(I45860) );
not I_2559 (I45877,I45860);
or I_2560 (I45894,I45877,I45798);
DFFARX1 I_2561  ( .D(I45894), .CLK(I2350), .RSTB(I45340), .Q(I45323) );
nand I_2562 (I45332,I45877,I45603);
DFFARX1 I_2563  ( .D(I45877), .CLK(I2350), .RSTB(I45340), .Q(I45302) );
not I_2564 (I45986,I2357);
not I_2565 (I46003,I326072);
nor I_2566 (I46020,I326057,I326084);
nand I_2567 (I46037,I46020,I326060);
DFFARX1 I_2568  ( .D(I46037), .CLK(I2350), .RSTB(I45986), .Q(I45960) );
nor I_2569 (I46068,I46003,I326057);
nand I_2570 (I46085,I46068,I326075);
not I_2571 (I45975,I46085);
DFFARX1 I_2572  ( .D(I46085), .CLK(I2350), .RSTB(I45986), .Q(I45957) );
not I_2573 (I46130,I326057);
not I_2574 (I46147,I46130);
not I_2575 (I46164,I326087);
nor I_2576 (I46181,I46164,I326069);
and I_2577 (I46198,I46181,I326078);
or I_2578 (I46215,I46198,I326063);
DFFARX1 I_2579  ( .D(I46215), .CLK(I2350), .RSTB(I45986), .Q(I46232) );
nor I_2580 (I46249,I46232,I46085);
nor I_2581 (I46266,I46232,I46147);
nand I_2582 (I45972,I46037,I46266);
nand I_2583 (I46297,I46003,I326087);
nand I_2584 (I46314,I46297,I46232);
and I_2585 (I46331,I46297,I46314);
DFFARX1 I_2586  ( .D(I46331), .CLK(I2350), .RSTB(I45986), .Q(I45954) );
DFFARX1 I_2587  ( .D(I46297), .CLK(I2350), .RSTB(I45986), .Q(I46362) );
and I_2588 (I45951,I46130,I46362);
DFFARX1 I_2589  ( .D(I326066), .CLK(I2350), .RSTB(I45986), .Q(I46393) );
not I_2590 (I46410,I46393);
nor I_2591 (I46427,I46085,I46410);
and I_2592 (I46444,I46393,I46427);
nand I_2593 (I45966,I46393,I46147);
DFFARX1 I_2594  ( .D(I46393), .CLK(I2350), .RSTB(I45986), .Q(I46475) );
not I_2595 (I45963,I46475);
DFFARX1 I_2596  ( .D(I326081), .CLK(I2350), .RSTB(I45986), .Q(I46506) );
not I_2597 (I46523,I46506);
or I_2598 (I46540,I46523,I46444);
DFFARX1 I_2599  ( .D(I46540), .CLK(I2350), .RSTB(I45986), .Q(I45969) );
nand I_2600 (I45978,I46523,I46249);
DFFARX1 I_2601  ( .D(I46523), .CLK(I2350), .RSTB(I45986), .Q(I45948) );
not I_2602 (I46632,I2357);
not I_2603 (I46649,I385668);
nor I_2604 (I46666,I385665,I385662);
nand I_2605 (I46683,I46666,I385683);
DFFARX1 I_2606  ( .D(I46683), .CLK(I2350), .RSTB(I46632), .Q(I46606) );
nor I_2607 (I46714,I46649,I385665);
nand I_2608 (I46731,I46714,I385686);
not I_2609 (I46621,I46731);
DFFARX1 I_2610  ( .D(I46731), .CLK(I2350), .RSTB(I46632), .Q(I46603) );
not I_2611 (I46776,I385665);
not I_2612 (I46793,I46776);
not I_2613 (I46810,I385659);
nor I_2614 (I46827,I46810,I385671);
and I_2615 (I46844,I46827,I385680);
or I_2616 (I46861,I46844,I385674);
DFFARX1 I_2617  ( .D(I46861), .CLK(I2350), .RSTB(I46632), .Q(I46878) );
nor I_2618 (I46895,I46878,I46731);
nor I_2619 (I46912,I46878,I46793);
nand I_2620 (I46618,I46683,I46912);
nand I_2621 (I46943,I46649,I385659);
nand I_2622 (I46960,I46943,I46878);
and I_2623 (I46977,I46943,I46960);
DFFARX1 I_2624  ( .D(I46977), .CLK(I2350), .RSTB(I46632), .Q(I46600) );
DFFARX1 I_2625  ( .D(I46943), .CLK(I2350), .RSTB(I46632), .Q(I47008) );
and I_2626 (I46597,I46776,I47008);
DFFARX1 I_2627  ( .D(I385689), .CLK(I2350), .RSTB(I46632), .Q(I47039) );
not I_2628 (I47056,I47039);
nor I_2629 (I47073,I46731,I47056);
and I_2630 (I47090,I47039,I47073);
nand I_2631 (I46612,I47039,I46793);
DFFARX1 I_2632  ( .D(I47039), .CLK(I2350), .RSTB(I46632), .Q(I47121) );
not I_2633 (I46609,I47121);
DFFARX1 I_2634  ( .D(I385677), .CLK(I2350), .RSTB(I46632), .Q(I47152) );
not I_2635 (I47169,I47152);
or I_2636 (I47186,I47169,I47090);
DFFARX1 I_2637  ( .D(I47186), .CLK(I2350), .RSTB(I46632), .Q(I46615) );
nand I_2638 (I46624,I47169,I46895);
DFFARX1 I_2639  ( .D(I47169), .CLK(I2350), .RSTB(I46632), .Q(I46594) );
not I_2640 (I47278,I2357);
not I_2641 (I47295,I144328);
nor I_2642 (I47312,I144325,I144313);
nand I_2643 (I47329,I47312,I144316);
DFFARX1 I_2644  ( .D(I47329), .CLK(I2350), .RSTB(I47278), .Q(I47252) );
nor I_2645 (I47360,I47295,I144325);
nand I_2646 (I47377,I47360,I144322);
not I_2647 (I47267,I47377);
DFFARX1 I_2648  ( .D(I47377), .CLK(I2350), .RSTB(I47278), .Q(I47249) );
not I_2649 (I47422,I144325);
not I_2650 (I47439,I47422);
not I_2651 (I47456,I144334);
nor I_2652 (I47473,I47456,I144310);
and I_2653 (I47490,I47473,I144331);
or I_2654 (I47507,I47490,I144319);
DFFARX1 I_2655  ( .D(I47507), .CLK(I2350), .RSTB(I47278), .Q(I47524) );
nor I_2656 (I47541,I47524,I47377);
nor I_2657 (I47558,I47524,I47439);
nand I_2658 (I47264,I47329,I47558);
nand I_2659 (I47589,I47295,I144334);
nand I_2660 (I47606,I47589,I47524);
and I_2661 (I47623,I47589,I47606);
DFFARX1 I_2662  ( .D(I47623), .CLK(I2350), .RSTB(I47278), .Q(I47246) );
DFFARX1 I_2663  ( .D(I47589), .CLK(I2350), .RSTB(I47278), .Q(I47654) );
and I_2664 (I47243,I47422,I47654);
DFFARX1 I_2665  ( .D(I144340), .CLK(I2350), .RSTB(I47278), .Q(I47685) );
not I_2666 (I47702,I47685);
nor I_2667 (I47719,I47377,I47702);
and I_2668 (I47736,I47685,I47719);
nand I_2669 (I47258,I47685,I47439);
DFFARX1 I_2670  ( .D(I47685), .CLK(I2350), .RSTB(I47278), .Q(I47767) );
not I_2671 (I47255,I47767);
DFFARX1 I_2672  ( .D(I144337), .CLK(I2350), .RSTB(I47278), .Q(I47798) );
not I_2673 (I47815,I47798);
or I_2674 (I47832,I47815,I47736);
DFFARX1 I_2675  ( .D(I47832), .CLK(I2350), .RSTB(I47278), .Q(I47261) );
nand I_2676 (I47270,I47815,I47541);
DFFARX1 I_2677  ( .D(I47815), .CLK(I2350), .RSTB(I47278), .Q(I47240) );
not I_2678 (I47924,I2357);
not I_2679 (I47941,I359649);
nor I_2680 (I47958,I359664,I359679);
nand I_2681 (I47975,I47958,I359667);
DFFARX1 I_2682  ( .D(I47975), .CLK(I2350), .RSTB(I47924), .Q(I47898) );
nor I_2683 (I48006,I47941,I359664);
nand I_2684 (I48023,I48006,I359670);
not I_2685 (I47913,I48023);
DFFARX1 I_2686  ( .D(I48023), .CLK(I2350), .RSTB(I47924), .Q(I47895) );
not I_2687 (I48068,I359664);
not I_2688 (I48085,I48068);
not I_2689 (I48102,I359676);
nor I_2690 (I48119,I48102,I359673);
and I_2691 (I48136,I48119,I359652);
or I_2692 (I48153,I48136,I359661);
DFFARX1 I_2693  ( .D(I48153), .CLK(I2350), .RSTB(I47924), .Q(I48170) );
nor I_2694 (I48187,I48170,I48023);
nor I_2695 (I48204,I48170,I48085);
nand I_2696 (I47910,I47975,I48204);
nand I_2697 (I48235,I47941,I359676);
nand I_2698 (I48252,I48235,I48170);
and I_2699 (I48269,I48235,I48252);
DFFARX1 I_2700  ( .D(I48269), .CLK(I2350), .RSTB(I47924), .Q(I47892) );
DFFARX1 I_2701  ( .D(I48235), .CLK(I2350), .RSTB(I47924), .Q(I48300) );
and I_2702 (I47889,I48068,I48300);
DFFARX1 I_2703  ( .D(I359658), .CLK(I2350), .RSTB(I47924), .Q(I48331) );
not I_2704 (I48348,I48331);
nor I_2705 (I48365,I48023,I48348);
and I_2706 (I48382,I48331,I48365);
nand I_2707 (I47904,I48331,I48085);
DFFARX1 I_2708  ( .D(I48331), .CLK(I2350), .RSTB(I47924), .Q(I48413) );
not I_2709 (I47901,I48413);
DFFARX1 I_2710  ( .D(I359655), .CLK(I2350), .RSTB(I47924), .Q(I48444) );
not I_2711 (I48461,I48444);
or I_2712 (I48478,I48461,I48382);
DFFARX1 I_2713  ( .D(I48478), .CLK(I2350), .RSTB(I47924), .Q(I47907) );
nand I_2714 (I47916,I48461,I48187);
DFFARX1 I_2715  ( .D(I48461), .CLK(I2350), .RSTB(I47924), .Q(I47886) );
not I_2716 (I48570,I2357);
not I_2717 (I48587,I184108);
nor I_2718 (I48604,I184105,I184093);
nand I_2719 (I48621,I48604,I184096);
DFFARX1 I_2720  ( .D(I48621), .CLK(I2350), .RSTB(I48570), .Q(I48544) );
nor I_2721 (I48652,I48587,I184105);
nand I_2722 (I48669,I48652,I184102);
not I_2723 (I48559,I48669);
DFFARX1 I_2724  ( .D(I48669), .CLK(I2350), .RSTB(I48570), .Q(I48541) );
not I_2725 (I48714,I184105);
not I_2726 (I48731,I48714);
not I_2727 (I48748,I184114);
nor I_2728 (I48765,I48748,I184090);
and I_2729 (I48782,I48765,I184111);
or I_2730 (I48799,I48782,I184099);
DFFARX1 I_2731  ( .D(I48799), .CLK(I2350), .RSTB(I48570), .Q(I48816) );
nor I_2732 (I48833,I48816,I48669);
nor I_2733 (I48850,I48816,I48731);
nand I_2734 (I48556,I48621,I48850);
nand I_2735 (I48881,I48587,I184114);
nand I_2736 (I48898,I48881,I48816);
and I_2737 (I48915,I48881,I48898);
DFFARX1 I_2738  ( .D(I48915), .CLK(I2350), .RSTB(I48570), .Q(I48538) );
DFFARX1 I_2739  ( .D(I48881), .CLK(I2350), .RSTB(I48570), .Q(I48946) );
and I_2740 (I48535,I48714,I48946);
DFFARX1 I_2741  ( .D(I184120), .CLK(I2350), .RSTB(I48570), .Q(I48977) );
not I_2742 (I48994,I48977);
nor I_2743 (I49011,I48669,I48994);
and I_2744 (I49028,I48977,I49011);
nand I_2745 (I48550,I48977,I48731);
DFFARX1 I_2746  ( .D(I48977), .CLK(I2350), .RSTB(I48570), .Q(I49059) );
not I_2747 (I48547,I49059);
DFFARX1 I_2748  ( .D(I184117), .CLK(I2350), .RSTB(I48570), .Q(I49090) );
not I_2749 (I49107,I49090);
or I_2750 (I49124,I49107,I49028);
DFFARX1 I_2751  ( .D(I49124), .CLK(I2350), .RSTB(I48570), .Q(I48553) );
nand I_2752 (I48562,I49107,I48833);
DFFARX1 I_2753  ( .D(I49107), .CLK(I2350), .RSTB(I48570), .Q(I48532) );
not I_2754 (I49216,I2357);
not I_2755 (I49233,I89367);
nor I_2756 (I49250,I89355,I89361);
nand I_2757 (I49267,I49250,I89370);
DFFARX1 I_2758  ( .D(I49267), .CLK(I2350), .RSTB(I49216), .Q(I49190) );
nor I_2759 (I49298,I49233,I89355);
nand I_2760 (I49315,I49298,I89358);
not I_2761 (I49205,I49315);
DFFARX1 I_2762  ( .D(I49315), .CLK(I2350), .RSTB(I49216), .Q(I49187) );
not I_2763 (I49360,I89355);
not I_2764 (I49377,I49360);
not I_2765 (I49394,I89379);
nor I_2766 (I49411,I49394,I89352);
and I_2767 (I49428,I49411,I89373);
or I_2768 (I49445,I49428,I89364);
DFFARX1 I_2769  ( .D(I49445), .CLK(I2350), .RSTB(I49216), .Q(I49462) );
nor I_2770 (I49479,I49462,I49315);
nor I_2771 (I49496,I49462,I49377);
nand I_2772 (I49202,I49267,I49496);
nand I_2773 (I49527,I49233,I89379);
nand I_2774 (I49544,I49527,I49462);
and I_2775 (I49561,I49527,I49544);
DFFARX1 I_2776  ( .D(I49561), .CLK(I2350), .RSTB(I49216), .Q(I49184) );
DFFARX1 I_2777  ( .D(I49527), .CLK(I2350), .RSTB(I49216), .Q(I49592) );
and I_2778 (I49181,I49360,I49592);
DFFARX1 I_2779  ( .D(I89349), .CLK(I2350), .RSTB(I49216), .Q(I49623) );
not I_2780 (I49640,I49623);
nor I_2781 (I49657,I49315,I49640);
and I_2782 (I49674,I49623,I49657);
nand I_2783 (I49196,I49623,I49377);
DFFARX1 I_2784  ( .D(I49623), .CLK(I2350), .RSTB(I49216), .Q(I49705) );
not I_2785 (I49193,I49705);
DFFARX1 I_2786  ( .D(I89376), .CLK(I2350), .RSTB(I49216), .Q(I49736) );
not I_2787 (I49753,I49736);
or I_2788 (I49770,I49753,I49674);
DFFARX1 I_2789  ( .D(I49770), .CLK(I2350), .RSTB(I49216), .Q(I49199) );
nand I_2790 (I49208,I49753,I49479);
DFFARX1 I_2791  ( .D(I49753), .CLK(I2350), .RSTB(I49216), .Q(I49178) );
not I_2792 (I49862,I2357);
not I_2793 (I49879,I247566);
nor I_2794 (I49896,I247554,I247560);
nand I_2795 (I49913,I49896,I247551);
DFFARX1 I_2796  ( .D(I49913), .CLK(I2350), .RSTB(I49862), .Q(I49836) );
nor I_2797 (I49944,I49879,I247554);
nand I_2798 (I49961,I49944,I247557);
not I_2799 (I49851,I49961);
DFFARX1 I_2800  ( .D(I49961), .CLK(I2350), .RSTB(I49862), .Q(I49833) );
not I_2801 (I50006,I247554);
not I_2802 (I50023,I50006);
not I_2803 (I50040,I247569);
nor I_2804 (I50057,I50040,I247581);
and I_2805 (I50074,I50057,I247563);
or I_2806 (I50091,I50074,I247578);
DFFARX1 I_2807  ( .D(I50091), .CLK(I2350), .RSTB(I49862), .Q(I50108) );
nor I_2808 (I50125,I50108,I49961);
nor I_2809 (I50142,I50108,I50023);
nand I_2810 (I49848,I49913,I50142);
nand I_2811 (I50173,I49879,I247569);
nand I_2812 (I50190,I50173,I50108);
and I_2813 (I50207,I50173,I50190);
DFFARX1 I_2814  ( .D(I50207), .CLK(I2350), .RSTB(I49862), .Q(I49830) );
DFFARX1 I_2815  ( .D(I50173), .CLK(I2350), .RSTB(I49862), .Q(I50238) );
and I_2816 (I49827,I50006,I50238);
DFFARX1 I_2817  ( .D(I247572), .CLK(I2350), .RSTB(I49862), .Q(I50269) );
not I_2818 (I50286,I50269);
nor I_2819 (I50303,I49961,I50286);
and I_2820 (I50320,I50269,I50303);
nand I_2821 (I49842,I50269,I50023);
DFFARX1 I_2822  ( .D(I50269), .CLK(I2350), .RSTB(I49862), .Q(I50351) );
not I_2823 (I49839,I50351);
DFFARX1 I_2824  ( .D(I247575), .CLK(I2350), .RSTB(I49862), .Q(I50382) );
not I_2825 (I50399,I50382);
or I_2826 (I50416,I50399,I50320);
DFFARX1 I_2827  ( .D(I50416), .CLK(I2350), .RSTB(I49862), .Q(I49845) );
nand I_2828 (I49854,I50399,I50125);
DFFARX1 I_2829  ( .D(I50399), .CLK(I2350), .RSTB(I49862), .Q(I49824) );
not I_2830 (I50508,I2357);
not I_2831 (I50525,I244098);
nor I_2832 (I50542,I244086,I244092);
nand I_2833 (I50559,I50542,I244083);
DFFARX1 I_2834  ( .D(I50559), .CLK(I2350), .RSTB(I50508), .Q(I50482) );
nor I_2835 (I50590,I50525,I244086);
nand I_2836 (I50607,I50590,I244089);
not I_2837 (I50497,I50607);
DFFARX1 I_2838  ( .D(I50607), .CLK(I2350), .RSTB(I50508), .Q(I50479) );
not I_2839 (I50652,I244086);
not I_2840 (I50669,I50652);
not I_2841 (I50686,I244101);
nor I_2842 (I50703,I50686,I244113);
and I_2843 (I50720,I50703,I244095);
or I_2844 (I50737,I50720,I244110);
DFFARX1 I_2845  ( .D(I50737), .CLK(I2350), .RSTB(I50508), .Q(I50754) );
nor I_2846 (I50771,I50754,I50607);
nor I_2847 (I50788,I50754,I50669);
nand I_2848 (I50494,I50559,I50788);
nand I_2849 (I50819,I50525,I244101);
nand I_2850 (I50836,I50819,I50754);
and I_2851 (I50853,I50819,I50836);
DFFARX1 I_2852  ( .D(I50853), .CLK(I2350), .RSTB(I50508), .Q(I50476) );
DFFARX1 I_2853  ( .D(I50819), .CLK(I2350), .RSTB(I50508), .Q(I50884) );
and I_2854 (I50473,I50652,I50884);
DFFARX1 I_2855  ( .D(I244104), .CLK(I2350), .RSTB(I50508), .Q(I50915) );
not I_2856 (I50932,I50915);
nor I_2857 (I50949,I50607,I50932);
and I_2858 (I50966,I50915,I50949);
nand I_2859 (I50488,I50915,I50669);
DFFARX1 I_2860  ( .D(I50915), .CLK(I2350), .RSTB(I50508), .Q(I50997) );
not I_2861 (I50485,I50997);
DFFARX1 I_2862  ( .D(I244107), .CLK(I2350), .RSTB(I50508), .Q(I51028) );
not I_2863 (I51045,I51028);
or I_2864 (I51062,I51045,I50966);
DFFARX1 I_2865  ( .D(I51062), .CLK(I2350), .RSTB(I50508), .Q(I50491) );
nand I_2866 (I50500,I51045,I50771);
DFFARX1 I_2867  ( .D(I51045), .CLK(I2350), .RSTB(I50508), .Q(I50470) );
not I_2868 (I51154,I2357);
not I_2869 (I51171,I396072);
nor I_2870 (I51188,I396069,I396066);
nand I_2871 (I51205,I51188,I396087);
DFFARX1 I_2872  ( .D(I51205), .CLK(I2350), .RSTB(I51154), .Q(I51128) );
nor I_2873 (I51236,I51171,I396069);
nand I_2874 (I51253,I51236,I396090);
not I_2875 (I51143,I51253);
DFFARX1 I_2876  ( .D(I51253), .CLK(I2350), .RSTB(I51154), .Q(I51125) );
not I_2877 (I51298,I396069);
not I_2878 (I51315,I51298);
not I_2879 (I51332,I396063);
nor I_2880 (I51349,I51332,I396075);
and I_2881 (I51366,I51349,I396084);
or I_2882 (I51383,I51366,I396078);
DFFARX1 I_2883  ( .D(I51383), .CLK(I2350), .RSTB(I51154), .Q(I51400) );
nor I_2884 (I51417,I51400,I51253);
nor I_2885 (I51434,I51400,I51315);
nand I_2886 (I51140,I51205,I51434);
nand I_2887 (I51465,I51171,I396063);
nand I_2888 (I51482,I51465,I51400);
and I_2889 (I51499,I51465,I51482);
DFFARX1 I_2890  ( .D(I51499), .CLK(I2350), .RSTB(I51154), .Q(I51122) );
DFFARX1 I_2891  ( .D(I51465), .CLK(I2350), .RSTB(I51154), .Q(I51530) );
and I_2892 (I51119,I51298,I51530);
DFFARX1 I_2893  ( .D(I396093), .CLK(I2350), .RSTB(I51154), .Q(I51561) );
not I_2894 (I51578,I51561);
nor I_2895 (I51595,I51253,I51578);
and I_2896 (I51612,I51561,I51595);
nand I_2897 (I51134,I51561,I51315);
DFFARX1 I_2898  ( .D(I51561), .CLK(I2350), .RSTB(I51154), .Q(I51643) );
not I_2899 (I51131,I51643);
DFFARX1 I_2900  ( .D(I396081), .CLK(I2350), .RSTB(I51154), .Q(I51674) );
not I_2901 (I51691,I51674);
or I_2902 (I51708,I51691,I51612);
DFFARX1 I_2903  ( .D(I51708), .CLK(I2350), .RSTB(I51154), .Q(I51137) );
nand I_2904 (I51146,I51691,I51417);
DFFARX1 I_2905  ( .D(I51691), .CLK(I2350), .RSTB(I51154), .Q(I51116) );
not I_2906 (I51800,I2357);
not I_2907 (I51817,I144991);
nor I_2908 (I51834,I144988,I144976);
nand I_2909 (I51851,I51834,I144979);
DFFARX1 I_2910  ( .D(I51851), .CLK(I2350), .RSTB(I51800), .Q(I51774) );
nor I_2911 (I51882,I51817,I144988);
nand I_2912 (I51899,I51882,I144985);
not I_2913 (I51789,I51899);
DFFARX1 I_2914  ( .D(I51899), .CLK(I2350), .RSTB(I51800), .Q(I51771) );
not I_2915 (I51944,I144988);
not I_2916 (I51961,I51944);
not I_2917 (I51978,I144997);
nor I_2918 (I51995,I51978,I144973);
and I_2919 (I52012,I51995,I144994);
or I_2920 (I52029,I52012,I144982);
DFFARX1 I_2921  ( .D(I52029), .CLK(I2350), .RSTB(I51800), .Q(I52046) );
nor I_2922 (I52063,I52046,I51899);
nor I_2923 (I52080,I52046,I51961);
nand I_2924 (I51786,I51851,I52080);
nand I_2925 (I52111,I51817,I144997);
nand I_2926 (I52128,I52111,I52046);
and I_2927 (I52145,I52111,I52128);
DFFARX1 I_2928  ( .D(I52145), .CLK(I2350), .RSTB(I51800), .Q(I51768) );
DFFARX1 I_2929  ( .D(I52111), .CLK(I2350), .RSTB(I51800), .Q(I52176) );
and I_2930 (I51765,I51944,I52176);
DFFARX1 I_2931  ( .D(I145003), .CLK(I2350), .RSTB(I51800), .Q(I52207) );
not I_2932 (I52224,I52207);
nor I_2933 (I52241,I51899,I52224);
and I_2934 (I52258,I52207,I52241);
nand I_2935 (I51780,I52207,I51961);
DFFARX1 I_2936  ( .D(I52207), .CLK(I2350), .RSTB(I51800), .Q(I52289) );
not I_2937 (I51777,I52289);
DFFARX1 I_2938  ( .D(I145000), .CLK(I2350), .RSTB(I51800), .Q(I52320) );
not I_2939 (I52337,I52320);
or I_2940 (I52354,I52337,I52258);
DFFARX1 I_2941  ( .D(I52354), .CLK(I2350), .RSTB(I51800), .Q(I51783) );
nand I_2942 (I51792,I52337,I52063);
DFFARX1 I_2943  ( .D(I52337), .CLK(I2350), .RSTB(I51800), .Q(I51762) );
not I_2944 (I52446,I2357);
not I_2945 (I52463,I248722);
nor I_2946 (I52480,I248710,I248716);
nand I_2947 (I52497,I52480,I248707);
DFFARX1 I_2948  ( .D(I52497), .CLK(I2350), .RSTB(I52446), .Q(I52420) );
nor I_2949 (I52528,I52463,I248710);
nand I_2950 (I52545,I52528,I248713);
not I_2951 (I52435,I52545);
DFFARX1 I_2952  ( .D(I52545), .CLK(I2350), .RSTB(I52446), .Q(I52417) );
not I_2953 (I52590,I248710);
not I_2954 (I52607,I52590);
not I_2955 (I52624,I248725);
nor I_2956 (I52641,I52624,I248737);
and I_2957 (I52658,I52641,I248719);
or I_2958 (I52675,I52658,I248734);
DFFARX1 I_2959  ( .D(I52675), .CLK(I2350), .RSTB(I52446), .Q(I52692) );
nor I_2960 (I52709,I52692,I52545);
nor I_2961 (I52726,I52692,I52607);
nand I_2962 (I52432,I52497,I52726);
nand I_2963 (I52757,I52463,I248725);
nand I_2964 (I52774,I52757,I52692);
and I_2965 (I52791,I52757,I52774);
DFFARX1 I_2966  ( .D(I52791), .CLK(I2350), .RSTB(I52446), .Q(I52414) );
DFFARX1 I_2967  ( .D(I52757), .CLK(I2350), .RSTB(I52446), .Q(I52822) );
and I_2968 (I52411,I52590,I52822);
DFFARX1 I_2969  ( .D(I248728), .CLK(I2350), .RSTB(I52446), .Q(I52853) );
not I_2970 (I52870,I52853);
nor I_2971 (I52887,I52545,I52870);
and I_2972 (I52904,I52853,I52887);
nand I_2973 (I52426,I52853,I52607);
DFFARX1 I_2974  ( .D(I52853), .CLK(I2350), .RSTB(I52446), .Q(I52935) );
not I_2975 (I52423,I52935);
DFFARX1 I_2976  ( .D(I248731), .CLK(I2350), .RSTB(I52446), .Q(I52966) );
not I_2977 (I52983,I52966);
or I_2978 (I53000,I52983,I52904);
DFFARX1 I_2979  ( .D(I53000), .CLK(I2350), .RSTB(I52446), .Q(I52429) );
nand I_2980 (I52438,I52983,I52709);
DFFARX1 I_2981  ( .D(I52983), .CLK(I2350), .RSTB(I52446), .Q(I52408) );
not I_2982 (I53092,I2357);
not I_2983 (I53109,I271539);
nor I_2984 (I53126,I271551,I271533);
nand I_2985 (I53143,I53126,I271542);
DFFARX1 I_2986  ( .D(I53143), .CLK(I2350), .RSTB(I53092), .Q(I53066) );
nor I_2987 (I53174,I53109,I271551);
nand I_2988 (I53191,I53174,I271548);
not I_2989 (I53081,I53191);
DFFARX1 I_2990  ( .D(I53191), .CLK(I2350), .RSTB(I53092), .Q(I53063) );
not I_2991 (I53236,I271551);
not I_2992 (I53253,I53236);
not I_2993 (I53270,I271521);
nor I_2994 (I53287,I53270,I271524);
and I_2995 (I53304,I53287,I271530);
or I_2996 (I53321,I53304,I271545);
DFFARX1 I_2997  ( .D(I53321), .CLK(I2350), .RSTB(I53092), .Q(I53338) );
nor I_2998 (I53355,I53338,I53191);
nor I_2999 (I53372,I53338,I53253);
nand I_3000 (I53078,I53143,I53372);
nand I_3001 (I53403,I53109,I271521);
nand I_3002 (I53420,I53403,I53338);
and I_3003 (I53437,I53403,I53420);
DFFARX1 I_3004  ( .D(I53437), .CLK(I2350), .RSTB(I53092), .Q(I53060) );
DFFARX1 I_3005  ( .D(I53403), .CLK(I2350), .RSTB(I53092), .Q(I53468) );
and I_3006 (I53057,I53236,I53468);
DFFARX1 I_3007  ( .D(I271527), .CLK(I2350), .RSTB(I53092), .Q(I53499) );
not I_3008 (I53516,I53499);
nor I_3009 (I53533,I53191,I53516);
and I_3010 (I53550,I53499,I53533);
nand I_3011 (I53072,I53499,I53253);
DFFARX1 I_3012  ( .D(I53499), .CLK(I2350), .RSTB(I53092), .Q(I53581) );
not I_3013 (I53069,I53581);
DFFARX1 I_3014  ( .D(I271536), .CLK(I2350), .RSTB(I53092), .Q(I53612) );
not I_3015 (I53629,I53612);
or I_3016 (I53646,I53629,I53550);
DFFARX1 I_3017  ( .D(I53646), .CLK(I2350), .RSTB(I53092), .Q(I53075) );
nand I_3018 (I53084,I53629,I53355);
DFFARX1 I_3019  ( .D(I53629), .CLK(I2350), .RSTB(I53092), .Q(I53054) );
not I_3020 (I53738,I2357);
not I_3021 (I53755,I240630);
nor I_3022 (I53772,I240618,I240624);
nand I_3023 (I53789,I53772,I240615);
DFFARX1 I_3024  ( .D(I53789), .CLK(I2350), .RSTB(I53738), .Q(I53712) );
nor I_3025 (I53820,I53755,I240618);
nand I_3026 (I53837,I53820,I240621);
not I_3027 (I53727,I53837);
DFFARX1 I_3028  ( .D(I53837), .CLK(I2350), .RSTB(I53738), .Q(I53709) );
not I_3029 (I53882,I240618);
not I_3030 (I53899,I53882);
not I_3031 (I53916,I240633);
nor I_3032 (I53933,I53916,I240645);
and I_3033 (I53950,I53933,I240627);
or I_3034 (I53967,I53950,I240642);
DFFARX1 I_3035  ( .D(I53967), .CLK(I2350), .RSTB(I53738), .Q(I53984) );
nor I_3036 (I54001,I53984,I53837);
nor I_3037 (I54018,I53984,I53899);
nand I_3038 (I53724,I53789,I54018);
nand I_3039 (I54049,I53755,I240633);
nand I_3040 (I54066,I54049,I53984);
and I_3041 (I54083,I54049,I54066);
DFFARX1 I_3042  ( .D(I54083), .CLK(I2350), .RSTB(I53738), .Q(I53706) );
DFFARX1 I_3043  ( .D(I54049), .CLK(I2350), .RSTB(I53738), .Q(I54114) );
and I_3044 (I53703,I53882,I54114);
DFFARX1 I_3045  ( .D(I240636), .CLK(I2350), .RSTB(I53738), .Q(I54145) );
not I_3046 (I54162,I54145);
nor I_3047 (I54179,I53837,I54162);
and I_3048 (I54196,I54145,I54179);
nand I_3049 (I53718,I54145,I53899);
DFFARX1 I_3050  ( .D(I54145), .CLK(I2350), .RSTB(I53738), .Q(I54227) );
not I_3051 (I53715,I54227);
DFFARX1 I_3052  ( .D(I240639), .CLK(I2350), .RSTB(I53738), .Q(I54258) );
not I_3053 (I54275,I54258);
or I_3054 (I54292,I54275,I54196);
DFFARX1 I_3055  ( .D(I54292), .CLK(I2350), .RSTB(I53738), .Q(I53721) );
nand I_3056 (I53730,I54275,I54001);
DFFARX1 I_3057  ( .D(I54275), .CLK(I2350), .RSTB(I53738), .Q(I53700) );
not I_3058 (I54384,I2357);
not I_3059 (I54401,I21437);
nor I_3060 (I54418,I21449,I21434);
nand I_3061 (I54435,I54418,I21446);
DFFARX1 I_3062  ( .D(I54435), .CLK(I2350), .RSTB(I54384), .Q(I54358) );
nor I_3063 (I54466,I54401,I21449);
nand I_3064 (I54483,I54466,I21464);
not I_3065 (I54373,I54483);
DFFARX1 I_3066  ( .D(I54483), .CLK(I2350), .RSTB(I54384), .Q(I54355) );
not I_3067 (I54528,I21449);
not I_3068 (I54545,I54528);
not I_3069 (I54562,I21440);
nor I_3070 (I54579,I54562,I21452);
and I_3071 (I54596,I54579,I21443);
or I_3072 (I54613,I54596,I21458);
DFFARX1 I_3073  ( .D(I54613), .CLK(I2350), .RSTB(I54384), .Q(I54630) );
nor I_3074 (I54647,I54630,I54483);
nor I_3075 (I54664,I54630,I54545);
nand I_3076 (I54370,I54435,I54664);
nand I_3077 (I54695,I54401,I21440);
nand I_3078 (I54712,I54695,I54630);
and I_3079 (I54729,I54695,I54712);
DFFARX1 I_3080  ( .D(I54729), .CLK(I2350), .RSTB(I54384), .Q(I54352) );
DFFARX1 I_3081  ( .D(I54695), .CLK(I2350), .RSTB(I54384), .Q(I54760) );
and I_3082 (I54349,I54528,I54760);
DFFARX1 I_3083  ( .D(I21461), .CLK(I2350), .RSTB(I54384), .Q(I54791) );
not I_3084 (I54808,I54791);
nor I_3085 (I54825,I54483,I54808);
and I_3086 (I54842,I54791,I54825);
nand I_3087 (I54364,I54791,I54545);
DFFARX1 I_3088  ( .D(I54791), .CLK(I2350), .RSTB(I54384), .Q(I54873) );
not I_3089 (I54361,I54873);
DFFARX1 I_3090  ( .D(I21455), .CLK(I2350), .RSTB(I54384), .Q(I54904) );
not I_3091 (I54921,I54904);
or I_3092 (I54938,I54921,I54842);
DFFARX1 I_3093  ( .D(I54938), .CLK(I2350), .RSTB(I54384), .Q(I54367) );
nand I_3094 (I54376,I54921,I54647);
DFFARX1 I_3095  ( .D(I54921), .CLK(I2350), .RSTB(I54384), .Q(I54346) );
not I_3096 (I55030,I2357);
not I_3097 (I55047,I252768);
nor I_3098 (I55064,I252756,I252762);
nand I_3099 (I55081,I55064,I252753);
DFFARX1 I_3100  ( .D(I55081), .CLK(I2350), .RSTB(I55030), .Q(I55004) );
nor I_3101 (I55112,I55047,I252756);
nand I_3102 (I55129,I55112,I252759);
not I_3103 (I55019,I55129);
DFFARX1 I_3104  ( .D(I55129), .CLK(I2350), .RSTB(I55030), .Q(I55001) );
not I_3105 (I55174,I252756);
not I_3106 (I55191,I55174);
not I_3107 (I55208,I252771);
nor I_3108 (I55225,I55208,I252783);
and I_3109 (I55242,I55225,I252765);
or I_3110 (I55259,I55242,I252780);
DFFARX1 I_3111  ( .D(I55259), .CLK(I2350), .RSTB(I55030), .Q(I55276) );
nor I_3112 (I55293,I55276,I55129);
nor I_3113 (I55310,I55276,I55191);
nand I_3114 (I55016,I55081,I55310);
nand I_3115 (I55341,I55047,I252771);
nand I_3116 (I55358,I55341,I55276);
and I_3117 (I55375,I55341,I55358);
DFFARX1 I_3118  ( .D(I55375), .CLK(I2350), .RSTB(I55030), .Q(I54998) );
DFFARX1 I_3119  ( .D(I55341), .CLK(I2350), .RSTB(I55030), .Q(I55406) );
and I_3120 (I54995,I55174,I55406);
DFFARX1 I_3121  ( .D(I252774), .CLK(I2350), .RSTB(I55030), .Q(I55437) );
not I_3122 (I55454,I55437);
nor I_3123 (I55471,I55129,I55454);
and I_3124 (I55488,I55437,I55471);
nand I_3125 (I55010,I55437,I55191);
DFFARX1 I_3126  ( .D(I55437), .CLK(I2350), .RSTB(I55030), .Q(I55519) );
not I_3127 (I55007,I55519);
DFFARX1 I_3128  ( .D(I252777), .CLK(I2350), .RSTB(I55030), .Q(I55550) );
not I_3129 (I55567,I55550);
or I_3130 (I55584,I55567,I55488);
DFFARX1 I_3131  ( .D(I55584), .CLK(I2350), .RSTB(I55030), .Q(I55013) );
nand I_3132 (I55022,I55567,I55293);
DFFARX1 I_3133  ( .D(I55567), .CLK(I2350), .RSTB(I55030), .Q(I54992) );
not I_3134 (I55676,I2357);
not I_3135 (I55693,I340150);
nor I_3136 (I55710,I340165,I340180);
nand I_3137 (I55727,I55710,I340168);
DFFARX1 I_3138  ( .D(I55727), .CLK(I2350), .RSTB(I55676), .Q(I55650) );
nor I_3139 (I55758,I55693,I340165);
nand I_3140 (I55775,I55758,I340171);
not I_3141 (I55665,I55775);
DFFARX1 I_3142  ( .D(I55775), .CLK(I2350), .RSTB(I55676), .Q(I55647) );
not I_3143 (I55820,I340165);
not I_3144 (I55837,I55820);
not I_3145 (I55854,I340177);
nor I_3146 (I55871,I55854,I340174);
and I_3147 (I55888,I55871,I340153);
or I_3148 (I55905,I55888,I340162);
DFFARX1 I_3149  ( .D(I55905), .CLK(I2350), .RSTB(I55676), .Q(I55922) );
nor I_3150 (I55939,I55922,I55775);
nor I_3151 (I55956,I55922,I55837);
nand I_3152 (I55662,I55727,I55956);
nand I_3153 (I55987,I55693,I340177);
nand I_3154 (I56004,I55987,I55922);
and I_3155 (I56021,I55987,I56004);
DFFARX1 I_3156  ( .D(I56021), .CLK(I2350), .RSTB(I55676), .Q(I55644) );
DFFARX1 I_3157  ( .D(I55987), .CLK(I2350), .RSTB(I55676), .Q(I56052) );
and I_3158 (I55641,I55820,I56052);
DFFARX1 I_3159  ( .D(I340159), .CLK(I2350), .RSTB(I55676), .Q(I56083) );
not I_3160 (I56100,I56083);
nor I_3161 (I56117,I55775,I56100);
and I_3162 (I56134,I56083,I56117);
nand I_3163 (I55656,I56083,I55837);
DFFARX1 I_3164  ( .D(I56083), .CLK(I2350), .RSTB(I55676), .Q(I56165) );
not I_3165 (I55653,I56165);
DFFARX1 I_3166  ( .D(I340156), .CLK(I2350), .RSTB(I55676), .Q(I56196) );
not I_3167 (I56213,I56196);
or I_3168 (I56230,I56213,I56134);
DFFARX1 I_3169  ( .D(I56230), .CLK(I2350), .RSTB(I55676), .Q(I55659) );
nand I_3170 (I55668,I56213,I55939);
DFFARX1 I_3171  ( .D(I56213), .CLK(I2350), .RSTB(I55676), .Q(I55638) );
not I_3172 (I56322,I2357);
not I_3173 (I56339,I267261);
nor I_3174 (I56356,I267243,I267252);
nand I_3175 (I56373,I56356,I267264);
DFFARX1 I_3176  ( .D(I56373), .CLK(I2350), .RSTB(I56322), .Q(I56296) );
nor I_3177 (I56404,I56339,I267243);
nand I_3178 (I56421,I56404,I267249);
not I_3179 (I56311,I56421);
DFFARX1 I_3180  ( .D(I56421), .CLK(I2350), .RSTB(I56322), .Q(I56293) );
not I_3181 (I56466,I267243);
not I_3182 (I56483,I56466);
not I_3183 (I56500,I267240);
nor I_3184 (I56517,I56500,I267258);
and I_3185 (I56534,I56517,I267246);
or I_3186 (I56551,I56534,I267267);
DFFARX1 I_3187  ( .D(I56551), .CLK(I2350), .RSTB(I56322), .Q(I56568) );
nor I_3188 (I56585,I56568,I56421);
nor I_3189 (I56602,I56568,I56483);
nand I_3190 (I56308,I56373,I56602);
nand I_3191 (I56633,I56339,I267240);
nand I_3192 (I56650,I56633,I56568);
and I_3193 (I56667,I56633,I56650);
DFFARX1 I_3194  ( .D(I56667), .CLK(I2350), .RSTB(I56322), .Q(I56290) );
DFFARX1 I_3195  ( .D(I56633), .CLK(I2350), .RSTB(I56322), .Q(I56698) );
and I_3196 (I56287,I56466,I56698);
DFFARX1 I_3197  ( .D(I267255), .CLK(I2350), .RSTB(I56322), .Q(I56729) );
not I_3198 (I56746,I56729);
nor I_3199 (I56763,I56421,I56746);
and I_3200 (I56780,I56729,I56763);
nand I_3201 (I56302,I56729,I56483);
DFFARX1 I_3202  ( .D(I56729), .CLK(I2350), .RSTB(I56322), .Q(I56811) );
not I_3203 (I56299,I56811);
DFFARX1 I_3204  ( .D(I267237), .CLK(I2350), .RSTB(I56322), .Q(I56842) );
not I_3205 (I56859,I56842);
or I_3206 (I56876,I56859,I56780);
DFFARX1 I_3207  ( .D(I56876), .CLK(I2350), .RSTB(I56322), .Q(I56305) );
nand I_3208 (I56314,I56859,I56585);
DFFARX1 I_3209  ( .D(I56859), .CLK(I2350), .RSTB(I56322), .Q(I56284) );
not I_3210 (I56968,I2357);
not I_3211 (I56985,I103290);
nor I_3212 (I57002,I103278,I103284);
nand I_3213 (I57019,I57002,I103293);
DFFARX1 I_3214  ( .D(I57019), .CLK(I2350), .RSTB(I56968), .Q(I56942) );
nor I_3215 (I57050,I56985,I103278);
nand I_3216 (I57067,I57050,I103281);
not I_3217 (I56957,I57067);
DFFARX1 I_3218  ( .D(I57067), .CLK(I2350), .RSTB(I56968), .Q(I56939) );
not I_3219 (I57112,I103278);
not I_3220 (I57129,I57112);
not I_3221 (I57146,I103302);
nor I_3222 (I57163,I57146,I103275);
and I_3223 (I57180,I57163,I103296);
or I_3224 (I57197,I57180,I103287);
DFFARX1 I_3225  ( .D(I57197), .CLK(I2350), .RSTB(I56968), .Q(I57214) );
nor I_3226 (I57231,I57214,I57067);
nor I_3227 (I57248,I57214,I57129);
nand I_3228 (I56954,I57019,I57248);
nand I_3229 (I57279,I56985,I103302);
nand I_3230 (I57296,I57279,I57214);
and I_3231 (I57313,I57279,I57296);
DFFARX1 I_3232  ( .D(I57313), .CLK(I2350), .RSTB(I56968), .Q(I56936) );
DFFARX1 I_3233  ( .D(I57279), .CLK(I2350), .RSTB(I56968), .Q(I57344) );
and I_3234 (I56933,I57112,I57344);
DFFARX1 I_3235  ( .D(I103272), .CLK(I2350), .RSTB(I56968), .Q(I57375) );
not I_3236 (I57392,I57375);
nor I_3237 (I57409,I57067,I57392);
and I_3238 (I57426,I57375,I57409);
nand I_3239 (I56948,I57375,I57129);
DFFARX1 I_3240  ( .D(I57375), .CLK(I2350), .RSTB(I56968), .Q(I57457) );
not I_3241 (I56945,I57457);
DFFARX1 I_3242  ( .D(I103299), .CLK(I2350), .RSTB(I56968), .Q(I57488) );
not I_3243 (I57505,I57488);
or I_3244 (I57522,I57505,I57426);
DFFARX1 I_3245  ( .D(I57522), .CLK(I2350), .RSTB(I56968), .Q(I56951) );
nand I_3246 (I56960,I57505,I57231);
DFFARX1 I_3247  ( .D(I57505), .CLK(I2350), .RSTB(I56968), .Q(I56930) );
not I_3248 (I57614,I2357);
not I_3249 (I57631,I329047);
nor I_3250 (I57648,I329032,I329059);
nand I_3251 (I57665,I57648,I329035);
DFFARX1 I_3252  ( .D(I57665), .CLK(I2350), .RSTB(I57614), .Q(I57588) );
nor I_3253 (I57696,I57631,I329032);
nand I_3254 (I57713,I57696,I329050);
not I_3255 (I57603,I57713);
DFFARX1 I_3256  ( .D(I57713), .CLK(I2350), .RSTB(I57614), .Q(I57585) );
not I_3257 (I57758,I329032);
not I_3258 (I57775,I57758);
not I_3259 (I57792,I329062);
nor I_3260 (I57809,I57792,I329044);
and I_3261 (I57826,I57809,I329053);
or I_3262 (I57843,I57826,I329038);
DFFARX1 I_3263  ( .D(I57843), .CLK(I2350), .RSTB(I57614), .Q(I57860) );
nor I_3264 (I57877,I57860,I57713);
nor I_3265 (I57894,I57860,I57775);
nand I_3266 (I57600,I57665,I57894);
nand I_3267 (I57925,I57631,I329062);
nand I_3268 (I57942,I57925,I57860);
and I_3269 (I57959,I57925,I57942);
DFFARX1 I_3270  ( .D(I57959), .CLK(I2350), .RSTB(I57614), .Q(I57582) );
DFFARX1 I_3271  ( .D(I57925), .CLK(I2350), .RSTB(I57614), .Q(I57990) );
and I_3272 (I57579,I57758,I57990);
DFFARX1 I_3273  ( .D(I329041), .CLK(I2350), .RSTB(I57614), .Q(I58021) );
not I_3274 (I58038,I58021);
nor I_3275 (I58055,I57713,I58038);
and I_3276 (I58072,I58021,I58055);
nand I_3277 (I57594,I58021,I57775);
DFFARX1 I_3278  ( .D(I58021), .CLK(I2350), .RSTB(I57614), .Q(I58103) );
not I_3279 (I57591,I58103);
DFFARX1 I_3280  ( .D(I329056), .CLK(I2350), .RSTB(I57614), .Q(I58134) );
not I_3281 (I58151,I58134);
or I_3282 (I58168,I58151,I58072);
DFFARX1 I_3283  ( .D(I58168), .CLK(I2350), .RSTB(I57614), .Q(I57597) );
nand I_3284 (I57606,I58151,I57877);
DFFARX1 I_3285  ( .D(I58151), .CLK(I2350), .RSTB(I57614), .Q(I57576) );
not I_3286 (I58260,I2357);
not I_3287 (I58277,I99312);
nor I_3288 (I58294,I99300,I99306);
nand I_3289 (I58311,I58294,I99315);
DFFARX1 I_3290  ( .D(I58311), .CLK(I2350), .RSTB(I58260), .Q(I58234) );
nor I_3291 (I58342,I58277,I99300);
nand I_3292 (I58359,I58342,I99303);
not I_3293 (I58249,I58359);
DFFARX1 I_3294  ( .D(I58359), .CLK(I2350), .RSTB(I58260), .Q(I58231) );
not I_3295 (I58404,I99300);
not I_3296 (I58421,I58404);
not I_3297 (I58438,I99324);
nor I_3298 (I58455,I58438,I99297);
and I_3299 (I58472,I58455,I99318);
or I_3300 (I58489,I58472,I99309);
DFFARX1 I_3301  ( .D(I58489), .CLK(I2350), .RSTB(I58260), .Q(I58506) );
nor I_3302 (I58523,I58506,I58359);
nor I_3303 (I58540,I58506,I58421);
nand I_3304 (I58246,I58311,I58540);
nand I_3305 (I58571,I58277,I99324);
nand I_3306 (I58588,I58571,I58506);
and I_3307 (I58605,I58571,I58588);
DFFARX1 I_3308  ( .D(I58605), .CLK(I2350), .RSTB(I58260), .Q(I58228) );
DFFARX1 I_3309  ( .D(I58571), .CLK(I2350), .RSTB(I58260), .Q(I58636) );
and I_3310 (I58225,I58404,I58636);
DFFARX1 I_3311  ( .D(I99294), .CLK(I2350), .RSTB(I58260), .Q(I58667) );
not I_3312 (I58684,I58667);
nor I_3313 (I58701,I58359,I58684);
and I_3314 (I58718,I58667,I58701);
nand I_3315 (I58240,I58667,I58421);
DFFARX1 I_3316  ( .D(I58667), .CLK(I2350), .RSTB(I58260), .Q(I58749) );
not I_3317 (I58237,I58749);
DFFARX1 I_3318  ( .D(I99321), .CLK(I2350), .RSTB(I58260), .Q(I58780) );
not I_3319 (I58797,I58780);
or I_3320 (I58814,I58797,I58718);
DFFARX1 I_3321  ( .D(I58814), .CLK(I2350), .RSTB(I58260), .Q(I58243) );
nand I_3322 (I58252,I58797,I58523);
DFFARX1 I_3323  ( .D(I58797), .CLK(I2350), .RSTB(I58260), .Q(I58222) );
not I_3324 (I58906,I2357);
not I_3325 (I58923,I370971);
nor I_3326 (I58940,I370986,I371001);
nand I_3327 (I58957,I58940,I370989);
DFFARX1 I_3328  ( .D(I58957), .CLK(I2350), .RSTB(I58906), .Q(I58880) );
nor I_3329 (I58988,I58923,I370986);
nand I_3330 (I59005,I58988,I370992);
not I_3331 (I58895,I59005);
DFFARX1 I_3332  ( .D(I59005), .CLK(I2350), .RSTB(I58906), .Q(I58877) );
not I_3333 (I59050,I370986);
not I_3334 (I59067,I59050);
not I_3335 (I59084,I370998);
nor I_3336 (I59101,I59084,I370995);
and I_3337 (I59118,I59101,I370974);
or I_3338 (I59135,I59118,I370983);
DFFARX1 I_3339  ( .D(I59135), .CLK(I2350), .RSTB(I58906), .Q(I59152) );
nor I_3340 (I59169,I59152,I59005);
nor I_3341 (I59186,I59152,I59067);
nand I_3342 (I58892,I58957,I59186);
nand I_3343 (I59217,I58923,I370998);
nand I_3344 (I59234,I59217,I59152);
and I_3345 (I59251,I59217,I59234);
DFFARX1 I_3346  ( .D(I59251), .CLK(I2350), .RSTB(I58906), .Q(I58874) );
DFFARX1 I_3347  ( .D(I59217), .CLK(I2350), .RSTB(I58906), .Q(I59282) );
and I_3348 (I58871,I59050,I59282);
DFFARX1 I_3349  ( .D(I370980), .CLK(I2350), .RSTB(I58906), .Q(I59313) );
not I_3350 (I59330,I59313);
nor I_3351 (I59347,I59005,I59330);
and I_3352 (I59364,I59313,I59347);
nand I_3353 (I58886,I59313,I59067);
DFFARX1 I_3354  ( .D(I59313), .CLK(I2350), .RSTB(I58906), .Q(I59395) );
not I_3355 (I58883,I59395);
DFFARX1 I_3356  ( .D(I370977), .CLK(I2350), .RSTB(I58906), .Q(I59426) );
not I_3357 (I59443,I59426);
or I_3358 (I59460,I59443,I59364);
DFFARX1 I_3359  ( .D(I59460), .CLK(I2350), .RSTB(I58906), .Q(I58889) );
nand I_3360 (I58898,I59443,I59169);
DFFARX1 I_3361  ( .D(I59443), .CLK(I2350), .RSTB(I58906), .Q(I58868) );
not I_3362 (I59552,I2357);
not I_3363 (I59569,I387980);
nor I_3364 (I59586,I387977,I387974);
nand I_3365 (I59603,I59586,I387995);
DFFARX1 I_3366  ( .D(I59603), .CLK(I2350), .RSTB(I59552), .Q(I59526) );
nor I_3367 (I59634,I59569,I387977);
nand I_3368 (I59651,I59634,I387998);
not I_3369 (I59541,I59651);
DFFARX1 I_3370  ( .D(I59651), .CLK(I2350), .RSTB(I59552), .Q(I59523) );
not I_3371 (I59696,I387977);
not I_3372 (I59713,I59696);
not I_3373 (I59730,I387971);
nor I_3374 (I59747,I59730,I387983);
and I_3375 (I59764,I59747,I387992);
or I_3376 (I59781,I59764,I387986);
DFFARX1 I_3377  ( .D(I59781), .CLK(I2350), .RSTB(I59552), .Q(I59798) );
nor I_3378 (I59815,I59798,I59651);
nor I_3379 (I59832,I59798,I59713);
nand I_3380 (I59538,I59603,I59832);
nand I_3381 (I59863,I59569,I387971);
nand I_3382 (I59880,I59863,I59798);
and I_3383 (I59897,I59863,I59880);
DFFARX1 I_3384  ( .D(I59897), .CLK(I2350), .RSTB(I59552), .Q(I59520) );
DFFARX1 I_3385  ( .D(I59863), .CLK(I2350), .RSTB(I59552), .Q(I59928) );
and I_3386 (I59517,I59696,I59928);
DFFARX1 I_3387  ( .D(I388001), .CLK(I2350), .RSTB(I59552), .Q(I59959) );
not I_3388 (I59976,I59959);
nor I_3389 (I59993,I59651,I59976);
and I_3390 (I60010,I59959,I59993);
nand I_3391 (I59532,I59959,I59713);
DFFARX1 I_3392  ( .D(I59959), .CLK(I2350), .RSTB(I59552), .Q(I60041) );
not I_3393 (I59529,I60041);
DFFARX1 I_3394  ( .D(I387989), .CLK(I2350), .RSTB(I59552), .Q(I60072) );
not I_3395 (I60089,I60072);
or I_3396 (I60106,I60089,I60010);
DFFARX1 I_3397  ( .D(I60106), .CLK(I2350), .RSTB(I59552), .Q(I59535) );
nand I_3398 (I59544,I60089,I59815);
DFFARX1 I_3399  ( .D(I60089), .CLK(I2350), .RSTB(I59552), .Q(I59514) );
not I_3400 (I60198,I2357);
not I_3401 (I60215,I251612);
nor I_3402 (I60232,I251600,I251606);
nand I_3403 (I60249,I60232,I251597);
DFFARX1 I_3404  ( .D(I60249), .CLK(I2350), .RSTB(I60198), .Q(I60172) );
nor I_3405 (I60280,I60215,I251600);
nand I_3406 (I60297,I60280,I251603);
not I_3407 (I60187,I60297);
DFFARX1 I_3408  ( .D(I60297), .CLK(I2350), .RSTB(I60198), .Q(I60169) );
not I_3409 (I60342,I251600);
not I_3410 (I60359,I60342);
not I_3411 (I60376,I251615);
nor I_3412 (I60393,I60376,I251627);
and I_3413 (I60410,I60393,I251609);
or I_3414 (I60427,I60410,I251624);
DFFARX1 I_3415  ( .D(I60427), .CLK(I2350), .RSTB(I60198), .Q(I60444) );
nor I_3416 (I60461,I60444,I60297);
nor I_3417 (I60478,I60444,I60359);
nand I_3418 (I60184,I60249,I60478);
nand I_3419 (I60509,I60215,I251615);
nand I_3420 (I60526,I60509,I60444);
and I_3421 (I60543,I60509,I60526);
DFFARX1 I_3422  ( .D(I60543), .CLK(I2350), .RSTB(I60198), .Q(I60166) );
DFFARX1 I_3423  ( .D(I60509), .CLK(I2350), .RSTB(I60198), .Q(I60574) );
and I_3424 (I60163,I60342,I60574);
DFFARX1 I_3425  ( .D(I251618), .CLK(I2350), .RSTB(I60198), .Q(I60605) );
not I_3426 (I60622,I60605);
nor I_3427 (I60639,I60297,I60622);
and I_3428 (I60656,I60605,I60639);
nand I_3429 (I60178,I60605,I60359);
DFFARX1 I_3430  ( .D(I60605), .CLK(I2350), .RSTB(I60198), .Q(I60687) );
not I_3431 (I60175,I60687);
DFFARX1 I_3432  ( .D(I251621), .CLK(I2350), .RSTB(I60198), .Q(I60718) );
not I_3433 (I60735,I60718);
or I_3434 (I60752,I60735,I60656);
DFFARX1 I_3435  ( .D(I60752), .CLK(I2350), .RSTB(I60198), .Q(I60181) );
nand I_3436 (I60190,I60735,I60461);
DFFARX1 I_3437  ( .D(I60735), .CLK(I2350), .RSTB(I60198), .Q(I60160) );
not I_3438 (I60844,I2357);
not I_3439 (I60861,I2103);
nor I_3440 (I60878,I1295,I1543);
nand I_3441 (I60895,I60878,I1839);
DFFARX1 I_3442  ( .D(I60895), .CLK(I2350), .RSTB(I60844), .Q(I60818) );
nor I_3443 (I60926,I60861,I1295);
nand I_3444 (I60943,I60926,I1255);
not I_3445 (I60833,I60943);
DFFARX1 I_3446  ( .D(I60943), .CLK(I2350), .RSTB(I60844), .Q(I60815) );
not I_3447 (I60988,I1295);
not I_3448 (I61005,I60988);
not I_3449 (I61022,I2303);
nor I_3450 (I61039,I61022,I2031);
and I_3451 (I61056,I61039,I1815);
or I_3452 (I61073,I61056,I1911);
DFFARX1 I_3453  ( .D(I61073), .CLK(I2350), .RSTB(I60844), .Q(I61090) );
nor I_3454 (I61107,I61090,I60943);
nor I_3455 (I61124,I61090,I61005);
nand I_3456 (I60830,I60895,I61124);
nand I_3457 (I61155,I60861,I2303);
nand I_3458 (I61172,I61155,I61090);
and I_3459 (I61189,I61155,I61172);
DFFARX1 I_3460  ( .D(I61189), .CLK(I2350), .RSTB(I60844), .Q(I60812) );
DFFARX1 I_3461  ( .D(I61155), .CLK(I2350), .RSTB(I60844), .Q(I61220) );
and I_3462 (I60809,I60988,I61220);
DFFARX1 I_3463  ( .D(I1919), .CLK(I2350), .RSTB(I60844), .Q(I61251) );
not I_3464 (I61268,I61251);
nor I_3465 (I61285,I60943,I61268);
and I_3466 (I61302,I61251,I61285);
nand I_3467 (I60824,I61251,I61005);
DFFARX1 I_3468  ( .D(I61251), .CLK(I2350), .RSTB(I60844), .Q(I61333) );
not I_3469 (I60821,I61333);
DFFARX1 I_3470  ( .D(I1631), .CLK(I2350), .RSTB(I60844), .Q(I61364) );
not I_3471 (I61381,I61364);
or I_3472 (I61398,I61381,I61302);
DFFARX1 I_3473  ( .D(I61398), .CLK(I2350), .RSTB(I60844), .Q(I60827) );
nand I_3474 (I60836,I61381,I61107);
DFFARX1 I_3475  ( .D(I61381), .CLK(I2350), .RSTB(I60844), .Q(I60806) );
not I_3476 (I61490,I2357);
not I_3477 (I61507,I172837);
nor I_3478 (I61524,I172834,I172822);
nand I_3479 (I61541,I61524,I172825);
DFFARX1 I_3480  ( .D(I61541), .CLK(I2350), .RSTB(I61490), .Q(I61464) );
nor I_3481 (I61572,I61507,I172834);
nand I_3482 (I61589,I61572,I172831);
not I_3483 (I61479,I61589);
DFFARX1 I_3484  ( .D(I61589), .CLK(I2350), .RSTB(I61490), .Q(I61461) );
not I_3485 (I61634,I172834);
not I_3486 (I61651,I61634);
not I_3487 (I61668,I172843);
nor I_3488 (I61685,I61668,I172819);
and I_3489 (I61702,I61685,I172840);
or I_3490 (I61719,I61702,I172828);
DFFARX1 I_3491  ( .D(I61719), .CLK(I2350), .RSTB(I61490), .Q(I61736) );
nor I_3492 (I61753,I61736,I61589);
nor I_3493 (I61770,I61736,I61651);
nand I_3494 (I61476,I61541,I61770);
nand I_3495 (I61801,I61507,I172843);
nand I_3496 (I61818,I61801,I61736);
and I_3497 (I61835,I61801,I61818);
DFFARX1 I_3498  ( .D(I61835), .CLK(I2350), .RSTB(I61490), .Q(I61458) );
DFFARX1 I_3499  ( .D(I61801), .CLK(I2350), .RSTB(I61490), .Q(I61866) );
and I_3500 (I61455,I61634,I61866);
DFFARX1 I_3501  ( .D(I172849), .CLK(I2350), .RSTB(I61490), .Q(I61897) );
not I_3502 (I61914,I61897);
nor I_3503 (I61931,I61589,I61914);
and I_3504 (I61948,I61897,I61931);
nand I_3505 (I61470,I61897,I61651);
DFFARX1 I_3506  ( .D(I61897), .CLK(I2350), .RSTB(I61490), .Q(I61979) );
not I_3507 (I61467,I61979);
DFFARX1 I_3508  ( .D(I172846), .CLK(I2350), .RSTB(I61490), .Q(I62010) );
not I_3509 (I62027,I62010);
or I_3510 (I62044,I62027,I61948);
DFFARX1 I_3511  ( .D(I62044), .CLK(I2350), .RSTB(I61490), .Q(I61473) );
nand I_3512 (I61482,I62027,I61753);
DFFARX1 I_3513  ( .D(I62027), .CLK(I2350), .RSTB(I61490), .Q(I61452) );
not I_3514 (I62136,I2357);
not I_3515 (I62153,I206293);
nor I_3516 (I62170,I206305,I206287);
nand I_3517 (I62187,I62170,I206302);
DFFARX1 I_3518  ( .D(I62187), .CLK(I2350), .RSTB(I62136), .Q(I62110) );
nor I_3519 (I62218,I62153,I206305);
nand I_3520 (I62235,I62218,I206290);
not I_3521 (I62125,I62235);
DFFARX1 I_3522  ( .D(I62235), .CLK(I2350), .RSTB(I62136), .Q(I62107) );
not I_3523 (I62280,I206305);
not I_3524 (I62297,I62280);
not I_3525 (I62314,I206299);
nor I_3526 (I62331,I62314,I206278);
and I_3527 (I62348,I62331,I206281);
or I_3528 (I62365,I62348,I206284);
DFFARX1 I_3529  ( .D(I62365), .CLK(I2350), .RSTB(I62136), .Q(I62382) );
nor I_3530 (I62399,I62382,I62235);
nor I_3531 (I62416,I62382,I62297);
nand I_3532 (I62122,I62187,I62416);
nand I_3533 (I62447,I62153,I206299);
nand I_3534 (I62464,I62447,I62382);
and I_3535 (I62481,I62447,I62464);
DFFARX1 I_3536  ( .D(I62481), .CLK(I2350), .RSTB(I62136), .Q(I62104) );
DFFARX1 I_3537  ( .D(I62447), .CLK(I2350), .RSTB(I62136), .Q(I62512) );
and I_3538 (I62101,I62280,I62512);
DFFARX1 I_3539  ( .D(I206275), .CLK(I2350), .RSTB(I62136), .Q(I62543) );
not I_3540 (I62560,I62543);
nor I_3541 (I62577,I62235,I62560);
and I_3542 (I62594,I62543,I62577);
nand I_3543 (I62116,I62543,I62297);
DFFARX1 I_3544  ( .D(I62543), .CLK(I2350), .RSTB(I62136), .Q(I62625) );
not I_3545 (I62113,I62625);
DFFARX1 I_3546  ( .D(I206296), .CLK(I2350), .RSTB(I62136), .Q(I62656) );
not I_3547 (I62673,I62656);
or I_3548 (I62690,I62673,I62594);
DFFARX1 I_3549  ( .D(I62690), .CLK(I2350), .RSTB(I62136), .Q(I62119) );
nand I_3550 (I62128,I62673,I62399);
DFFARX1 I_3551  ( .D(I62673), .CLK(I2350), .RSTB(I62136), .Q(I62098) );
not I_3552 (I62782,I2357);
not I_3553 (I62799,I239474);
nor I_3554 (I62816,I239462,I239468);
nand I_3555 (I62833,I62816,I239459);
DFFARX1 I_3556  ( .D(I62833), .CLK(I2350), .RSTB(I62782), .Q(I62756) );
nor I_3557 (I62864,I62799,I239462);
nand I_3558 (I62881,I62864,I239465);
not I_3559 (I62771,I62881);
DFFARX1 I_3560  ( .D(I62881), .CLK(I2350), .RSTB(I62782), .Q(I62753) );
not I_3561 (I62926,I239462);
not I_3562 (I62943,I62926);
not I_3563 (I62960,I239477);
nor I_3564 (I62977,I62960,I239489);
and I_3565 (I62994,I62977,I239471);
or I_3566 (I63011,I62994,I239486);
DFFARX1 I_3567  ( .D(I63011), .CLK(I2350), .RSTB(I62782), .Q(I63028) );
nor I_3568 (I63045,I63028,I62881);
nor I_3569 (I63062,I63028,I62943);
nand I_3570 (I62768,I62833,I63062);
nand I_3571 (I63093,I62799,I239477);
nand I_3572 (I63110,I63093,I63028);
and I_3573 (I63127,I63093,I63110);
DFFARX1 I_3574  ( .D(I63127), .CLK(I2350), .RSTB(I62782), .Q(I62750) );
DFFARX1 I_3575  ( .D(I63093), .CLK(I2350), .RSTB(I62782), .Q(I63158) );
and I_3576 (I62747,I62926,I63158);
DFFARX1 I_3577  ( .D(I239480), .CLK(I2350), .RSTB(I62782), .Q(I63189) );
not I_3578 (I63206,I63189);
nor I_3579 (I63223,I62881,I63206);
and I_3580 (I63240,I63189,I63223);
nand I_3581 (I62762,I63189,I62943);
DFFARX1 I_3582  ( .D(I63189), .CLK(I2350), .RSTB(I62782), .Q(I63271) );
not I_3583 (I62759,I63271);
DFFARX1 I_3584  ( .D(I239483), .CLK(I2350), .RSTB(I62782), .Q(I63302) );
not I_3585 (I63319,I63302);
or I_3586 (I63336,I63319,I63240);
DFFARX1 I_3587  ( .D(I63336), .CLK(I2350), .RSTB(I62782), .Q(I62765) );
nand I_3588 (I62774,I63319,I63045);
DFFARX1 I_3589  ( .D(I63319), .CLK(I2350), .RSTB(I62782), .Q(I62744) );
not I_3590 (I63428,I2357);
not I_3591 (I63445,I241786);
nor I_3592 (I63462,I241774,I241780);
nand I_3593 (I63479,I63462,I241771);
DFFARX1 I_3594  ( .D(I63479), .CLK(I2350), .RSTB(I63428), .Q(I63402) );
nor I_3595 (I63510,I63445,I241774);
nand I_3596 (I63527,I63510,I241777);
not I_3597 (I63417,I63527);
DFFARX1 I_3598  ( .D(I63527), .CLK(I2350), .RSTB(I63428), .Q(I63399) );
not I_3599 (I63572,I241774);
not I_3600 (I63589,I63572);
not I_3601 (I63606,I241789);
nor I_3602 (I63623,I63606,I241801);
and I_3603 (I63640,I63623,I241783);
or I_3604 (I63657,I63640,I241798);
DFFARX1 I_3605  ( .D(I63657), .CLK(I2350), .RSTB(I63428), .Q(I63674) );
nor I_3606 (I63691,I63674,I63527);
nor I_3607 (I63708,I63674,I63589);
nand I_3608 (I63414,I63479,I63708);
nand I_3609 (I63739,I63445,I241789);
nand I_3610 (I63756,I63739,I63674);
and I_3611 (I63773,I63739,I63756);
DFFARX1 I_3612  ( .D(I63773), .CLK(I2350), .RSTB(I63428), .Q(I63396) );
DFFARX1 I_3613  ( .D(I63739), .CLK(I2350), .RSTB(I63428), .Q(I63804) );
and I_3614 (I63393,I63572,I63804);
DFFARX1 I_3615  ( .D(I241792), .CLK(I2350), .RSTB(I63428), .Q(I63835) );
not I_3616 (I63852,I63835);
nor I_3617 (I63869,I63527,I63852);
and I_3618 (I63886,I63835,I63869);
nand I_3619 (I63408,I63835,I63589);
DFFARX1 I_3620  ( .D(I63835), .CLK(I2350), .RSTB(I63428), .Q(I63917) );
not I_3621 (I63405,I63917);
DFFARX1 I_3622  ( .D(I241795), .CLK(I2350), .RSTB(I63428), .Q(I63948) );
not I_3623 (I63965,I63948);
or I_3624 (I63982,I63965,I63886);
DFFARX1 I_3625  ( .D(I63982), .CLK(I2350), .RSTB(I63428), .Q(I63411) );
nand I_3626 (I63420,I63965,I63691);
DFFARX1 I_3627  ( .D(I63965), .CLK(I2350), .RSTB(I63428), .Q(I63390) );
not I_3628 (I64074,I2357);
not I_3629 (I64091,I296929);
nor I_3630 (I64108,I296905,I296911);
nand I_3631 (I64125,I64108,I296914);
DFFARX1 I_3632  ( .D(I64125), .CLK(I2350), .RSTB(I64074), .Q(I64048) );
nor I_3633 (I64156,I64091,I296905);
nand I_3634 (I64173,I64156,I296923);
not I_3635 (I64063,I64173);
DFFARX1 I_3636  ( .D(I64173), .CLK(I2350), .RSTB(I64074), .Q(I64045) );
not I_3637 (I64218,I296905);
not I_3638 (I64235,I64218);
not I_3639 (I64252,I296902);
nor I_3640 (I64269,I64252,I296917);
and I_3641 (I64286,I64269,I296908);
or I_3642 (I64303,I64286,I296920);
DFFARX1 I_3643  ( .D(I64303), .CLK(I2350), .RSTB(I64074), .Q(I64320) );
nor I_3644 (I64337,I64320,I64173);
nor I_3645 (I64354,I64320,I64235);
nand I_3646 (I64060,I64125,I64354);
nand I_3647 (I64385,I64091,I296902);
nand I_3648 (I64402,I64385,I64320);
and I_3649 (I64419,I64385,I64402);
DFFARX1 I_3650  ( .D(I64419), .CLK(I2350), .RSTB(I64074), .Q(I64042) );
DFFARX1 I_3651  ( .D(I64385), .CLK(I2350), .RSTB(I64074), .Q(I64450) );
and I_3652 (I64039,I64218,I64450);
DFFARX1 I_3653  ( .D(I296932), .CLK(I2350), .RSTB(I64074), .Q(I64481) );
not I_3654 (I64498,I64481);
nor I_3655 (I64515,I64173,I64498);
and I_3656 (I64532,I64481,I64515);
nand I_3657 (I64054,I64481,I64235);
DFFARX1 I_3658  ( .D(I64481), .CLK(I2350), .RSTB(I64074), .Q(I64563) );
not I_3659 (I64051,I64563);
DFFARX1 I_3660  ( .D(I296926), .CLK(I2350), .RSTB(I64074), .Q(I64594) );
not I_3661 (I64611,I64594);
or I_3662 (I64628,I64611,I64532);
DFFARX1 I_3663  ( .D(I64628), .CLK(I2350), .RSTB(I64074), .Q(I64057) );
nand I_3664 (I64066,I64611,I64337);
DFFARX1 I_3665  ( .D(I64611), .CLK(I2350), .RSTB(I64074), .Q(I64036) );
not I_3666 (I64720,I2357);
not I_3667 (I64737,I392026);
nor I_3668 (I64754,I392023,I392020);
nand I_3669 (I64771,I64754,I392041);
DFFARX1 I_3670  ( .D(I64771), .CLK(I2350), .RSTB(I64720), .Q(I64694) );
nor I_3671 (I64802,I64737,I392023);
nand I_3672 (I64819,I64802,I392044);
not I_3673 (I64709,I64819);
DFFARX1 I_3674  ( .D(I64819), .CLK(I2350), .RSTB(I64720), .Q(I64691) );
not I_3675 (I64864,I392023);
not I_3676 (I64881,I64864);
not I_3677 (I64898,I392017);
nor I_3678 (I64915,I64898,I392029);
and I_3679 (I64932,I64915,I392038);
or I_3680 (I64949,I64932,I392032);
DFFARX1 I_3681  ( .D(I64949), .CLK(I2350), .RSTB(I64720), .Q(I64966) );
nor I_3682 (I64983,I64966,I64819);
nor I_3683 (I65000,I64966,I64881);
nand I_3684 (I64706,I64771,I65000);
nand I_3685 (I65031,I64737,I392017);
nand I_3686 (I65048,I65031,I64966);
and I_3687 (I65065,I65031,I65048);
DFFARX1 I_3688  ( .D(I65065), .CLK(I2350), .RSTB(I64720), .Q(I64688) );
DFFARX1 I_3689  ( .D(I65031), .CLK(I2350), .RSTB(I64720), .Q(I65096) );
and I_3690 (I64685,I64864,I65096);
DFFARX1 I_3691  ( .D(I392047), .CLK(I2350), .RSTB(I64720), .Q(I65127) );
not I_3692 (I65144,I65127);
nor I_3693 (I65161,I64819,I65144);
and I_3694 (I65178,I65127,I65161);
nand I_3695 (I64700,I65127,I64881);
DFFARX1 I_3696  ( .D(I65127), .CLK(I2350), .RSTB(I64720), .Q(I65209) );
not I_3697 (I64697,I65209);
DFFARX1 I_3698  ( .D(I392035), .CLK(I2350), .RSTB(I64720), .Q(I65240) );
not I_3699 (I65257,I65240);
or I_3700 (I65274,I65257,I65178);
DFFARX1 I_3701  ( .D(I65274), .CLK(I2350), .RSTB(I64720), .Q(I64703) );
nand I_3702 (I64712,I65257,I64983);
DFFARX1 I_3703  ( .D(I65257), .CLK(I2350), .RSTB(I64720), .Q(I64682) );
not I_3704 (I65366,I2357);
not I_3705 (I65383,I233391);
nor I_3706 (I65400,I233373,I233388);
nand I_3707 (I65417,I65400,I233397);
DFFARX1 I_3708  ( .D(I65417), .CLK(I2350), .RSTB(I65366), .Q(I65340) );
nor I_3709 (I65448,I65383,I233373);
nand I_3710 (I65465,I65448,I233400);
not I_3711 (I65355,I65465);
DFFARX1 I_3712  ( .D(I65465), .CLK(I2350), .RSTB(I65366), .Q(I65337) );
not I_3713 (I65510,I233373);
not I_3714 (I65527,I65510);
not I_3715 (I65544,I233403);
nor I_3716 (I65561,I65544,I233379);
and I_3717 (I65578,I65561,I233382);
or I_3718 (I65595,I65578,I233376);
DFFARX1 I_3719  ( .D(I65595), .CLK(I2350), .RSTB(I65366), .Q(I65612) );
nor I_3720 (I65629,I65612,I65465);
nor I_3721 (I65646,I65612,I65527);
nand I_3722 (I65352,I65417,I65646);
nand I_3723 (I65677,I65383,I233403);
nand I_3724 (I65694,I65677,I65612);
and I_3725 (I65711,I65677,I65694);
DFFARX1 I_3726  ( .D(I65711), .CLK(I2350), .RSTB(I65366), .Q(I65334) );
DFFARX1 I_3727  ( .D(I65677), .CLK(I2350), .RSTB(I65366), .Q(I65742) );
and I_3728 (I65331,I65510,I65742);
DFFARX1 I_3729  ( .D(I233385), .CLK(I2350), .RSTB(I65366), .Q(I65773) );
not I_3730 (I65790,I65773);
nor I_3731 (I65807,I65465,I65790);
and I_3732 (I65824,I65773,I65807);
nand I_3733 (I65346,I65773,I65527);
DFFARX1 I_3734  ( .D(I65773), .CLK(I2350), .RSTB(I65366), .Q(I65855) );
not I_3735 (I65343,I65855);
DFFARX1 I_3736  ( .D(I233394), .CLK(I2350), .RSTB(I65366), .Q(I65886) );
not I_3737 (I65903,I65886);
or I_3738 (I65920,I65903,I65824);
DFFARX1 I_3739  ( .D(I65920), .CLK(I2350), .RSTB(I65366), .Q(I65349) );
nand I_3740 (I65358,I65903,I65629);
DFFARX1 I_3741  ( .D(I65903), .CLK(I2350), .RSTB(I65366), .Q(I65328) );
not I_3742 (I66012,I2357);
not I_3743 (I66029,I1727);
nor I_3744 (I66046,I1671,I1479);
nand I_3745 (I66063,I66046,I2167);
DFFARX1 I_3746  ( .D(I66063), .CLK(I2350), .RSTB(I66012), .Q(I65986) );
nor I_3747 (I66094,I66029,I1671);
nand I_3748 (I66111,I66094,I2047);
not I_3749 (I66001,I66111);
DFFARX1 I_3750  ( .D(I66111), .CLK(I2350), .RSTB(I66012), .Q(I65983) );
not I_3751 (I66156,I1671);
not I_3752 (I66173,I66156);
not I_3753 (I66190,I1863);
nor I_3754 (I66207,I66190,I2343);
and I_3755 (I66224,I66207,I2079);
or I_3756 (I66241,I66224,I1247);
DFFARX1 I_3757  ( .D(I66241), .CLK(I2350), .RSTB(I66012), .Q(I66258) );
nor I_3758 (I66275,I66258,I66111);
nor I_3759 (I66292,I66258,I66173);
nand I_3760 (I65998,I66063,I66292);
nand I_3761 (I66323,I66029,I1863);
nand I_3762 (I66340,I66323,I66258);
and I_3763 (I66357,I66323,I66340);
DFFARX1 I_3764  ( .D(I66357), .CLK(I2350), .RSTB(I66012), .Q(I65980) );
DFFARX1 I_3765  ( .D(I66323), .CLK(I2350), .RSTB(I66012), .Q(I66388) );
and I_3766 (I65977,I66156,I66388);
DFFARX1 I_3767  ( .D(I2247), .CLK(I2350), .RSTB(I66012), .Q(I66419) );
not I_3768 (I66436,I66419);
nor I_3769 (I66453,I66111,I66436);
and I_3770 (I66470,I66419,I66453);
nand I_3771 (I65992,I66419,I66173);
DFFARX1 I_3772  ( .D(I66419), .CLK(I2350), .RSTB(I66012), .Q(I66501) );
not I_3773 (I65989,I66501);
DFFARX1 I_3774  ( .D(I1487), .CLK(I2350), .RSTB(I66012), .Q(I66532) );
not I_3775 (I66549,I66532);
or I_3776 (I66566,I66549,I66470);
DFFARX1 I_3777  ( .D(I66566), .CLK(I2350), .RSTB(I66012), .Q(I65995) );
nand I_3778 (I66004,I66549,I66275);
DFFARX1 I_3779  ( .D(I66549), .CLK(I2350), .RSTB(I66012), .Q(I65974) );
not I_3780 (I66658,I2357);
not I_3781 (I66675,I211461);
nor I_3782 (I66692,I211473,I211455);
nand I_3783 (I66709,I66692,I211470);
DFFARX1 I_3784  ( .D(I66709), .CLK(I2350), .RSTB(I66658), .Q(I66632) );
nor I_3785 (I66740,I66675,I211473);
nand I_3786 (I66757,I66740,I211458);
not I_3787 (I66647,I66757);
DFFARX1 I_3788  ( .D(I66757), .CLK(I2350), .RSTB(I66658), .Q(I66629) );
not I_3789 (I66802,I211473);
not I_3790 (I66819,I66802);
not I_3791 (I66836,I211467);
nor I_3792 (I66853,I66836,I211446);
and I_3793 (I66870,I66853,I211449);
or I_3794 (I66887,I66870,I211452);
DFFARX1 I_3795  ( .D(I66887), .CLK(I2350), .RSTB(I66658), .Q(I66904) );
nor I_3796 (I66921,I66904,I66757);
nor I_3797 (I66938,I66904,I66819);
nand I_3798 (I66644,I66709,I66938);
nand I_3799 (I66969,I66675,I211467);
nand I_3800 (I66986,I66969,I66904);
and I_3801 (I67003,I66969,I66986);
DFFARX1 I_3802  ( .D(I67003), .CLK(I2350), .RSTB(I66658), .Q(I66626) );
DFFARX1 I_3803  ( .D(I66969), .CLK(I2350), .RSTB(I66658), .Q(I67034) );
and I_3804 (I66623,I66802,I67034);
DFFARX1 I_3805  ( .D(I211443), .CLK(I2350), .RSTB(I66658), .Q(I67065) );
not I_3806 (I67082,I67065);
nor I_3807 (I67099,I66757,I67082);
and I_3808 (I67116,I67065,I67099);
nand I_3809 (I66638,I67065,I66819);
DFFARX1 I_3810  ( .D(I67065), .CLK(I2350), .RSTB(I66658), .Q(I67147) );
not I_3811 (I66635,I67147);
DFFARX1 I_3812  ( .D(I211464), .CLK(I2350), .RSTB(I66658), .Q(I67178) );
not I_3813 (I67195,I67178);
or I_3814 (I67212,I67195,I67116);
DFFARX1 I_3815  ( .D(I67212), .CLK(I2350), .RSTB(I66658), .Q(I66641) );
nand I_3816 (I66650,I67195,I66921);
DFFARX1 I_3817  ( .D(I67195), .CLK(I2350), .RSTB(I66658), .Q(I66620) );
not I_3818 (I67304,I2357);
not I_3819 (I67321,I160240);
nor I_3820 (I67338,I160237,I160225);
nand I_3821 (I67355,I67338,I160228);
DFFARX1 I_3822  ( .D(I67355), .CLK(I2350), .RSTB(I67304), .Q(I67278) );
nor I_3823 (I67386,I67321,I160237);
nand I_3824 (I67403,I67386,I160234);
not I_3825 (I67293,I67403);
DFFARX1 I_3826  ( .D(I67403), .CLK(I2350), .RSTB(I67304), .Q(I67275) );
not I_3827 (I67448,I160237);
not I_3828 (I67465,I67448);
not I_3829 (I67482,I160246);
nor I_3830 (I67499,I67482,I160222);
and I_3831 (I67516,I67499,I160243);
or I_3832 (I67533,I67516,I160231);
DFFARX1 I_3833  ( .D(I67533), .CLK(I2350), .RSTB(I67304), .Q(I67550) );
nor I_3834 (I67567,I67550,I67403);
nor I_3835 (I67584,I67550,I67465);
nand I_3836 (I67290,I67355,I67584);
nand I_3837 (I67615,I67321,I160246);
nand I_3838 (I67632,I67615,I67550);
and I_3839 (I67649,I67615,I67632);
DFFARX1 I_3840  ( .D(I67649), .CLK(I2350), .RSTB(I67304), .Q(I67272) );
DFFARX1 I_3841  ( .D(I67615), .CLK(I2350), .RSTB(I67304), .Q(I67680) );
and I_3842 (I67269,I67448,I67680);
DFFARX1 I_3843  ( .D(I160252), .CLK(I2350), .RSTB(I67304), .Q(I67711) );
not I_3844 (I67728,I67711);
nor I_3845 (I67745,I67403,I67728);
and I_3846 (I67762,I67711,I67745);
nand I_3847 (I67284,I67711,I67465);
DFFARX1 I_3848  ( .D(I67711), .CLK(I2350), .RSTB(I67304), .Q(I67793) );
not I_3849 (I67281,I67793);
DFFARX1 I_3850  ( .D(I160249), .CLK(I2350), .RSTB(I67304), .Q(I67824) );
not I_3851 (I67841,I67824);
or I_3852 (I67858,I67841,I67762);
DFFARX1 I_3853  ( .D(I67858), .CLK(I2350), .RSTB(I67304), .Q(I67287) );
nand I_3854 (I67296,I67841,I67567);
DFFARX1 I_3855  ( .D(I67841), .CLK(I2350), .RSTB(I67304), .Q(I67266) );
not I_3856 (I67950,I2357);
not I_3857 (I67967,I86715);
nor I_3858 (I67984,I86703,I86709);
nand I_3859 (I68001,I67984,I86718);
DFFARX1 I_3860  ( .D(I68001), .CLK(I2350), .RSTB(I67950), .Q(I67924) );
nor I_3861 (I68032,I67967,I86703);
nand I_3862 (I68049,I68032,I86706);
not I_3863 (I67939,I68049);
DFFARX1 I_3864  ( .D(I68049), .CLK(I2350), .RSTB(I67950), .Q(I67921) );
not I_3865 (I68094,I86703);
not I_3866 (I68111,I68094);
not I_3867 (I68128,I86727);
nor I_3868 (I68145,I68128,I86700);
and I_3869 (I68162,I68145,I86721);
or I_3870 (I68179,I68162,I86712);
DFFARX1 I_3871  ( .D(I68179), .CLK(I2350), .RSTB(I67950), .Q(I68196) );
nor I_3872 (I68213,I68196,I68049);
nor I_3873 (I68230,I68196,I68111);
nand I_3874 (I67936,I68001,I68230);
nand I_3875 (I68261,I67967,I86727);
nand I_3876 (I68278,I68261,I68196);
and I_3877 (I68295,I68261,I68278);
DFFARX1 I_3878  ( .D(I68295), .CLK(I2350), .RSTB(I67950), .Q(I67918) );
DFFARX1 I_3879  ( .D(I68261), .CLK(I2350), .RSTB(I67950), .Q(I68326) );
and I_3880 (I67915,I68094,I68326);
DFFARX1 I_3881  ( .D(I86697), .CLK(I2350), .RSTB(I67950), .Q(I68357) );
not I_3882 (I68374,I68357);
nor I_3883 (I68391,I68049,I68374);
and I_3884 (I68408,I68357,I68391);
nand I_3885 (I67930,I68357,I68111);
DFFARX1 I_3886  ( .D(I68357), .CLK(I2350), .RSTB(I67950), .Q(I68439) );
not I_3887 (I67927,I68439);
DFFARX1 I_3888  ( .D(I86724), .CLK(I2350), .RSTB(I67950), .Q(I68470) );
not I_3889 (I68487,I68470);
or I_3890 (I68504,I68487,I68408);
DFFARX1 I_3891  ( .D(I68504), .CLK(I2350), .RSTB(I67950), .Q(I67933) );
nand I_3892 (I67942,I68487,I68213);
DFFARX1 I_3893  ( .D(I68487), .CLK(I2350), .RSTB(I67950), .Q(I67912) );
not I_3894 (I68596,I2357);
not I_3895 (I68613,I290979);
nor I_3896 (I68630,I290955,I290961);
nand I_3897 (I68647,I68630,I290964);
DFFARX1 I_3898  ( .D(I68647), .CLK(I2350), .RSTB(I68596), .Q(I68570) );
nor I_3899 (I68678,I68613,I290955);
nand I_3900 (I68695,I68678,I290973);
not I_3901 (I68585,I68695);
DFFARX1 I_3902  ( .D(I68695), .CLK(I2350), .RSTB(I68596), .Q(I68567) );
not I_3903 (I68740,I290955);
not I_3904 (I68757,I68740);
not I_3905 (I68774,I290952);
nor I_3906 (I68791,I68774,I290967);
and I_3907 (I68808,I68791,I290958);
or I_3908 (I68825,I68808,I290970);
DFFARX1 I_3909  ( .D(I68825), .CLK(I2350), .RSTB(I68596), .Q(I68842) );
nor I_3910 (I68859,I68842,I68695);
nor I_3911 (I68876,I68842,I68757);
nand I_3912 (I68582,I68647,I68876);
nand I_3913 (I68907,I68613,I290952);
nand I_3914 (I68924,I68907,I68842);
and I_3915 (I68941,I68907,I68924);
DFFARX1 I_3916  ( .D(I68941), .CLK(I2350), .RSTB(I68596), .Q(I68564) );
DFFARX1 I_3917  ( .D(I68907), .CLK(I2350), .RSTB(I68596), .Q(I68972) );
and I_3918 (I68561,I68740,I68972);
DFFARX1 I_3919  ( .D(I290982), .CLK(I2350), .RSTB(I68596), .Q(I69003) );
not I_3920 (I69020,I69003);
nor I_3921 (I69037,I68695,I69020);
and I_3922 (I69054,I69003,I69037);
nand I_3923 (I68576,I69003,I68757);
DFFARX1 I_3924  ( .D(I69003), .CLK(I2350), .RSTB(I68596), .Q(I69085) );
not I_3925 (I68573,I69085);
DFFARX1 I_3926  ( .D(I290976), .CLK(I2350), .RSTB(I68596), .Q(I69116) );
not I_3927 (I69133,I69116);
or I_3928 (I69150,I69133,I69054);
DFFARX1 I_3929  ( .D(I69150), .CLK(I2350), .RSTB(I68596), .Q(I68579) );
nand I_3930 (I68588,I69133,I68859);
DFFARX1 I_3931  ( .D(I69133), .CLK(I2350), .RSTB(I68596), .Q(I68558) );
not I_3932 (I69242,I2357);
not I_3933 (I69259,I355246);
nor I_3934 (I69276,I355261,I355276);
nand I_3935 (I69293,I69276,I355264);
DFFARX1 I_3936  ( .D(I69293), .CLK(I2350), .RSTB(I69242), .Q(I69216) );
nor I_3937 (I69324,I69259,I355261);
nand I_3938 (I69341,I69324,I355267);
not I_3939 (I69231,I69341);
DFFARX1 I_3940  ( .D(I69341), .CLK(I2350), .RSTB(I69242), .Q(I69213) );
not I_3941 (I69386,I355261);
not I_3942 (I69403,I69386);
not I_3943 (I69420,I355273);
nor I_3944 (I69437,I69420,I355270);
and I_3945 (I69454,I69437,I355249);
or I_3946 (I69471,I69454,I355258);
DFFARX1 I_3947  ( .D(I69471), .CLK(I2350), .RSTB(I69242), .Q(I69488) );
nor I_3948 (I69505,I69488,I69341);
nor I_3949 (I69522,I69488,I69403);
nand I_3950 (I69228,I69293,I69522);
nand I_3951 (I69553,I69259,I355273);
nand I_3952 (I69570,I69553,I69488);
and I_3953 (I69587,I69553,I69570);
DFFARX1 I_3954  ( .D(I69587), .CLK(I2350), .RSTB(I69242), .Q(I69210) );
DFFARX1 I_3955  ( .D(I69553), .CLK(I2350), .RSTB(I69242), .Q(I69618) );
and I_3956 (I69207,I69386,I69618);
DFFARX1 I_3957  ( .D(I355255), .CLK(I2350), .RSTB(I69242), .Q(I69649) );
not I_3958 (I69666,I69649);
nor I_3959 (I69683,I69341,I69666);
and I_3960 (I69700,I69649,I69683);
nand I_3961 (I69222,I69649,I69403);
DFFARX1 I_3962  ( .D(I69649), .CLK(I2350), .RSTB(I69242), .Q(I69731) );
not I_3963 (I69219,I69731);
DFFARX1 I_3964  ( .D(I355252), .CLK(I2350), .RSTB(I69242), .Q(I69762) );
not I_3965 (I69779,I69762);
or I_3966 (I69796,I69779,I69700);
DFFARX1 I_3967  ( .D(I69796), .CLK(I2350), .RSTB(I69242), .Q(I69225) );
nand I_3968 (I69234,I69779,I69505);
DFFARX1 I_3969  ( .D(I69779), .CLK(I2350), .RSTB(I69242), .Q(I69204) );
not I_3970 (I69888,I2357);
not I_3971 (I69905,I294549);
nor I_3972 (I69922,I294525,I294531);
nand I_3973 (I69939,I69922,I294534);
DFFARX1 I_3974  ( .D(I69939), .CLK(I2350), .RSTB(I69888), .Q(I69862) );
nor I_3975 (I69970,I69905,I294525);
nand I_3976 (I69987,I69970,I294543);
not I_3977 (I69877,I69987);
DFFARX1 I_3978  ( .D(I69987), .CLK(I2350), .RSTB(I69888), .Q(I69859) );
not I_3979 (I70032,I294525);
not I_3980 (I70049,I70032);
not I_3981 (I70066,I294522);
nor I_3982 (I70083,I70066,I294537);
and I_3983 (I70100,I70083,I294528);
or I_3984 (I70117,I70100,I294540);
DFFARX1 I_3985  ( .D(I70117), .CLK(I2350), .RSTB(I69888), .Q(I70134) );
nor I_3986 (I70151,I70134,I69987);
nor I_3987 (I70168,I70134,I70049);
nand I_3988 (I69874,I69939,I70168);
nand I_3989 (I70199,I69905,I294522);
nand I_3990 (I70216,I70199,I70134);
and I_3991 (I70233,I70199,I70216);
DFFARX1 I_3992  ( .D(I70233), .CLK(I2350), .RSTB(I69888), .Q(I69856) );
DFFARX1 I_3993  ( .D(I70199), .CLK(I2350), .RSTB(I69888), .Q(I70264) );
and I_3994 (I69853,I70032,I70264);
DFFARX1 I_3995  ( .D(I294552), .CLK(I2350), .RSTB(I69888), .Q(I70295) );
not I_3996 (I70312,I70295);
nor I_3997 (I70329,I69987,I70312);
and I_3998 (I70346,I70295,I70329);
nand I_3999 (I69868,I70295,I70049);
DFFARX1 I_4000  ( .D(I70295), .CLK(I2350), .RSTB(I69888), .Q(I70377) );
not I_4001 (I69865,I70377);
DFFARX1 I_4002  ( .D(I294546), .CLK(I2350), .RSTB(I69888), .Q(I70408) );
not I_4003 (I70425,I70408);
or I_4004 (I70442,I70425,I70346);
DFFARX1 I_4005  ( .D(I70442), .CLK(I2350), .RSTB(I69888), .Q(I69871) );
nand I_4006 (I69880,I70425,I70151);
DFFARX1 I_4007  ( .D(I70425), .CLK(I2350), .RSTB(I69888), .Q(I69850) );
not I_4008 (I70534,I2357);
not I_4009 (I70551,I328452);
nor I_4010 (I70568,I328437,I328464);
nand I_4011 (I70585,I70568,I328440);
DFFARX1 I_4012  ( .D(I70585), .CLK(I2350), .RSTB(I70534), .Q(I70508) );
nor I_4013 (I70616,I70551,I328437);
nand I_4014 (I70633,I70616,I328455);
not I_4015 (I70523,I70633);
DFFARX1 I_4016  ( .D(I70633), .CLK(I2350), .RSTB(I70534), .Q(I70505) );
not I_4017 (I70678,I328437);
not I_4018 (I70695,I70678);
not I_4019 (I70712,I328467);
nor I_4020 (I70729,I70712,I328449);
and I_4021 (I70746,I70729,I328458);
or I_4022 (I70763,I70746,I328443);
DFFARX1 I_4023  ( .D(I70763), .CLK(I2350), .RSTB(I70534), .Q(I70780) );
nor I_4024 (I70797,I70780,I70633);
nor I_4025 (I70814,I70780,I70695);
nand I_4026 (I70520,I70585,I70814);
nand I_4027 (I70845,I70551,I328467);
nand I_4028 (I70862,I70845,I70780);
and I_4029 (I70879,I70845,I70862);
DFFARX1 I_4030  ( .D(I70879), .CLK(I2350), .RSTB(I70534), .Q(I70502) );
DFFARX1 I_4031  ( .D(I70845), .CLK(I2350), .RSTB(I70534), .Q(I70910) );
and I_4032 (I70499,I70678,I70910);
DFFARX1 I_4033  ( .D(I328446), .CLK(I2350), .RSTB(I70534), .Q(I70941) );
not I_4034 (I70958,I70941);
nor I_4035 (I70975,I70633,I70958);
and I_4036 (I70992,I70941,I70975);
nand I_4037 (I70514,I70941,I70695);
DFFARX1 I_4038  ( .D(I70941), .CLK(I2350), .RSTB(I70534), .Q(I71023) );
not I_4039 (I70511,I71023);
DFFARX1 I_4040  ( .D(I328461), .CLK(I2350), .RSTB(I70534), .Q(I71054) );
not I_4041 (I71071,I71054);
or I_4042 (I71088,I71071,I70992);
DFFARX1 I_4043  ( .D(I71088), .CLK(I2350), .RSTB(I70534), .Q(I70517) );
nand I_4044 (I70526,I71071,I70797);
DFFARX1 I_4045  ( .D(I71071), .CLK(I2350), .RSTB(I70534), .Q(I70496) );
not I_4046 (I71180,I2357);
not I_4047 (I71197,I1775);
nor I_4048 (I71214,I2175,I1567);
nand I_4049 (I71231,I71214,I2287);
DFFARX1 I_4050  ( .D(I71231), .CLK(I2350), .RSTB(I71180), .Q(I71154) );
nor I_4051 (I71262,I71197,I2175);
nand I_4052 (I71279,I71262,I1591);
not I_4053 (I71169,I71279);
DFFARX1 I_4054  ( .D(I71279), .CLK(I2350), .RSTB(I71180), .Q(I71151) );
not I_4055 (I71324,I2175);
not I_4056 (I71341,I71324);
not I_4057 (I71358,I2095);
nor I_4058 (I71375,I71358,I1807);
and I_4059 (I71392,I71375,I2295);
or I_4060 (I71409,I71392,I1391);
DFFARX1 I_4061  ( .D(I71409), .CLK(I2350), .RSTB(I71180), .Q(I71426) );
nor I_4062 (I71443,I71426,I71279);
nor I_4063 (I71460,I71426,I71341);
nand I_4064 (I71166,I71231,I71460);
nand I_4065 (I71491,I71197,I2095);
nand I_4066 (I71508,I71491,I71426);
and I_4067 (I71525,I71491,I71508);
DFFARX1 I_4068  ( .D(I71525), .CLK(I2350), .RSTB(I71180), .Q(I71148) );
DFFARX1 I_4069  ( .D(I71491), .CLK(I2350), .RSTB(I71180), .Q(I71556) );
and I_4070 (I71145,I71324,I71556);
DFFARX1 I_4071  ( .D(I1999), .CLK(I2350), .RSTB(I71180), .Q(I71587) );
not I_4072 (I71604,I71587);
nor I_4073 (I71621,I71279,I71604);
and I_4074 (I71638,I71587,I71621);
nand I_4075 (I71160,I71587,I71341);
DFFARX1 I_4076  ( .D(I71587), .CLK(I2350), .RSTB(I71180), .Q(I71669) );
not I_4077 (I71157,I71669);
DFFARX1 I_4078  ( .D(I2063), .CLK(I2350), .RSTB(I71180), .Q(I71700) );
not I_4079 (I71717,I71700);
or I_4080 (I71734,I71717,I71638);
DFFARX1 I_4081  ( .D(I71734), .CLK(I2350), .RSTB(I71180), .Q(I71163) );
nand I_4082 (I71172,I71717,I71443);
DFFARX1 I_4083  ( .D(I71717), .CLK(I2350), .RSTB(I71180), .Q(I71142) );
not I_4084 (I71826,I2357);
not I_4085 (I71843,I352730);
nor I_4086 (I71860,I352745,I352760);
nand I_4087 (I71877,I71860,I352748);
DFFARX1 I_4088  ( .D(I71877), .CLK(I2350), .RSTB(I71826), .Q(I71800) );
nor I_4089 (I71908,I71843,I352745);
nand I_4090 (I71925,I71908,I352751);
not I_4091 (I71815,I71925);
DFFARX1 I_4092  ( .D(I71925), .CLK(I2350), .RSTB(I71826), .Q(I71797) );
not I_4093 (I71970,I352745);
not I_4094 (I71987,I71970);
not I_4095 (I72004,I352757);
nor I_4096 (I72021,I72004,I352754);
and I_4097 (I72038,I72021,I352733);
or I_4098 (I72055,I72038,I352742);
DFFARX1 I_4099  ( .D(I72055), .CLK(I2350), .RSTB(I71826), .Q(I72072) );
nor I_4100 (I72089,I72072,I71925);
nor I_4101 (I72106,I72072,I71987);
nand I_4102 (I71812,I71877,I72106);
nand I_4103 (I72137,I71843,I352757);
nand I_4104 (I72154,I72137,I72072);
and I_4105 (I72171,I72137,I72154);
DFFARX1 I_4106  ( .D(I72171), .CLK(I2350), .RSTB(I71826), .Q(I71794) );
DFFARX1 I_4107  ( .D(I72137), .CLK(I2350), .RSTB(I71826), .Q(I72202) );
and I_4108 (I71791,I71970,I72202);
DFFARX1 I_4109  ( .D(I352739), .CLK(I2350), .RSTB(I71826), .Q(I72233) );
not I_4110 (I72250,I72233);
nor I_4111 (I72267,I71925,I72250);
and I_4112 (I72284,I72233,I72267);
nand I_4113 (I71806,I72233,I71987);
DFFARX1 I_4114  ( .D(I72233), .CLK(I2350), .RSTB(I71826), .Q(I72315) );
not I_4115 (I71803,I72315);
DFFARX1 I_4116  ( .D(I352736), .CLK(I2350), .RSTB(I71826), .Q(I72346) );
not I_4117 (I72363,I72346);
or I_4118 (I72380,I72363,I72284);
DFFARX1 I_4119  ( .D(I72380), .CLK(I2350), .RSTB(I71826), .Q(I71809) );
nand I_4120 (I71818,I72363,I72089);
DFFARX1 I_4121  ( .D(I72363), .CLK(I2350), .RSTB(I71826), .Q(I71788) );
not I_4122 (I72472,I2357);
not I_4123 (I72489,I298714);
nor I_4124 (I72506,I298690,I298696);
nand I_4125 (I72523,I72506,I298699);
DFFARX1 I_4126  ( .D(I72523), .CLK(I2350), .RSTB(I72472), .Q(I72446) );
nor I_4127 (I72554,I72489,I298690);
nand I_4128 (I72571,I72554,I298708);
not I_4129 (I72461,I72571);
DFFARX1 I_4130  ( .D(I72571), .CLK(I2350), .RSTB(I72472), .Q(I72443) );
not I_4131 (I72616,I298690);
not I_4132 (I72633,I72616);
not I_4133 (I72650,I298687);
nor I_4134 (I72667,I72650,I298702);
and I_4135 (I72684,I72667,I298693);
or I_4136 (I72701,I72684,I298705);
DFFARX1 I_4137  ( .D(I72701), .CLK(I2350), .RSTB(I72472), .Q(I72718) );
nor I_4138 (I72735,I72718,I72571);
nor I_4139 (I72752,I72718,I72633);
nand I_4140 (I72458,I72523,I72752);
nand I_4141 (I72783,I72489,I298687);
nand I_4142 (I72800,I72783,I72718);
and I_4143 (I72817,I72783,I72800);
DFFARX1 I_4144  ( .D(I72817), .CLK(I2350), .RSTB(I72472), .Q(I72440) );
DFFARX1 I_4145  ( .D(I72783), .CLK(I2350), .RSTB(I72472), .Q(I72848) );
and I_4146 (I72437,I72616,I72848);
DFFARX1 I_4147  ( .D(I298717), .CLK(I2350), .RSTB(I72472), .Q(I72879) );
not I_4148 (I72896,I72879);
nor I_4149 (I72913,I72571,I72896);
and I_4150 (I72930,I72879,I72913);
nand I_4151 (I72452,I72879,I72633);
DFFARX1 I_4152  ( .D(I72879), .CLK(I2350), .RSTB(I72472), .Q(I72961) );
not I_4153 (I72449,I72961);
DFFARX1 I_4154  ( .D(I298711), .CLK(I2350), .RSTB(I72472), .Q(I72992) );
not I_4155 (I73009,I72992);
or I_4156 (I73026,I73009,I72930);
DFFARX1 I_4157  ( .D(I73026), .CLK(I2350), .RSTB(I72472), .Q(I72455) );
nand I_4158 (I72464,I73009,I72735);
DFFARX1 I_4159  ( .D(I73009), .CLK(I2350), .RSTB(I72472), .Q(I72434) );
not I_4160 (I73118,I2357);
not I_4161 (I73135,I257392);
nor I_4162 (I73152,I257380,I257386);
nand I_4163 (I73169,I73152,I257377);
DFFARX1 I_4164  ( .D(I73169), .CLK(I2350), .RSTB(I73118), .Q(I73092) );
nor I_4165 (I73200,I73135,I257380);
nand I_4166 (I73217,I73200,I257383);
not I_4167 (I73107,I73217);
DFFARX1 I_4168  ( .D(I73217), .CLK(I2350), .RSTB(I73118), .Q(I73089) );
not I_4169 (I73262,I257380);
not I_4170 (I73279,I73262);
not I_4171 (I73296,I257395);
nor I_4172 (I73313,I73296,I257407);
and I_4173 (I73330,I73313,I257389);
or I_4174 (I73347,I73330,I257404);
DFFARX1 I_4175  ( .D(I73347), .CLK(I2350), .RSTB(I73118), .Q(I73364) );
nor I_4176 (I73381,I73364,I73217);
nor I_4177 (I73398,I73364,I73279);
nand I_4178 (I73104,I73169,I73398);
nand I_4179 (I73429,I73135,I257395);
nand I_4180 (I73446,I73429,I73364);
and I_4181 (I73463,I73429,I73446);
DFFARX1 I_4182  ( .D(I73463), .CLK(I2350), .RSTB(I73118), .Q(I73086) );
DFFARX1 I_4183  ( .D(I73429), .CLK(I2350), .RSTB(I73118), .Q(I73494) );
and I_4184 (I73083,I73262,I73494);
DFFARX1 I_4185  ( .D(I257398), .CLK(I2350), .RSTB(I73118), .Q(I73525) );
not I_4186 (I73542,I73525);
nor I_4187 (I73559,I73217,I73542);
and I_4188 (I73576,I73525,I73559);
nand I_4189 (I73098,I73525,I73279);
DFFARX1 I_4190  ( .D(I73525), .CLK(I2350), .RSTB(I73118), .Q(I73607) );
not I_4191 (I73095,I73607);
DFFARX1 I_4192  ( .D(I257401), .CLK(I2350), .RSTB(I73118), .Q(I73638) );
not I_4193 (I73655,I73638);
or I_4194 (I73672,I73655,I73576);
DFFARX1 I_4195  ( .D(I73672), .CLK(I2350), .RSTB(I73118), .Q(I73101) );
nand I_4196 (I73110,I73655,I73381);
DFFARX1 I_4197  ( .D(I73655), .CLK(I2350), .RSTB(I73118), .Q(I73080) );
not I_4198 (I73764,I2357);
not I_4199 (I73781,I180793);
nor I_4200 (I73798,I180790,I180778);
nand I_4201 (I73815,I73798,I180781);
DFFARX1 I_4202  ( .D(I73815), .CLK(I2350), .RSTB(I73764), .Q(I73738) );
nor I_4203 (I73846,I73781,I180790);
nand I_4204 (I73863,I73846,I180787);
not I_4205 (I73753,I73863);
DFFARX1 I_4206  ( .D(I73863), .CLK(I2350), .RSTB(I73764), .Q(I73735) );
not I_4207 (I73908,I180790);
not I_4208 (I73925,I73908);
not I_4209 (I73942,I180799);
nor I_4210 (I73959,I73942,I180775);
and I_4211 (I73976,I73959,I180796);
or I_4212 (I73993,I73976,I180784);
DFFARX1 I_4213  ( .D(I73993), .CLK(I2350), .RSTB(I73764), .Q(I74010) );
nor I_4214 (I74027,I74010,I73863);
nor I_4215 (I74044,I74010,I73925);
nand I_4216 (I73750,I73815,I74044);
nand I_4217 (I74075,I73781,I180799);
nand I_4218 (I74092,I74075,I74010);
and I_4219 (I74109,I74075,I74092);
DFFARX1 I_4220  ( .D(I74109), .CLK(I2350), .RSTB(I73764), .Q(I73732) );
DFFARX1 I_4221  ( .D(I74075), .CLK(I2350), .RSTB(I73764), .Q(I74140) );
and I_4222 (I73729,I73908,I74140);
DFFARX1 I_4223  ( .D(I180805), .CLK(I2350), .RSTB(I73764), .Q(I74171) );
not I_4224 (I74188,I74171);
nor I_4225 (I74205,I73863,I74188);
and I_4226 (I74222,I74171,I74205);
nand I_4227 (I73744,I74171,I73925);
DFFARX1 I_4228  ( .D(I74171), .CLK(I2350), .RSTB(I73764), .Q(I74253) );
not I_4229 (I73741,I74253);
DFFARX1 I_4230  ( .D(I180802), .CLK(I2350), .RSTB(I73764), .Q(I74284) );
not I_4231 (I74301,I74284);
or I_4232 (I74318,I74301,I74222);
DFFARX1 I_4233  ( .D(I74318), .CLK(I2350), .RSTB(I73764), .Q(I73747) );
nand I_4234 (I73756,I74301,I74027);
DFFARX1 I_4235  ( .D(I74301), .CLK(I2350), .RSTB(I73764), .Q(I73726) );
not I_4236 (I74410,I2357);
not I_4237 (I74427,I178804);
nor I_4238 (I74444,I178801,I178789);
nand I_4239 (I74461,I74444,I178792);
DFFARX1 I_4240  ( .D(I74461), .CLK(I2350), .RSTB(I74410), .Q(I74384) );
nor I_4241 (I74492,I74427,I178801);
nand I_4242 (I74509,I74492,I178798);
not I_4243 (I74399,I74509);
DFFARX1 I_4244  ( .D(I74509), .CLK(I2350), .RSTB(I74410), .Q(I74381) );
not I_4245 (I74554,I178801);
not I_4246 (I74571,I74554);
not I_4247 (I74588,I178810);
nor I_4248 (I74605,I74588,I178786);
and I_4249 (I74622,I74605,I178807);
or I_4250 (I74639,I74622,I178795);
DFFARX1 I_4251  ( .D(I74639), .CLK(I2350), .RSTB(I74410), .Q(I74656) );
nor I_4252 (I74673,I74656,I74509);
nor I_4253 (I74690,I74656,I74571);
nand I_4254 (I74396,I74461,I74690);
nand I_4255 (I74721,I74427,I178810);
nand I_4256 (I74738,I74721,I74656);
and I_4257 (I74755,I74721,I74738);
DFFARX1 I_4258  ( .D(I74755), .CLK(I2350), .RSTB(I74410), .Q(I74378) );
DFFARX1 I_4259  ( .D(I74721), .CLK(I2350), .RSTB(I74410), .Q(I74786) );
and I_4260 (I74375,I74554,I74786);
DFFARX1 I_4261  ( .D(I178816), .CLK(I2350), .RSTB(I74410), .Q(I74817) );
not I_4262 (I74834,I74817);
nor I_4263 (I74851,I74509,I74834);
and I_4264 (I74868,I74817,I74851);
nand I_4265 (I74390,I74817,I74571);
DFFARX1 I_4266  ( .D(I74817), .CLK(I2350), .RSTB(I74410), .Q(I74899) );
not I_4267 (I74387,I74899);
DFFARX1 I_4268  ( .D(I178813), .CLK(I2350), .RSTB(I74410), .Q(I74930) );
not I_4269 (I74947,I74930);
or I_4270 (I74964,I74947,I74868);
DFFARX1 I_4271  ( .D(I74964), .CLK(I2350), .RSTB(I74410), .Q(I74393) );
nand I_4272 (I74402,I74947,I74673);
DFFARX1 I_4273  ( .D(I74947), .CLK(I2350), .RSTB(I74410), .Q(I74372) );
not I_4274 (I75056,I2357);
not I_4275 (I75073,I150958);
nor I_4276 (I75090,I150955,I150943);
nand I_4277 (I75107,I75090,I150946);
DFFARX1 I_4278  ( .D(I75107), .CLK(I2350), .RSTB(I75056), .Q(I75030) );
nor I_4279 (I75138,I75073,I150955);
nand I_4280 (I75155,I75138,I150952);
not I_4281 (I75045,I75155);
DFFARX1 I_4282  ( .D(I75155), .CLK(I2350), .RSTB(I75056), .Q(I75027) );
not I_4283 (I75200,I150955);
not I_4284 (I75217,I75200);
not I_4285 (I75234,I150964);
nor I_4286 (I75251,I75234,I150940);
and I_4287 (I75268,I75251,I150961);
or I_4288 (I75285,I75268,I150949);
DFFARX1 I_4289  ( .D(I75285), .CLK(I2350), .RSTB(I75056), .Q(I75302) );
nor I_4290 (I75319,I75302,I75155);
nor I_4291 (I75336,I75302,I75217);
nand I_4292 (I75042,I75107,I75336);
nand I_4293 (I75367,I75073,I150964);
nand I_4294 (I75384,I75367,I75302);
and I_4295 (I75401,I75367,I75384);
DFFARX1 I_4296  ( .D(I75401), .CLK(I2350), .RSTB(I75056), .Q(I75024) );
DFFARX1 I_4297  ( .D(I75367), .CLK(I2350), .RSTB(I75056), .Q(I75432) );
and I_4298 (I75021,I75200,I75432);
DFFARX1 I_4299  ( .D(I150970), .CLK(I2350), .RSTB(I75056), .Q(I75463) );
not I_4300 (I75480,I75463);
nor I_4301 (I75497,I75155,I75480);
and I_4302 (I75514,I75463,I75497);
nand I_4303 (I75036,I75463,I75217);
DFFARX1 I_4304  ( .D(I75463), .CLK(I2350), .RSTB(I75056), .Q(I75545) );
not I_4305 (I75033,I75545);
DFFARX1 I_4306  ( .D(I150967), .CLK(I2350), .RSTB(I75056), .Q(I75576) );
not I_4307 (I75593,I75576);
or I_4308 (I75610,I75593,I75514);
DFFARX1 I_4309  ( .D(I75610), .CLK(I2350), .RSTB(I75056), .Q(I75039) );
nand I_4310 (I75048,I75593,I75319);
DFFARX1 I_4311  ( .D(I75593), .CLK(I2350), .RSTB(I75056), .Q(I75018) );
not I_4312 (I75702,I2357);
not I_4313 (I75719,I305259);
nor I_4314 (I75736,I305235,I305241);
nand I_4315 (I75753,I75736,I305244);
DFFARX1 I_4316  ( .D(I75753), .CLK(I2350), .RSTB(I75702), .Q(I75676) );
nor I_4317 (I75784,I75719,I305235);
nand I_4318 (I75801,I75784,I305253);
not I_4319 (I75691,I75801);
DFFARX1 I_4320  ( .D(I75801), .CLK(I2350), .RSTB(I75702), .Q(I75673) );
not I_4321 (I75846,I305235);
not I_4322 (I75863,I75846);
not I_4323 (I75880,I305232);
nor I_4324 (I75897,I75880,I305247);
and I_4325 (I75914,I75897,I305238);
or I_4326 (I75931,I75914,I305250);
DFFARX1 I_4327  ( .D(I75931), .CLK(I2350), .RSTB(I75702), .Q(I75948) );
nor I_4328 (I75965,I75948,I75801);
nor I_4329 (I75982,I75948,I75863);
nand I_4330 (I75688,I75753,I75982);
nand I_4331 (I76013,I75719,I305232);
nand I_4332 (I76030,I76013,I75948);
and I_4333 (I76047,I76013,I76030);
DFFARX1 I_4334  ( .D(I76047), .CLK(I2350), .RSTB(I75702), .Q(I75670) );
DFFARX1 I_4335  ( .D(I76013), .CLK(I2350), .RSTB(I75702), .Q(I76078) );
and I_4336 (I75667,I75846,I76078);
DFFARX1 I_4337  ( .D(I305262), .CLK(I2350), .RSTB(I75702), .Q(I76109) );
not I_4338 (I76126,I76109);
nor I_4339 (I76143,I75801,I76126);
and I_4340 (I76160,I76109,I76143);
nand I_4341 (I75682,I76109,I75863);
DFFARX1 I_4342  ( .D(I76109), .CLK(I2350), .RSTB(I75702), .Q(I76191) );
not I_4343 (I75679,I76191);
DFFARX1 I_4344  ( .D(I305256), .CLK(I2350), .RSTB(I75702), .Q(I76222) );
not I_4345 (I76239,I76222);
or I_4346 (I76256,I76239,I76160);
DFFARX1 I_4347  ( .D(I76256), .CLK(I2350), .RSTB(I75702), .Q(I75685) );
nand I_4348 (I75694,I76239,I75965);
DFFARX1 I_4349  ( .D(I76239), .CLK(I2350), .RSTB(I75702), .Q(I75664) );
not I_4350 (I76348,I2357);
not I_4351 (I76365,I145654);
nor I_4352 (I76382,I145651,I145639);
nand I_4353 (I76399,I76382,I145642);
DFFARX1 I_4354  ( .D(I76399), .CLK(I2350), .RSTB(I76348), .Q(I76322) );
nor I_4355 (I76430,I76365,I145651);
nand I_4356 (I76447,I76430,I145648);
not I_4357 (I76337,I76447);
DFFARX1 I_4358  ( .D(I76447), .CLK(I2350), .RSTB(I76348), .Q(I76319) );
not I_4359 (I76492,I145651);
not I_4360 (I76509,I76492);
not I_4361 (I76526,I145660);
nor I_4362 (I76543,I76526,I145636);
and I_4363 (I76560,I76543,I145657);
or I_4364 (I76577,I76560,I145645);
DFFARX1 I_4365  ( .D(I76577), .CLK(I2350), .RSTB(I76348), .Q(I76594) );
nor I_4366 (I76611,I76594,I76447);
nor I_4367 (I76628,I76594,I76509);
nand I_4368 (I76334,I76399,I76628);
nand I_4369 (I76659,I76365,I145660);
nand I_4370 (I76676,I76659,I76594);
and I_4371 (I76693,I76659,I76676);
DFFARX1 I_4372  ( .D(I76693), .CLK(I2350), .RSTB(I76348), .Q(I76316) );
DFFARX1 I_4373  ( .D(I76659), .CLK(I2350), .RSTB(I76348), .Q(I76724) );
and I_4374 (I76313,I76492,I76724);
DFFARX1 I_4375  ( .D(I145666), .CLK(I2350), .RSTB(I76348), .Q(I76755) );
not I_4376 (I76772,I76755);
nor I_4377 (I76789,I76447,I76772);
and I_4378 (I76806,I76755,I76789);
nand I_4379 (I76328,I76755,I76509);
DFFARX1 I_4380  ( .D(I76755), .CLK(I2350), .RSTB(I76348), .Q(I76837) );
not I_4381 (I76325,I76837);
DFFARX1 I_4382  ( .D(I145663), .CLK(I2350), .RSTB(I76348), .Q(I76868) );
not I_4383 (I76885,I76868);
or I_4384 (I76902,I76885,I76806);
DFFARX1 I_4385  ( .D(I76902), .CLK(I2350), .RSTB(I76348), .Q(I76331) );
nand I_4386 (I76340,I76885,I76611);
DFFARX1 I_4387  ( .D(I76885), .CLK(I2350), .RSTB(I76348), .Q(I76310) );
not I_4388 (I76994,I2357);
not I_4389 (I77011,I295739);
nor I_4390 (I77028,I295715,I295721);
nand I_4391 (I77045,I77028,I295724);
DFFARX1 I_4392  ( .D(I77045), .CLK(I2350), .RSTB(I76994), .Q(I76968) );
nor I_4393 (I77076,I77011,I295715);
nand I_4394 (I77093,I77076,I295733);
not I_4395 (I76983,I77093);
DFFARX1 I_4396  ( .D(I77093), .CLK(I2350), .RSTB(I76994), .Q(I76965) );
not I_4397 (I77138,I295715);
not I_4398 (I77155,I77138);
not I_4399 (I77172,I295712);
nor I_4400 (I77189,I77172,I295727);
and I_4401 (I77206,I77189,I295718);
or I_4402 (I77223,I77206,I295730);
DFFARX1 I_4403  ( .D(I77223), .CLK(I2350), .RSTB(I76994), .Q(I77240) );
nor I_4404 (I77257,I77240,I77093);
nor I_4405 (I77274,I77240,I77155);
nand I_4406 (I76980,I77045,I77274);
nand I_4407 (I77305,I77011,I295712);
nand I_4408 (I77322,I77305,I77240);
and I_4409 (I77339,I77305,I77322);
DFFARX1 I_4410  ( .D(I77339), .CLK(I2350), .RSTB(I76994), .Q(I76962) );
DFFARX1 I_4411  ( .D(I77305), .CLK(I2350), .RSTB(I76994), .Q(I77370) );
and I_4412 (I76959,I77138,I77370);
DFFARX1 I_4413  ( .D(I295742), .CLK(I2350), .RSTB(I76994), .Q(I77401) );
not I_4414 (I77418,I77401);
nor I_4415 (I77435,I77093,I77418);
and I_4416 (I77452,I77401,I77435);
nand I_4417 (I76974,I77401,I77155);
DFFARX1 I_4418  ( .D(I77401), .CLK(I2350), .RSTB(I76994), .Q(I77483) );
not I_4419 (I76971,I77483);
DFFARX1 I_4420  ( .D(I295736), .CLK(I2350), .RSTB(I76994), .Q(I77514) );
not I_4421 (I77531,I77514);
or I_4422 (I77548,I77531,I77452);
DFFARX1 I_4423  ( .D(I77548), .CLK(I2350), .RSTB(I76994), .Q(I76977) );
nand I_4424 (I76986,I77531,I77257);
DFFARX1 I_4425  ( .D(I77531), .CLK(I2350), .RSTB(I76994), .Q(I76956) );
not I_4426 (I77640,I2357);
not I_4427 (I77657,I18071);
nor I_4428 (I77674,I18083,I18068);
nand I_4429 (I77691,I77674,I18080);
DFFARX1 I_4430  ( .D(I77691), .CLK(I2350), .RSTB(I77640), .Q(I77614) );
nor I_4431 (I77722,I77657,I18083);
nand I_4432 (I77739,I77722,I18098);
not I_4433 (I77629,I77739);
DFFARX1 I_4434  ( .D(I77739), .CLK(I2350), .RSTB(I77640), .Q(I77611) );
not I_4435 (I77784,I18083);
not I_4436 (I77801,I77784);
not I_4437 (I77818,I18074);
nor I_4438 (I77835,I77818,I18086);
and I_4439 (I77852,I77835,I18077);
or I_4440 (I77869,I77852,I18092);
DFFARX1 I_4441  ( .D(I77869), .CLK(I2350), .RSTB(I77640), .Q(I77886) );
nor I_4442 (I77903,I77886,I77739);
nor I_4443 (I77920,I77886,I77801);
nand I_4444 (I77626,I77691,I77920);
nand I_4445 (I77951,I77657,I18074);
nand I_4446 (I77968,I77951,I77886);
and I_4447 (I77985,I77951,I77968);
DFFARX1 I_4448  ( .D(I77985), .CLK(I2350), .RSTB(I77640), .Q(I77608) );
DFFARX1 I_4449  ( .D(I77951), .CLK(I2350), .RSTB(I77640), .Q(I78016) );
and I_4450 (I77605,I77784,I78016);
DFFARX1 I_4451  ( .D(I18095), .CLK(I2350), .RSTB(I77640), .Q(I78047) );
not I_4452 (I78064,I78047);
nor I_4453 (I78081,I77739,I78064);
and I_4454 (I78098,I78047,I78081);
nand I_4455 (I77620,I78047,I77801);
DFFARX1 I_4456  ( .D(I78047), .CLK(I2350), .RSTB(I77640), .Q(I78129) );
not I_4457 (I77617,I78129);
DFFARX1 I_4458  ( .D(I18089), .CLK(I2350), .RSTB(I77640), .Q(I78160) );
not I_4459 (I78177,I78160);
or I_4460 (I78194,I78177,I78098);
DFFARX1 I_4461  ( .D(I78194), .CLK(I2350), .RSTB(I77640), .Q(I77623) );
nand I_4462 (I77632,I78177,I77903);
DFFARX1 I_4463  ( .D(I78177), .CLK(I2350), .RSTB(I77640), .Q(I77602) );
not I_4464 (I78286,I2357);
not I_4465 (I78303,I1527);
nor I_4466 (I78320,I1415,I1887);
nand I_4467 (I78337,I78320,I2327);
DFFARX1 I_4468  ( .D(I78337), .CLK(I2350), .RSTB(I78286), .Q(I78260) );
nor I_4469 (I78368,I78303,I1415);
nand I_4470 (I78385,I78368,I2023);
not I_4471 (I78275,I78385);
DFFARX1 I_4472  ( .D(I78385), .CLK(I2350), .RSTB(I78286), .Q(I78257) );
not I_4473 (I78430,I1415);
not I_4474 (I78447,I78430);
not I_4475 (I78464,I1983);
nor I_4476 (I78481,I78464,I1791);
and I_4477 (I78498,I78481,I1663);
or I_4478 (I78515,I78498,I1511);
DFFARX1 I_4479  ( .D(I78515), .CLK(I2350), .RSTB(I78286), .Q(I78532) );
nor I_4480 (I78549,I78532,I78385);
nor I_4481 (I78566,I78532,I78447);
nand I_4482 (I78272,I78337,I78566);
nand I_4483 (I78597,I78303,I1983);
nand I_4484 (I78614,I78597,I78532);
and I_4485 (I78631,I78597,I78614);
DFFARX1 I_4486  ( .D(I78631), .CLK(I2350), .RSTB(I78286), .Q(I78254) );
DFFARX1 I_4487  ( .D(I78597), .CLK(I2350), .RSTB(I78286), .Q(I78662) );
and I_4488 (I78251,I78430,I78662);
DFFARX1 I_4489  ( .D(I1927), .CLK(I2350), .RSTB(I78286), .Q(I78693) );
not I_4490 (I78710,I78693);
nor I_4491 (I78727,I78385,I78710);
and I_4492 (I78744,I78693,I78727);
nand I_4493 (I78266,I78693,I78447);
DFFARX1 I_4494  ( .D(I78693), .CLK(I2350), .RSTB(I78286), .Q(I78775) );
not I_4495 (I78263,I78775);
DFFARX1 I_4496  ( .D(I2191), .CLK(I2350), .RSTB(I78286), .Q(I78806) );
not I_4497 (I78823,I78806);
or I_4498 (I78840,I78823,I78744);
DFFARX1 I_4499  ( .D(I78840), .CLK(I2350), .RSTB(I78286), .Q(I78269) );
nand I_4500 (I78278,I78823,I78549);
DFFARX1 I_4501  ( .D(I78823), .CLK(I2350), .RSTB(I78286), .Q(I78248) );
not I_4502 (I78932,I2357);
not I_4503 (I78949,I122210);
nor I_4504 (I78966,I122240,I122219);
nand I_4505 (I78983,I78966,I122231);
DFFARX1 I_4506  ( .D(I78983), .CLK(I2350), .RSTB(I78932), .Q(I78906) );
nor I_4507 (I79014,I78949,I122240);
nand I_4508 (I79031,I79014,I122213);
not I_4509 (I78921,I79031);
DFFARX1 I_4510  ( .D(I79031), .CLK(I2350), .RSTB(I78932), .Q(I78903) );
not I_4511 (I79076,I122240);
not I_4512 (I79093,I79076);
not I_4513 (I79110,I122216);
nor I_4514 (I79127,I79110,I122234);
and I_4515 (I79144,I79127,I122225);
or I_4516 (I79161,I79144,I122222);
DFFARX1 I_4517  ( .D(I79161), .CLK(I2350), .RSTB(I78932), .Q(I79178) );
nor I_4518 (I79195,I79178,I79031);
nor I_4519 (I79212,I79178,I79093);
nand I_4520 (I78918,I78983,I79212);
nand I_4521 (I79243,I78949,I122216);
nand I_4522 (I79260,I79243,I79178);
and I_4523 (I79277,I79243,I79260);
DFFARX1 I_4524  ( .D(I79277), .CLK(I2350), .RSTB(I78932), .Q(I78900) );
DFFARX1 I_4525  ( .D(I79243), .CLK(I2350), .RSTB(I78932), .Q(I79308) );
and I_4526 (I78897,I79076,I79308);
DFFARX1 I_4527  ( .D(I122228), .CLK(I2350), .RSTB(I78932), .Q(I79339) );
not I_4528 (I79356,I79339);
nor I_4529 (I79373,I79031,I79356);
and I_4530 (I79390,I79339,I79373);
nand I_4531 (I78912,I79339,I79093);
DFFARX1 I_4532  ( .D(I79339), .CLK(I2350), .RSTB(I78932), .Q(I79421) );
not I_4533 (I78909,I79421);
DFFARX1 I_4534  ( .D(I122237), .CLK(I2350), .RSTB(I78932), .Q(I79452) );
not I_4535 (I79469,I79452);
or I_4536 (I79486,I79469,I79390);
DFFARX1 I_4537  ( .D(I79486), .CLK(I2350), .RSTB(I78932), .Q(I78915) );
nand I_4538 (I78924,I79469,I79195);
DFFARX1 I_4539  ( .D(I79469), .CLK(I2350), .RSTB(I78932), .Q(I78894) );
not I_4540 (I79578,I2357);
not I_4541 (I79595,I194665);
nor I_4542 (I79612,I194677,I194659);
nand I_4543 (I79629,I79612,I194674);
DFFARX1 I_4544  ( .D(I79629), .CLK(I2350), .RSTB(I79578), .Q(I79552) );
nor I_4545 (I79660,I79595,I194677);
nand I_4546 (I79677,I79660,I194662);
not I_4547 (I79567,I79677);
DFFARX1 I_4548  ( .D(I79677), .CLK(I2350), .RSTB(I79578), .Q(I79549) );
not I_4549 (I79722,I194677);
not I_4550 (I79739,I79722);
not I_4551 (I79756,I194671);
nor I_4552 (I79773,I79756,I194650);
and I_4553 (I79790,I79773,I194653);
or I_4554 (I79807,I79790,I194656);
DFFARX1 I_4555  ( .D(I79807), .CLK(I2350), .RSTB(I79578), .Q(I79824) );
nor I_4556 (I79841,I79824,I79677);
nor I_4557 (I79858,I79824,I79739);
nand I_4558 (I79564,I79629,I79858);
nand I_4559 (I79889,I79595,I194671);
nand I_4560 (I79906,I79889,I79824);
and I_4561 (I79923,I79889,I79906);
DFFARX1 I_4562  ( .D(I79923), .CLK(I2350), .RSTB(I79578), .Q(I79546) );
DFFARX1 I_4563  ( .D(I79889), .CLK(I2350), .RSTB(I79578), .Q(I79954) );
and I_4564 (I79543,I79722,I79954);
DFFARX1 I_4565  ( .D(I194647), .CLK(I2350), .RSTB(I79578), .Q(I79985) );
not I_4566 (I80002,I79985);
nor I_4567 (I80019,I79677,I80002);
and I_4568 (I80036,I79985,I80019);
nand I_4569 (I79558,I79985,I79739);
DFFARX1 I_4570  ( .D(I79985), .CLK(I2350), .RSTB(I79578), .Q(I80067) );
not I_4571 (I79555,I80067);
DFFARX1 I_4572  ( .D(I194668), .CLK(I2350), .RSTB(I79578), .Q(I80098) );
not I_4573 (I80115,I80098);
or I_4574 (I80132,I80115,I80036);
DFFARX1 I_4575  ( .D(I80132), .CLK(I2350), .RSTB(I79578), .Q(I79561) );
nand I_4576 (I79570,I80115,I79841);
DFFARX1 I_4577  ( .D(I80115), .CLK(I2350), .RSTB(I79578), .Q(I79540) );
not I_4578 (I80224,I2357);
not I_4579 (I80241,I258548);
nor I_4580 (I80258,I258536,I258542);
nand I_4581 (I80275,I80258,I258533);
DFFARX1 I_4582  ( .D(I80275), .CLK(I2350), .RSTB(I80224), .Q(I80198) );
nor I_4583 (I80306,I80241,I258536);
nand I_4584 (I80323,I80306,I258539);
not I_4585 (I80213,I80323);
DFFARX1 I_4586  ( .D(I80323), .CLK(I2350), .RSTB(I80224), .Q(I80195) );
not I_4587 (I80368,I258536);
not I_4588 (I80385,I80368);
not I_4589 (I80402,I258551);
nor I_4590 (I80419,I80402,I258563);
and I_4591 (I80436,I80419,I258545);
or I_4592 (I80453,I80436,I258560);
DFFARX1 I_4593  ( .D(I80453), .CLK(I2350), .RSTB(I80224), .Q(I80470) );
nor I_4594 (I80487,I80470,I80323);
nor I_4595 (I80504,I80470,I80385);
nand I_4596 (I80210,I80275,I80504);
nand I_4597 (I80535,I80241,I258551);
nand I_4598 (I80552,I80535,I80470);
and I_4599 (I80569,I80535,I80552);
DFFARX1 I_4600  ( .D(I80569), .CLK(I2350), .RSTB(I80224), .Q(I80192) );
DFFARX1 I_4601  ( .D(I80535), .CLK(I2350), .RSTB(I80224), .Q(I80600) );
and I_4602 (I80189,I80368,I80600);
DFFARX1 I_4603  ( .D(I258554), .CLK(I2350), .RSTB(I80224), .Q(I80631) );
not I_4604 (I80648,I80631);
nor I_4605 (I80665,I80323,I80648);
and I_4606 (I80682,I80631,I80665);
nand I_4607 (I80204,I80631,I80385);
DFFARX1 I_4608  ( .D(I80631), .CLK(I2350), .RSTB(I80224), .Q(I80713) );
not I_4609 (I80201,I80713);
DFFARX1 I_4610  ( .D(I258557), .CLK(I2350), .RSTB(I80224), .Q(I80744) );
not I_4611 (I80761,I80744);
or I_4612 (I80778,I80761,I80682);
DFFARX1 I_4613  ( .D(I80778), .CLK(I2350), .RSTB(I80224), .Q(I80207) );
nand I_4614 (I80216,I80761,I80487);
DFFARX1 I_4615  ( .D(I80761), .CLK(I2350), .RSTB(I80224), .Q(I80186) );
not I_4616 (I80870,I2357);
not I_4617 (I80887,I299309);
nor I_4618 (I80904,I299285,I299291);
nand I_4619 (I80921,I80904,I299294);
DFFARX1 I_4620  ( .D(I80921), .CLK(I2350), .RSTB(I80870), .Q(I80844) );
nor I_4621 (I80952,I80887,I299285);
nand I_4622 (I80969,I80952,I299303);
not I_4623 (I80859,I80969);
DFFARX1 I_4624  ( .D(I80969), .CLK(I2350), .RSTB(I80870), .Q(I80841) );
not I_4625 (I81014,I299285);
not I_4626 (I81031,I81014);
not I_4627 (I81048,I299282);
nor I_4628 (I81065,I81048,I299297);
and I_4629 (I81082,I81065,I299288);
or I_4630 (I81099,I81082,I299300);
DFFARX1 I_4631  ( .D(I81099), .CLK(I2350), .RSTB(I80870), .Q(I81116) );
nor I_4632 (I81133,I81116,I80969);
nor I_4633 (I81150,I81116,I81031);
nand I_4634 (I80856,I80921,I81150);
nand I_4635 (I81181,I80887,I299282);
nand I_4636 (I81198,I81181,I81116);
and I_4637 (I81215,I81181,I81198);
DFFARX1 I_4638  ( .D(I81215), .CLK(I2350), .RSTB(I80870), .Q(I80838) );
DFFARX1 I_4639  ( .D(I81181), .CLK(I2350), .RSTB(I80870), .Q(I81246) );
and I_4640 (I80835,I81014,I81246);
DFFARX1 I_4641  ( .D(I299312), .CLK(I2350), .RSTB(I80870), .Q(I81277) );
not I_4642 (I81294,I81277);
nor I_4643 (I81311,I80969,I81294);
and I_4644 (I81328,I81277,I81311);
nand I_4645 (I80850,I81277,I81031);
DFFARX1 I_4646  ( .D(I81277), .CLK(I2350), .RSTB(I80870), .Q(I81359) );
not I_4647 (I80847,I81359);
DFFARX1 I_4648  ( .D(I299306), .CLK(I2350), .RSTB(I80870), .Q(I81390) );
not I_4649 (I81407,I81390);
or I_4650 (I81424,I81407,I81328);
DFFARX1 I_4651  ( .D(I81424), .CLK(I2350), .RSTB(I80870), .Q(I80853) );
nand I_4652 (I80862,I81407,I81133);
DFFARX1 I_4653  ( .D(I81407), .CLK(I2350), .RSTB(I80870), .Q(I80832) );
not I_4654 (I81516,I2357);
not I_4655 (I81533,I146317);
nor I_4656 (I81550,I146314,I146302);
nand I_4657 (I81567,I81550,I146305);
DFFARX1 I_4658  ( .D(I81567), .CLK(I2350), .RSTB(I81516), .Q(I81490) );
nor I_4659 (I81598,I81533,I146314);
nand I_4660 (I81615,I81598,I146311);
not I_4661 (I81505,I81615);
DFFARX1 I_4662  ( .D(I81615), .CLK(I2350), .RSTB(I81516), .Q(I81487) );
not I_4663 (I81660,I146314);
not I_4664 (I81677,I81660);
not I_4665 (I81694,I146323);
nor I_4666 (I81711,I81694,I146299);
and I_4667 (I81728,I81711,I146320);
or I_4668 (I81745,I81728,I146308);
DFFARX1 I_4669  ( .D(I81745), .CLK(I2350), .RSTB(I81516), .Q(I81762) );
nor I_4670 (I81779,I81762,I81615);
nor I_4671 (I81796,I81762,I81677);
nand I_4672 (I81502,I81567,I81796);
nand I_4673 (I81827,I81533,I146323);
nand I_4674 (I81844,I81827,I81762);
and I_4675 (I81861,I81827,I81844);
DFFARX1 I_4676  ( .D(I81861), .CLK(I2350), .RSTB(I81516), .Q(I81484) );
DFFARX1 I_4677  ( .D(I81827), .CLK(I2350), .RSTB(I81516), .Q(I81892) );
and I_4678 (I81481,I81660,I81892);
DFFARX1 I_4679  ( .D(I146329), .CLK(I2350), .RSTB(I81516), .Q(I81923) );
not I_4680 (I81940,I81923);
nor I_4681 (I81957,I81615,I81940);
and I_4682 (I81974,I81923,I81957);
nand I_4683 (I81496,I81923,I81677);
DFFARX1 I_4684  ( .D(I81923), .CLK(I2350), .RSTB(I81516), .Q(I82005) );
not I_4685 (I81493,I82005);
DFFARX1 I_4686  ( .D(I146326), .CLK(I2350), .RSTB(I81516), .Q(I82036) );
not I_4687 (I82053,I82036);
or I_4688 (I82070,I82053,I81974);
DFFARX1 I_4689  ( .D(I82070), .CLK(I2350), .RSTB(I81516), .Q(I81499) );
nand I_4690 (I81508,I82053,I81779);
DFFARX1 I_4691  ( .D(I82053), .CLK(I2350), .RSTB(I81516), .Q(I81478) );
not I_4692 (I82162,I2357);
not I_4693 (I82179,I312994);
nor I_4694 (I82196,I312970,I312976);
nand I_4695 (I82213,I82196,I312979);
DFFARX1 I_4696  ( .D(I82213), .CLK(I2350), .RSTB(I82162), .Q(I82136) );
nor I_4697 (I82244,I82179,I312970);
nand I_4698 (I82261,I82244,I312988);
not I_4699 (I82151,I82261);
DFFARX1 I_4700  ( .D(I82261), .CLK(I2350), .RSTB(I82162), .Q(I82133) );
not I_4701 (I82306,I312970);
not I_4702 (I82323,I82306);
not I_4703 (I82340,I312967);
nor I_4704 (I82357,I82340,I312982);
and I_4705 (I82374,I82357,I312973);
or I_4706 (I82391,I82374,I312985);
DFFARX1 I_4707  ( .D(I82391), .CLK(I2350), .RSTB(I82162), .Q(I82408) );
nor I_4708 (I82425,I82408,I82261);
nor I_4709 (I82442,I82408,I82323);
nand I_4710 (I82148,I82213,I82442);
nand I_4711 (I82473,I82179,I312967);
nand I_4712 (I82490,I82473,I82408);
and I_4713 (I82507,I82473,I82490);
DFFARX1 I_4714  ( .D(I82507), .CLK(I2350), .RSTB(I82162), .Q(I82130) );
DFFARX1 I_4715  ( .D(I82473), .CLK(I2350), .RSTB(I82162), .Q(I82538) );
and I_4716 (I82127,I82306,I82538);
DFFARX1 I_4717  ( .D(I312997), .CLK(I2350), .RSTB(I82162), .Q(I82569) );
not I_4718 (I82586,I82569);
nor I_4719 (I82603,I82261,I82586);
and I_4720 (I82620,I82569,I82603);
nand I_4721 (I82142,I82569,I82323);
DFFARX1 I_4722  ( .D(I82569), .CLK(I2350), .RSTB(I82162), .Q(I82651) );
not I_4723 (I82139,I82651);
DFFARX1 I_4724  ( .D(I312991), .CLK(I2350), .RSTB(I82162), .Q(I82682) );
not I_4725 (I82699,I82682);
or I_4726 (I82716,I82699,I82620);
DFFARX1 I_4727  ( .D(I82716), .CLK(I2350), .RSTB(I82162), .Q(I82145) );
nand I_4728 (I82154,I82699,I82425);
DFFARX1 I_4729  ( .D(I82699), .CLK(I2350), .RSTB(I82162), .Q(I82124) );
not I_4730 (I82808,I2357);
not I_4731 (I82825,I214691);
nor I_4732 (I82842,I214703,I214685);
nand I_4733 (I82859,I82842,I214700);
DFFARX1 I_4734  ( .D(I82859), .CLK(I2350), .RSTB(I82808), .Q(I82782) );
nor I_4735 (I82890,I82825,I214703);
nand I_4736 (I82907,I82890,I214688);
not I_4737 (I82797,I82907);
DFFARX1 I_4738  ( .D(I82907), .CLK(I2350), .RSTB(I82808), .Q(I82779) );
not I_4739 (I82952,I214703);
not I_4740 (I82969,I82952);
not I_4741 (I82986,I214697);
nor I_4742 (I83003,I82986,I214676);
and I_4743 (I83020,I83003,I214679);
or I_4744 (I83037,I83020,I214682);
DFFARX1 I_4745  ( .D(I83037), .CLK(I2350), .RSTB(I82808), .Q(I83054) );
nor I_4746 (I83071,I83054,I82907);
nor I_4747 (I83088,I83054,I82969);
nand I_4748 (I82794,I82859,I83088);
nand I_4749 (I83119,I82825,I214697);
nand I_4750 (I83136,I83119,I83054);
and I_4751 (I83153,I83119,I83136);
DFFARX1 I_4752  ( .D(I83153), .CLK(I2350), .RSTB(I82808), .Q(I82776) );
DFFARX1 I_4753  ( .D(I83119), .CLK(I2350), .RSTB(I82808), .Q(I83184) );
and I_4754 (I82773,I82952,I83184);
DFFARX1 I_4755  ( .D(I214673), .CLK(I2350), .RSTB(I82808), .Q(I83215) );
not I_4756 (I83232,I83215);
nor I_4757 (I83249,I82907,I83232);
and I_4758 (I83266,I83215,I83249);
nand I_4759 (I82788,I83215,I82969);
DFFARX1 I_4760  ( .D(I83215), .CLK(I2350), .RSTB(I82808), .Q(I83297) );
not I_4761 (I82785,I83297);
DFFARX1 I_4762  ( .D(I214694), .CLK(I2350), .RSTB(I82808), .Q(I83328) );
not I_4763 (I83345,I83328);
or I_4764 (I83362,I83345,I83266);
DFFARX1 I_4765  ( .D(I83362), .CLK(I2350), .RSTB(I82808), .Q(I82791) );
nand I_4766 (I82800,I83345,I83071);
DFFARX1 I_4767  ( .D(I83345), .CLK(I2350), .RSTB(I82808), .Q(I82770) );
not I_4768 (I83454,I2357);
not I_4769 (I83471,I323097);
nor I_4770 (I83488,I323082,I323109);
nand I_4771 (I83505,I83488,I323085);
DFFARX1 I_4772  ( .D(I83505), .CLK(I2350), .RSTB(I83454), .Q(I83428) );
nor I_4773 (I83536,I83471,I323082);
nand I_4774 (I83553,I83536,I323100);
not I_4775 (I83443,I83553);
DFFARX1 I_4776  ( .D(I83553), .CLK(I2350), .RSTB(I83454), .Q(I83425) );
not I_4777 (I83598,I323082);
not I_4778 (I83615,I83598);
not I_4779 (I83632,I323112);
nor I_4780 (I83649,I83632,I323094);
and I_4781 (I83666,I83649,I323103);
or I_4782 (I83683,I83666,I323088);
DFFARX1 I_4783  ( .D(I83683), .CLK(I2350), .RSTB(I83454), .Q(I83700) );
nor I_4784 (I83717,I83700,I83553);
nor I_4785 (I83734,I83700,I83615);
nand I_4786 (I83440,I83505,I83734);
nand I_4787 (I83765,I83471,I323112);
nand I_4788 (I83782,I83765,I83700);
and I_4789 (I83799,I83765,I83782);
DFFARX1 I_4790  ( .D(I83799), .CLK(I2350), .RSTB(I83454), .Q(I83422) );
DFFARX1 I_4791  ( .D(I83765), .CLK(I2350), .RSTB(I83454), .Q(I83830) );
and I_4792 (I83419,I83598,I83830);
DFFARX1 I_4793  ( .D(I323091), .CLK(I2350), .RSTB(I83454), .Q(I83861) );
not I_4794 (I83878,I83861);
nor I_4795 (I83895,I83553,I83878);
and I_4796 (I83912,I83861,I83895);
nand I_4797 (I83434,I83861,I83615);
DFFARX1 I_4798  ( .D(I83861), .CLK(I2350), .RSTB(I83454), .Q(I83943) );
not I_4799 (I83431,I83943);
DFFARX1 I_4800  ( .D(I323106), .CLK(I2350), .RSTB(I83454), .Q(I83974) );
not I_4801 (I83991,I83974);
or I_4802 (I84008,I83991,I83912);
DFFARX1 I_4803  ( .D(I84008), .CLK(I2350), .RSTB(I83454), .Q(I83437) );
nand I_4804 (I83446,I83991,I83717);
DFFARX1 I_4805  ( .D(I83991), .CLK(I2350), .RSTB(I83454), .Q(I83416) );
not I_4806 (I84100,I2357);
not I_4807 (I84117,I186760);
nor I_4808 (I84134,I186757,I186745);
nand I_4809 (I84151,I84134,I186748);
DFFARX1 I_4810  ( .D(I84151), .CLK(I2350), .RSTB(I84100), .Q(I84074) );
nor I_4811 (I84182,I84117,I186757);
nand I_4812 (I84199,I84182,I186754);
not I_4813 (I84089,I84199);
DFFARX1 I_4814  ( .D(I84199), .CLK(I2350), .RSTB(I84100), .Q(I84071) );
not I_4815 (I84244,I186757);
not I_4816 (I84261,I84244);
not I_4817 (I84278,I186766);
nor I_4818 (I84295,I84278,I186742);
and I_4819 (I84312,I84295,I186763);
or I_4820 (I84329,I84312,I186751);
DFFARX1 I_4821  ( .D(I84329), .CLK(I2350), .RSTB(I84100), .Q(I84346) );
nor I_4822 (I84363,I84346,I84199);
nor I_4823 (I84380,I84346,I84261);
nand I_4824 (I84086,I84151,I84380);
nand I_4825 (I84411,I84117,I186766);
nand I_4826 (I84428,I84411,I84346);
and I_4827 (I84445,I84411,I84428);
DFFARX1 I_4828  ( .D(I84445), .CLK(I2350), .RSTB(I84100), .Q(I84068) );
DFFARX1 I_4829  ( .D(I84411), .CLK(I2350), .RSTB(I84100), .Q(I84476) );
and I_4830 (I84065,I84244,I84476);
DFFARX1 I_4831  ( .D(I186772), .CLK(I2350), .RSTB(I84100), .Q(I84507) );
not I_4832 (I84524,I84507);
nor I_4833 (I84541,I84199,I84524);
and I_4834 (I84558,I84507,I84541);
nand I_4835 (I84080,I84507,I84261);
DFFARX1 I_4836  ( .D(I84507), .CLK(I2350), .RSTB(I84100), .Q(I84589) );
not I_4837 (I84077,I84589);
DFFARX1 I_4838  ( .D(I186769), .CLK(I2350), .RSTB(I84100), .Q(I84620) );
not I_4839 (I84637,I84620);
or I_4840 (I84654,I84637,I84558);
DFFARX1 I_4841  ( .D(I84654), .CLK(I2350), .RSTB(I84100), .Q(I84083) );
nand I_4842 (I84092,I84637,I84363);
DFFARX1 I_4843  ( .D(I84637), .CLK(I2350), .RSTB(I84100), .Q(I84062) );
not I_4844 (I84746,I2357);
not I_4845 (I84763,I345823);
nor I_4846 (I84780,I345829,I345841);
nand I_4847 (I84797,I84780,I345832);
DFFARX1 I_4848  ( .D(I84797), .CLK(I2350), .RSTB(I84746), .Q(I84717) );
nor I_4849 (I84828,I84763,I345829);
nand I_4850 (I84845,I84828,I345811);
nand I_4851 (I84862,I84845,I84797);
not I_4852 (I84879,I345829);
not I_4853 (I84896,I345826);
nor I_4854 (I84913,I84896,I345814);
and I_4855 (I84930,I84913,I345835);
or I_4856 (I84947,I84930,I345817);
DFFARX1 I_4857  ( .D(I84947), .CLK(I2350), .RSTB(I84746), .Q(I84964) );
nor I_4858 (I84981,I84964,I84845);
nand I_4859 (I84732,I84879,I84981);
not I_4860 (I84729,I84964);
and I_4861 (I85026,I84964,I84862);
DFFARX1 I_4862  ( .D(I85026), .CLK(I2350), .RSTB(I84746), .Q(I84714) );
DFFARX1 I_4863  ( .D(I84964), .CLK(I2350), .RSTB(I84746), .Q(I85057) );
and I_4864 (I84711,I84879,I85057);
nand I_4865 (I85088,I84763,I345826);
not I_4866 (I85105,I85088);
nor I_4867 (I85122,I84964,I85105);
DFFARX1 I_4868  ( .D(I345838), .CLK(I2350), .RSTB(I84746), .Q(I85139) );
nand I_4869 (I85156,I85139,I85088);
and I_4870 (I85173,I84879,I85156);
DFFARX1 I_4871  ( .D(I85173), .CLK(I2350), .RSTB(I84746), .Q(I84738) );
not I_4872 (I85204,I85139);
nand I_4873 (I84726,I85139,I85122);
nand I_4874 (I84720,I85139,I85105);
DFFARX1 I_4875  ( .D(I345820), .CLK(I2350), .RSTB(I84746), .Q(I85249) );
not I_4876 (I85266,I85249);
nor I_4877 (I84735,I85139,I85266);
nor I_4878 (I85297,I85266,I85204);
and I_4879 (I85314,I84845,I85297);
or I_4880 (I85331,I85088,I85314);
DFFARX1 I_4881  ( .D(I85331), .CLK(I2350), .RSTB(I84746), .Q(I84723) );
DFFARX1 I_4882  ( .D(I85266), .CLK(I2350), .RSTB(I84746), .Q(I84708) );
not I_4883 (I85409,I2357);
not I_4884 (I85426,I165526);
nor I_4885 (I85443,I165535,I165547);
nand I_4886 (I85460,I85443,I165538);
DFFARX1 I_4887  ( .D(I85460), .CLK(I2350), .RSTB(I85409), .Q(I85380) );
nor I_4888 (I85491,I85426,I165535);
nand I_4889 (I85508,I85491,I165550);
nand I_4890 (I85525,I85508,I85460);
not I_4891 (I85542,I165535);
not I_4892 (I85559,I165556);
nor I_4893 (I85576,I85559,I165532);
and I_4894 (I85593,I85576,I165541);
or I_4895 (I85610,I85593,I165529);
DFFARX1 I_4896  ( .D(I85610), .CLK(I2350), .RSTB(I85409), .Q(I85627) );
nor I_4897 (I85644,I85627,I85508);
nand I_4898 (I85395,I85542,I85644);
not I_4899 (I85392,I85627);
and I_4900 (I85689,I85627,I85525);
DFFARX1 I_4901  ( .D(I85689), .CLK(I2350), .RSTB(I85409), .Q(I85377) );
DFFARX1 I_4902  ( .D(I85627), .CLK(I2350), .RSTB(I85409), .Q(I85720) );
and I_4903 (I85374,I85542,I85720);
nand I_4904 (I85751,I85426,I165556);
not I_4905 (I85768,I85751);
nor I_4906 (I85785,I85627,I85768);
DFFARX1 I_4907  ( .D(I165553), .CLK(I2350), .RSTB(I85409), .Q(I85802) );
nand I_4908 (I85819,I85802,I85751);
and I_4909 (I85836,I85542,I85819);
DFFARX1 I_4910  ( .D(I85836), .CLK(I2350), .RSTB(I85409), .Q(I85401) );
not I_4911 (I85867,I85802);
nand I_4912 (I85389,I85802,I85785);
nand I_4913 (I85383,I85802,I85768);
DFFARX1 I_4914  ( .D(I165544), .CLK(I2350), .RSTB(I85409), .Q(I85912) );
not I_4915 (I85929,I85912);
nor I_4916 (I85398,I85802,I85929);
nor I_4917 (I85960,I85929,I85867);
and I_4918 (I85977,I85508,I85960);
or I_4919 (I85994,I85751,I85977);
DFFARX1 I_4920  ( .D(I85994), .CLK(I2350), .RSTB(I85409), .Q(I85386) );
DFFARX1 I_4921  ( .D(I85929), .CLK(I2350), .RSTB(I85409), .Q(I85371) );
not I_4922 (I86072,I2357);
not I_4923 (I86089,I190720);
nor I_4924 (I86106,I190729,I190741);
nand I_4925 (I86123,I86106,I190732);
DFFARX1 I_4926  ( .D(I86123), .CLK(I2350), .RSTB(I86072), .Q(I86043) );
nor I_4927 (I86154,I86089,I190729);
nand I_4928 (I86171,I86154,I190744);
nand I_4929 (I86188,I86171,I86123);
not I_4930 (I86205,I190729);
not I_4931 (I86222,I190750);
nor I_4932 (I86239,I86222,I190726);
and I_4933 (I86256,I86239,I190735);
or I_4934 (I86273,I86256,I190723);
DFFARX1 I_4935  ( .D(I86273), .CLK(I2350), .RSTB(I86072), .Q(I86290) );
nor I_4936 (I86307,I86290,I86171);
nand I_4937 (I86058,I86205,I86307);
not I_4938 (I86055,I86290);
and I_4939 (I86352,I86290,I86188);
DFFARX1 I_4940  ( .D(I86352), .CLK(I2350), .RSTB(I86072), .Q(I86040) );
DFFARX1 I_4941  ( .D(I86290), .CLK(I2350), .RSTB(I86072), .Q(I86383) );
and I_4942 (I86037,I86205,I86383);
nand I_4943 (I86414,I86089,I190750);
not I_4944 (I86431,I86414);
nor I_4945 (I86448,I86290,I86431);
DFFARX1 I_4946  ( .D(I190747), .CLK(I2350), .RSTB(I86072), .Q(I86465) );
nand I_4947 (I86482,I86465,I86414);
and I_4948 (I86499,I86205,I86482);
DFFARX1 I_4949  ( .D(I86499), .CLK(I2350), .RSTB(I86072), .Q(I86064) );
not I_4950 (I86530,I86465);
nand I_4951 (I86052,I86465,I86448);
nand I_4952 (I86046,I86465,I86431);
DFFARX1 I_4953  ( .D(I190738), .CLK(I2350), .RSTB(I86072), .Q(I86575) );
not I_4954 (I86592,I86575);
nor I_4955 (I86061,I86465,I86592);
nor I_4956 (I86623,I86592,I86530);
and I_4957 (I86640,I86171,I86623);
or I_4958 (I86657,I86414,I86640);
DFFARX1 I_4959  ( .D(I86657), .CLK(I2350), .RSTB(I86072), .Q(I86049) );
DFFARX1 I_4960  ( .D(I86592), .CLK(I2350), .RSTB(I86072), .Q(I86034) );
not I_4961 (I86735,I2357);
not I_4962 (I86752,I199187);
nor I_4963 (I86769,I199196,I199169);
nand I_4964 (I86786,I86769,I199181);
DFFARX1 I_4965  ( .D(I86786), .CLK(I2350), .RSTB(I86735), .Q(I86706) );
nor I_4966 (I86817,I86752,I199196);
nand I_4967 (I86834,I86817,I199193);
nand I_4968 (I86851,I86834,I86786);
not I_4969 (I86868,I199196);
not I_4970 (I86885,I199172);
nor I_4971 (I86902,I86885,I199178);
and I_4972 (I86919,I86902,I199190);
or I_4973 (I86936,I86919,I199175);
DFFARX1 I_4974  ( .D(I86936), .CLK(I2350), .RSTB(I86735), .Q(I86953) );
nor I_4975 (I86970,I86953,I86834);
nand I_4976 (I86721,I86868,I86970);
not I_4977 (I86718,I86953);
and I_4978 (I87015,I86953,I86851);
DFFARX1 I_4979  ( .D(I87015), .CLK(I2350), .RSTB(I86735), .Q(I86703) );
DFFARX1 I_4980  ( .D(I86953), .CLK(I2350), .RSTB(I86735), .Q(I87046) );
and I_4981 (I86700,I86868,I87046);
nand I_4982 (I87077,I86752,I199172);
not I_4983 (I87094,I87077);
nor I_4984 (I87111,I86953,I87094);
DFFARX1 I_4985  ( .D(I199199), .CLK(I2350), .RSTB(I86735), .Q(I87128) );
nand I_4986 (I87145,I87128,I87077);
and I_4987 (I87162,I86868,I87145);
DFFARX1 I_4988  ( .D(I87162), .CLK(I2350), .RSTB(I86735), .Q(I86727) );
not I_4989 (I87193,I87128);
nand I_4990 (I86715,I87128,I87111);
nand I_4991 (I86709,I87128,I87094);
DFFARX1 I_4992  ( .D(I199184), .CLK(I2350), .RSTB(I86735), .Q(I87238) );
not I_4993 (I87255,I87238);
nor I_4994 (I86724,I87128,I87255);
nor I_4995 (I87286,I87255,I87193);
and I_4996 (I87303,I86834,I87286);
or I_4997 (I87320,I87077,I87303);
DFFARX1 I_4998  ( .D(I87320), .CLK(I2350), .RSTB(I86735), .Q(I86712) );
DFFARX1 I_4999  ( .D(I87255), .CLK(I2350), .RSTB(I86735), .Q(I86697) );
not I_5000 (I87398,I2357);
not I_5001 (I87415,I230195);
nor I_5002 (I87432,I230204,I230177);
nand I_5003 (I87449,I87432,I230189);
DFFARX1 I_5004  ( .D(I87449), .CLK(I2350), .RSTB(I87398), .Q(I87369) );
nor I_5005 (I87480,I87415,I230204);
nand I_5006 (I87497,I87480,I230201);
nand I_5007 (I87514,I87497,I87449);
not I_5008 (I87531,I230204);
not I_5009 (I87548,I230180);
nor I_5010 (I87565,I87548,I230186);
and I_5011 (I87582,I87565,I230198);
or I_5012 (I87599,I87582,I230183);
DFFARX1 I_5013  ( .D(I87599), .CLK(I2350), .RSTB(I87398), .Q(I87616) );
nor I_5014 (I87633,I87616,I87497);
nand I_5015 (I87384,I87531,I87633);
not I_5016 (I87381,I87616);
and I_5017 (I87678,I87616,I87514);
DFFARX1 I_5018  ( .D(I87678), .CLK(I2350), .RSTB(I87398), .Q(I87366) );
DFFARX1 I_5019  ( .D(I87616), .CLK(I2350), .RSTB(I87398), .Q(I87709) );
and I_5020 (I87363,I87531,I87709);
nand I_5021 (I87740,I87415,I230180);
not I_5022 (I87757,I87740);
nor I_5023 (I87774,I87616,I87757);
DFFARX1 I_5024  ( .D(I230207), .CLK(I2350), .RSTB(I87398), .Q(I87791) );
nand I_5025 (I87808,I87791,I87740);
and I_5026 (I87825,I87531,I87808);
DFFARX1 I_5027  ( .D(I87825), .CLK(I2350), .RSTB(I87398), .Q(I87390) );
not I_5028 (I87856,I87791);
nand I_5029 (I87378,I87791,I87774);
nand I_5030 (I87372,I87791,I87757);
DFFARX1 I_5031  ( .D(I230192), .CLK(I2350), .RSTB(I87398), .Q(I87901) );
not I_5032 (I87918,I87901);
nor I_5033 (I87387,I87791,I87918);
nor I_5034 (I87949,I87918,I87856);
and I_5035 (I87966,I87497,I87949);
or I_5036 (I87983,I87740,I87966);
DFFARX1 I_5037  ( .D(I87983), .CLK(I2350), .RSTB(I87398), .Q(I87375) );
DFFARX1 I_5038  ( .D(I87918), .CLK(I2350), .RSTB(I87398), .Q(I87360) );
not I_5039 (I88061,I2357);
not I_5040 (I88078,I266047);
nor I_5041 (I88095,I266053,I266050);
nand I_5042 (I88112,I88095,I266068);
DFFARX1 I_5043  ( .D(I88112), .CLK(I2350), .RSTB(I88061), .Q(I88032) );
nor I_5044 (I88143,I88078,I266053);
nand I_5045 (I88160,I88143,I266077);
nand I_5046 (I88177,I88160,I88112);
not I_5047 (I88194,I266053);
not I_5048 (I88211,I266071);
nor I_5049 (I88228,I88211,I266062);
and I_5050 (I88245,I88228,I266065);
or I_5051 (I88262,I88245,I266056);
DFFARX1 I_5052  ( .D(I88262), .CLK(I2350), .RSTB(I88061), .Q(I88279) );
nor I_5053 (I88296,I88279,I88160);
nand I_5054 (I88047,I88194,I88296);
not I_5055 (I88044,I88279);
and I_5056 (I88341,I88279,I88177);
DFFARX1 I_5057  ( .D(I88341), .CLK(I2350), .RSTB(I88061), .Q(I88029) );
DFFARX1 I_5058  ( .D(I88279), .CLK(I2350), .RSTB(I88061), .Q(I88372) );
and I_5059 (I88026,I88194,I88372);
nand I_5060 (I88403,I88078,I266071);
not I_5061 (I88420,I88403);
nor I_5062 (I88437,I88279,I88420);
DFFARX1 I_5063  ( .D(I266074), .CLK(I2350), .RSTB(I88061), .Q(I88454) );
nand I_5064 (I88471,I88454,I88403);
and I_5065 (I88488,I88194,I88471);
DFFARX1 I_5066  ( .D(I88488), .CLK(I2350), .RSTB(I88061), .Q(I88053) );
not I_5067 (I88519,I88454);
nand I_5068 (I88041,I88454,I88437);
nand I_5069 (I88035,I88454,I88420);
DFFARX1 I_5070  ( .D(I266059), .CLK(I2350), .RSTB(I88061), .Q(I88564) );
not I_5071 (I88581,I88564);
nor I_5072 (I88050,I88454,I88581);
nor I_5073 (I88612,I88581,I88519);
and I_5074 (I88629,I88160,I88612);
or I_5075 (I88646,I88403,I88629);
DFFARX1 I_5076  ( .D(I88646), .CLK(I2350), .RSTB(I88061), .Q(I88038) );
DFFARX1 I_5077  ( .D(I88581), .CLK(I2350), .RSTB(I88061), .Q(I88023) );
not I_5078 (I88724,I2357);
not I_5079 (I88741,I352113);
nor I_5080 (I88758,I352119,I352131);
nand I_5081 (I88775,I88758,I352122);
DFFARX1 I_5082  ( .D(I88775), .CLK(I2350), .RSTB(I88724), .Q(I88695) );
nor I_5083 (I88806,I88741,I352119);
nand I_5084 (I88823,I88806,I352101);
nand I_5085 (I88840,I88823,I88775);
not I_5086 (I88857,I352119);
not I_5087 (I88874,I352116);
nor I_5088 (I88891,I88874,I352104);
and I_5089 (I88908,I88891,I352125);
or I_5090 (I88925,I88908,I352107);
DFFARX1 I_5091  ( .D(I88925), .CLK(I2350), .RSTB(I88724), .Q(I88942) );
nor I_5092 (I88959,I88942,I88823);
nand I_5093 (I88710,I88857,I88959);
not I_5094 (I88707,I88942);
and I_5095 (I89004,I88942,I88840);
DFFARX1 I_5096  ( .D(I89004), .CLK(I2350), .RSTB(I88724), .Q(I88692) );
DFFARX1 I_5097  ( .D(I88942), .CLK(I2350), .RSTB(I88724), .Q(I89035) );
and I_5098 (I88689,I88857,I89035);
nand I_5099 (I89066,I88741,I352116);
not I_5100 (I89083,I89066);
nor I_5101 (I89100,I88942,I89083);
DFFARX1 I_5102  ( .D(I352128), .CLK(I2350), .RSTB(I88724), .Q(I89117) );
nand I_5103 (I89134,I89117,I89066);
and I_5104 (I89151,I88857,I89134);
DFFARX1 I_5105  ( .D(I89151), .CLK(I2350), .RSTB(I88724), .Q(I88716) );
not I_5106 (I89182,I89117);
nand I_5107 (I88704,I89117,I89100);
nand I_5108 (I88698,I89117,I89083);
DFFARX1 I_5109  ( .D(I352110), .CLK(I2350), .RSTB(I88724), .Q(I89227) );
not I_5110 (I89244,I89227);
nor I_5111 (I88713,I89117,I89244);
nor I_5112 (I89275,I89244,I89182);
and I_5113 (I89292,I88823,I89275);
or I_5114 (I89309,I89066,I89292);
DFFARX1 I_5115  ( .D(I89309), .CLK(I2350), .RSTB(I88724), .Q(I88701) );
DFFARX1 I_5116  ( .D(I89244), .CLK(I2350), .RSTB(I88724), .Q(I88686) );
not I_5117 (I89387,I2357);
not I_5118 (I89404,I338275);
nor I_5119 (I89421,I338281,I338293);
nand I_5120 (I89438,I89421,I338284);
DFFARX1 I_5121  ( .D(I89438), .CLK(I2350), .RSTB(I89387), .Q(I89358) );
nor I_5122 (I89469,I89404,I338281);
nand I_5123 (I89486,I89469,I338263);
nand I_5124 (I89503,I89486,I89438);
not I_5125 (I89520,I338281);
not I_5126 (I89537,I338278);
nor I_5127 (I89554,I89537,I338266);
and I_5128 (I89571,I89554,I338287);
or I_5129 (I89588,I89571,I338269);
DFFARX1 I_5130  ( .D(I89588), .CLK(I2350), .RSTB(I89387), .Q(I89605) );
nor I_5131 (I89622,I89605,I89486);
nand I_5132 (I89373,I89520,I89622);
not I_5133 (I89370,I89605);
and I_5134 (I89667,I89605,I89503);
DFFARX1 I_5135  ( .D(I89667), .CLK(I2350), .RSTB(I89387), .Q(I89355) );
DFFARX1 I_5136  ( .D(I89605), .CLK(I2350), .RSTB(I89387), .Q(I89698) );
and I_5137 (I89352,I89520,I89698);
nand I_5138 (I89729,I89404,I338278);
not I_5139 (I89746,I89729);
nor I_5140 (I89763,I89605,I89746);
DFFARX1 I_5141  ( .D(I338290), .CLK(I2350), .RSTB(I89387), .Q(I89780) );
nand I_5142 (I89797,I89780,I89729);
and I_5143 (I89814,I89520,I89797);
DFFARX1 I_5144  ( .D(I89814), .CLK(I2350), .RSTB(I89387), .Q(I89379) );
not I_5145 (I89845,I89780);
nand I_5146 (I89367,I89780,I89763);
nand I_5147 (I89361,I89780,I89746);
DFFARX1 I_5148  ( .D(I338272), .CLK(I2350), .RSTB(I89387), .Q(I89890) );
not I_5149 (I89907,I89890);
nor I_5150 (I89376,I89780,I89907);
nor I_5151 (I89938,I89907,I89845);
and I_5152 (I89955,I89486,I89938);
or I_5153 (I89972,I89729,I89955);
DFFARX1 I_5154  ( .D(I89972), .CLK(I2350), .RSTB(I89387), .Q(I89364) );
DFFARX1 I_5155  ( .D(I89907), .CLK(I2350), .RSTB(I89387), .Q(I89349) );
not I_5156 (I90050,I2357);
not I_5157 (I90067,I47901);
nor I_5158 (I90084,I47889,I47913);
nand I_5159 (I90101,I90084,I47898);
DFFARX1 I_5160  ( .D(I90101), .CLK(I2350), .RSTB(I90050), .Q(I90021) );
nor I_5161 (I90132,I90067,I47889);
nand I_5162 (I90149,I90132,I47916);
nand I_5163 (I90166,I90149,I90101);
not I_5164 (I90183,I47889);
not I_5165 (I90200,I47886);
nor I_5166 (I90217,I90200,I47895);
and I_5167 (I90234,I90217,I47910);
or I_5168 (I90251,I90234,I47892);
DFFARX1 I_5169  ( .D(I90251), .CLK(I2350), .RSTB(I90050), .Q(I90268) );
nor I_5170 (I90285,I90268,I90149);
nand I_5171 (I90036,I90183,I90285);
not I_5172 (I90033,I90268);
and I_5173 (I90330,I90268,I90166);
DFFARX1 I_5174  ( .D(I90330), .CLK(I2350), .RSTB(I90050), .Q(I90018) );
DFFARX1 I_5175  ( .D(I90268), .CLK(I2350), .RSTB(I90050), .Q(I90361) );
and I_5176 (I90015,I90183,I90361);
nand I_5177 (I90392,I90067,I47886);
not I_5178 (I90409,I90392);
nor I_5179 (I90426,I90268,I90409);
DFFARX1 I_5180  ( .D(I47907), .CLK(I2350), .RSTB(I90050), .Q(I90443) );
nand I_5181 (I90460,I90443,I90392);
and I_5182 (I90477,I90183,I90460);
DFFARX1 I_5183  ( .D(I90477), .CLK(I2350), .RSTB(I90050), .Q(I90042) );
not I_5184 (I90508,I90443);
nand I_5185 (I90030,I90443,I90426);
nand I_5186 (I90024,I90443,I90409);
DFFARX1 I_5187  ( .D(I47904), .CLK(I2350), .RSTB(I90050), .Q(I90553) );
not I_5188 (I90570,I90553);
nor I_5189 (I90039,I90443,I90570);
nor I_5190 (I90601,I90570,I90508);
and I_5191 (I90618,I90149,I90601);
or I_5192 (I90635,I90392,I90618);
DFFARX1 I_5193  ( .D(I90635), .CLK(I2350), .RSTB(I90050), .Q(I90027) );
DFFARX1 I_5194  ( .D(I90570), .CLK(I2350), .RSTB(I90050), .Q(I90012) );
not I_5195 (I90713,I2357);
not I_5196 (I90730,I127589);
nor I_5197 (I90747,I127571,I127565);
nand I_5198 (I90764,I90747,I127568);
DFFARX1 I_5199  ( .D(I90764), .CLK(I2350), .RSTB(I90713), .Q(I90684) );
nor I_5200 (I90795,I90730,I127571);
nand I_5201 (I90812,I90795,I127577);
nand I_5202 (I90829,I90812,I90764);
not I_5203 (I90846,I127571);
not I_5204 (I90863,I127586);
nor I_5205 (I90880,I90863,I127574);
and I_5206 (I90897,I90880,I127580);
or I_5207 (I90914,I90897,I127595);
DFFARX1 I_5208  ( .D(I90914), .CLK(I2350), .RSTB(I90713), .Q(I90931) );
nor I_5209 (I90948,I90931,I90812);
nand I_5210 (I90699,I90846,I90948);
not I_5211 (I90696,I90931);
and I_5212 (I90993,I90931,I90829);
DFFARX1 I_5213  ( .D(I90993), .CLK(I2350), .RSTB(I90713), .Q(I90681) );
DFFARX1 I_5214  ( .D(I90931), .CLK(I2350), .RSTB(I90713), .Q(I91024) );
and I_5215 (I90678,I90846,I91024);
nand I_5216 (I91055,I90730,I127586);
not I_5217 (I91072,I91055);
nor I_5218 (I91089,I90931,I91072);
DFFARX1 I_5219  ( .D(I127583), .CLK(I2350), .RSTB(I90713), .Q(I91106) );
nand I_5220 (I91123,I91106,I91055);
and I_5221 (I91140,I90846,I91123);
DFFARX1 I_5222  ( .D(I91140), .CLK(I2350), .RSTB(I90713), .Q(I90705) );
not I_5223 (I91171,I91106);
nand I_5224 (I90693,I91106,I91089);
nand I_5225 (I90687,I91106,I91072);
DFFARX1 I_5226  ( .D(I127592), .CLK(I2350), .RSTB(I90713), .Q(I91216) );
not I_5227 (I91233,I91216);
nor I_5228 (I90702,I91106,I91233);
nor I_5229 (I91264,I91233,I91171);
and I_5230 (I91281,I90812,I91264);
or I_5231 (I91298,I91055,I91281);
DFFARX1 I_5232  ( .D(I91298), .CLK(I2350), .RSTB(I90713), .Q(I90690) );
DFFARX1 I_5233  ( .D(I91233), .CLK(I2350), .RSTB(I90713), .Q(I90675) );
not I_5234 (I91376,I2357);
not I_5235 (I91393,I146962);
nor I_5236 (I91410,I146971,I146983);
nand I_5237 (I91427,I91410,I146974);
DFFARX1 I_5238  ( .D(I91427), .CLK(I2350), .RSTB(I91376), .Q(I91347) );
nor I_5239 (I91458,I91393,I146971);
nand I_5240 (I91475,I91458,I146986);
nand I_5241 (I91492,I91475,I91427);
not I_5242 (I91509,I146971);
not I_5243 (I91526,I146992);
nor I_5244 (I91543,I91526,I146968);
and I_5245 (I91560,I91543,I146977);
or I_5246 (I91577,I91560,I146965);
DFFARX1 I_5247  ( .D(I91577), .CLK(I2350), .RSTB(I91376), .Q(I91594) );
nor I_5248 (I91611,I91594,I91475);
nand I_5249 (I91362,I91509,I91611);
not I_5250 (I91359,I91594);
and I_5251 (I91656,I91594,I91492);
DFFARX1 I_5252  ( .D(I91656), .CLK(I2350), .RSTB(I91376), .Q(I91344) );
DFFARX1 I_5253  ( .D(I91594), .CLK(I2350), .RSTB(I91376), .Q(I91687) );
and I_5254 (I91341,I91509,I91687);
nand I_5255 (I91718,I91393,I146992);
not I_5256 (I91735,I91718);
nor I_5257 (I91752,I91594,I91735);
DFFARX1 I_5258  ( .D(I146989), .CLK(I2350), .RSTB(I91376), .Q(I91769) );
nand I_5259 (I91786,I91769,I91718);
and I_5260 (I91803,I91509,I91786);
DFFARX1 I_5261  ( .D(I91803), .CLK(I2350), .RSTB(I91376), .Q(I91368) );
not I_5262 (I91834,I91769);
nand I_5263 (I91356,I91769,I91752);
nand I_5264 (I91350,I91769,I91735);
DFFARX1 I_5265  ( .D(I146980), .CLK(I2350), .RSTB(I91376), .Q(I91879) );
not I_5266 (I91896,I91879);
nor I_5267 (I91365,I91769,I91896);
nor I_5268 (I91927,I91896,I91834);
and I_5269 (I91944,I91475,I91927);
or I_5270 (I91961,I91718,I91944);
DFFARX1 I_5271  ( .D(I91961), .CLK(I2350), .RSTB(I91376), .Q(I91353) );
DFFARX1 I_5272  ( .D(I91896), .CLK(I2350), .RSTB(I91376), .Q(I91338) );
not I_5273 (I92039,I2357);
not I_5274 (I92056,I333243);
nor I_5275 (I92073,I333249,I333261);
nand I_5276 (I92090,I92073,I333252);
DFFARX1 I_5277  ( .D(I92090), .CLK(I2350), .RSTB(I92039), .Q(I92010) );
nor I_5278 (I92121,I92056,I333249);
nand I_5279 (I92138,I92121,I333231);
nand I_5280 (I92155,I92138,I92090);
not I_5281 (I92172,I333249);
not I_5282 (I92189,I333246);
nor I_5283 (I92206,I92189,I333234);
and I_5284 (I92223,I92206,I333255);
or I_5285 (I92240,I92223,I333237);
DFFARX1 I_5286  ( .D(I92240), .CLK(I2350), .RSTB(I92039), .Q(I92257) );
nor I_5287 (I92274,I92257,I92138);
nand I_5288 (I92025,I92172,I92274);
not I_5289 (I92022,I92257);
and I_5290 (I92319,I92257,I92155);
DFFARX1 I_5291  ( .D(I92319), .CLK(I2350), .RSTB(I92039), .Q(I92007) );
DFFARX1 I_5292  ( .D(I92257), .CLK(I2350), .RSTB(I92039), .Q(I92350) );
and I_5293 (I92004,I92172,I92350);
nand I_5294 (I92381,I92056,I333246);
not I_5295 (I92398,I92381);
nor I_5296 (I92415,I92257,I92398);
DFFARX1 I_5297  ( .D(I333258), .CLK(I2350), .RSTB(I92039), .Q(I92432) );
nand I_5298 (I92449,I92432,I92381);
and I_5299 (I92466,I92172,I92449);
DFFARX1 I_5300  ( .D(I92466), .CLK(I2350), .RSTB(I92039), .Q(I92031) );
not I_5301 (I92497,I92432);
nand I_5302 (I92019,I92432,I92415);
nand I_5303 (I92013,I92432,I92398);
DFFARX1 I_5304  ( .D(I333240), .CLK(I2350), .RSTB(I92039), .Q(I92542) );
not I_5305 (I92559,I92542);
nor I_5306 (I92028,I92432,I92559);
nor I_5307 (I92590,I92559,I92497);
and I_5308 (I92607,I92138,I92590);
or I_5309 (I92624,I92381,I92607);
DFFARX1 I_5310  ( .D(I92624), .CLK(I2350), .RSTB(I92039), .Q(I92016) );
DFFARX1 I_5311  ( .D(I92559), .CLK(I2350), .RSTB(I92039), .Q(I92001) );
not I_5312 (I92702,I2357);
not I_5313 (I92719,I343936);
nor I_5314 (I92736,I343942,I343954);
nand I_5315 (I92753,I92736,I343945);
DFFARX1 I_5316  ( .D(I92753), .CLK(I2350), .RSTB(I92702), .Q(I92673) );
nor I_5317 (I92784,I92719,I343942);
nand I_5318 (I92801,I92784,I343924);
nand I_5319 (I92818,I92801,I92753);
not I_5320 (I92835,I343942);
not I_5321 (I92852,I343939);
nor I_5322 (I92869,I92852,I343927);
and I_5323 (I92886,I92869,I343948);
or I_5324 (I92903,I92886,I343930);
DFFARX1 I_5325  ( .D(I92903), .CLK(I2350), .RSTB(I92702), .Q(I92920) );
nor I_5326 (I92937,I92920,I92801);
nand I_5327 (I92688,I92835,I92937);
not I_5328 (I92685,I92920);
and I_5329 (I92982,I92920,I92818);
DFFARX1 I_5330  ( .D(I92982), .CLK(I2350), .RSTB(I92702), .Q(I92670) );
DFFARX1 I_5331  ( .D(I92920), .CLK(I2350), .RSTB(I92702), .Q(I93013) );
and I_5332 (I92667,I92835,I93013);
nand I_5333 (I93044,I92719,I343939);
not I_5334 (I93061,I93044);
nor I_5335 (I93078,I92920,I93061);
DFFARX1 I_5336  ( .D(I343951), .CLK(I2350), .RSTB(I92702), .Q(I93095) );
nand I_5337 (I93112,I93095,I93044);
and I_5338 (I93129,I92835,I93112);
DFFARX1 I_5339  ( .D(I93129), .CLK(I2350), .RSTB(I92702), .Q(I92694) );
not I_5340 (I93160,I93095);
nand I_5341 (I92682,I93095,I93078);
nand I_5342 (I92676,I93095,I93061);
DFFARX1 I_5343  ( .D(I343933), .CLK(I2350), .RSTB(I92702), .Q(I93205) );
not I_5344 (I93222,I93205);
nor I_5345 (I92691,I93095,I93222);
nor I_5346 (I93253,I93222,I93160);
and I_5347 (I93270,I92801,I93253);
or I_5348 (I93287,I93044,I93270);
DFFARX1 I_5349  ( .D(I93287), .CLK(I2350), .RSTB(I92702), .Q(I92679) );
DFFARX1 I_5350  ( .D(I93222), .CLK(I2350), .RSTB(I92702), .Q(I92664) );
not I_5351 (I93365,I2357);
not I_5352 (I93382,I259111);
nor I_5353 (I93399,I259117,I259114);
nand I_5354 (I93416,I93399,I259132);
DFFARX1 I_5355  ( .D(I93416), .CLK(I2350), .RSTB(I93365), .Q(I93336) );
nor I_5356 (I93447,I93382,I259117);
nand I_5357 (I93464,I93447,I259141);
nand I_5358 (I93481,I93464,I93416);
not I_5359 (I93498,I259117);
not I_5360 (I93515,I259135);
nor I_5361 (I93532,I93515,I259126);
and I_5362 (I93549,I93532,I259129);
or I_5363 (I93566,I93549,I259120);
DFFARX1 I_5364  ( .D(I93566), .CLK(I2350), .RSTB(I93365), .Q(I93583) );
nor I_5365 (I93600,I93583,I93464);
nand I_5366 (I93351,I93498,I93600);
not I_5367 (I93348,I93583);
and I_5368 (I93645,I93583,I93481);
DFFARX1 I_5369  ( .D(I93645), .CLK(I2350), .RSTB(I93365), .Q(I93333) );
DFFARX1 I_5370  ( .D(I93583), .CLK(I2350), .RSTB(I93365), .Q(I93676) );
and I_5371 (I93330,I93498,I93676);
nand I_5372 (I93707,I93382,I259135);
not I_5373 (I93724,I93707);
nor I_5374 (I93741,I93583,I93724);
DFFARX1 I_5375  ( .D(I259138), .CLK(I2350), .RSTB(I93365), .Q(I93758) );
nand I_5376 (I93775,I93758,I93707);
and I_5377 (I93792,I93498,I93775);
DFFARX1 I_5378  ( .D(I93792), .CLK(I2350), .RSTB(I93365), .Q(I93357) );
not I_5379 (I93823,I93758);
nand I_5380 (I93345,I93758,I93741);
nand I_5381 (I93339,I93758,I93724);
DFFARX1 I_5382  ( .D(I259123), .CLK(I2350), .RSTB(I93365), .Q(I93868) );
not I_5383 (I93885,I93868);
nor I_5384 (I93354,I93758,I93885);
nor I_5385 (I93916,I93885,I93823);
and I_5386 (I93933,I93464,I93916);
or I_5387 (I93950,I93707,I93933);
DFFARX1 I_5388  ( .D(I93950), .CLK(I2350), .RSTB(I93365), .Q(I93342) );
DFFARX1 I_5389  ( .D(I93885), .CLK(I2350), .RSTB(I93365), .Q(I93327) );
not I_5390 (I94028,I2357);
not I_5391 (I94045,I354629);
nor I_5392 (I94062,I354635,I354647);
nand I_5393 (I94079,I94062,I354638);
DFFARX1 I_5394  ( .D(I94079), .CLK(I2350), .RSTB(I94028), .Q(I93999) );
nor I_5395 (I94110,I94045,I354635);
nand I_5396 (I94127,I94110,I354617);
nand I_5397 (I94144,I94127,I94079);
not I_5398 (I94161,I354635);
not I_5399 (I94178,I354632);
nor I_5400 (I94195,I94178,I354620);
and I_5401 (I94212,I94195,I354641);
or I_5402 (I94229,I94212,I354623);
DFFARX1 I_5403  ( .D(I94229), .CLK(I2350), .RSTB(I94028), .Q(I94246) );
nor I_5404 (I94263,I94246,I94127);
nand I_5405 (I94014,I94161,I94263);
not I_5406 (I94011,I94246);
and I_5407 (I94308,I94246,I94144);
DFFARX1 I_5408  ( .D(I94308), .CLK(I2350), .RSTB(I94028), .Q(I93996) );
DFFARX1 I_5409  ( .D(I94246), .CLK(I2350), .RSTB(I94028), .Q(I94339) );
and I_5410 (I93993,I94161,I94339);
nand I_5411 (I94370,I94045,I354632);
not I_5412 (I94387,I94370);
nor I_5413 (I94404,I94246,I94387);
DFFARX1 I_5414  ( .D(I354644), .CLK(I2350), .RSTB(I94028), .Q(I94421) );
nand I_5415 (I94438,I94421,I94370);
and I_5416 (I94455,I94161,I94438);
DFFARX1 I_5417  ( .D(I94455), .CLK(I2350), .RSTB(I94028), .Q(I94020) );
not I_5418 (I94486,I94421);
nand I_5419 (I94008,I94421,I94404);
nand I_5420 (I94002,I94421,I94387);
DFFARX1 I_5421  ( .D(I354626), .CLK(I2350), .RSTB(I94028), .Q(I94531) );
not I_5422 (I94548,I94531);
nor I_5423 (I94017,I94421,I94548);
nor I_5424 (I94579,I94548,I94486);
and I_5425 (I94596,I94127,I94579);
or I_5426 (I94613,I94370,I94596);
DFFARX1 I_5427  ( .D(I94613), .CLK(I2350), .RSTB(I94028), .Q(I94005) );
DFFARX1 I_5428  ( .D(I94548), .CLK(I2350), .RSTB(I94028), .Q(I93990) );
not I_5429 (I94691,I2357);
not I_5430 (I94708,I44671);
nor I_5431 (I94725,I44659,I44683);
nand I_5432 (I94742,I94725,I44668);
DFFARX1 I_5433  ( .D(I94742), .CLK(I2350), .RSTB(I94691), .Q(I94662) );
nor I_5434 (I94773,I94708,I44659);
nand I_5435 (I94790,I94773,I44686);
nand I_5436 (I94807,I94790,I94742);
not I_5437 (I94824,I44659);
not I_5438 (I94841,I44656);
nor I_5439 (I94858,I94841,I44665);
and I_5440 (I94875,I94858,I44680);
or I_5441 (I94892,I94875,I44662);
DFFARX1 I_5442  ( .D(I94892), .CLK(I2350), .RSTB(I94691), .Q(I94909) );
nor I_5443 (I94926,I94909,I94790);
nand I_5444 (I94677,I94824,I94926);
not I_5445 (I94674,I94909);
and I_5446 (I94971,I94909,I94807);
DFFARX1 I_5447  ( .D(I94971), .CLK(I2350), .RSTB(I94691), .Q(I94659) );
DFFARX1 I_5448  ( .D(I94909), .CLK(I2350), .RSTB(I94691), .Q(I95002) );
and I_5449 (I94656,I94824,I95002);
nand I_5450 (I95033,I94708,I44656);
not I_5451 (I95050,I95033);
nor I_5452 (I95067,I94909,I95050);
DFFARX1 I_5453  ( .D(I44677), .CLK(I2350), .RSTB(I94691), .Q(I95084) );
nand I_5454 (I95101,I95084,I95033);
and I_5455 (I95118,I94824,I95101);
DFFARX1 I_5456  ( .D(I95118), .CLK(I2350), .RSTB(I94691), .Q(I94683) );
not I_5457 (I95149,I95084);
nand I_5458 (I94671,I95084,I95067);
nand I_5459 (I94665,I95084,I95050);
DFFARX1 I_5460  ( .D(I44674), .CLK(I2350), .RSTB(I94691), .Q(I95194) );
not I_5461 (I95211,I95194);
nor I_5462 (I94680,I95084,I95211);
nor I_5463 (I95242,I95211,I95149);
and I_5464 (I95259,I94790,I95242);
or I_5465 (I95276,I95033,I95259);
DFFARX1 I_5466  ( .D(I95276), .CLK(I2350), .RSTB(I94691), .Q(I94668) );
DFFARX1 I_5467  ( .D(I95211), .CLK(I2350), .RSTB(I94691), .Q(I94653) );
not I_5468 (I95354,I2357);
not I_5469 (I95371,I273255);
nor I_5470 (I95388,I273267,I273270);
nand I_5471 (I95405,I95388,I273276);
DFFARX1 I_5472  ( .D(I95405), .CLK(I2350), .RSTB(I95354), .Q(I95325) );
nor I_5473 (I95436,I95371,I273267);
nand I_5474 (I95453,I95436,I273279);
nand I_5475 (I95470,I95453,I95405);
not I_5476 (I95487,I273267);
not I_5477 (I95504,I273258);
nor I_5478 (I95521,I95504,I273273);
and I_5479 (I95538,I95521,I273282);
or I_5480 (I95555,I95538,I273285);
DFFARX1 I_5481  ( .D(I95555), .CLK(I2350), .RSTB(I95354), .Q(I95572) );
nor I_5482 (I95589,I95572,I95453);
nand I_5483 (I95340,I95487,I95589);
not I_5484 (I95337,I95572);
and I_5485 (I95634,I95572,I95470);
DFFARX1 I_5486  ( .D(I95634), .CLK(I2350), .RSTB(I95354), .Q(I95322) );
DFFARX1 I_5487  ( .D(I95572), .CLK(I2350), .RSTB(I95354), .Q(I95665) );
and I_5488 (I95319,I95487,I95665);
nand I_5489 (I95696,I95371,I273258);
not I_5490 (I95713,I95696);
nor I_5491 (I95730,I95572,I95713);
DFFARX1 I_5492  ( .D(I273261), .CLK(I2350), .RSTB(I95354), .Q(I95747) );
nand I_5493 (I95764,I95747,I95696);
and I_5494 (I95781,I95487,I95764);
DFFARX1 I_5495  ( .D(I95781), .CLK(I2350), .RSTB(I95354), .Q(I95346) );
not I_5496 (I95812,I95747);
nand I_5497 (I95334,I95747,I95730);
nand I_5498 (I95328,I95747,I95713);
DFFARX1 I_5499  ( .D(I273264), .CLK(I2350), .RSTB(I95354), .Q(I95857) );
not I_5500 (I95874,I95857);
nor I_5501 (I95343,I95747,I95874);
nor I_5502 (I95905,I95874,I95812);
and I_5503 (I95922,I95453,I95905);
or I_5504 (I95939,I95696,I95922);
DFFARX1 I_5505  ( .D(I95939), .CLK(I2350), .RSTB(I95354), .Q(I95331) );
DFFARX1 I_5506  ( .D(I95874), .CLK(I2350), .RSTB(I95354), .Q(I95316) );
not I_5507 (I96017,I2357);
not I_5508 (I96034,I53069);
nor I_5509 (I96051,I53057,I53081);
nand I_5510 (I96068,I96051,I53066);
DFFARX1 I_5511  ( .D(I96068), .CLK(I2350), .RSTB(I96017), .Q(I95988) );
nor I_5512 (I96099,I96034,I53057);
nand I_5513 (I96116,I96099,I53084);
nand I_5514 (I96133,I96116,I96068);
not I_5515 (I96150,I53057);
not I_5516 (I96167,I53054);
nor I_5517 (I96184,I96167,I53063);
and I_5518 (I96201,I96184,I53078);
or I_5519 (I96218,I96201,I53060);
DFFARX1 I_5520  ( .D(I96218), .CLK(I2350), .RSTB(I96017), .Q(I96235) );
nor I_5521 (I96252,I96235,I96116);
nand I_5522 (I96003,I96150,I96252);
not I_5523 (I96000,I96235);
and I_5524 (I96297,I96235,I96133);
DFFARX1 I_5525  ( .D(I96297), .CLK(I2350), .RSTB(I96017), .Q(I95985) );
DFFARX1 I_5526  ( .D(I96235), .CLK(I2350), .RSTB(I96017), .Q(I96328) );
and I_5527 (I95982,I96150,I96328);
nand I_5528 (I96359,I96034,I53054);
not I_5529 (I96376,I96359);
nor I_5530 (I96393,I96235,I96376);
DFFARX1 I_5531  ( .D(I53075), .CLK(I2350), .RSTB(I96017), .Q(I96410) );
nand I_5532 (I96427,I96410,I96359);
and I_5533 (I96444,I96150,I96427);
DFFARX1 I_5534  ( .D(I96444), .CLK(I2350), .RSTB(I96017), .Q(I96009) );
not I_5535 (I96475,I96410);
nand I_5536 (I95997,I96410,I96393);
nand I_5537 (I95991,I96410,I96376);
DFFARX1 I_5538  ( .D(I53072), .CLK(I2350), .RSTB(I96017), .Q(I96520) );
not I_5539 (I96537,I96520);
nor I_5540 (I96006,I96410,I96537);
nor I_5541 (I96568,I96537,I96475);
and I_5542 (I96585,I96116,I96568);
or I_5543 (I96602,I96359,I96585);
DFFARX1 I_5544  ( .D(I96602), .CLK(I2350), .RSTB(I96017), .Q(I95994) );
DFFARX1 I_5545  ( .D(I96537), .CLK(I2350), .RSTB(I96017), .Q(I95979) );
not I_5546 (I96680,I2357);
not I_5547 (I96697,I324278);
nor I_5548 (I96714,I324293,I324275);
nand I_5549 (I96731,I96714,I324287);
DFFARX1 I_5550  ( .D(I96731), .CLK(I2350), .RSTB(I96680), .Q(I96651) );
nor I_5551 (I96762,I96697,I324293);
nand I_5552 (I96779,I96762,I324284);
nand I_5553 (I96796,I96779,I96731);
not I_5554 (I96813,I324293);
not I_5555 (I96830,I324302);
nor I_5556 (I96847,I96830,I324272);
and I_5557 (I96864,I96847,I324281);
or I_5558 (I96881,I96864,I324299);
DFFARX1 I_5559  ( .D(I96881), .CLK(I2350), .RSTB(I96680), .Q(I96898) );
nor I_5560 (I96915,I96898,I96779);
nand I_5561 (I96666,I96813,I96915);
not I_5562 (I96663,I96898);
and I_5563 (I96960,I96898,I96796);
DFFARX1 I_5564  ( .D(I96960), .CLK(I2350), .RSTB(I96680), .Q(I96648) );
DFFARX1 I_5565  ( .D(I96898), .CLK(I2350), .RSTB(I96680), .Q(I96991) );
and I_5566 (I96645,I96813,I96991);
nand I_5567 (I97022,I96697,I324302);
not I_5568 (I97039,I97022);
nor I_5569 (I97056,I96898,I97039);
DFFARX1 I_5570  ( .D(I324290), .CLK(I2350), .RSTB(I96680), .Q(I97073) );
nand I_5571 (I97090,I97073,I97022);
and I_5572 (I97107,I96813,I97090);
DFFARX1 I_5573  ( .D(I97107), .CLK(I2350), .RSTB(I96680), .Q(I96672) );
not I_5574 (I97138,I97073);
nand I_5575 (I96660,I97073,I97056);
nand I_5576 (I96654,I97073,I97039);
DFFARX1 I_5577  ( .D(I324296), .CLK(I2350), .RSTB(I96680), .Q(I97183) );
not I_5578 (I97200,I97183);
nor I_5579 (I96669,I97073,I97200);
nor I_5580 (I97231,I97200,I97138);
and I_5581 (I97248,I96779,I97231);
or I_5582 (I97265,I97022,I97248);
DFFARX1 I_5583  ( .D(I97265), .CLK(I2350), .RSTB(I96680), .Q(I96657) );
DFFARX1 I_5584  ( .D(I97200), .CLK(I2350), .RSTB(I96680), .Q(I96642) );
not I_5585 (I97343,I2357);
not I_5586 (I97360,I51131);
nor I_5587 (I97377,I51119,I51143);
nand I_5588 (I97394,I97377,I51128);
DFFARX1 I_5589  ( .D(I97394), .CLK(I2350), .RSTB(I97343), .Q(I97314) );
nor I_5590 (I97425,I97360,I51119);
nand I_5591 (I97442,I97425,I51146);
nand I_5592 (I97459,I97442,I97394);
not I_5593 (I97476,I51119);
not I_5594 (I97493,I51116);
nor I_5595 (I97510,I97493,I51125);
and I_5596 (I97527,I97510,I51140);
or I_5597 (I97544,I97527,I51122);
DFFARX1 I_5598  ( .D(I97544), .CLK(I2350), .RSTB(I97343), .Q(I97561) );
nor I_5599 (I97578,I97561,I97442);
nand I_5600 (I97329,I97476,I97578);
not I_5601 (I97326,I97561);
and I_5602 (I97623,I97561,I97459);
DFFARX1 I_5603  ( .D(I97623), .CLK(I2350), .RSTB(I97343), .Q(I97311) );
DFFARX1 I_5604  ( .D(I97561), .CLK(I2350), .RSTB(I97343), .Q(I97654) );
and I_5605 (I97308,I97476,I97654);
nand I_5606 (I97685,I97360,I51116);
not I_5607 (I97702,I97685);
nor I_5608 (I97719,I97561,I97702);
DFFARX1 I_5609  ( .D(I51137), .CLK(I2350), .RSTB(I97343), .Q(I97736) );
nand I_5610 (I97753,I97736,I97685);
and I_5611 (I97770,I97476,I97753);
DFFARX1 I_5612  ( .D(I97770), .CLK(I2350), .RSTB(I97343), .Q(I97335) );
not I_5613 (I97801,I97736);
nand I_5614 (I97323,I97736,I97719);
nand I_5615 (I97317,I97736,I97702);
DFFARX1 I_5616  ( .D(I51134), .CLK(I2350), .RSTB(I97343), .Q(I97846) );
not I_5617 (I97863,I97846);
nor I_5618 (I97332,I97736,I97863);
nor I_5619 (I97894,I97863,I97801);
and I_5620 (I97911,I97442,I97894);
or I_5621 (I97928,I97685,I97911);
DFFARX1 I_5622  ( .D(I97928), .CLK(I2350), .RSTB(I97343), .Q(I97320) );
DFFARX1 I_5623  ( .D(I97863), .CLK(I2350), .RSTB(I97343), .Q(I97305) );
not I_5624 (I98006,I2357);
not I_5625 (I98023,I209523);
nor I_5626 (I98040,I209532,I209505);
nand I_5627 (I98057,I98040,I209517);
DFFARX1 I_5628  ( .D(I98057), .CLK(I2350), .RSTB(I98006), .Q(I97977) );
nor I_5629 (I98088,I98023,I209532);
nand I_5630 (I98105,I98088,I209529);
nand I_5631 (I98122,I98105,I98057);
not I_5632 (I98139,I209532);
not I_5633 (I98156,I209508);
nor I_5634 (I98173,I98156,I209514);
and I_5635 (I98190,I98173,I209526);
or I_5636 (I98207,I98190,I209511);
DFFARX1 I_5637  ( .D(I98207), .CLK(I2350), .RSTB(I98006), .Q(I98224) );
nor I_5638 (I98241,I98224,I98105);
nand I_5639 (I97992,I98139,I98241);
not I_5640 (I97989,I98224);
and I_5641 (I98286,I98224,I98122);
DFFARX1 I_5642  ( .D(I98286), .CLK(I2350), .RSTB(I98006), .Q(I97974) );
DFFARX1 I_5643  ( .D(I98224), .CLK(I2350), .RSTB(I98006), .Q(I98317) );
and I_5644 (I97971,I98139,I98317);
nand I_5645 (I98348,I98023,I209508);
not I_5646 (I98365,I98348);
nor I_5647 (I98382,I98224,I98365);
DFFARX1 I_5648  ( .D(I209535), .CLK(I2350), .RSTB(I98006), .Q(I98399) );
nand I_5649 (I98416,I98399,I98348);
and I_5650 (I98433,I98139,I98416);
DFFARX1 I_5651  ( .D(I98433), .CLK(I2350), .RSTB(I98006), .Q(I97998) );
not I_5652 (I98464,I98399);
nand I_5653 (I97986,I98399,I98382);
nand I_5654 (I97980,I98399,I98365);
DFFARX1 I_5655  ( .D(I209520), .CLK(I2350), .RSTB(I98006), .Q(I98509) );
not I_5656 (I98526,I98509);
nor I_5657 (I97995,I98399,I98526);
nor I_5658 (I98557,I98526,I98464);
and I_5659 (I98574,I98105,I98557);
or I_5660 (I98591,I98348,I98574);
DFFARX1 I_5661  ( .D(I98591), .CLK(I2350), .RSTB(I98006), .Q(I97983) );
DFFARX1 I_5662  ( .D(I98526), .CLK(I2350), .RSTB(I98006), .Q(I97968) );
not I_5663 (I98669,I2357);
not I_5664 (I98686,I233997);
nor I_5665 (I98703,I234015,I234003);
nand I_5666 (I98720,I98703,I234009);
DFFARX1 I_5667  ( .D(I98720), .CLK(I2350), .RSTB(I98669), .Q(I98640) );
nor I_5668 (I98751,I98686,I234015);
nand I_5669 (I98768,I98751,I234012);
nand I_5670 (I98785,I98768,I98720);
not I_5671 (I98802,I234015);
not I_5672 (I98819,I233991);
nor I_5673 (I98836,I98819,I233985);
and I_5674 (I98853,I98836,I233994);
or I_5675 (I98870,I98853,I234006);
DFFARX1 I_5676  ( .D(I98870), .CLK(I2350), .RSTB(I98669), .Q(I98887) );
nor I_5677 (I98904,I98887,I98768);
nand I_5678 (I98655,I98802,I98904);
not I_5679 (I98652,I98887);
and I_5680 (I98949,I98887,I98785);
DFFARX1 I_5681  ( .D(I98949), .CLK(I2350), .RSTB(I98669), .Q(I98637) );
DFFARX1 I_5682  ( .D(I98887), .CLK(I2350), .RSTB(I98669), .Q(I98980) );
and I_5683 (I98634,I98802,I98980);
nand I_5684 (I99011,I98686,I233991);
not I_5685 (I99028,I99011);
nor I_5686 (I99045,I98887,I99028);
DFFARX1 I_5687  ( .D(I234000), .CLK(I2350), .RSTB(I98669), .Q(I99062) );
nand I_5688 (I99079,I99062,I99011);
and I_5689 (I99096,I98802,I99079);
DFFARX1 I_5690  ( .D(I99096), .CLK(I2350), .RSTB(I98669), .Q(I98661) );
not I_5691 (I99127,I99062);
nand I_5692 (I98649,I99062,I99045);
nand I_5693 (I98643,I99062,I99028);
DFFARX1 I_5694  ( .D(I233988), .CLK(I2350), .RSTB(I98669), .Q(I99172) );
not I_5695 (I99189,I99172);
nor I_5696 (I98658,I99062,I99189);
nor I_5697 (I99220,I99189,I99127);
and I_5698 (I99237,I98768,I99220);
or I_5699 (I99254,I99011,I99237);
DFFARX1 I_5700  ( .D(I99254), .CLK(I2350), .RSTB(I98669), .Q(I98646) );
DFFARX1 I_5701  ( .D(I99189), .CLK(I2350), .RSTB(I98669), .Q(I98631) );
not I_5702 (I99332,I2357);
not I_5703 (I99349,I301082);
nor I_5704 (I99366,I301094,I301097);
nand I_5705 (I99383,I99366,I301085);
DFFARX1 I_5706  ( .D(I99383), .CLK(I2350), .RSTB(I99332), .Q(I99303) );
nor I_5707 (I99414,I99349,I301094);
nand I_5708 (I99431,I99414,I301070);
nand I_5709 (I99448,I99431,I99383);
not I_5710 (I99465,I301094);
not I_5711 (I99482,I301073);
nor I_5712 (I99499,I99482,I301076);
and I_5713 (I99516,I99499,I301079);
or I_5714 (I99533,I99516,I301088);
DFFARX1 I_5715  ( .D(I99533), .CLK(I2350), .RSTB(I99332), .Q(I99550) );
nor I_5716 (I99567,I99550,I99431);
nand I_5717 (I99318,I99465,I99567);
not I_5718 (I99315,I99550);
and I_5719 (I99612,I99550,I99448);
DFFARX1 I_5720  ( .D(I99612), .CLK(I2350), .RSTB(I99332), .Q(I99300) );
DFFARX1 I_5721  ( .D(I99550), .CLK(I2350), .RSTB(I99332), .Q(I99643) );
and I_5722 (I99297,I99465,I99643);
nand I_5723 (I99674,I99349,I301073);
not I_5724 (I99691,I99674);
nor I_5725 (I99708,I99550,I99691);
DFFARX1 I_5726  ( .D(I301091), .CLK(I2350), .RSTB(I99332), .Q(I99725) );
nand I_5727 (I99742,I99725,I99674);
and I_5728 (I99759,I99465,I99742);
DFFARX1 I_5729  ( .D(I99759), .CLK(I2350), .RSTB(I99332), .Q(I99324) );
not I_5730 (I99790,I99725);
nand I_5731 (I99312,I99725,I99708);
nand I_5732 (I99306,I99725,I99691);
DFFARX1 I_5733  ( .D(I301067), .CLK(I2350), .RSTB(I99332), .Q(I99835) );
not I_5734 (I99852,I99835);
nor I_5735 (I99321,I99725,I99852);
nor I_5736 (I99883,I99852,I99790);
and I_5737 (I99900,I99431,I99883);
or I_5738 (I99917,I99674,I99900);
DFFARX1 I_5739  ( .D(I99917), .CLK(I2350), .RSTB(I99332), .Q(I99309) );
DFFARX1 I_5740  ( .D(I99852), .CLK(I2350), .RSTB(I99332), .Q(I99294) );
not I_5741 (I99995,I2357);
not I_5742 (I100012,I253909);
nor I_5743 (I100029,I253915,I253912);
nand I_5744 (I100046,I100029,I253930);
DFFARX1 I_5745  ( .D(I100046), .CLK(I2350), .RSTB(I99995), .Q(I99966) );
nor I_5746 (I100077,I100012,I253915);
nand I_5747 (I100094,I100077,I253939);
nand I_5748 (I100111,I100094,I100046);
not I_5749 (I100128,I253915);
not I_5750 (I100145,I253933);
nor I_5751 (I100162,I100145,I253924);
and I_5752 (I100179,I100162,I253927);
or I_5753 (I100196,I100179,I253918);
DFFARX1 I_5754  ( .D(I100196), .CLK(I2350), .RSTB(I99995), .Q(I100213) );
nor I_5755 (I100230,I100213,I100094);
nand I_5756 (I99981,I100128,I100230);
not I_5757 (I99978,I100213);
and I_5758 (I100275,I100213,I100111);
DFFARX1 I_5759  ( .D(I100275), .CLK(I2350), .RSTB(I99995), .Q(I99963) );
DFFARX1 I_5760  ( .D(I100213), .CLK(I2350), .RSTB(I99995), .Q(I100306) );
and I_5761 (I99960,I100128,I100306);
nand I_5762 (I100337,I100012,I253933);
not I_5763 (I100354,I100337);
nor I_5764 (I100371,I100213,I100354);
DFFARX1 I_5765  ( .D(I253936), .CLK(I2350), .RSTB(I99995), .Q(I100388) );
nand I_5766 (I100405,I100388,I100337);
and I_5767 (I100422,I100128,I100405);
DFFARX1 I_5768  ( .D(I100422), .CLK(I2350), .RSTB(I99995), .Q(I99987) );
not I_5769 (I100453,I100388);
nand I_5770 (I99975,I100388,I100371);
nand I_5771 (I99969,I100388,I100354);
DFFARX1 I_5772  ( .D(I253921), .CLK(I2350), .RSTB(I99995), .Q(I100498) );
not I_5773 (I100515,I100498);
nor I_5774 (I99984,I100388,I100515);
nor I_5775 (I100546,I100515,I100453);
and I_5776 (I100563,I100094,I100546);
or I_5777 (I100580,I100337,I100563);
DFFARX1 I_5778  ( .D(I100580), .CLK(I2350), .RSTB(I99995), .Q(I99972) );
DFFARX1 I_5779  ( .D(I100515), .CLK(I2350), .RSTB(I99995), .Q(I99957) );
not I_5780 (I100658,I2357);
not I_5781 (I100675,I58883);
nor I_5782 (I100692,I58871,I58895);
nand I_5783 (I100709,I100692,I58880);
DFFARX1 I_5784  ( .D(I100709), .CLK(I2350), .RSTB(I100658), .Q(I100629) );
nor I_5785 (I100740,I100675,I58871);
nand I_5786 (I100757,I100740,I58898);
nand I_5787 (I100774,I100757,I100709);
not I_5788 (I100791,I58871);
not I_5789 (I100808,I58868);
nor I_5790 (I100825,I100808,I58877);
and I_5791 (I100842,I100825,I58892);
or I_5792 (I100859,I100842,I58874);
DFFARX1 I_5793  ( .D(I100859), .CLK(I2350), .RSTB(I100658), .Q(I100876) );
nor I_5794 (I100893,I100876,I100757);
nand I_5795 (I100644,I100791,I100893);
not I_5796 (I100641,I100876);
and I_5797 (I100938,I100876,I100774);
DFFARX1 I_5798  ( .D(I100938), .CLK(I2350), .RSTB(I100658), .Q(I100626) );
DFFARX1 I_5799  ( .D(I100876), .CLK(I2350), .RSTB(I100658), .Q(I100969) );
and I_5800 (I100623,I100791,I100969);
nand I_5801 (I101000,I100675,I58868);
not I_5802 (I101017,I101000);
nor I_5803 (I101034,I100876,I101017);
DFFARX1 I_5804  ( .D(I58889), .CLK(I2350), .RSTB(I100658), .Q(I101051) );
nand I_5805 (I101068,I101051,I101000);
and I_5806 (I101085,I100791,I101068);
DFFARX1 I_5807  ( .D(I101085), .CLK(I2350), .RSTB(I100658), .Q(I100650) );
not I_5808 (I101116,I101051);
nand I_5809 (I100638,I101051,I101034);
nand I_5810 (I100632,I101051,I101017);
DFFARX1 I_5811  ( .D(I58886), .CLK(I2350), .RSTB(I100658), .Q(I101161) );
not I_5812 (I101178,I101161);
nor I_5813 (I100647,I101051,I101178);
nor I_5814 (I101209,I101178,I101116);
and I_5815 (I101226,I100757,I101209);
or I_5816 (I101243,I101000,I101226);
DFFARX1 I_5817  ( .D(I101243), .CLK(I2350), .RSTB(I100658), .Q(I100635) );
DFFARX1 I_5818  ( .D(I101178), .CLK(I2350), .RSTB(I100658), .Q(I100620) );
not I_5819 (I101321,I2357);
not I_5820 (I101338,I56299);
nor I_5821 (I101355,I56287,I56311);
nand I_5822 (I101372,I101355,I56296);
DFFARX1 I_5823  ( .D(I101372), .CLK(I2350), .RSTB(I101321), .Q(I101292) );
nor I_5824 (I101403,I101338,I56287);
nand I_5825 (I101420,I101403,I56314);
nand I_5826 (I101437,I101420,I101372);
not I_5827 (I101454,I56287);
not I_5828 (I101471,I56284);
nor I_5829 (I101488,I101471,I56293);
and I_5830 (I101505,I101488,I56308);
or I_5831 (I101522,I101505,I56290);
DFFARX1 I_5832  ( .D(I101522), .CLK(I2350), .RSTB(I101321), .Q(I101539) );
nor I_5833 (I101556,I101539,I101420);
nand I_5834 (I101307,I101454,I101556);
not I_5835 (I101304,I101539);
and I_5836 (I101601,I101539,I101437);
DFFARX1 I_5837  ( .D(I101601), .CLK(I2350), .RSTB(I101321), .Q(I101289) );
DFFARX1 I_5838  ( .D(I101539), .CLK(I2350), .RSTB(I101321), .Q(I101632) );
and I_5839 (I101286,I101454,I101632);
nand I_5840 (I101663,I101338,I56284);
not I_5841 (I101680,I101663);
nor I_5842 (I101697,I101539,I101680);
DFFARX1 I_5843  ( .D(I56305), .CLK(I2350), .RSTB(I101321), .Q(I101714) );
nand I_5844 (I101731,I101714,I101663);
and I_5845 (I101748,I101454,I101731);
DFFARX1 I_5846  ( .D(I101748), .CLK(I2350), .RSTB(I101321), .Q(I101313) );
not I_5847 (I101779,I101714);
nand I_5848 (I101301,I101714,I101697);
nand I_5849 (I101295,I101714,I101680);
DFFARX1 I_5850  ( .D(I56302), .CLK(I2350), .RSTB(I101321), .Q(I101824) );
not I_5851 (I101841,I101824);
nor I_5852 (I101310,I101714,I101841);
nor I_5853 (I101872,I101841,I101779);
and I_5854 (I101889,I101420,I101872);
or I_5855 (I101906,I101663,I101889);
DFFARX1 I_5856  ( .D(I101906), .CLK(I2350), .RSTB(I101321), .Q(I101298) );
DFFARX1 I_5857  ( .D(I101841), .CLK(I2350), .RSTB(I101321), .Q(I101283) );
not I_5858 (I101984,I2357);
not I_5859 (I102001,I385105);
nor I_5860 (I102018,I385084,I385096);
nand I_5861 (I102035,I102018,I385090);
DFFARX1 I_5862  ( .D(I102035), .CLK(I2350), .RSTB(I101984), .Q(I101955) );
nor I_5863 (I102066,I102001,I385084);
nand I_5864 (I102083,I102066,I385111);
nand I_5865 (I102100,I102083,I102035);
not I_5866 (I102117,I385084);
not I_5867 (I102134,I385087);
nor I_5868 (I102151,I102134,I385099);
and I_5869 (I102168,I102151,I385102);
or I_5870 (I102185,I102168,I385108);
DFFARX1 I_5871  ( .D(I102185), .CLK(I2350), .RSTB(I101984), .Q(I102202) );
nor I_5872 (I102219,I102202,I102083);
nand I_5873 (I101970,I102117,I102219);
not I_5874 (I101967,I102202);
and I_5875 (I102264,I102202,I102100);
DFFARX1 I_5876  ( .D(I102264), .CLK(I2350), .RSTB(I101984), .Q(I101952) );
DFFARX1 I_5877  ( .D(I102202), .CLK(I2350), .RSTB(I101984), .Q(I102295) );
and I_5878 (I101949,I102117,I102295);
nand I_5879 (I102326,I102001,I385087);
not I_5880 (I102343,I102326);
nor I_5881 (I102360,I102202,I102343);
DFFARX1 I_5882  ( .D(I385081), .CLK(I2350), .RSTB(I101984), .Q(I102377) );
nand I_5883 (I102394,I102377,I102326);
and I_5884 (I102411,I102117,I102394);
DFFARX1 I_5885  ( .D(I102411), .CLK(I2350), .RSTB(I101984), .Q(I101976) );
not I_5886 (I102442,I102377);
nand I_5887 (I101964,I102377,I102360);
nand I_5888 (I101958,I102377,I102343);
DFFARX1 I_5889  ( .D(I385093), .CLK(I2350), .RSTB(I101984), .Q(I102487) );
not I_5890 (I102504,I102487);
nor I_5891 (I101973,I102377,I102504);
nor I_5892 (I102535,I102504,I102442);
and I_5893 (I102552,I102083,I102535);
or I_5894 (I102569,I102326,I102552);
DFFARX1 I_5895  ( .D(I102569), .CLK(I2350), .RSTB(I101984), .Q(I101961) );
DFFARX1 I_5896  ( .D(I102504), .CLK(I2350), .RSTB(I101984), .Q(I101946) );
not I_5897 (I102647,I2357);
not I_5898 (I102664,I161548);
nor I_5899 (I102681,I161557,I161569);
nand I_5900 (I102698,I102681,I161560);
DFFARX1 I_5901  ( .D(I102698), .CLK(I2350), .RSTB(I102647), .Q(I102618) );
nor I_5902 (I102729,I102664,I161557);
nand I_5903 (I102746,I102729,I161572);
nand I_5904 (I102763,I102746,I102698);
not I_5905 (I102780,I161557);
not I_5906 (I102797,I161578);
nor I_5907 (I102814,I102797,I161554);
and I_5908 (I102831,I102814,I161563);
or I_5909 (I102848,I102831,I161551);
DFFARX1 I_5910  ( .D(I102848), .CLK(I2350), .RSTB(I102647), .Q(I102865) );
nor I_5911 (I102882,I102865,I102746);
nand I_5912 (I102633,I102780,I102882);
not I_5913 (I102630,I102865);
and I_5914 (I102927,I102865,I102763);
DFFARX1 I_5915  ( .D(I102927), .CLK(I2350), .RSTB(I102647), .Q(I102615) );
DFFARX1 I_5916  ( .D(I102865), .CLK(I2350), .RSTB(I102647), .Q(I102958) );
and I_5917 (I102612,I102780,I102958);
nand I_5918 (I102989,I102664,I161578);
not I_5919 (I103006,I102989);
nor I_5920 (I103023,I102865,I103006);
DFFARX1 I_5921  ( .D(I161575), .CLK(I2350), .RSTB(I102647), .Q(I103040) );
nand I_5922 (I103057,I103040,I102989);
and I_5923 (I103074,I102780,I103057);
DFFARX1 I_5924  ( .D(I103074), .CLK(I2350), .RSTB(I102647), .Q(I102639) );
not I_5925 (I103105,I103040);
nand I_5926 (I102627,I103040,I103023);
nand I_5927 (I102621,I103040,I103006);
DFFARX1 I_5928  ( .D(I161566), .CLK(I2350), .RSTB(I102647), .Q(I103150) );
not I_5929 (I103167,I103150);
nor I_5930 (I102636,I103040,I103167);
nor I_5931 (I103198,I103167,I103105);
and I_5932 (I103215,I102746,I103198);
or I_5933 (I103232,I102989,I103215);
DFFARX1 I_5934  ( .D(I103232), .CLK(I2350), .RSTB(I102647), .Q(I102624) );
DFFARX1 I_5935  ( .D(I103167), .CLK(I2350), .RSTB(I102647), .Q(I102609) );
not I_5936 (I103310,I2357);
not I_5937 (I103327,I254487);
nor I_5938 (I103344,I254493,I254490);
nand I_5939 (I103361,I103344,I254508);
DFFARX1 I_5940  ( .D(I103361), .CLK(I2350), .RSTB(I103310), .Q(I103281) );
nor I_5941 (I103392,I103327,I254493);
nand I_5942 (I103409,I103392,I254517);
nand I_5943 (I103426,I103409,I103361);
not I_5944 (I103443,I254493);
not I_5945 (I103460,I254511);
nor I_5946 (I103477,I103460,I254502);
and I_5947 (I103494,I103477,I254505);
or I_5948 (I103511,I103494,I254496);
DFFARX1 I_5949  ( .D(I103511), .CLK(I2350), .RSTB(I103310), .Q(I103528) );
nor I_5950 (I103545,I103528,I103409);
nand I_5951 (I103296,I103443,I103545);
not I_5952 (I103293,I103528);
and I_5953 (I103590,I103528,I103426);
DFFARX1 I_5954  ( .D(I103590), .CLK(I2350), .RSTB(I103310), .Q(I103278) );
DFFARX1 I_5955  ( .D(I103528), .CLK(I2350), .RSTB(I103310), .Q(I103621) );
and I_5956 (I103275,I103443,I103621);
nand I_5957 (I103652,I103327,I254511);
not I_5958 (I103669,I103652);
nor I_5959 (I103686,I103528,I103669);
DFFARX1 I_5960  ( .D(I254514), .CLK(I2350), .RSTB(I103310), .Q(I103703) );
nand I_5961 (I103720,I103703,I103652);
and I_5962 (I103737,I103443,I103720);
DFFARX1 I_5963  ( .D(I103737), .CLK(I2350), .RSTB(I103310), .Q(I103302) );
not I_5964 (I103768,I103703);
nand I_5965 (I103290,I103703,I103686);
nand I_5966 (I103284,I103703,I103669);
DFFARX1 I_5967  ( .D(I254499), .CLK(I2350), .RSTB(I103310), .Q(I103813) );
not I_5968 (I103830,I103813);
nor I_5969 (I103299,I103703,I103830);
nor I_5970 (I103861,I103830,I103768);
and I_5971 (I103878,I103409,I103861);
or I_5972 (I103895,I103652,I103878);
DFFARX1 I_5973  ( .D(I103895), .CLK(I2350), .RSTB(I103310), .Q(I103287) );
DFFARX1 I_5974  ( .D(I103830), .CLK(I2350), .RSTB(I103310), .Q(I103272) );
not I_5975 (I103973,I2357);
not I_5976 (I103990,I316543);
nor I_5977 (I104007,I316558,I316540);
nand I_5978 (I104024,I104007,I316552);
DFFARX1 I_5979  ( .D(I104024), .CLK(I2350), .RSTB(I103973), .Q(I103944) );
nor I_5980 (I104055,I103990,I316558);
nand I_5981 (I104072,I104055,I316549);
nand I_5982 (I104089,I104072,I104024);
not I_5983 (I104106,I316558);
not I_5984 (I104123,I316567);
nor I_5985 (I104140,I104123,I316537);
and I_5986 (I104157,I104140,I316546);
or I_5987 (I104174,I104157,I316564);
DFFARX1 I_5988  ( .D(I104174), .CLK(I2350), .RSTB(I103973), .Q(I104191) );
nor I_5989 (I104208,I104191,I104072);
nand I_5990 (I103959,I104106,I104208);
not I_5991 (I103956,I104191);
and I_5992 (I104253,I104191,I104089);
DFFARX1 I_5993  ( .D(I104253), .CLK(I2350), .RSTB(I103973), .Q(I103941) );
DFFARX1 I_5994  ( .D(I104191), .CLK(I2350), .RSTB(I103973), .Q(I104284) );
and I_5995 (I103938,I104106,I104284);
nand I_5996 (I104315,I103990,I316567);
not I_5997 (I104332,I104315);
nor I_5998 (I104349,I104191,I104332);
DFFARX1 I_5999  ( .D(I316555), .CLK(I2350), .RSTB(I103973), .Q(I104366) );
nand I_6000 (I104383,I104366,I104315);
and I_6001 (I104400,I104106,I104383);
DFFARX1 I_6002  ( .D(I104400), .CLK(I2350), .RSTB(I103973), .Q(I103965) );
not I_6003 (I104431,I104366);
nand I_6004 (I103953,I104366,I104349);
nand I_6005 (I103947,I104366,I104332);
DFFARX1 I_6006  ( .D(I316561), .CLK(I2350), .RSTB(I103973), .Q(I104476) );
not I_6007 (I104493,I104476);
nor I_6008 (I103962,I104366,I104493);
nor I_6009 (I104524,I104493,I104431);
and I_6010 (I104541,I104072,I104524);
or I_6011 (I104558,I104315,I104541);
DFFARX1 I_6012  ( .D(I104558), .CLK(I2350), .RSTB(I103973), .Q(I103950) );
DFFARX1 I_6013  ( .D(I104493), .CLK(I2350), .RSTB(I103973), .Q(I103935) );
not I_6014 (I104636,I2357);
not I_6015 (I104653,I266631);
nor I_6016 (I104670,I266637,I266628);
nand I_6017 (I104687,I104670,I266646);
DFFARX1 I_6018  ( .D(I104687), .CLK(I2350), .RSTB(I104636), .Q(I104607) );
nor I_6019 (I104718,I104653,I266637);
nand I_6020 (I104735,I104718,I266625);
nand I_6021 (I104752,I104735,I104687);
not I_6022 (I104769,I266637);
not I_6023 (I104786,I266655);
nor I_6024 (I104803,I104786,I266634);
and I_6025 (I104820,I104803,I266643);
or I_6026 (I104837,I104820,I266649);
DFFARX1 I_6027  ( .D(I104837), .CLK(I2350), .RSTB(I104636), .Q(I104854) );
nor I_6028 (I104871,I104854,I104735);
nand I_6029 (I104622,I104769,I104871);
not I_6030 (I104619,I104854);
and I_6031 (I104916,I104854,I104752);
DFFARX1 I_6032  ( .D(I104916), .CLK(I2350), .RSTB(I104636), .Q(I104604) );
DFFARX1 I_6033  ( .D(I104854), .CLK(I2350), .RSTB(I104636), .Q(I104947) );
and I_6034 (I104601,I104769,I104947);
nand I_6035 (I104978,I104653,I266655);
not I_6036 (I104995,I104978);
nor I_6037 (I105012,I104854,I104995);
DFFARX1 I_6038  ( .D(I266640), .CLK(I2350), .RSTB(I104636), .Q(I105029) );
nand I_6039 (I105046,I105029,I104978);
and I_6040 (I105063,I104769,I105046);
DFFARX1 I_6041  ( .D(I105063), .CLK(I2350), .RSTB(I104636), .Q(I104628) );
not I_6042 (I105094,I105029);
nand I_6043 (I104616,I105029,I105012);
nand I_6044 (I104610,I105029,I104995);
DFFARX1 I_6045  ( .D(I266652), .CLK(I2350), .RSTB(I104636), .Q(I105139) );
not I_6046 (I105156,I105139);
nor I_6047 (I104625,I105029,I105156);
nor I_6048 (I105187,I105156,I105094);
and I_6049 (I105204,I104735,I105187);
or I_6050 (I105221,I104978,I105204);
DFFARX1 I_6051  ( .D(I105221), .CLK(I2350), .RSTB(I104636), .Q(I104613) );
DFFARX1 I_6052  ( .D(I105156), .CLK(I2350), .RSTB(I104636), .Q(I104598) );
not I_6053 (I105299,I2357);
not I_6054 (I105316,I33043);
nor I_6055 (I105333,I33031,I33055);
nand I_6056 (I105350,I105333,I33040);
DFFARX1 I_6057  ( .D(I105350), .CLK(I2350), .RSTB(I105299), .Q(I105270) );
nor I_6058 (I105381,I105316,I33031);
nand I_6059 (I105398,I105381,I33058);
nand I_6060 (I105415,I105398,I105350);
not I_6061 (I105432,I33031);
not I_6062 (I105449,I33028);
nor I_6063 (I105466,I105449,I33037);
and I_6064 (I105483,I105466,I33052);
or I_6065 (I105500,I105483,I33034);
DFFARX1 I_6066  ( .D(I105500), .CLK(I2350), .RSTB(I105299), .Q(I105517) );
nor I_6067 (I105534,I105517,I105398);
nand I_6068 (I105285,I105432,I105534);
not I_6069 (I105282,I105517);
and I_6070 (I105579,I105517,I105415);
DFFARX1 I_6071  ( .D(I105579), .CLK(I2350), .RSTB(I105299), .Q(I105267) );
DFFARX1 I_6072  ( .D(I105517), .CLK(I2350), .RSTB(I105299), .Q(I105610) );
and I_6073 (I105264,I105432,I105610);
nand I_6074 (I105641,I105316,I33028);
not I_6075 (I105658,I105641);
nor I_6076 (I105675,I105517,I105658);
DFFARX1 I_6077  ( .D(I33049), .CLK(I2350), .RSTB(I105299), .Q(I105692) );
nand I_6078 (I105709,I105692,I105641);
and I_6079 (I105726,I105432,I105709);
DFFARX1 I_6080  ( .D(I105726), .CLK(I2350), .RSTB(I105299), .Q(I105291) );
not I_6081 (I105757,I105692);
nand I_6082 (I105279,I105692,I105675);
nand I_6083 (I105273,I105692,I105658);
DFFARX1 I_6084  ( .D(I33046), .CLK(I2350), .RSTB(I105299), .Q(I105802) );
not I_6085 (I105819,I105802);
nor I_6086 (I105288,I105692,I105819);
nor I_6087 (I105850,I105819,I105757);
and I_6088 (I105867,I105398,I105850);
or I_6089 (I105884,I105641,I105867);
DFFARX1 I_6090  ( .D(I105884), .CLK(I2350), .RSTB(I105299), .Q(I105276) );
DFFARX1 I_6091  ( .D(I105819), .CLK(I2350), .RSTB(I105299), .Q(I105261) );
not I_6092 (I105962,I2357);
not I_6093 (I105979,I320708);
nor I_6094 (I105996,I320723,I320705);
nand I_6095 (I106013,I105996,I320717);
DFFARX1 I_6096  ( .D(I106013), .CLK(I2350), .RSTB(I105962), .Q(I105933) );
nor I_6097 (I106044,I105979,I320723);
nand I_6098 (I106061,I106044,I320714);
nand I_6099 (I106078,I106061,I106013);
not I_6100 (I106095,I320723);
not I_6101 (I106112,I320732);
nor I_6102 (I106129,I106112,I320702);
and I_6103 (I106146,I106129,I320711);
or I_6104 (I106163,I106146,I320729);
DFFARX1 I_6105  ( .D(I106163), .CLK(I2350), .RSTB(I105962), .Q(I106180) );
nor I_6106 (I106197,I106180,I106061);
nand I_6107 (I105948,I106095,I106197);
not I_6108 (I105945,I106180);
and I_6109 (I106242,I106180,I106078);
DFFARX1 I_6110  ( .D(I106242), .CLK(I2350), .RSTB(I105962), .Q(I105930) );
DFFARX1 I_6111  ( .D(I106180), .CLK(I2350), .RSTB(I105962), .Q(I106273) );
and I_6112 (I105927,I106095,I106273);
nand I_6113 (I106304,I105979,I320732);
not I_6114 (I106321,I106304);
nor I_6115 (I106338,I106180,I106321);
DFFARX1 I_6116  ( .D(I320720), .CLK(I2350), .RSTB(I105962), .Q(I106355) );
nand I_6117 (I106372,I106355,I106304);
and I_6118 (I106389,I106095,I106372);
DFFARX1 I_6119  ( .D(I106389), .CLK(I2350), .RSTB(I105962), .Q(I105954) );
not I_6120 (I106420,I106355);
nand I_6121 (I105942,I106355,I106338);
nand I_6122 (I105936,I106355,I106321);
DFFARX1 I_6123  ( .D(I320726), .CLK(I2350), .RSTB(I105962), .Q(I106465) );
not I_6124 (I106482,I106465);
nor I_6125 (I105951,I106355,I106482);
nor I_6126 (I106513,I106482,I106420);
and I_6127 (I106530,I106061,I106513);
or I_6128 (I106547,I106304,I106530);
DFFARX1 I_6129  ( .D(I106547), .CLK(I2350), .RSTB(I105962), .Q(I105939) );
DFFARX1 I_6130  ( .D(I106482), .CLK(I2350), .RSTB(I105962), .Q(I105924) );
not I_6131 (I106625,I2357);
not I_6132 (I106642,I19205);
nor I_6133 (I106659,I19193,I19196);
nand I_6134 (I106676,I106659,I19211);
DFFARX1 I_6135  ( .D(I106676), .CLK(I2350), .RSTB(I106625), .Q(I106596) );
nor I_6136 (I106707,I106642,I19193);
nand I_6137 (I106724,I106707,I19202);
nand I_6138 (I106741,I106724,I106676);
not I_6139 (I106758,I19193);
not I_6140 (I106775,I19214);
nor I_6141 (I106792,I106775,I19190);
and I_6142 (I106809,I106792,I19199);
or I_6143 (I106826,I106809,I19208);
DFFARX1 I_6144  ( .D(I106826), .CLK(I2350), .RSTB(I106625), .Q(I106843) );
nor I_6145 (I106860,I106843,I106724);
nand I_6146 (I106611,I106758,I106860);
not I_6147 (I106608,I106843);
and I_6148 (I106905,I106843,I106741);
DFFARX1 I_6149  ( .D(I106905), .CLK(I2350), .RSTB(I106625), .Q(I106593) );
DFFARX1 I_6150  ( .D(I106843), .CLK(I2350), .RSTB(I106625), .Q(I106936) );
and I_6151 (I106590,I106758,I106936);
nand I_6152 (I106967,I106642,I19214);
not I_6153 (I106984,I106967);
nor I_6154 (I107001,I106843,I106984);
DFFARX1 I_6155  ( .D(I19220), .CLK(I2350), .RSTB(I106625), .Q(I107018) );
nand I_6156 (I107035,I107018,I106967);
and I_6157 (I107052,I106758,I107035);
DFFARX1 I_6158  ( .D(I107052), .CLK(I2350), .RSTB(I106625), .Q(I106617) );
not I_6159 (I107083,I107018);
nand I_6160 (I106605,I107018,I107001);
nand I_6161 (I106599,I107018,I106984);
DFFARX1 I_6162  ( .D(I19217), .CLK(I2350), .RSTB(I106625), .Q(I107128) );
not I_6163 (I107145,I107128);
nor I_6164 (I106614,I107018,I107145);
nor I_6165 (I107176,I107145,I107083);
and I_6166 (I107193,I106724,I107176);
or I_6167 (I107210,I106967,I107193);
DFFARX1 I_6168  ( .D(I107210), .CLK(I2350), .RSTB(I106625), .Q(I106602) );
DFFARX1 I_6169  ( .D(I107145), .CLK(I2350), .RSTB(I106625), .Q(I106587) );
not I_6170 (I107288,I2357);
not I_6171 (I107305,I8546);
nor I_6172 (I107322,I8534,I8537);
nand I_6173 (I107339,I107322,I8552);
DFFARX1 I_6174  ( .D(I107339), .CLK(I2350), .RSTB(I107288), .Q(I107259) );
nor I_6175 (I107370,I107305,I8534);
nand I_6176 (I107387,I107370,I8543);
nand I_6177 (I107404,I107387,I107339);
not I_6178 (I107421,I8534);
not I_6179 (I107438,I8555);
nor I_6180 (I107455,I107438,I8531);
and I_6181 (I107472,I107455,I8540);
or I_6182 (I107489,I107472,I8549);
DFFARX1 I_6183  ( .D(I107489), .CLK(I2350), .RSTB(I107288), .Q(I107506) );
nor I_6184 (I107523,I107506,I107387);
nand I_6185 (I107274,I107421,I107523);
not I_6186 (I107271,I107506);
and I_6187 (I107568,I107506,I107404);
DFFARX1 I_6188  ( .D(I107568), .CLK(I2350), .RSTB(I107288), .Q(I107256) );
DFFARX1 I_6189  ( .D(I107506), .CLK(I2350), .RSTB(I107288), .Q(I107599) );
and I_6190 (I107253,I107421,I107599);
nand I_6191 (I107630,I107305,I8555);
not I_6192 (I107647,I107630);
nor I_6193 (I107664,I107506,I107647);
DFFARX1 I_6194  ( .D(I8561), .CLK(I2350), .RSTB(I107288), .Q(I107681) );
nand I_6195 (I107698,I107681,I107630);
and I_6196 (I107715,I107421,I107698);
DFFARX1 I_6197  ( .D(I107715), .CLK(I2350), .RSTB(I107288), .Q(I107280) );
not I_6198 (I107746,I107681);
nand I_6199 (I107268,I107681,I107664);
nand I_6200 (I107262,I107681,I107647);
DFFARX1 I_6201  ( .D(I8558), .CLK(I2350), .RSTB(I107288), .Q(I107791) );
not I_6202 (I107808,I107791);
nor I_6203 (I107277,I107681,I107808);
nor I_6204 (I107839,I107808,I107746);
and I_6205 (I107856,I107387,I107839);
or I_6206 (I107873,I107630,I107856);
DFFARX1 I_6207  ( .D(I107873), .CLK(I2350), .RSTB(I107288), .Q(I107265) );
DFFARX1 I_6208  ( .D(I107808), .CLK(I2350), .RSTB(I107288), .Q(I107250) );
not I_6209 (I107951,I2357);
not I_6210 (I107968,I73095);
nor I_6211 (I107985,I73083,I73107);
nand I_6212 (I108002,I107985,I73092);
DFFARX1 I_6213  ( .D(I108002), .CLK(I2350), .RSTB(I107951), .Q(I107922) );
nor I_6214 (I108033,I107968,I73083);
nand I_6215 (I108050,I108033,I73110);
nand I_6216 (I108067,I108050,I108002);
not I_6217 (I108084,I73083);
not I_6218 (I108101,I73080);
nor I_6219 (I108118,I108101,I73089);
and I_6220 (I108135,I108118,I73104);
or I_6221 (I108152,I108135,I73086);
DFFARX1 I_6222  ( .D(I108152), .CLK(I2350), .RSTB(I107951), .Q(I108169) );
nor I_6223 (I108186,I108169,I108050);
nand I_6224 (I107937,I108084,I108186);
not I_6225 (I107934,I108169);
and I_6226 (I108231,I108169,I108067);
DFFARX1 I_6227  ( .D(I108231), .CLK(I2350), .RSTB(I107951), .Q(I107919) );
DFFARX1 I_6228  ( .D(I108169), .CLK(I2350), .RSTB(I107951), .Q(I108262) );
and I_6229 (I107916,I108084,I108262);
nand I_6230 (I108293,I107968,I73080);
not I_6231 (I108310,I108293);
nor I_6232 (I108327,I108169,I108310);
DFFARX1 I_6233  ( .D(I73101), .CLK(I2350), .RSTB(I107951), .Q(I108344) );
nand I_6234 (I108361,I108344,I108293);
and I_6235 (I108378,I108084,I108361);
DFFARX1 I_6236  ( .D(I108378), .CLK(I2350), .RSTB(I107951), .Q(I107943) );
not I_6237 (I108409,I108344);
nand I_6238 (I107931,I108344,I108327);
nand I_6239 (I107925,I108344,I108310);
DFFARX1 I_6240  ( .D(I73098), .CLK(I2350), .RSTB(I107951), .Q(I108454) );
not I_6241 (I108471,I108454);
nor I_6242 (I107940,I108344,I108471);
nor I_6243 (I108502,I108471,I108409);
and I_6244 (I108519,I108050,I108502);
or I_6245 (I108536,I108293,I108519);
DFFARX1 I_6246  ( .D(I108536), .CLK(I2350), .RSTB(I107951), .Q(I107928) );
DFFARX1 I_6247  ( .D(I108471), .CLK(I2350), .RSTB(I107951), .Q(I107913) );
not I_6248 (I108614,I2357);
not I_6249 (I108631,I51777);
nor I_6250 (I108648,I51765,I51789);
nand I_6251 (I108665,I108648,I51774);
DFFARX1 I_6252  ( .D(I108665), .CLK(I2350), .RSTB(I108614), .Q(I108585) );
nor I_6253 (I108696,I108631,I51765);
nand I_6254 (I108713,I108696,I51792);
nand I_6255 (I108730,I108713,I108665);
not I_6256 (I108747,I51765);
not I_6257 (I108764,I51762);
nor I_6258 (I108781,I108764,I51771);
and I_6259 (I108798,I108781,I51786);
or I_6260 (I108815,I108798,I51768);
DFFARX1 I_6261  ( .D(I108815), .CLK(I2350), .RSTB(I108614), .Q(I108832) );
nor I_6262 (I108849,I108832,I108713);
nand I_6263 (I108600,I108747,I108849);
not I_6264 (I108597,I108832);
and I_6265 (I108894,I108832,I108730);
DFFARX1 I_6266  ( .D(I108894), .CLK(I2350), .RSTB(I108614), .Q(I108582) );
DFFARX1 I_6267  ( .D(I108832), .CLK(I2350), .RSTB(I108614), .Q(I108925) );
and I_6268 (I108579,I108747,I108925);
nand I_6269 (I108956,I108631,I51762);
not I_6270 (I108973,I108956);
nor I_6271 (I108990,I108832,I108973);
DFFARX1 I_6272  ( .D(I51783), .CLK(I2350), .RSTB(I108614), .Q(I109007) );
nand I_6273 (I109024,I109007,I108956);
and I_6274 (I109041,I108747,I109024);
DFFARX1 I_6275  ( .D(I109041), .CLK(I2350), .RSTB(I108614), .Q(I108606) );
not I_6276 (I109072,I109007);
nand I_6277 (I108594,I109007,I108990);
nand I_6278 (I108588,I109007,I108973);
DFFARX1 I_6279  ( .D(I51780), .CLK(I2350), .RSTB(I108614), .Q(I109117) );
not I_6280 (I109134,I109117);
nor I_6281 (I108603,I109007,I109134);
nor I_6282 (I109165,I109134,I109072);
and I_6283 (I109182,I108713,I109165);
or I_6284 (I109199,I108956,I109182);
DFFARX1 I_6285  ( .D(I109199), .CLK(I2350), .RSTB(I108614), .Q(I108591) );
DFFARX1 I_6286  ( .D(I109134), .CLK(I2350), .RSTB(I108614), .Q(I108576) );
not I_6287 (I109277,I2357);
not I_6288 (I109294,I310007);
nor I_6289 (I109311,I310019,I310022);
nand I_6290 (I109328,I109311,I310010);
DFFARX1 I_6291  ( .D(I109328), .CLK(I2350), .RSTB(I109277), .Q(I109248) );
nor I_6292 (I109359,I109294,I310019);
nand I_6293 (I109376,I109359,I309995);
nand I_6294 (I109393,I109376,I109328);
not I_6295 (I109410,I310019);
not I_6296 (I109427,I309998);
nor I_6297 (I109444,I109427,I310001);
and I_6298 (I109461,I109444,I310004);
or I_6299 (I109478,I109461,I310013);
DFFARX1 I_6300  ( .D(I109478), .CLK(I2350), .RSTB(I109277), .Q(I109495) );
nor I_6301 (I109512,I109495,I109376);
nand I_6302 (I109263,I109410,I109512);
not I_6303 (I109260,I109495);
and I_6304 (I109557,I109495,I109393);
DFFARX1 I_6305  ( .D(I109557), .CLK(I2350), .RSTB(I109277), .Q(I109245) );
DFFARX1 I_6306  ( .D(I109495), .CLK(I2350), .RSTB(I109277), .Q(I109588) );
and I_6307 (I109242,I109410,I109588);
nand I_6308 (I109619,I109294,I309998);
not I_6309 (I109636,I109619);
nor I_6310 (I109653,I109495,I109636);
DFFARX1 I_6311  ( .D(I310016), .CLK(I2350), .RSTB(I109277), .Q(I109670) );
nand I_6312 (I109687,I109670,I109619);
and I_6313 (I109704,I109410,I109687);
DFFARX1 I_6314  ( .D(I109704), .CLK(I2350), .RSTB(I109277), .Q(I109269) );
not I_6315 (I109735,I109670);
nand I_6316 (I109257,I109670,I109653);
nand I_6317 (I109251,I109670,I109636);
DFFARX1 I_6318  ( .D(I309992), .CLK(I2350), .RSTB(I109277), .Q(I109780) );
not I_6319 (I109797,I109780);
nor I_6320 (I109266,I109670,I109797);
nor I_6321 (I109828,I109797,I109735);
and I_6322 (I109845,I109376,I109828);
or I_6323 (I109862,I109619,I109845);
DFFARX1 I_6324  ( .D(I109862), .CLK(I2350), .RSTB(I109277), .Q(I109254) );
DFFARX1 I_6325  ( .D(I109797), .CLK(I2350), .RSTB(I109277), .Q(I109239) );
not I_6326 (I109940,I2357);
not I_6327 (I109957,I393197);
nor I_6328 (I109974,I393176,I393188);
nand I_6329 (I109991,I109974,I393182);
DFFARX1 I_6330  ( .D(I109991), .CLK(I2350), .RSTB(I109940), .Q(I109911) );
nor I_6331 (I110022,I109957,I393176);
nand I_6332 (I110039,I110022,I393203);
nand I_6333 (I110056,I110039,I109991);
not I_6334 (I110073,I393176);
not I_6335 (I110090,I393179);
nor I_6336 (I110107,I110090,I393191);
and I_6337 (I110124,I110107,I393194);
or I_6338 (I110141,I110124,I393200);
DFFARX1 I_6339  ( .D(I110141), .CLK(I2350), .RSTB(I109940), .Q(I110158) );
nor I_6340 (I110175,I110158,I110039);
nand I_6341 (I109926,I110073,I110175);
not I_6342 (I109923,I110158);
and I_6343 (I110220,I110158,I110056);
DFFARX1 I_6344  ( .D(I110220), .CLK(I2350), .RSTB(I109940), .Q(I109908) );
DFFARX1 I_6345  ( .D(I110158), .CLK(I2350), .RSTB(I109940), .Q(I110251) );
and I_6346 (I109905,I110073,I110251);
nand I_6347 (I110282,I109957,I393179);
not I_6348 (I110299,I110282);
nor I_6349 (I110316,I110158,I110299);
DFFARX1 I_6350  ( .D(I393173), .CLK(I2350), .RSTB(I109940), .Q(I110333) );
nand I_6351 (I110350,I110333,I110282);
and I_6352 (I110367,I110073,I110350);
DFFARX1 I_6353  ( .D(I110367), .CLK(I2350), .RSTB(I109940), .Q(I109932) );
not I_6354 (I110398,I110333);
nand I_6355 (I109920,I110333,I110316);
nand I_6356 (I109914,I110333,I110299);
DFFARX1 I_6357  ( .D(I393185), .CLK(I2350), .RSTB(I109940), .Q(I110443) );
not I_6358 (I110460,I110443);
nor I_6359 (I109929,I110333,I110460);
nor I_6360 (I110491,I110460,I110398);
and I_6361 (I110508,I110039,I110491);
or I_6362 (I110525,I110282,I110508);
DFFARX1 I_6363  ( .D(I110525), .CLK(I2350), .RSTB(I109940), .Q(I109917) );
DFFARX1 I_6364  ( .D(I110460), .CLK(I2350), .RSTB(I109940), .Q(I109902) );
not I_6365 (I110603,I2357);
not I_6366 (I110620,I286207);
nor I_6367 (I110637,I286219,I286222);
nand I_6368 (I110654,I110637,I286210);
DFFARX1 I_6369  ( .D(I110654), .CLK(I2350), .RSTB(I110603), .Q(I110574) );
nor I_6370 (I110685,I110620,I286219);
nand I_6371 (I110702,I110685,I286195);
nand I_6372 (I110719,I110702,I110654);
not I_6373 (I110736,I286219);
not I_6374 (I110753,I286198);
nor I_6375 (I110770,I110753,I286201);
and I_6376 (I110787,I110770,I286204);
or I_6377 (I110804,I110787,I286213);
DFFARX1 I_6378  ( .D(I110804), .CLK(I2350), .RSTB(I110603), .Q(I110821) );
nor I_6379 (I110838,I110821,I110702);
nand I_6380 (I110589,I110736,I110838);
not I_6381 (I110586,I110821);
and I_6382 (I110883,I110821,I110719);
DFFARX1 I_6383  ( .D(I110883), .CLK(I2350), .RSTB(I110603), .Q(I110571) );
DFFARX1 I_6384  ( .D(I110821), .CLK(I2350), .RSTB(I110603), .Q(I110914) );
and I_6385 (I110568,I110736,I110914);
nand I_6386 (I110945,I110620,I286198);
not I_6387 (I110962,I110945);
nor I_6388 (I110979,I110821,I110962);
DFFARX1 I_6389  ( .D(I286216), .CLK(I2350), .RSTB(I110603), .Q(I110996) );
nand I_6390 (I111013,I110996,I110945);
and I_6391 (I111030,I110736,I111013);
DFFARX1 I_6392  ( .D(I111030), .CLK(I2350), .RSTB(I110603), .Q(I110595) );
not I_6393 (I111061,I110996);
nand I_6394 (I110583,I110996,I110979);
nand I_6395 (I110577,I110996,I110962);
DFFARX1 I_6396  ( .D(I286192), .CLK(I2350), .RSTB(I110603), .Q(I111106) );
not I_6397 (I111123,I111106);
nor I_6398 (I110592,I110996,I111123);
nor I_6399 (I111154,I111123,I111061);
and I_6400 (I111171,I110702,I111154);
or I_6401 (I111188,I110945,I111171);
DFFARX1 I_6402  ( .D(I111188), .CLK(I2350), .RSTB(I110603), .Q(I110580) );
DFFARX1 I_6403  ( .D(I111123), .CLK(I2350), .RSTB(I110603), .Q(I110565) );
not I_6404 (I111266,I2357);
not I_6405 (I111283,I20327);
nor I_6406 (I111300,I20315,I20318);
nand I_6407 (I111317,I111300,I20333);
DFFARX1 I_6408  ( .D(I111317), .CLK(I2350), .RSTB(I111266), .Q(I111237) );
nor I_6409 (I111348,I111283,I20315);
nand I_6410 (I111365,I111348,I20324);
nand I_6411 (I111382,I111365,I111317);
not I_6412 (I111399,I20315);
not I_6413 (I111416,I20336);
nor I_6414 (I111433,I111416,I20312);
and I_6415 (I111450,I111433,I20321);
or I_6416 (I111467,I111450,I20330);
DFFARX1 I_6417  ( .D(I111467), .CLK(I2350), .RSTB(I111266), .Q(I111484) );
nor I_6418 (I111501,I111484,I111365);
nand I_6419 (I111252,I111399,I111501);
not I_6420 (I111249,I111484);
and I_6421 (I111546,I111484,I111382);
DFFARX1 I_6422  ( .D(I111546), .CLK(I2350), .RSTB(I111266), .Q(I111234) );
DFFARX1 I_6423  ( .D(I111484), .CLK(I2350), .RSTB(I111266), .Q(I111577) );
and I_6424 (I111231,I111399,I111577);
nand I_6425 (I111608,I111283,I20336);
not I_6426 (I111625,I111608);
nor I_6427 (I111642,I111484,I111625);
DFFARX1 I_6428  ( .D(I20342), .CLK(I2350), .RSTB(I111266), .Q(I111659) );
nand I_6429 (I111676,I111659,I111608);
and I_6430 (I111693,I111399,I111676);
DFFARX1 I_6431  ( .D(I111693), .CLK(I2350), .RSTB(I111266), .Q(I111258) );
not I_6432 (I111724,I111659);
nand I_6433 (I111246,I111659,I111642);
nand I_6434 (I111240,I111659,I111625);
DFFARX1 I_6435  ( .D(I20339), .CLK(I2350), .RSTB(I111266), .Q(I111769) );
not I_6436 (I111786,I111769);
nor I_6437 (I111255,I111659,I111786);
nor I_6438 (I111817,I111786,I111724);
and I_6439 (I111834,I111365,I111817);
or I_6440 (I111851,I111608,I111834);
DFFARX1 I_6441  ( .D(I111851), .CLK(I2350), .RSTB(I111266), .Q(I111243) );
DFFARX1 I_6442  ( .D(I111786), .CLK(I2350), .RSTB(I111266), .Q(I111228) );
not I_6443 (I111929,I2357);
not I_6444 (I111946,I126994);
nor I_6445 (I111963,I126976,I126970);
nand I_6446 (I111980,I111963,I126973);
DFFARX1 I_6447  ( .D(I111980), .CLK(I2350), .RSTB(I111929), .Q(I111900) );
nor I_6448 (I112011,I111946,I126976);
nand I_6449 (I112028,I112011,I126982);
nand I_6450 (I112045,I112028,I111980);
not I_6451 (I112062,I126976);
not I_6452 (I112079,I126991);
nor I_6453 (I112096,I112079,I126979);
and I_6454 (I112113,I112096,I126985);
or I_6455 (I112130,I112113,I127000);
DFFARX1 I_6456  ( .D(I112130), .CLK(I2350), .RSTB(I111929), .Q(I112147) );
nor I_6457 (I112164,I112147,I112028);
nand I_6458 (I111915,I112062,I112164);
not I_6459 (I111912,I112147);
and I_6460 (I112209,I112147,I112045);
DFFARX1 I_6461  ( .D(I112209), .CLK(I2350), .RSTB(I111929), .Q(I111897) );
DFFARX1 I_6462  ( .D(I112147), .CLK(I2350), .RSTB(I111929), .Q(I112240) );
and I_6463 (I111894,I112062,I112240);
nand I_6464 (I112271,I111946,I126991);
not I_6465 (I112288,I112271);
nor I_6466 (I112305,I112147,I112288);
DFFARX1 I_6467  ( .D(I126988), .CLK(I2350), .RSTB(I111929), .Q(I112322) );
nand I_6468 (I112339,I112322,I112271);
and I_6469 (I112356,I112062,I112339);
DFFARX1 I_6470  ( .D(I112356), .CLK(I2350), .RSTB(I111929), .Q(I111921) );
not I_6471 (I112387,I112322);
nand I_6472 (I111909,I112322,I112305);
nand I_6473 (I111903,I112322,I112288);
DFFARX1 I_6474  ( .D(I126997), .CLK(I2350), .RSTB(I111929), .Q(I112432) );
not I_6475 (I112449,I112432);
nor I_6476 (I111918,I112322,I112449);
nor I_6477 (I112480,I112449,I112387);
and I_6478 (I112497,I112028,I112480);
or I_6479 (I112514,I112271,I112497);
DFFARX1 I_6480  ( .D(I112514), .CLK(I2350), .RSTB(I111929), .Q(I111906) );
DFFARX1 I_6481  ( .D(I112449), .CLK(I2350), .RSTB(I111929), .Q(I111891) );
not I_6482 (I112592,I2357);
not I_6483 (I112609,I71157);
nor I_6484 (I112626,I71145,I71169);
nand I_6485 (I112643,I112626,I71154);
DFFARX1 I_6486  ( .D(I112643), .CLK(I2350), .RSTB(I112592), .Q(I112563) );
nor I_6487 (I112674,I112609,I71145);
nand I_6488 (I112691,I112674,I71172);
nand I_6489 (I112708,I112691,I112643);
not I_6490 (I112725,I71145);
not I_6491 (I112742,I71142);
nor I_6492 (I112759,I112742,I71151);
and I_6493 (I112776,I112759,I71166);
or I_6494 (I112793,I112776,I71148);
DFFARX1 I_6495  ( .D(I112793), .CLK(I2350), .RSTB(I112592), .Q(I112810) );
nor I_6496 (I112827,I112810,I112691);
nand I_6497 (I112578,I112725,I112827);
not I_6498 (I112575,I112810);
and I_6499 (I112872,I112810,I112708);
DFFARX1 I_6500  ( .D(I112872), .CLK(I2350), .RSTB(I112592), .Q(I112560) );
DFFARX1 I_6501  ( .D(I112810), .CLK(I2350), .RSTB(I112592), .Q(I112903) );
and I_6502 (I112557,I112725,I112903);
nand I_6503 (I112934,I112609,I71142);
not I_6504 (I112951,I112934);
nor I_6505 (I112968,I112810,I112951);
DFFARX1 I_6506  ( .D(I71163), .CLK(I2350), .RSTB(I112592), .Q(I112985) );
nand I_6507 (I113002,I112985,I112934);
and I_6508 (I113019,I112725,I113002);
DFFARX1 I_6509  ( .D(I113019), .CLK(I2350), .RSTB(I112592), .Q(I112584) );
not I_6510 (I113050,I112985);
nand I_6511 (I112572,I112985,I112968);
nand I_6512 (I112566,I112985,I112951);
DFFARX1 I_6513  ( .D(I71160), .CLK(I2350), .RSTB(I112592), .Q(I113095) );
not I_6514 (I113112,I113095);
nor I_6515 (I112581,I112985,I113112);
nor I_6516 (I113143,I113112,I113050);
and I_6517 (I113160,I112691,I113143);
or I_6518 (I113177,I112934,I113160);
DFFARX1 I_6519  ( .D(I113177), .CLK(I2350), .RSTB(I112592), .Q(I112569) );
DFFARX1 I_6520  ( .D(I113112), .CLK(I2350), .RSTB(I112592), .Q(I112554) );
not I_6521 (I113255,I2357);
not I_6522 (I113272,I16400);
nor I_6523 (I113289,I16388,I16391);
nand I_6524 (I113306,I113289,I16406);
DFFARX1 I_6525  ( .D(I113306), .CLK(I2350), .RSTB(I113255), .Q(I113226) );
nor I_6526 (I113337,I113272,I16388);
nand I_6527 (I113354,I113337,I16397);
nand I_6528 (I113371,I113354,I113306);
not I_6529 (I113388,I16388);
not I_6530 (I113405,I16409);
nor I_6531 (I113422,I113405,I16385);
and I_6532 (I113439,I113422,I16394);
or I_6533 (I113456,I113439,I16403);
DFFARX1 I_6534  ( .D(I113456), .CLK(I2350), .RSTB(I113255), .Q(I113473) );
nor I_6535 (I113490,I113473,I113354);
nand I_6536 (I113241,I113388,I113490);
not I_6537 (I113238,I113473);
and I_6538 (I113535,I113473,I113371);
DFFARX1 I_6539  ( .D(I113535), .CLK(I2350), .RSTB(I113255), .Q(I113223) );
DFFARX1 I_6540  ( .D(I113473), .CLK(I2350), .RSTB(I113255), .Q(I113566) );
and I_6541 (I113220,I113388,I113566);
nand I_6542 (I113597,I113272,I16409);
not I_6543 (I113614,I113597);
nor I_6544 (I113631,I113473,I113614);
DFFARX1 I_6545  ( .D(I16415), .CLK(I2350), .RSTB(I113255), .Q(I113648) );
nand I_6546 (I113665,I113648,I113597);
and I_6547 (I113682,I113388,I113665);
DFFARX1 I_6548  ( .D(I113682), .CLK(I2350), .RSTB(I113255), .Q(I113247) );
not I_6549 (I113713,I113648);
nand I_6550 (I113235,I113648,I113631);
nand I_6551 (I113229,I113648,I113614);
DFFARX1 I_6552  ( .D(I16412), .CLK(I2350), .RSTB(I113255), .Q(I113758) );
not I_6553 (I113775,I113758);
nor I_6554 (I113244,I113648,I113775);
nor I_6555 (I113806,I113775,I113713);
and I_6556 (I113823,I113354,I113806);
or I_6557 (I113840,I113597,I113823);
DFFARX1 I_6558  ( .D(I113840), .CLK(I2350), .RSTB(I113255), .Q(I113232) );
DFFARX1 I_6559  ( .D(I113775), .CLK(I2350), .RSTB(I113255), .Q(I113217) );
not I_6560 (I113918,I2357);
or I_6561 (I113935,I217275,I217272);
or I_6562 (I113952,I217257,I217275);
DFFARX1 I_6563  ( .D(I113952), .CLK(I2350), .RSTB(I113918), .Q(I113892) );
nor I_6564 (I113983,I217266,I217269);
not I_6565 (I114000,I113983);
not I_6566 (I114017,I217266);
and I_6567 (I114034,I114017,I217281);
nor I_6568 (I114051,I114034,I217272);
nor I_6569 (I114068,I217287,I217263);
DFFARX1 I_6570  ( .D(I114068), .CLK(I2350), .RSTB(I113918), .Q(I114085) );
nand I_6571 (I114102,I114085,I113935);
and I_6572 (I114119,I114051,I114102);
DFFARX1 I_6573  ( .D(I114119), .CLK(I2350), .RSTB(I113918), .Q(I113886) );
nor I_6574 (I114150,I217287,I217257);
DFFARX1 I_6575  ( .D(I114150), .CLK(I2350), .RSTB(I113918), .Q(I114167) );
and I_6576 (I113883,I113983,I114167);
DFFARX1 I_6577  ( .D(I217278), .CLK(I2350), .RSTB(I113918), .Q(I114198) );
and I_6578 (I114215,I114198,I217284);
DFFARX1 I_6579  ( .D(I114215), .CLK(I2350), .RSTB(I113918), .Q(I114232) );
not I_6580 (I113895,I114232);
DFFARX1 I_6581  ( .D(I114215), .CLK(I2350), .RSTB(I113918), .Q(I113880) );
DFFARX1 I_6582  ( .D(I217260), .CLK(I2350), .RSTB(I113918), .Q(I114277) );
not I_6583 (I114294,I114277);
nor I_6584 (I114311,I113952,I114294);
and I_6585 (I114328,I114215,I114311);
or I_6586 (I114345,I113935,I114328);
DFFARX1 I_6587  ( .D(I114345), .CLK(I2350), .RSTB(I113918), .Q(I113901) );
nor I_6588 (I114376,I114277,I114085);
nand I_6589 (I113910,I114051,I114376);
nor I_6590 (I114407,I114277,I114000);
nand I_6591 (I113904,I114150,I114407);
not I_6592 (I113907,I114277);
nand I_6593 (I113898,I114277,I114000);
DFFARX1 I_6594  ( .D(I114277), .CLK(I2350), .RSTB(I113918), .Q(I113889) );
not I_6595 (I114513,I2357);
or I_6596 (I114530,I75039,I75033);
or I_6597 (I114547,I75027,I75039);
DFFARX1 I_6598  ( .D(I114547), .CLK(I2350), .RSTB(I114513), .Q(I114487) );
nor I_6599 (I114578,I75045,I75036);
not I_6600 (I114595,I114578);
not I_6601 (I114612,I75045);
and I_6602 (I114629,I114612,I75042);
nor I_6603 (I114646,I114629,I75033);
nor I_6604 (I114663,I75018,I75024);
DFFARX1 I_6605  ( .D(I114663), .CLK(I2350), .RSTB(I114513), .Q(I114680) );
nand I_6606 (I114697,I114680,I114530);
and I_6607 (I114714,I114646,I114697);
DFFARX1 I_6608  ( .D(I114714), .CLK(I2350), .RSTB(I114513), .Q(I114481) );
nor I_6609 (I114745,I75018,I75027);
DFFARX1 I_6610  ( .D(I114745), .CLK(I2350), .RSTB(I114513), .Q(I114762) );
and I_6611 (I114478,I114578,I114762);
DFFARX1 I_6612  ( .D(I75030), .CLK(I2350), .RSTB(I114513), .Q(I114793) );
and I_6613 (I114810,I114793,I75048);
DFFARX1 I_6614  ( .D(I114810), .CLK(I2350), .RSTB(I114513), .Q(I114827) );
not I_6615 (I114490,I114827);
DFFARX1 I_6616  ( .D(I114810), .CLK(I2350), .RSTB(I114513), .Q(I114475) );
DFFARX1 I_6617  ( .D(I75021), .CLK(I2350), .RSTB(I114513), .Q(I114872) );
not I_6618 (I114889,I114872);
nor I_6619 (I114906,I114547,I114889);
and I_6620 (I114923,I114810,I114906);
or I_6621 (I114940,I114530,I114923);
DFFARX1 I_6622  ( .D(I114940), .CLK(I2350), .RSTB(I114513), .Q(I114496) );
nor I_6623 (I114971,I114872,I114680);
nand I_6624 (I114505,I114646,I114971);
nor I_6625 (I115002,I114872,I114595);
nand I_6626 (I114499,I114745,I115002);
not I_6627 (I114502,I114872);
nand I_6628 (I114493,I114872,I114595);
DFFARX1 I_6629  ( .D(I114872), .CLK(I2350), .RSTB(I114513), .Q(I114484) );
not I_6630 (I115108,I2357);
or I_6631 (I115125,I39509,I39503);
or I_6632 (I115142,I39497,I39509);
DFFARX1 I_6633  ( .D(I115142), .CLK(I2350), .RSTB(I115108), .Q(I115082) );
nor I_6634 (I115173,I39515,I39506);
not I_6635 (I115190,I115173);
not I_6636 (I115207,I39515);
and I_6637 (I115224,I115207,I39512);
nor I_6638 (I115241,I115224,I39503);
nor I_6639 (I115258,I39488,I39494);
DFFARX1 I_6640  ( .D(I115258), .CLK(I2350), .RSTB(I115108), .Q(I115275) );
nand I_6641 (I115292,I115275,I115125);
and I_6642 (I115309,I115241,I115292);
DFFARX1 I_6643  ( .D(I115309), .CLK(I2350), .RSTB(I115108), .Q(I115076) );
nor I_6644 (I115340,I39488,I39497);
DFFARX1 I_6645  ( .D(I115340), .CLK(I2350), .RSTB(I115108), .Q(I115357) );
and I_6646 (I115073,I115173,I115357);
DFFARX1 I_6647  ( .D(I39500), .CLK(I2350), .RSTB(I115108), .Q(I115388) );
and I_6648 (I115405,I115388,I39518);
DFFARX1 I_6649  ( .D(I115405), .CLK(I2350), .RSTB(I115108), .Q(I115422) );
not I_6650 (I115085,I115422);
DFFARX1 I_6651  ( .D(I115405), .CLK(I2350), .RSTB(I115108), .Q(I115070) );
DFFARX1 I_6652  ( .D(I39491), .CLK(I2350), .RSTB(I115108), .Q(I115467) );
not I_6653 (I115484,I115467);
nor I_6654 (I115501,I115142,I115484);
and I_6655 (I115518,I115405,I115501);
or I_6656 (I115535,I115125,I115518);
DFFARX1 I_6657  ( .D(I115535), .CLK(I2350), .RSTB(I115108), .Q(I115091) );
nor I_6658 (I115566,I115467,I115275);
nand I_6659 (I115100,I115241,I115566);
nor I_6660 (I115597,I115467,I115190);
nand I_6661 (I115094,I115340,I115597);
not I_6662 (I115097,I115467);
nand I_6663 (I115088,I115467,I115190);
DFFARX1 I_6664  ( .D(I115467), .CLK(I2350), .RSTB(I115108), .Q(I115079) );
not I_6665 (I115703,I2357);
or I_6666 (I115720,I143647,I143662);
or I_6667 (I115737,I143650,I143647);
DFFARX1 I_6668  ( .D(I115737), .CLK(I2350), .RSTB(I115703), .Q(I115677) );
nor I_6669 (I115768,I143653,I143668);
not I_6670 (I115785,I115768);
not I_6671 (I115802,I143653);
and I_6672 (I115819,I115802,I143656);
nor I_6673 (I115836,I115819,I143662);
nor I_6674 (I115853,I143659,I143677);
DFFARX1 I_6675  ( .D(I115853), .CLK(I2350), .RSTB(I115703), .Q(I115870) );
nand I_6676 (I115887,I115870,I115720);
and I_6677 (I115904,I115836,I115887);
DFFARX1 I_6678  ( .D(I115904), .CLK(I2350), .RSTB(I115703), .Q(I115671) );
nor I_6679 (I115935,I143659,I143650);
DFFARX1 I_6680  ( .D(I115935), .CLK(I2350), .RSTB(I115703), .Q(I115952) );
and I_6681 (I115668,I115768,I115952);
DFFARX1 I_6682  ( .D(I143674), .CLK(I2350), .RSTB(I115703), .Q(I115983) );
and I_6683 (I116000,I115983,I143665);
DFFARX1 I_6684  ( .D(I116000), .CLK(I2350), .RSTB(I115703), .Q(I116017) );
not I_6685 (I115680,I116017);
DFFARX1 I_6686  ( .D(I116000), .CLK(I2350), .RSTB(I115703), .Q(I115665) );
DFFARX1 I_6687  ( .D(I143671), .CLK(I2350), .RSTB(I115703), .Q(I116062) );
not I_6688 (I116079,I116062);
nor I_6689 (I116096,I115737,I116079);
and I_6690 (I116113,I116000,I116096);
or I_6691 (I116130,I115720,I116113);
DFFARX1 I_6692  ( .D(I116130), .CLK(I2350), .RSTB(I115703), .Q(I115686) );
nor I_6693 (I116161,I116062,I115870);
nand I_6694 (I115695,I115836,I116161);
nor I_6695 (I116192,I116062,I115785);
nand I_6696 (I115689,I115935,I116192);
not I_6697 (I115692,I116062);
nand I_6698 (I115683,I116062,I115785);
DFFARX1 I_6699  ( .D(I116062), .CLK(I2350), .RSTB(I115703), .Q(I115674) );
not I_6700 (I116298,I2357);
or I_6701 (I116315,I253361,I253346);
or I_6702 (I116332,I253358,I253361);
DFFARX1 I_6703  ( .D(I116332), .CLK(I2350), .RSTB(I116298), .Q(I116272) );
nor I_6704 (I116363,I253340,I253331);
not I_6705 (I116380,I116363);
not I_6706 (I116397,I253340);
and I_6707 (I116414,I116397,I253355);
nor I_6708 (I116431,I116414,I253346);
nor I_6709 (I116448,I253334,I253352);
DFFARX1 I_6710  ( .D(I116448), .CLK(I2350), .RSTB(I116298), .Q(I116465) );
nand I_6711 (I116482,I116465,I116315);
and I_6712 (I116499,I116431,I116482);
DFFARX1 I_6713  ( .D(I116499), .CLK(I2350), .RSTB(I116298), .Q(I116266) );
nor I_6714 (I116530,I253334,I253358);
DFFARX1 I_6715  ( .D(I116530), .CLK(I2350), .RSTB(I116298), .Q(I116547) );
and I_6716 (I116263,I116363,I116547);
DFFARX1 I_6717  ( .D(I253343), .CLK(I2350), .RSTB(I116298), .Q(I116578) );
and I_6718 (I116595,I116578,I253337);
DFFARX1 I_6719  ( .D(I116595), .CLK(I2350), .RSTB(I116298), .Q(I116612) );
not I_6720 (I116275,I116612);
DFFARX1 I_6721  ( .D(I116595), .CLK(I2350), .RSTB(I116298), .Q(I116260) );
DFFARX1 I_6722  ( .D(I253349), .CLK(I2350), .RSTB(I116298), .Q(I116657) );
not I_6723 (I116674,I116657);
nor I_6724 (I116691,I116332,I116674);
and I_6725 (I116708,I116595,I116691);
or I_6726 (I116725,I116315,I116708);
DFFARX1 I_6727  ( .D(I116725), .CLK(I2350), .RSTB(I116298), .Q(I116281) );
nor I_6728 (I116756,I116657,I116465);
nand I_6729 (I116290,I116431,I116756);
nor I_6730 (I116787,I116657,I116380);
nand I_6731 (I116284,I116530,I116787);
not I_6732 (I116287,I116657);
nand I_6733 (I116278,I116657,I116380);
DFFARX1 I_6734  ( .D(I116657), .CLK(I2350), .RSTB(I116298), .Q(I116269) );
not I_6735 (I116893,I2357);
or I_6736 (I116910,I2159,I1559);
or I_6737 (I116927,I1711,I2159);
DFFARX1 I_6738  ( .D(I116927), .CLK(I2350), .RSTB(I116893), .Q(I116867) );
nor I_6739 (I116958,I1687,I1735);
not I_6740 (I116975,I116958);
not I_6741 (I116992,I1687);
and I_6742 (I117009,I116992,I1455);
nor I_6743 (I117026,I117009,I1559);
nor I_6744 (I117043,I1583,I1759);
DFFARX1 I_6745  ( .D(I117043), .CLK(I2350), .RSTB(I116893), .Q(I117060) );
nand I_6746 (I117077,I117060,I116910);
and I_6747 (I117094,I117026,I117077);
DFFARX1 I_6748  ( .D(I117094), .CLK(I2350), .RSTB(I116893), .Q(I116861) );
nor I_6749 (I117125,I1583,I1711);
DFFARX1 I_6750  ( .D(I117125), .CLK(I2350), .RSTB(I116893), .Q(I117142) );
and I_6751 (I116858,I116958,I117142);
DFFARX1 I_6752  ( .D(I1303), .CLK(I2350), .RSTB(I116893), .Q(I117173) );
and I_6753 (I117190,I117173,I1943);
DFFARX1 I_6754  ( .D(I117190), .CLK(I2350), .RSTB(I116893), .Q(I117207) );
not I_6755 (I116870,I117207);
DFFARX1 I_6756  ( .D(I117190), .CLK(I2350), .RSTB(I116893), .Q(I116855) );
DFFARX1 I_6757  ( .D(I1743), .CLK(I2350), .RSTB(I116893), .Q(I117252) );
not I_6758 (I117269,I117252);
nor I_6759 (I117286,I116927,I117269);
and I_6760 (I117303,I117190,I117286);
or I_6761 (I117320,I116910,I117303);
DFFARX1 I_6762  ( .D(I117320), .CLK(I2350), .RSTB(I116893), .Q(I116876) );
nor I_6763 (I117351,I117252,I117060);
nand I_6764 (I116885,I117026,I117351);
nor I_6765 (I117382,I117252,I116975);
nand I_6766 (I116879,I117125,I117382);
not I_6767 (I116882,I117252);
nand I_6768 (I116873,I117252,I116975);
DFFARX1 I_6769  ( .D(I117252), .CLK(I2350), .RSTB(I116893), .Q(I116864) );
not I_6770 (I117488,I2357);
or I_6771 (I117505,I2119,I1895);
or I_6772 (I117522,I2111,I2119);
DFFARX1 I_6773  ( .D(I117522), .CLK(I2350), .RSTB(I117488), .Q(I117462) );
nor I_6774 (I117553,I2319,I1823);
not I_6775 (I117570,I117553);
not I_6776 (I117587,I2319);
and I_6777 (I117604,I117587,I1903);
nor I_6778 (I117621,I117604,I1895);
nor I_6779 (I117638,I1615,I1439);
DFFARX1 I_6780  ( .D(I117638), .CLK(I2350), .RSTB(I117488), .Q(I117655) );
nand I_6781 (I117672,I117655,I117505);
and I_6782 (I117689,I117621,I117672);
DFFARX1 I_6783  ( .D(I117689), .CLK(I2350), .RSTB(I117488), .Q(I117456) );
nor I_6784 (I117720,I1615,I2111);
DFFARX1 I_6785  ( .D(I117720), .CLK(I2350), .RSTB(I117488), .Q(I117737) );
and I_6786 (I117453,I117553,I117737);
DFFARX1 I_6787  ( .D(I2207), .CLK(I2350), .RSTB(I117488), .Q(I117768) );
and I_6788 (I117785,I117768,I2143);
DFFARX1 I_6789  ( .D(I117785), .CLK(I2350), .RSTB(I117488), .Q(I117802) );
not I_6790 (I117465,I117802);
DFFARX1 I_6791  ( .D(I117785), .CLK(I2350), .RSTB(I117488), .Q(I117450) );
DFFARX1 I_6792  ( .D(I1959), .CLK(I2350), .RSTB(I117488), .Q(I117847) );
not I_6793 (I117864,I117847);
nor I_6794 (I117881,I117522,I117864);
and I_6795 (I117898,I117785,I117881);
or I_6796 (I117915,I117505,I117898);
DFFARX1 I_6797  ( .D(I117915), .CLK(I2350), .RSTB(I117488), .Q(I117471) );
nor I_6798 (I117946,I117847,I117655);
nand I_6799 (I117480,I117621,I117946);
nor I_6800 (I117977,I117847,I117570);
nand I_6801 (I117474,I117720,I117977);
not I_6802 (I117477,I117847);
nand I_6803 (I117468,I117847,I117570);
DFFARX1 I_6804  ( .D(I117847), .CLK(I2350), .RSTB(I117488), .Q(I117459) );
not I_6805 (I118083,I2357);
or I_6806 (I118100,I315359,I315353);
or I_6807 (I118117,I315347,I315359);
DFFARX1 I_6808  ( .D(I118117), .CLK(I2350), .RSTB(I118083), .Q(I118057) );
nor I_6809 (I118148,I315350,I315356);
not I_6810 (I118165,I118148);
not I_6811 (I118182,I315350);
and I_6812 (I118199,I118182,I315374);
nor I_6813 (I118216,I118199,I315353);
nor I_6814 (I118233,I315377,I315368);
DFFARX1 I_6815  ( .D(I118233), .CLK(I2350), .RSTB(I118083), .Q(I118250) );
nand I_6816 (I118267,I118250,I118100);
and I_6817 (I118284,I118216,I118267);
DFFARX1 I_6818  ( .D(I118284), .CLK(I2350), .RSTB(I118083), .Q(I118051) );
nor I_6819 (I118315,I315377,I315347);
DFFARX1 I_6820  ( .D(I118315), .CLK(I2350), .RSTB(I118083), .Q(I118332) );
and I_6821 (I118048,I118148,I118332);
DFFARX1 I_6822  ( .D(I315365), .CLK(I2350), .RSTB(I118083), .Q(I118363) );
and I_6823 (I118380,I118363,I315362);
DFFARX1 I_6824  ( .D(I118380), .CLK(I2350), .RSTB(I118083), .Q(I118397) );
not I_6825 (I118060,I118397);
DFFARX1 I_6826  ( .D(I118380), .CLK(I2350), .RSTB(I118083), .Q(I118045) );
DFFARX1 I_6827  ( .D(I315371), .CLK(I2350), .RSTB(I118083), .Q(I118442) );
not I_6828 (I118459,I118442);
nor I_6829 (I118476,I118117,I118459);
and I_6830 (I118493,I118380,I118476);
or I_6831 (I118510,I118100,I118493);
DFFARX1 I_6832  ( .D(I118510), .CLK(I2350), .RSTB(I118083), .Q(I118066) );
nor I_6833 (I118541,I118442,I118250);
nand I_6834 (I118075,I118216,I118541);
nor I_6835 (I118572,I118442,I118165);
nand I_6836 (I118069,I118315,I118572);
not I_6837 (I118072,I118442);
nand I_6838 (I118063,I118442,I118165);
DFFARX1 I_6839  ( .D(I118442), .CLK(I2350), .RSTB(I118083), .Q(I118054) );
not I_6840 (I118678,I2357);
or I_6841 (I118695,I222443,I222440);
or I_6842 (I118712,I222425,I222443);
DFFARX1 I_6843  ( .D(I118712), .CLK(I2350), .RSTB(I118678), .Q(I118652) );
nor I_6844 (I118743,I222434,I222437);
not I_6845 (I118760,I118743);
not I_6846 (I118777,I222434);
and I_6847 (I118794,I118777,I222449);
nor I_6848 (I118811,I118794,I222440);
nor I_6849 (I118828,I222455,I222431);
DFFARX1 I_6850  ( .D(I118828), .CLK(I2350), .RSTB(I118678), .Q(I118845) );
nand I_6851 (I118862,I118845,I118695);
and I_6852 (I118879,I118811,I118862);
DFFARX1 I_6853  ( .D(I118879), .CLK(I2350), .RSTB(I118678), .Q(I118646) );
nor I_6854 (I118910,I222455,I222425);
DFFARX1 I_6855  ( .D(I118910), .CLK(I2350), .RSTB(I118678), .Q(I118927) );
and I_6856 (I118643,I118743,I118927);
DFFARX1 I_6857  ( .D(I222446), .CLK(I2350), .RSTB(I118678), .Q(I118958) );
and I_6858 (I118975,I118958,I222452);
DFFARX1 I_6859  ( .D(I118975), .CLK(I2350), .RSTB(I118678), .Q(I118992) );
not I_6860 (I118655,I118992);
DFFARX1 I_6861  ( .D(I118975), .CLK(I2350), .RSTB(I118678), .Q(I118640) );
DFFARX1 I_6862  ( .D(I222428), .CLK(I2350), .RSTB(I118678), .Q(I119037) );
not I_6863 (I119054,I119037);
nor I_6864 (I119071,I118712,I119054);
and I_6865 (I119088,I118975,I119071);
or I_6866 (I119105,I118695,I119088);
DFFARX1 I_6867  ( .D(I119105), .CLK(I2350), .RSTB(I118678), .Q(I118661) );
nor I_6868 (I119136,I119037,I118845);
nand I_6869 (I118670,I118811,I119136);
nor I_6870 (I119167,I119037,I118760);
nand I_6871 (I118664,I118910,I119167);
not I_6872 (I118667,I119037);
nand I_6873 (I118658,I119037,I118760);
DFFARX1 I_6874  ( .D(I119037), .CLK(I2350), .RSTB(I118678), .Q(I118649) );
not I_6875 (I119273,I2357);
or I_6876 (I119290,I18650,I18659);
or I_6877 (I119307,I18653,I18650);
DFFARX1 I_6878  ( .D(I119307), .CLK(I2350), .RSTB(I119273), .Q(I119247) );
nor I_6879 (I119338,I18629,I18632);
not I_6880 (I119355,I119338);
not I_6881 (I119372,I18629);
and I_6882 (I119389,I119372,I18641);
nor I_6883 (I119406,I119389,I18659);
nor I_6884 (I119423,I18647,I18638);
DFFARX1 I_6885  ( .D(I119423), .CLK(I2350), .RSTB(I119273), .Q(I119440) );
nand I_6886 (I119457,I119440,I119290);
and I_6887 (I119474,I119406,I119457);
DFFARX1 I_6888  ( .D(I119474), .CLK(I2350), .RSTB(I119273), .Q(I119241) );
nor I_6889 (I119505,I18647,I18653);
DFFARX1 I_6890  ( .D(I119505), .CLK(I2350), .RSTB(I119273), .Q(I119522) );
and I_6891 (I119238,I119338,I119522);
DFFARX1 I_6892  ( .D(I18644), .CLK(I2350), .RSTB(I119273), .Q(I119553) );
and I_6893 (I119570,I119553,I18635);
DFFARX1 I_6894  ( .D(I119570), .CLK(I2350), .RSTB(I119273), .Q(I119587) );
not I_6895 (I119250,I119587);
DFFARX1 I_6896  ( .D(I119570), .CLK(I2350), .RSTB(I119273), .Q(I119235) );
DFFARX1 I_6897  ( .D(I18656), .CLK(I2350), .RSTB(I119273), .Q(I119632) );
not I_6898 (I119649,I119632);
nor I_6899 (I119666,I119307,I119649);
and I_6900 (I119683,I119570,I119666);
or I_6901 (I119700,I119290,I119683);
DFFARX1 I_6902  ( .D(I119700), .CLK(I2350), .RSTB(I119273), .Q(I119256) );
nor I_6903 (I119731,I119632,I119440);
nand I_6904 (I119265,I119406,I119731);
nor I_6905 (I119762,I119632,I119355);
nand I_6906 (I119259,I119505,I119762);
not I_6907 (I119262,I119632);
nand I_6908 (I119253,I119632,I119355);
DFFARX1 I_6909  ( .D(I119632), .CLK(I2350), .RSTB(I119273), .Q(I119244) );
not I_6910 (I119868,I2357);
or I_6911 (I119885,I83437,I83431);
or I_6912 (I119902,I83425,I83437);
DFFARX1 I_6913  ( .D(I119902), .CLK(I2350), .RSTB(I119868), .Q(I119842) );
nor I_6914 (I119933,I83443,I83434);
not I_6915 (I119950,I119933);
not I_6916 (I119967,I83443);
and I_6917 (I119984,I119967,I83440);
nor I_6918 (I120001,I119984,I83431);
nor I_6919 (I120018,I83416,I83422);
DFFARX1 I_6920  ( .D(I120018), .CLK(I2350), .RSTB(I119868), .Q(I120035) );
nand I_6921 (I120052,I120035,I119885);
and I_6922 (I120069,I120001,I120052);
DFFARX1 I_6923  ( .D(I120069), .CLK(I2350), .RSTB(I119868), .Q(I119836) );
nor I_6924 (I120100,I83416,I83425);
DFFARX1 I_6925  ( .D(I120100), .CLK(I2350), .RSTB(I119868), .Q(I120117) );
and I_6926 (I119833,I119933,I120117);
DFFARX1 I_6927  ( .D(I83428), .CLK(I2350), .RSTB(I119868), .Q(I120148) );
and I_6928 (I120165,I120148,I83446);
DFFARX1 I_6929  ( .D(I120165), .CLK(I2350), .RSTB(I119868), .Q(I120182) );
not I_6930 (I119845,I120182);
DFFARX1 I_6931  ( .D(I120165), .CLK(I2350), .RSTB(I119868), .Q(I119830) );
DFFARX1 I_6932  ( .D(I83419), .CLK(I2350), .RSTB(I119868), .Q(I120227) );
not I_6933 (I120244,I120227);
nor I_6934 (I120261,I119902,I120244);
and I_6935 (I120278,I120165,I120261);
or I_6936 (I120295,I119885,I120278);
DFFARX1 I_6937  ( .D(I120295), .CLK(I2350), .RSTB(I119868), .Q(I119851) );
nor I_6938 (I120326,I120227,I120035);
nand I_6939 (I119860,I120001,I120326);
nor I_6940 (I120357,I120227,I119950);
nand I_6941 (I119854,I120100,I120357);
not I_6942 (I119857,I120227);
nand I_6943 (I119848,I120227,I119950);
DFFARX1 I_6944  ( .D(I120227), .CLK(I2350), .RSTB(I119868), .Q(I119839) );
not I_6945 (I120463,I2357);
or I_6946 (I120480,I152266,I152281);
or I_6947 (I120497,I152269,I152266);
DFFARX1 I_6948  ( .D(I120497), .CLK(I2350), .RSTB(I120463), .Q(I120437) );
nor I_6949 (I120528,I152272,I152287);
not I_6950 (I120545,I120528);
not I_6951 (I120562,I152272);
and I_6952 (I120579,I120562,I152275);
nor I_6953 (I120596,I120579,I152281);
nor I_6954 (I120613,I152278,I152296);
DFFARX1 I_6955  ( .D(I120613), .CLK(I2350), .RSTB(I120463), .Q(I120630) );
nand I_6956 (I120647,I120630,I120480);
and I_6957 (I120664,I120596,I120647);
DFFARX1 I_6958  ( .D(I120664), .CLK(I2350), .RSTB(I120463), .Q(I120431) );
nor I_6959 (I120695,I152278,I152269);
DFFARX1 I_6960  ( .D(I120695), .CLK(I2350), .RSTB(I120463), .Q(I120712) );
and I_6961 (I120428,I120528,I120712);
DFFARX1 I_6962  ( .D(I152293), .CLK(I2350), .RSTB(I120463), .Q(I120743) );
and I_6963 (I120760,I120743,I152284);
DFFARX1 I_6964  ( .D(I120760), .CLK(I2350), .RSTB(I120463), .Q(I120777) );
not I_6965 (I120440,I120777);
DFFARX1 I_6966  ( .D(I120760), .CLK(I2350), .RSTB(I120463), .Q(I120425) );
DFFARX1 I_6967  ( .D(I152290), .CLK(I2350), .RSTB(I120463), .Q(I120822) );
not I_6968 (I120839,I120822);
nor I_6969 (I120856,I120497,I120839);
and I_6970 (I120873,I120760,I120856);
or I_6971 (I120890,I120480,I120873);
DFFARX1 I_6972  ( .D(I120890), .CLK(I2350), .RSTB(I120463), .Q(I120446) );
nor I_6973 (I120921,I120822,I120630);
nand I_6974 (I120455,I120596,I120921);
nor I_6975 (I120952,I120822,I120545);
nand I_6976 (I120449,I120695,I120952);
not I_6977 (I120452,I120822);
nand I_6978 (I120443,I120822,I120545);
DFFARX1 I_6979  ( .D(I120822), .CLK(I2350), .RSTB(I120463), .Q(I120434) );
not I_6980 (I121058,I2357);
or I_6981 (I121075,I347701,I347698);
or I_6982 (I121092,I347728,I347701);
DFFARX1 I_6983  ( .D(I121092), .CLK(I2350), .RSTB(I121058), .Q(I121032) );
nor I_6984 (I121123,I347707,I347713);
not I_6985 (I121140,I121123);
not I_6986 (I121157,I347707);
and I_6987 (I121174,I121157,I347704);
nor I_6988 (I121191,I121174,I347698);
nor I_6989 (I121208,I347716,I347725);
DFFARX1 I_6990  ( .D(I121208), .CLK(I2350), .RSTB(I121058), .Q(I121225) );
nand I_6991 (I121242,I121225,I121075);
and I_6992 (I121259,I121191,I121242);
DFFARX1 I_6993  ( .D(I121259), .CLK(I2350), .RSTB(I121058), .Q(I121026) );
nor I_6994 (I121290,I347716,I347728);
DFFARX1 I_6995  ( .D(I121290), .CLK(I2350), .RSTB(I121058), .Q(I121307) );
and I_6996 (I121023,I121123,I121307);
DFFARX1 I_6997  ( .D(I347719), .CLK(I2350), .RSTB(I121058), .Q(I121338) );
and I_6998 (I121355,I121338,I347710);
DFFARX1 I_6999  ( .D(I121355), .CLK(I2350), .RSTB(I121058), .Q(I121372) );
not I_7000 (I121035,I121372);
DFFARX1 I_7001  ( .D(I121355), .CLK(I2350), .RSTB(I121058), .Q(I121020) );
DFFARX1 I_7002  ( .D(I347722), .CLK(I2350), .RSTB(I121058), .Q(I121417) );
not I_7003 (I121434,I121417);
nor I_7004 (I121451,I121092,I121434);
and I_7005 (I121468,I121355,I121451);
or I_7006 (I121485,I121075,I121468);
DFFARX1 I_7007  ( .D(I121485), .CLK(I2350), .RSTB(I121058), .Q(I121041) );
nor I_7008 (I121516,I121417,I121225);
nand I_7009 (I121050,I121191,I121516);
nor I_7010 (I121547,I121417,I121140);
nand I_7011 (I121044,I121290,I121547);
not I_7012 (I121047,I121417);
nand I_7013 (I121038,I121417,I121140);
DFFARX1 I_7014  ( .D(I121417), .CLK(I2350), .RSTB(I121058), .Q(I121029) );
not I_7015 (I121653,I2357);
or I_7016 (I121670,I327854,I327848);
or I_7017 (I121687,I327842,I327854);
DFFARX1 I_7018  ( .D(I121687), .CLK(I2350), .RSTB(I121653), .Q(I121627) );
nor I_7019 (I121718,I327845,I327851);
not I_7020 (I121735,I121718);
not I_7021 (I121752,I327845);
and I_7022 (I121769,I121752,I327869);
nor I_7023 (I121786,I121769,I327848);
nor I_7024 (I121803,I327872,I327863);
DFFARX1 I_7025  ( .D(I121803), .CLK(I2350), .RSTB(I121653), .Q(I121820) );
nand I_7026 (I121837,I121820,I121670);
and I_7027 (I121854,I121786,I121837);
DFFARX1 I_7028  ( .D(I121854), .CLK(I2350), .RSTB(I121653), .Q(I121621) );
nor I_7029 (I121885,I327872,I327842);
DFFARX1 I_7030  ( .D(I121885), .CLK(I2350), .RSTB(I121653), .Q(I121902) );
and I_7031 (I121618,I121718,I121902);
DFFARX1 I_7032  ( .D(I327860), .CLK(I2350), .RSTB(I121653), .Q(I121933) );
and I_7033 (I121950,I121933,I327857);
DFFARX1 I_7034  ( .D(I121950), .CLK(I2350), .RSTB(I121653), .Q(I121967) );
not I_7035 (I121630,I121967);
DFFARX1 I_7036  ( .D(I121950), .CLK(I2350), .RSTB(I121653), .Q(I121615) );
DFFARX1 I_7037  ( .D(I327866), .CLK(I2350), .RSTB(I121653), .Q(I122012) );
not I_7038 (I122029,I122012);
nor I_7039 (I122046,I121687,I122029);
and I_7040 (I122063,I121950,I122046);
or I_7041 (I122080,I121670,I122063);
DFFARX1 I_7042  ( .D(I122080), .CLK(I2350), .RSTB(I121653), .Q(I121636) );
nor I_7043 (I122111,I122012,I121820);
nand I_7044 (I121645,I121786,I122111);
nor I_7045 (I122142,I122012,I121735);
nand I_7046 (I121639,I121885,I122142);
not I_7047 (I121642,I122012);
nand I_7048 (I121633,I122012,I121735);
DFFARX1 I_7049  ( .D(I122012), .CLK(I2350), .RSTB(I121653), .Q(I121624) );
not I_7050 (I122248,I2357);
or I_7051 (I122265,I88053,I88038);
or I_7052 (I122282,I88035,I88053);
DFFARX1 I_7053  ( .D(I122282), .CLK(I2350), .RSTB(I122248), .Q(I122222) );
nor I_7054 (I122313,I88023,I88032);
not I_7055 (I122330,I122313);
not I_7056 (I122347,I88023);
and I_7057 (I122364,I122347,I88047);
nor I_7058 (I122381,I122364,I88038);
nor I_7059 (I122398,I88026,I88041);
DFFARX1 I_7060  ( .D(I122398), .CLK(I2350), .RSTB(I122248), .Q(I122415) );
nand I_7061 (I122432,I122415,I122265);
and I_7062 (I122449,I122381,I122432);
DFFARX1 I_7063  ( .D(I122449), .CLK(I2350), .RSTB(I122248), .Q(I122216) );
nor I_7064 (I122480,I88026,I88035);
DFFARX1 I_7065  ( .D(I122480), .CLK(I2350), .RSTB(I122248), .Q(I122497) );
and I_7066 (I122213,I122313,I122497);
DFFARX1 I_7067  ( .D(I88029), .CLK(I2350), .RSTB(I122248), .Q(I122528) );
and I_7068 (I122545,I122528,I88050);
DFFARX1 I_7069  ( .D(I122545), .CLK(I2350), .RSTB(I122248), .Q(I122562) );
not I_7070 (I122225,I122562);
DFFARX1 I_7071  ( .D(I122545), .CLK(I2350), .RSTB(I122248), .Q(I122210) );
DFFARX1 I_7072  ( .D(I88044), .CLK(I2350), .RSTB(I122248), .Q(I122607) );
not I_7073 (I122624,I122607);
nor I_7074 (I122641,I122282,I122624);
and I_7075 (I122658,I122545,I122641);
or I_7076 (I122675,I122265,I122658);
DFFARX1 I_7077  ( .D(I122675), .CLK(I2350), .RSTB(I122248), .Q(I122231) );
nor I_7078 (I122706,I122607,I122415);
nand I_7079 (I122240,I122381,I122706);
nor I_7080 (I122737,I122607,I122330);
nand I_7081 (I122234,I122480,I122737);
not I_7082 (I122237,I122607);
nand I_7083 (I122228,I122607,I122330);
DFFARX1 I_7084  ( .D(I122607), .CLK(I2350), .RSTB(I122248), .Q(I122219) );
not I_7085 (I122843,I2357);
or I_7086 (I122860,I225027,I225024);
or I_7087 (I122877,I225009,I225027);
DFFARX1 I_7088  ( .D(I122877), .CLK(I2350), .RSTB(I122843), .Q(I122817) );
nor I_7089 (I122908,I225018,I225021);
not I_7090 (I122925,I122908);
not I_7091 (I122942,I225018);
and I_7092 (I122959,I122942,I225033);
nor I_7093 (I122976,I122959,I225024);
nor I_7094 (I122993,I225039,I225015);
DFFARX1 I_7095  ( .D(I122993), .CLK(I2350), .RSTB(I122843), .Q(I123010) );
nand I_7096 (I123027,I123010,I122860);
and I_7097 (I123044,I122976,I123027);
DFFARX1 I_7098  ( .D(I123044), .CLK(I2350), .RSTB(I122843), .Q(I122811) );
nor I_7099 (I123075,I225039,I225009);
DFFARX1 I_7100  ( .D(I123075), .CLK(I2350), .RSTB(I122843), .Q(I123092) );
and I_7101 (I122808,I122908,I123092);
DFFARX1 I_7102  ( .D(I225030), .CLK(I2350), .RSTB(I122843), .Q(I123123) );
and I_7103 (I123140,I123123,I225036);
DFFARX1 I_7104  ( .D(I123140), .CLK(I2350), .RSTB(I122843), .Q(I123157) );
not I_7105 (I122820,I123157);
DFFARX1 I_7106  ( .D(I123140), .CLK(I2350), .RSTB(I122843), .Q(I122805) );
DFFARX1 I_7107  ( .D(I225012), .CLK(I2350), .RSTB(I122843), .Q(I123202) );
not I_7108 (I123219,I123202);
nor I_7109 (I123236,I122877,I123219);
and I_7110 (I123253,I123140,I123236);
or I_7111 (I123270,I122860,I123253);
DFFARX1 I_7112  ( .D(I123270), .CLK(I2350), .RSTB(I122843), .Q(I122826) );
nor I_7113 (I123301,I123202,I123010);
nand I_7114 (I122835,I122976,I123301);
nor I_7115 (I123332,I123202,I122925);
nand I_7116 (I122829,I123075,I123332);
not I_7117 (I122832,I123202);
nand I_7118 (I122823,I123202,I122925);
DFFARX1 I_7119  ( .D(I123202), .CLK(I2350), .RSTB(I122843), .Q(I122814) );
not I_7120 (I123438,I2357);
or I_7121 (I123455,I1599,I1383);
or I_7122 (I123472,I2271,I1599);
DFFARX1 I_7123  ( .D(I123472), .CLK(I2350), .RSTB(I123438), .Q(I123412) );
nor I_7124 (I123503,I1503,I1951);
not I_7125 (I123520,I123503);
not I_7126 (I123537,I1503);
and I_7127 (I123554,I123537,I2007);
nor I_7128 (I123571,I123554,I1383);
nor I_7129 (I123588,I1935,I1783);
DFFARX1 I_7130  ( .D(I123588), .CLK(I2350), .RSTB(I123438), .Q(I123605) );
nand I_7131 (I123622,I123605,I123455);
and I_7132 (I123639,I123571,I123622);
DFFARX1 I_7133  ( .D(I123639), .CLK(I2350), .RSTB(I123438), .Q(I123406) );
nor I_7134 (I123670,I1935,I2271);
DFFARX1 I_7135  ( .D(I123670), .CLK(I2350), .RSTB(I123438), .Q(I123687) );
and I_7136 (I123403,I123503,I123687);
DFFARX1 I_7137  ( .D(I1655), .CLK(I2350), .RSTB(I123438), .Q(I123718) );
and I_7138 (I123735,I123718,I1535);
DFFARX1 I_7139  ( .D(I123735), .CLK(I2350), .RSTB(I123438), .Q(I123752) );
not I_7140 (I123415,I123752);
DFFARX1 I_7141  ( .D(I123735), .CLK(I2350), .RSTB(I123438), .Q(I123400) );
DFFARX1 I_7142  ( .D(I2279), .CLK(I2350), .RSTB(I123438), .Q(I123797) );
not I_7143 (I123814,I123797);
nor I_7144 (I123831,I123472,I123814);
and I_7145 (I123848,I123735,I123831);
or I_7146 (I123865,I123455,I123848);
DFFARX1 I_7147  ( .D(I123865), .CLK(I2350), .RSTB(I123438), .Q(I123421) );
nor I_7148 (I123896,I123797,I123605);
nand I_7149 (I123430,I123571,I123896);
nor I_7150 (I123927,I123797,I123520);
nand I_7151 (I123424,I123670,I123927);
not I_7152 (I123427,I123797);
nand I_7153 (I123418,I123797,I123520);
DFFARX1 I_7154  ( .D(I123797), .CLK(I2350), .RSTB(I123438), .Q(I123409) );
not I_7155 (I124033,I2357);
or I_7156 (I124050,I73747,I73741);
or I_7157 (I124067,I73735,I73747);
DFFARX1 I_7158  ( .D(I124067), .CLK(I2350), .RSTB(I124033), .Q(I124007) );
nor I_7159 (I124098,I73753,I73744);
not I_7160 (I124115,I124098);
not I_7161 (I124132,I73753);
and I_7162 (I124149,I124132,I73750);
nor I_7163 (I124166,I124149,I73741);
nor I_7164 (I124183,I73726,I73732);
DFFARX1 I_7165  ( .D(I124183), .CLK(I2350), .RSTB(I124033), .Q(I124200) );
nand I_7166 (I124217,I124200,I124050);
and I_7167 (I124234,I124166,I124217);
DFFARX1 I_7168  ( .D(I124234), .CLK(I2350), .RSTB(I124033), .Q(I124001) );
nor I_7169 (I124265,I73726,I73735);
DFFARX1 I_7170  ( .D(I124265), .CLK(I2350), .RSTB(I124033), .Q(I124282) );
and I_7171 (I123998,I124098,I124282);
DFFARX1 I_7172  ( .D(I73738), .CLK(I2350), .RSTB(I124033), .Q(I124313) );
and I_7173 (I124330,I124313,I73756);
DFFARX1 I_7174  ( .D(I124330), .CLK(I2350), .RSTB(I124033), .Q(I124347) );
not I_7175 (I124010,I124347);
DFFARX1 I_7176  ( .D(I124330), .CLK(I2350), .RSTB(I124033), .Q(I123995) );
DFFARX1 I_7177  ( .D(I73729), .CLK(I2350), .RSTB(I124033), .Q(I124392) );
not I_7178 (I124409,I124392);
nor I_7179 (I124426,I124067,I124409);
and I_7180 (I124443,I124330,I124426);
or I_7181 (I124460,I124050,I124443);
DFFARX1 I_7182  ( .D(I124460), .CLK(I2350), .RSTB(I124033), .Q(I124016) );
nor I_7183 (I124491,I124392,I124200);
nand I_7184 (I124025,I124166,I124491);
nor I_7185 (I124522,I124392,I124115);
nand I_7186 (I124019,I124265,I124522);
not I_7187 (I124022,I124392);
nand I_7188 (I124013,I124392,I124115);
DFFARX1 I_7189  ( .D(I124392), .CLK(I2350), .RSTB(I124033), .Q(I124004) );
not I_7190 (I124628,I2357);
or I_7191 (I124645,I54367,I54361);
or I_7192 (I124662,I54355,I54367);
DFFARX1 I_7193  ( .D(I124662), .CLK(I2350), .RSTB(I124628), .Q(I124602) );
nor I_7194 (I124693,I54373,I54364);
not I_7195 (I124710,I124693);
not I_7196 (I124727,I54373);
and I_7197 (I124744,I124727,I54370);
nor I_7198 (I124761,I124744,I54361);
nor I_7199 (I124778,I54346,I54352);
DFFARX1 I_7200  ( .D(I124778), .CLK(I2350), .RSTB(I124628), .Q(I124795) );
nand I_7201 (I124812,I124795,I124645);
and I_7202 (I124829,I124761,I124812);
DFFARX1 I_7203  ( .D(I124829), .CLK(I2350), .RSTB(I124628), .Q(I124596) );
nor I_7204 (I124860,I54346,I54355);
DFFARX1 I_7205  ( .D(I124860), .CLK(I2350), .RSTB(I124628), .Q(I124877) );
and I_7206 (I124593,I124693,I124877);
DFFARX1 I_7207  ( .D(I54358), .CLK(I2350), .RSTB(I124628), .Q(I124908) );
and I_7208 (I124925,I124908,I54376);
DFFARX1 I_7209  ( .D(I124925), .CLK(I2350), .RSTB(I124628), .Q(I124942) );
not I_7210 (I124605,I124942);
DFFARX1 I_7211  ( .D(I124925), .CLK(I2350), .RSTB(I124628), .Q(I124590) );
DFFARX1 I_7212  ( .D(I54349), .CLK(I2350), .RSTB(I124628), .Q(I124987) );
not I_7213 (I125004,I124987);
nor I_7214 (I125021,I124662,I125004);
and I_7215 (I125038,I124925,I125021);
or I_7216 (I125055,I124645,I125038);
DFFARX1 I_7217  ( .D(I125055), .CLK(I2350), .RSTB(I124628), .Q(I124611) );
nor I_7218 (I125086,I124987,I124795);
nand I_7219 (I124620,I124761,I125086);
nor I_7220 (I125117,I124987,I124710);
nand I_7221 (I124614,I124860,I125117);
not I_7222 (I124617,I124987);
nand I_7223 (I124608,I124987,I124710);
DFFARX1 I_7224  ( .D(I124987), .CLK(I2350), .RSTB(I124628), .Q(I124599) );
not I_7225 (I125223,I2357);
or I_7226 (I125240,I380409,I380406);
or I_7227 (I125257,I380436,I380409);
DFFARX1 I_7228  ( .D(I125257), .CLK(I2350), .RSTB(I125223), .Q(I125197) );
nor I_7229 (I125288,I380415,I380421);
not I_7230 (I125305,I125288);
not I_7231 (I125322,I380415);
and I_7232 (I125339,I125322,I380412);
nor I_7233 (I125356,I125339,I380406);
nor I_7234 (I125373,I380424,I380433);
DFFARX1 I_7235  ( .D(I125373), .CLK(I2350), .RSTB(I125223), .Q(I125390) );
nand I_7236 (I125407,I125390,I125240);
and I_7237 (I125424,I125356,I125407);
DFFARX1 I_7238  ( .D(I125424), .CLK(I2350), .RSTB(I125223), .Q(I125191) );
nor I_7239 (I125455,I380424,I380436);
DFFARX1 I_7240  ( .D(I125455), .CLK(I2350), .RSTB(I125223), .Q(I125472) );
and I_7241 (I125188,I125288,I125472);
DFFARX1 I_7242  ( .D(I380427), .CLK(I2350), .RSTB(I125223), .Q(I125503) );
and I_7243 (I125520,I125503,I380418);
DFFARX1 I_7244  ( .D(I125520), .CLK(I2350), .RSTB(I125223), .Q(I125537) );
not I_7245 (I125200,I125537);
DFFARX1 I_7246  ( .D(I125520), .CLK(I2350), .RSTB(I125223), .Q(I125185) );
DFFARX1 I_7247  ( .D(I380430), .CLK(I2350), .RSTB(I125223), .Q(I125582) );
not I_7248 (I125599,I125582);
nor I_7249 (I125616,I125257,I125599);
and I_7250 (I125633,I125520,I125616);
or I_7251 (I125650,I125240,I125633);
DFFARX1 I_7252  ( .D(I125650), .CLK(I2350), .RSTB(I125223), .Q(I125206) );
nor I_7253 (I125681,I125582,I125390);
nand I_7254 (I125215,I125356,I125681);
nor I_7255 (I125712,I125582,I125305);
nand I_7256 (I125209,I125455,I125712);
not I_7257 (I125212,I125582);
nand I_7258 (I125203,I125582,I125305);
DFFARX1 I_7259  ( .D(I125582), .CLK(I2350), .RSTB(I125223), .Q(I125194) );
not I_7260 (I125818,I2357);
or I_7261 (I125835,I166852,I166867);
or I_7262 (I125852,I166855,I166852);
DFFARX1 I_7263  ( .D(I125852), .CLK(I2350), .RSTB(I125818), .Q(I125792) );
nor I_7264 (I125883,I166858,I166873);
not I_7265 (I125900,I125883);
not I_7266 (I125917,I166858);
and I_7267 (I125934,I125917,I166861);
nor I_7268 (I125951,I125934,I166867);
nor I_7269 (I125968,I166864,I166882);
DFFARX1 I_7270  ( .D(I125968), .CLK(I2350), .RSTB(I125818), .Q(I125985) );
nand I_7271 (I126002,I125985,I125835);
and I_7272 (I126019,I125951,I126002);
DFFARX1 I_7273  ( .D(I126019), .CLK(I2350), .RSTB(I125818), .Q(I125786) );
nor I_7274 (I126050,I166864,I166855);
DFFARX1 I_7275  ( .D(I126050), .CLK(I2350), .RSTB(I125818), .Q(I126067) );
and I_7276 (I125783,I125883,I126067);
DFFARX1 I_7277  ( .D(I166879), .CLK(I2350), .RSTB(I125818), .Q(I126098) );
and I_7278 (I126115,I126098,I166870);
DFFARX1 I_7279  ( .D(I126115), .CLK(I2350), .RSTB(I125818), .Q(I126132) );
not I_7280 (I125795,I126132);
DFFARX1 I_7281  ( .D(I126115), .CLK(I2350), .RSTB(I125818), .Q(I125780) );
DFFARX1 I_7282  ( .D(I166876), .CLK(I2350), .RSTB(I125818), .Q(I126177) );
not I_7283 (I126194,I126177);
nor I_7284 (I126211,I125852,I126194);
and I_7285 (I126228,I126115,I126211);
or I_7286 (I126245,I125835,I126228);
DFFARX1 I_7287  ( .D(I126245), .CLK(I2350), .RSTB(I125818), .Q(I125801) );
nor I_7288 (I126276,I126177,I125985);
nand I_7289 (I125810,I125951,I126276);
nor I_7290 (I126307,I126177,I125900);
nand I_7291 (I125804,I126050,I126307);
not I_7292 (I125807,I126177);
nand I_7293 (I125798,I126177,I125900);
DFFARX1 I_7294  ( .D(I126177), .CLK(I2350), .RSTB(I125818), .Q(I125789) );
not I_7295 (I126413,I2357);
or I_7296 (I126430,I377893,I377890);
or I_7297 (I126447,I377920,I377893);
DFFARX1 I_7298  ( .D(I126447), .CLK(I2350), .RSTB(I126413), .Q(I126387) );
nor I_7299 (I126478,I377899,I377905);
not I_7300 (I126495,I126478);
not I_7301 (I126512,I377899);
and I_7302 (I126529,I126512,I377896);
nor I_7303 (I126546,I126529,I377890);
nor I_7304 (I126563,I377908,I377917);
DFFARX1 I_7305  ( .D(I126563), .CLK(I2350), .RSTB(I126413), .Q(I126580) );
nand I_7306 (I126597,I126580,I126430);
and I_7307 (I126614,I126546,I126597);
DFFARX1 I_7308  ( .D(I126614), .CLK(I2350), .RSTB(I126413), .Q(I126381) );
nor I_7309 (I126645,I377908,I377920);
DFFARX1 I_7310  ( .D(I126645), .CLK(I2350), .RSTB(I126413), .Q(I126662) );
and I_7311 (I126378,I126478,I126662);
DFFARX1 I_7312  ( .D(I377911), .CLK(I2350), .RSTB(I126413), .Q(I126693) );
and I_7313 (I126710,I126693,I377902);
DFFARX1 I_7314  ( .D(I126710), .CLK(I2350), .RSTB(I126413), .Q(I126727) );
not I_7315 (I126390,I126727);
DFFARX1 I_7316  ( .D(I126710), .CLK(I2350), .RSTB(I126413), .Q(I126375) );
DFFARX1 I_7317  ( .D(I377914), .CLK(I2350), .RSTB(I126413), .Q(I126772) );
not I_7318 (I126789,I126772);
nor I_7319 (I126806,I126447,I126789);
and I_7320 (I126823,I126710,I126806);
or I_7321 (I126840,I126430,I126823);
DFFARX1 I_7322  ( .D(I126840), .CLK(I2350), .RSTB(I126413), .Q(I126396) );
nor I_7323 (I126871,I126772,I126580);
nand I_7324 (I126405,I126546,I126871);
nor I_7325 (I126902,I126772,I126495);
nand I_7326 (I126399,I126645,I126902);
not I_7327 (I126402,I126772);
nand I_7328 (I126393,I126772,I126495);
DFFARX1 I_7329  ( .D(I126772), .CLK(I2350), .RSTB(I126413), .Q(I126384) );
not I_7330 (I127008,I2357);
or I_7331 (I127025,I368458,I368455);
or I_7332 (I127042,I368485,I368458);
DFFARX1 I_7333  ( .D(I127042), .CLK(I2350), .RSTB(I127008), .Q(I126982) );
nor I_7334 (I127073,I368464,I368470);
not I_7335 (I127090,I127073);
not I_7336 (I127107,I368464);
and I_7337 (I127124,I127107,I368461);
nor I_7338 (I127141,I127124,I368455);
nor I_7339 (I127158,I368473,I368482);
DFFARX1 I_7340  ( .D(I127158), .CLK(I2350), .RSTB(I127008), .Q(I127175) );
nand I_7341 (I127192,I127175,I127025);
and I_7342 (I127209,I127141,I127192);
DFFARX1 I_7343  ( .D(I127209), .CLK(I2350), .RSTB(I127008), .Q(I126976) );
nor I_7344 (I127240,I368473,I368485);
DFFARX1 I_7345  ( .D(I127240), .CLK(I2350), .RSTB(I127008), .Q(I127257) );
and I_7346 (I126973,I127073,I127257);
DFFARX1 I_7347  ( .D(I368476), .CLK(I2350), .RSTB(I127008), .Q(I127288) );
and I_7348 (I127305,I127288,I368467);
DFFARX1 I_7349  ( .D(I127305), .CLK(I2350), .RSTB(I127008), .Q(I127322) );
not I_7350 (I126985,I127322);
DFFARX1 I_7351  ( .D(I127305), .CLK(I2350), .RSTB(I127008), .Q(I126970) );
DFFARX1 I_7352  ( .D(I368479), .CLK(I2350), .RSTB(I127008), .Q(I127367) );
not I_7353 (I127384,I127367);
nor I_7354 (I127401,I127042,I127384);
and I_7355 (I127418,I127305,I127401);
or I_7356 (I127435,I127025,I127418);
DFFARX1 I_7357  ( .D(I127435), .CLK(I2350), .RSTB(I127008), .Q(I126991) );
nor I_7358 (I127466,I127367,I127175);
nand I_7359 (I127000,I127141,I127466);
nor I_7360 (I127497,I127367,I127090);
nand I_7361 (I126994,I127240,I127497);
not I_7362 (I126997,I127367);
nand I_7363 (I126988,I127367,I127090);
DFFARX1 I_7364  ( .D(I127367), .CLK(I2350), .RSTB(I127008), .Q(I126979) );
not I_7365 (I127603,I2357);
or I_7366 (I127620,I177460,I177475);
or I_7367 (I127637,I177463,I177460);
DFFARX1 I_7368  ( .D(I127637), .CLK(I2350), .RSTB(I127603), .Q(I127577) );
nor I_7369 (I127668,I177466,I177481);
not I_7370 (I127685,I127668);
not I_7371 (I127702,I177466);
and I_7372 (I127719,I127702,I177469);
nor I_7373 (I127736,I127719,I177475);
nor I_7374 (I127753,I177472,I177490);
DFFARX1 I_7375  ( .D(I127753), .CLK(I2350), .RSTB(I127603), .Q(I127770) );
nand I_7376 (I127787,I127770,I127620);
and I_7377 (I127804,I127736,I127787);
DFFARX1 I_7378  ( .D(I127804), .CLK(I2350), .RSTB(I127603), .Q(I127571) );
nor I_7379 (I127835,I177472,I177463);
DFFARX1 I_7380  ( .D(I127835), .CLK(I2350), .RSTB(I127603), .Q(I127852) );
and I_7381 (I127568,I127668,I127852);
DFFARX1 I_7382  ( .D(I177487), .CLK(I2350), .RSTB(I127603), .Q(I127883) );
and I_7383 (I127900,I127883,I177478);
DFFARX1 I_7384  ( .D(I127900), .CLK(I2350), .RSTB(I127603), .Q(I127917) );
not I_7385 (I127580,I127917);
DFFARX1 I_7386  ( .D(I127900), .CLK(I2350), .RSTB(I127603), .Q(I127565) );
DFFARX1 I_7387  ( .D(I177484), .CLK(I2350), .RSTB(I127603), .Q(I127962) );
not I_7388 (I127979,I127962);
nor I_7389 (I127996,I127637,I127979);
and I_7390 (I128013,I127900,I127996);
or I_7391 (I128030,I127620,I128013);
DFFARX1 I_7392  ( .D(I128030), .CLK(I2350), .RSTB(I127603), .Q(I127586) );
nor I_7393 (I128061,I127962,I127770);
nand I_7394 (I127595,I127736,I128061);
nor I_7395 (I128092,I127962,I127685);
nand I_7396 (I127589,I127835,I128092);
not I_7397 (I127592,I127962);
nand I_7398 (I127583,I127962,I127685);
DFFARX1 I_7399  ( .D(I127962), .CLK(I2350), .RSTB(I127603), .Q(I127574) );
not I_7400 (I128198,I2357);
or I_7401 (I128215,I301677,I301662);
or I_7402 (I128232,I301683,I301677);
DFFARX1 I_7403  ( .D(I128232), .CLK(I2350), .RSTB(I128198), .Q(I128172) );
nor I_7404 (I128263,I301689,I301671);
not I_7405 (I128280,I128263);
not I_7406 (I128297,I301689);
and I_7407 (I128314,I128297,I301668);
nor I_7408 (I128331,I128314,I301662);
nor I_7409 (I128348,I301665,I301674);
DFFARX1 I_7410  ( .D(I128348), .CLK(I2350), .RSTB(I128198), .Q(I128365) );
nand I_7411 (I128382,I128365,I128215);
and I_7412 (I128399,I128331,I128382);
DFFARX1 I_7413  ( .D(I128399), .CLK(I2350), .RSTB(I128198), .Q(I128166) );
nor I_7414 (I128430,I301665,I301683);
DFFARX1 I_7415  ( .D(I128430), .CLK(I2350), .RSTB(I128198), .Q(I128447) );
and I_7416 (I128163,I128263,I128447);
DFFARX1 I_7417  ( .D(I301692), .CLK(I2350), .RSTB(I128198), .Q(I128478) );
and I_7418 (I128495,I128478,I301680);
DFFARX1 I_7419  ( .D(I128495), .CLK(I2350), .RSTB(I128198), .Q(I128512) );
not I_7420 (I128175,I128512);
DFFARX1 I_7421  ( .D(I128495), .CLK(I2350), .RSTB(I128198), .Q(I128160) );
DFFARX1 I_7422  ( .D(I301686), .CLK(I2350), .RSTB(I128198), .Q(I128557) );
not I_7423 (I128574,I128557);
nor I_7424 (I128591,I128232,I128574);
and I_7425 (I128608,I128495,I128591);
or I_7426 (I128625,I128215,I128608);
DFFARX1 I_7427  ( .D(I128625), .CLK(I2350), .RSTB(I128198), .Q(I128181) );
nor I_7428 (I128656,I128557,I128365);
nand I_7429 (I128190,I128331,I128656);
nor I_7430 (I128687,I128557,I128280);
nand I_7431 (I128184,I128430,I128687);
not I_7432 (I128187,I128557);
nand I_7433 (I128178,I128557,I128280);
DFFARX1 I_7434  ( .D(I128557), .CLK(I2350), .RSTB(I128198), .Q(I128169) );
not I_7435 (I128793,I2357);
or I_7436 (I128810,I314169,I314163);
or I_7437 (I128827,I314157,I314169);
DFFARX1 I_7438  ( .D(I128827), .CLK(I2350), .RSTB(I128793), .Q(I128767) );
nor I_7439 (I128858,I314160,I314166);
not I_7440 (I128875,I128858);
not I_7441 (I128892,I314160);
and I_7442 (I128909,I128892,I314184);
nor I_7443 (I128926,I128909,I314163);
nor I_7444 (I128943,I314187,I314178);
DFFARX1 I_7445  ( .D(I128943), .CLK(I2350), .RSTB(I128793), .Q(I128960) );
nand I_7446 (I128977,I128960,I128810);
and I_7447 (I128994,I128926,I128977);
DFFARX1 I_7448  ( .D(I128994), .CLK(I2350), .RSTB(I128793), .Q(I128761) );
nor I_7449 (I129025,I314187,I314157);
DFFARX1 I_7450  ( .D(I129025), .CLK(I2350), .RSTB(I128793), .Q(I129042) );
and I_7451 (I128758,I128858,I129042);
DFFARX1 I_7452  ( .D(I314175), .CLK(I2350), .RSTB(I128793), .Q(I129073) );
and I_7453 (I129090,I129073,I314172);
DFFARX1 I_7454  ( .D(I129090), .CLK(I2350), .RSTB(I128793), .Q(I129107) );
not I_7455 (I128770,I129107);
DFFARX1 I_7456  ( .D(I129090), .CLK(I2350), .RSTB(I128793), .Q(I128755) );
DFFARX1 I_7457  ( .D(I314181), .CLK(I2350), .RSTB(I128793), .Q(I129152) );
not I_7458 (I129169,I129152);
nor I_7459 (I129186,I128827,I129169);
and I_7460 (I129203,I129090,I129186);
or I_7461 (I129220,I128810,I129203);
DFFARX1 I_7462  ( .D(I129220), .CLK(I2350), .RSTB(I128793), .Q(I128776) );
nor I_7463 (I129251,I129152,I128960);
nand I_7464 (I128785,I128926,I129251);
nor I_7465 (I129282,I129152,I128875);
nand I_7466 (I128779,I129025,I129282);
not I_7467 (I128782,I129152);
nand I_7468 (I128773,I129152,I128875);
DFFARX1 I_7469  ( .D(I129152), .CLK(I2350), .RSTB(I128793), .Q(I128764) );
not I_7470 (I129388,I2357);
or I_7471 (I129405,I269706,I269715);
or I_7472 (I129422,I269709,I269706);
DFFARX1 I_7473  ( .D(I129422), .CLK(I2350), .RSTB(I129388), .Q(I129362) );
nor I_7474 (I129453,I269694,I269685);
not I_7475 (I129470,I129453);
not I_7476 (I129487,I269694);
and I_7477 (I129504,I129487,I269712);
nor I_7478 (I129521,I129504,I269715);
nor I_7479 (I129538,I269688,I269697);
DFFARX1 I_7480  ( .D(I129538), .CLK(I2350), .RSTB(I129388), .Q(I129555) );
nand I_7481 (I129572,I129555,I129405);
and I_7482 (I129589,I129521,I129572);
DFFARX1 I_7483  ( .D(I129589), .CLK(I2350), .RSTB(I129388), .Q(I129356) );
nor I_7484 (I129620,I269688,I269709);
DFFARX1 I_7485  ( .D(I129620), .CLK(I2350), .RSTB(I129388), .Q(I129637) );
and I_7486 (I129353,I129453,I129637);
DFFARX1 I_7487  ( .D(I269691), .CLK(I2350), .RSTB(I129388), .Q(I129668) );
and I_7488 (I129685,I129668,I269703);
DFFARX1 I_7489  ( .D(I129685), .CLK(I2350), .RSTB(I129388), .Q(I129702) );
not I_7490 (I129365,I129702);
DFFARX1 I_7491  ( .D(I129685), .CLK(I2350), .RSTB(I129388), .Q(I129350) );
DFFARX1 I_7492  ( .D(I269700), .CLK(I2350), .RSTB(I129388), .Q(I129747) );
not I_7493 (I129764,I129747);
nor I_7494 (I129781,I129422,I129764);
and I_7495 (I129798,I129685,I129781);
or I_7496 (I129815,I129405,I129798);
DFFARX1 I_7497  ( .D(I129815), .CLK(I2350), .RSTB(I129388), .Q(I129371) );
nor I_7498 (I129846,I129747,I129555);
nand I_7499 (I129380,I129521,I129846);
nor I_7500 (I129877,I129747,I129470);
nand I_7501 (I129374,I129620,I129877);
not I_7502 (I129377,I129747);
nand I_7503 (I129368,I129747,I129470);
DFFARX1 I_7504  ( .D(I129747), .CLK(I2350), .RSTB(I129388), .Q(I129359) );
not I_7505 (I129983,I2357);
or I_7506 (I130000,I170845,I170833);
not I_7507 (I129966,I130000);
DFFARX1 I_7508  ( .D(I130000), .CLK(I2350), .RSTB(I129983), .Q(I129945) );
or I_7509 (I130045,I170830,I170845);
nor I_7510 (I130062,I170860,I170851);
nor I_7511 (I130079,I130062,I130000);
not I_7512 (I130096,I170860);
and I_7513 (I130113,I130096,I170839);
nor I_7514 (I130130,I130113,I170833);
DFFARX1 I_7515  ( .D(I130130), .CLK(I2350), .RSTB(I129983), .Q(I130147) );
nor I_7516 (I130164,I170842,I170836);
DFFARX1 I_7517  ( .D(I130164), .CLK(I2350), .RSTB(I129983), .Q(I130181) );
nor I_7518 (I129972,I130181,I130130);
not I_7519 (I130212,I130181);
nor I_7520 (I130229,I170842,I170830);
nand I_7521 (I130246,I130130,I130229);
and I_7522 (I130263,I130045,I130246);
DFFARX1 I_7523  ( .D(I130263), .CLK(I2350), .RSTB(I129983), .Q(I129975) );
DFFARX1 I_7524  ( .D(I170857), .CLK(I2350), .RSTB(I129983), .Q(I130294) );
and I_7525 (I130311,I130294,I170854);
nor I_7526 (I130328,I130311,I130212);
and I_7527 (I130345,I130229,I130328);
or I_7528 (I130362,I130062,I130345);
DFFARX1 I_7529  ( .D(I130362), .CLK(I2350), .RSTB(I129983), .Q(I129960) );
not I_7530 (I130393,I130311);
nor I_7531 (I130410,I130000,I130393);
nand I_7532 (I129963,I130045,I130410);
nand I_7533 (I129957,I130181,I130393);
DFFARX1 I_7534  ( .D(I130311), .CLK(I2350), .RSTB(I129983), .Q(I129951) );
DFFARX1 I_7535  ( .D(I170848), .CLK(I2350), .RSTB(I129983), .Q(I130469) );
nand I_7536 (I129969,I130469,I130079);
DFFARX1 I_7537  ( .D(I130469), .CLK(I2350), .RSTB(I129983), .Q(I130500) );
not I_7538 (I129954,I130500);
and I_7539 (I129948,I130469,I130147);
not I_7540 (I130578,I2357);
or I_7541 (I130595,I31754,I31751);
not I_7542 (I130561,I130595);
DFFARX1 I_7543  ( .D(I130595), .CLK(I2350), .RSTB(I130578), .Q(I130540) );
or I_7544 (I130640,I31745,I31754);
nor I_7545 (I130657,I31763,I31736);
nor I_7546 (I130674,I130657,I130595);
not I_7547 (I130691,I31763);
and I_7548 (I130708,I130691,I31757);
nor I_7549 (I130725,I130708,I31751);
DFFARX1 I_7550  ( .D(I130725), .CLK(I2350), .RSTB(I130578), .Q(I130742) );
nor I_7551 (I130759,I31739,I31766);
DFFARX1 I_7552  ( .D(I130759), .CLK(I2350), .RSTB(I130578), .Q(I130776) );
nor I_7553 (I130567,I130776,I130725);
not I_7554 (I130807,I130776);
nor I_7555 (I130824,I31739,I31745);
nand I_7556 (I130841,I130725,I130824);
and I_7557 (I130858,I130640,I130841);
DFFARX1 I_7558  ( .D(I130858), .CLK(I2350), .RSTB(I130578), .Q(I130570) );
DFFARX1 I_7559  ( .D(I31742), .CLK(I2350), .RSTB(I130578), .Q(I130889) );
and I_7560 (I130906,I130889,I31748);
nor I_7561 (I130923,I130906,I130807);
and I_7562 (I130940,I130824,I130923);
or I_7563 (I130957,I130657,I130940);
DFFARX1 I_7564  ( .D(I130957), .CLK(I2350), .RSTB(I130578), .Q(I130555) );
not I_7565 (I130988,I130906);
nor I_7566 (I131005,I130595,I130988);
nand I_7567 (I130558,I130640,I131005);
nand I_7568 (I130552,I130776,I130988);
DFFARX1 I_7569  ( .D(I130906), .CLK(I2350), .RSTB(I130578), .Q(I130546) );
DFFARX1 I_7570  ( .D(I31760), .CLK(I2350), .RSTB(I130578), .Q(I131064) );
nand I_7571 (I130564,I131064,I130674);
DFFARX1 I_7572  ( .D(I131064), .CLK(I2350), .RSTB(I130578), .Q(I131095) );
not I_7573 (I130549,I131095);
and I_7574 (I130543,I131064,I130742);
not I_7575 (I131173,I2357);
or I_7576 (I131190,I125197,I125194);
not I_7577 (I131156,I131190);
DFFARX1 I_7578  ( .D(I131190), .CLK(I2350), .RSTB(I131173), .Q(I131135) );
or I_7579 (I131235,I125185,I125197);
nor I_7580 (I131252,I125212,I125191);
nor I_7581 (I131269,I131252,I131190);
not I_7582 (I131286,I125212);
and I_7583 (I131303,I131286,I125200);
nor I_7584 (I131320,I131303,I125194);
DFFARX1 I_7585  ( .D(I131320), .CLK(I2350), .RSTB(I131173), .Q(I131337) );
nor I_7586 (I131354,I125188,I125206);
DFFARX1 I_7587  ( .D(I131354), .CLK(I2350), .RSTB(I131173), .Q(I131371) );
nor I_7588 (I131162,I131371,I131320);
not I_7589 (I131402,I131371);
nor I_7590 (I131419,I125188,I125185);
nand I_7591 (I131436,I131320,I131419);
and I_7592 (I131453,I131235,I131436);
DFFARX1 I_7593  ( .D(I131453), .CLK(I2350), .RSTB(I131173), .Q(I131165) );
DFFARX1 I_7594  ( .D(I125203), .CLK(I2350), .RSTB(I131173), .Q(I131484) );
and I_7595 (I131501,I131484,I125215);
nor I_7596 (I131518,I131501,I131402);
and I_7597 (I131535,I131419,I131518);
or I_7598 (I131552,I131252,I131535);
DFFARX1 I_7599  ( .D(I131552), .CLK(I2350), .RSTB(I131173), .Q(I131150) );
not I_7600 (I131583,I131501);
nor I_7601 (I131600,I131190,I131583);
nand I_7602 (I131153,I131235,I131600);
nand I_7603 (I131147,I131371,I131583);
DFFARX1 I_7604  ( .D(I131501), .CLK(I2350), .RSTB(I131173), .Q(I131141) );
DFFARX1 I_7605  ( .D(I125209), .CLK(I2350), .RSTB(I131173), .Q(I131659) );
nand I_7606 (I131159,I131659,I131269);
DFFARX1 I_7607  ( .D(I131659), .CLK(I2350), .RSTB(I131173), .Q(I131690) );
not I_7608 (I131144,I131690);
and I_7609 (I131138,I131659,I131337);
not I_7610 (I131768,I2357);
or I_7611 (I131785,I183442,I183430);
not I_7612 (I131751,I131785);
DFFARX1 I_7613  ( .D(I131785), .CLK(I2350), .RSTB(I131768), .Q(I131730) );
or I_7614 (I131830,I183427,I183442);
nor I_7615 (I131847,I183457,I183448);
nor I_7616 (I131864,I131847,I131785);
not I_7617 (I131881,I183457);
and I_7618 (I131898,I131881,I183436);
nor I_7619 (I131915,I131898,I183430);
DFFARX1 I_7620  ( .D(I131915), .CLK(I2350), .RSTB(I131768), .Q(I131932) );
nor I_7621 (I131949,I183439,I183433);
DFFARX1 I_7622  ( .D(I131949), .CLK(I2350), .RSTB(I131768), .Q(I131966) );
nor I_7623 (I131757,I131966,I131915);
not I_7624 (I131997,I131966);
nor I_7625 (I132014,I183439,I183427);
nand I_7626 (I132031,I131915,I132014);
and I_7627 (I132048,I131830,I132031);
DFFARX1 I_7628  ( .D(I132048), .CLK(I2350), .RSTB(I131768), .Q(I131760) );
DFFARX1 I_7629  ( .D(I183454), .CLK(I2350), .RSTB(I131768), .Q(I132079) );
and I_7630 (I132096,I132079,I183451);
nor I_7631 (I132113,I132096,I131997);
and I_7632 (I132130,I132014,I132113);
or I_7633 (I132147,I131847,I132130);
DFFARX1 I_7634  ( .D(I132147), .CLK(I2350), .RSTB(I131768), .Q(I131745) );
not I_7635 (I132178,I132096);
nor I_7636 (I132195,I131785,I132178);
nand I_7637 (I131748,I131830,I132195);
nand I_7638 (I131742,I131966,I132178);
DFFARX1 I_7639  ( .D(I132096), .CLK(I2350), .RSTB(I131768), .Q(I131736) );
DFFARX1 I_7640  ( .D(I183445), .CLK(I2350), .RSTB(I131768), .Q(I132254) );
nand I_7641 (I131754,I132254,I131864);
DFFARX1 I_7642  ( .D(I132254), .CLK(I2350), .RSTB(I131768), .Q(I132285) );
not I_7643 (I131739,I132285);
and I_7644 (I131733,I132254,I131932);
not I_7645 (I132363,I2357);
or I_7646 (I132380,I50488,I50485);
not I_7647 (I132346,I132380);
DFFARX1 I_7648  ( .D(I132380), .CLK(I2350), .RSTB(I132363), .Q(I132325) );
or I_7649 (I132425,I50479,I50488);
nor I_7650 (I132442,I50497,I50470);
nor I_7651 (I132459,I132442,I132380);
not I_7652 (I132476,I50497);
and I_7653 (I132493,I132476,I50491);
nor I_7654 (I132510,I132493,I50485);
DFFARX1 I_7655  ( .D(I132510), .CLK(I2350), .RSTB(I132363), .Q(I132527) );
nor I_7656 (I132544,I50473,I50500);
DFFARX1 I_7657  ( .D(I132544), .CLK(I2350), .RSTB(I132363), .Q(I132561) );
nor I_7658 (I132352,I132561,I132510);
not I_7659 (I132592,I132561);
nor I_7660 (I132609,I50473,I50479);
nand I_7661 (I132626,I132510,I132609);
and I_7662 (I132643,I132425,I132626);
DFFARX1 I_7663  ( .D(I132643), .CLK(I2350), .RSTB(I132363), .Q(I132355) );
DFFARX1 I_7664  ( .D(I50476), .CLK(I2350), .RSTB(I132363), .Q(I132674) );
and I_7665 (I132691,I132674,I50482);
nor I_7666 (I132708,I132691,I132592);
and I_7667 (I132725,I132609,I132708);
or I_7668 (I132742,I132442,I132725);
DFFARX1 I_7669  ( .D(I132742), .CLK(I2350), .RSTB(I132363), .Q(I132340) );
not I_7670 (I132773,I132691);
nor I_7671 (I132790,I132380,I132773);
nand I_7672 (I132343,I132425,I132790);
nand I_7673 (I132337,I132561,I132773);
DFFARX1 I_7674  ( .D(I132691), .CLK(I2350), .RSTB(I132363), .Q(I132331) );
DFFARX1 I_7675  ( .D(I50494), .CLK(I2350), .RSTB(I132363), .Q(I132849) );
nand I_7676 (I132349,I132849,I132459);
DFFARX1 I_7677  ( .D(I132849), .CLK(I2350), .RSTB(I132363), .Q(I132880) );
not I_7678 (I132334,I132880);
and I_7679 (I132328,I132849,I132527);
not I_7680 (I132958,I2357);
or I_7681 (I132975,I245817,I245847);
not I_7682 (I132941,I132975);
DFFARX1 I_7683  ( .D(I132975), .CLK(I2350), .RSTB(I132958), .Q(I132920) );
or I_7684 (I133020,I245826,I245817);
nor I_7685 (I133037,I245832,I245829);
nor I_7686 (I133054,I133037,I132975);
not I_7687 (I133071,I245832);
and I_7688 (I133088,I133071,I245838);
nor I_7689 (I133105,I133088,I245847);
DFFARX1 I_7690  ( .D(I133105), .CLK(I2350), .RSTB(I132958), .Q(I133122) );
nor I_7691 (I133139,I245823,I245841);
DFFARX1 I_7692  ( .D(I133139), .CLK(I2350), .RSTB(I132958), .Q(I133156) );
nor I_7693 (I132947,I133156,I133105);
not I_7694 (I133187,I133156);
nor I_7695 (I133204,I245823,I245826);
nand I_7696 (I133221,I133105,I133204);
and I_7697 (I133238,I133020,I133221);
DFFARX1 I_7698  ( .D(I133238), .CLK(I2350), .RSTB(I132958), .Q(I132950) );
DFFARX1 I_7699  ( .D(I245844), .CLK(I2350), .RSTB(I132958), .Q(I133269) );
and I_7700 (I133286,I133269,I245835);
nor I_7701 (I133303,I133286,I133187);
and I_7702 (I133320,I133204,I133303);
or I_7703 (I133337,I133037,I133320);
DFFARX1 I_7704  ( .D(I133337), .CLK(I2350), .RSTB(I132958), .Q(I132935) );
not I_7705 (I133368,I133286);
nor I_7706 (I133385,I132975,I133368);
nand I_7707 (I132938,I133020,I133385);
nand I_7708 (I132932,I133156,I133368);
DFFARX1 I_7709  ( .D(I133286), .CLK(I2350), .RSTB(I132958), .Q(I132926) );
DFFARX1 I_7710  ( .D(I245820), .CLK(I2350), .RSTB(I132958), .Q(I133444) );
nand I_7711 (I132944,I133444,I133054);
DFFARX1 I_7712  ( .D(I133444), .CLK(I2350), .RSTB(I132958), .Q(I133475) );
not I_7713 (I132929,I133475);
and I_7714 (I132923,I133444,I133122);
not I_7715 (I133553,I2357);
or I_7716 (I133570,I84717,I84714);
not I_7717 (I133536,I133570);
DFFARX1 I_7718  ( .D(I133570), .CLK(I2350), .RSTB(I133553), .Q(I133515) );
or I_7719 (I133615,I84732,I84717);
nor I_7720 (I133632,I84723,I84708);
nor I_7721 (I133649,I133632,I133570);
not I_7722 (I133666,I84723);
and I_7723 (I133683,I133666,I84726);
nor I_7724 (I133700,I133683,I84714);
DFFARX1 I_7725  ( .D(I133700), .CLK(I2350), .RSTB(I133553), .Q(I133717) );
nor I_7726 (I133734,I84711,I84720);
DFFARX1 I_7727  ( .D(I133734), .CLK(I2350), .RSTB(I133553), .Q(I133751) );
nor I_7728 (I133542,I133751,I133700);
not I_7729 (I133782,I133751);
nor I_7730 (I133799,I84711,I84732);
nand I_7731 (I133816,I133700,I133799);
and I_7732 (I133833,I133615,I133816);
DFFARX1 I_7733  ( .D(I133833), .CLK(I2350), .RSTB(I133553), .Q(I133545) );
DFFARX1 I_7734  ( .D(I84729), .CLK(I2350), .RSTB(I133553), .Q(I133864) );
and I_7735 (I133881,I133864,I84738);
nor I_7736 (I133898,I133881,I133782);
and I_7737 (I133915,I133799,I133898);
or I_7738 (I133932,I133632,I133915);
DFFARX1 I_7739  ( .D(I133932), .CLK(I2350), .RSTB(I133553), .Q(I133530) );
not I_7740 (I133963,I133881);
nor I_7741 (I133980,I133570,I133963);
nand I_7742 (I133533,I133615,I133980);
nand I_7743 (I133527,I133751,I133963);
DFFARX1 I_7744  ( .D(I133881), .CLK(I2350), .RSTB(I133553), .Q(I133521) );
DFFARX1 I_7745  ( .D(I84735), .CLK(I2350), .RSTB(I133553), .Q(I134039) );
nand I_7746 (I133539,I134039,I133649);
DFFARX1 I_7747  ( .D(I134039), .CLK(I2350), .RSTB(I133553), .Q(I134070) );
not I_7748 (I133524,I134070);
and I_7749 (I133518,I134039,I133717);
not I_7750 (I134148,I2357);
or I_7751 (I134165,I152944,I152932);
not I_7752 (I134131,I134165);
DFFARX1 I_7753  ( .D(I134165), .CLK(I2350), .RSTB(I134148), .Q(I134110) );
or I_7754 (I134210,I152929,I152944);
nor I_7755 (I134227,I152959,I152950);
nor I_7756 (I134244,I134227,I134165);
not I_7757 (I134261,I152959);
and I_7758 (I134278,I134261,I152938);
nor I_7759 (I134295,I134278,I152932);
DFFARX1 I_7760  ( .D(I134295), .CLK(I2350), .RSTB(I134148), .Q(I134312) );
nor I_7761 (I134329,I152941,I152935);
DFFARX1 I_7762  ( .D(I134329), .CLK(I2350), .RSTB(I134148), .Q(I134346) );
nor I_7763 (I134137,I134346,I134295);
not I_7764 (I134377,I134346);
nor I_7765 (I134394,I152941,I152929);
nand I_7766 (I134411,I134295,I134394);
and I_7767 (I134428,I134210,I134411);
DFFARX1 I_7768  ( .D(I134428), .CLK(I2350), .RSTB(I134148), .Q(I134140) );
DFFARX1 I_7769  ( .D(I152956), .CLK(I2350), .RSTB(I134148), .Q(I134459) );
and I_7770 (I134476,I134459,I152953);
nor I_7771 (I134493,I134476,I134377);
and I_7772 (I134510,I134394,I134493);
or I_7773 (I134527,I134227,I134510);
DFFARX1 I_7774  ( .D(I134527), .CLK(I2350), .RSTB(I134148), .Q(I134125) );
not I_7775 (I134558,I134476);
nor I_7776 (I134575,I134165,I134558);
nand I_7777 (I134128,I134210,I134575);
nand I_7778 (I134122,I134346,I134558);
DFFARX1 I_7779  ( .D(I134476), .CLK(I2350), .RSTB(I134148), .Q(I134116) );
DFFARX1 I_7780  ( .D(I152947), .CLK(I2350), .RSTB(I134148), .Q(I134634) );
nand I_7781 (I134134,I134634,I134244);
DFFARX1 I_7782  ( .D(I134634), .CLK(I2350), .RSTB(I134148), .Q(I134665) );
not I_7783 (I134119,I134665);
and I_7784 (I134113,I134634,I134312);
not I_7785 (I134743,I2357);
or I_7786 (I134760,I348333,I348342);
not I_7787 (I134726,I134760);
DFFARX1 I_7788  ( .D(I134760), .CLK(I2350), .RSTB(I134743), .Q(I134705) );
or I_7789 (I134805,I348351,I348333);
nor I_7790 (I134822,I348345,I348339);
nor I_7791 (I134839,I134822,I134760);
not I_7792 (I134856,I348345);
and I_7793 (I134873,I134856,I348348);
nor I_7794 (I134890,I134873,I348342);
DFFARX1 I_7795  ( .D(I134890), .CLK(I2350), .RSTB(I134743), .Q(I134907) );
nor I_7796 (I134924,I348336,I348354);
DFFARX1 I_7797  ( .D(I134924), .CLK(I2350), .RSTB(I134743), .Q(I134941) );
nor I_7798 (I134732,I134941,I134890);
not I_7799 (I134972,I134941);
nor I_7800 (I134989,I348336,I348351);
nand I_7801 (I135006,I134890,I134989);
and I_7802 (I135023,I134805,I135006);
DFFARX1 I_7803  ( .D(I135023), .CLK(I2350), .RSTB(I134743), .Q(I134735) );
DFFARX1 I_7804  ( .D(I348357), .CLK(I2350), .RSTB(I134743), .Q(I135054) );
and I_7805 (I135071,I135054,I348330);
nor I_7806 (I135088,I135071,I134972);
and I_7807 (I135105,I134989,I135088);
or I_7808 (I135122,I134822,I135105);
DFFARX1 I_7809  ( .D(I135122), .CLK(I2350), .RSTB(I134743), .Q(I134720) );
not I_7810 (I135153,I135071);
nor I_7811 (I135170,I134760,I135153);
nand I_7812 (I134723,I134805,I135170);
nand I_7813 (I134717,I134941,I135153);
DFFARX1 I_7814  ( .D(I135071), .CLK(I2350), .RSTB(I134743), .Q(I134711) );
DFFARX1 I_7815  ( .D(I348327), .CLK(I2350), .RSTB(I134743), .Q(I135229) );
nand I_7816 (I134729,I135229,I134839);
DFFARX1 I_7817  ( .D(I135229), .CLK(I2350), .RSTB(I134743), .Q(I135260) );
not I_7818 (I134714,I135260);
and I_7819 (I134708,I135229,I134907);
not I_7820 (I135338,I2357);
or I_7821 (I135355,I90684,I90681);
not I_7822 (I135321,I135355);
DFFARX1 I_7823  ( .D(I135355), .CLK(I2350), .RSTB(I135338), .Q(I135300) );
or I_7824 (I135400,I90699,I90684);
nor I_7825 (I135417,I90690,I90675);
nor I_7826 (I135434,I135417,I135355);
not I_7827 (I135451,I90690);
and I_7828 (I135468,I135451,I90693);
nor I_7829 (I135485,I135468,I90681);
DFFARX1 I_7830  ( .D(I135485), .CLK(I2350), .RSTB(I135338), .Q(I135502) );
nor I_7831 (I135519,I90678,I90687);
DFFARX1 I_7832  ( .D(I135519), .CLK(I2350), .RSTB(I135338), .Q(I135536) );
nor I_7833 (I135327,I135536,I135485);
not I_7834 (I135567,I135536);
nor I_7835 (I135584,I90678,I90699);
nand I_7836 (I135601,I135485,I135584);
and I_7837 (I135618,I135400,I135601);
DFFARX1 I_7838  ( .D(I135618), .CLK(I2350), .RSTB(I135338), .Q(I135330) );
DFFARX1 I_7839  ( .D(I90696), .CLK(I2350), .RSTB(I135338), .Q(I135649) );
and I_7840 (I135666,I135649,I90705);
nor I_7841 (I135683,I135666,I135567);
and I_7842 (I135700,I135584,I135683);
or I_7843 (I135717,I135417,I135700);
DFFARX1 I_7844  ( .D(I135717), .CLK(I2350), .RSTB(I135338), .Q(I135315) );
not I_7845 (I135748,I135666);
nor I_7846 (I135765,I135355,I135748);
nand I_7847 (I135318,I135400,I135765);
nand I_7848 (I135312,I135536,I135748);
DFFARX1 I_7849  ( .D(I135666), .CLK(I2350), .RSTB(I135338), .Q(I135306) );
DFFARX1 I_7850  ( .D(I90702), .CLK(I2350), .RSTB(I135338), .Q(I135824) );
nand I_7851 (I135324,I135824,I135434);
DFFARX1 I_7852  ( .D(I135824), .CLK(I2350), .RSTB(I135338), .Q(I135855) );
not I_7853 (I135309,I135855);
and I_7854 (I135303,I135824,I135502);
not I_7855 (I135933,I2357);
or I_7856 (I135950,I9116,I9092);
not I_7857 (I135916,I135950);
DFFARX1 I_7858  ( .D(I135950), .CLK(I2350), .RSTB(I135933), .Q(I135895) );
or I_7859 (I135995,I9119,I9116);
nor I_7860 (I136012,I9101,I9107);
nor I_7861 (I136029,I136012,I135950);
not I_7862 (I136046,I9101);
and I_7863 (I136063,I136046,I9095);
nor I_7864 (I136080,I136063,I9092);
DFFARX1 I_7865  ( .D(I136080), .CLK(I2350), .RSTB(I135933), .Q(I136097) );
nor I_7866 (I136114,I9122,I9113);
DFFARX1 I_7867  ( .D(I136114), .CLK(I2350), .RSTB(I135933), .Q(I136131) );
nor I_7868 (I135922,I136131,I136080);
not I_7869 (I136162,I136131);
nor I_7870 (I136179,I9122,I9119);
nand I_7871 (I136196,I136080,I136179);
and I_7872 (I136213,I135995,I136196);
DFFARX1 I_7873  ( .D(I136213), .CLK(I2350), .RSTB(I135933), .Q(I135925) );
DFFARX1 I_7874  ( .D(I9098), .CLK(I2350), .RSTB(I135933), .Q(I136244) );
and I_7875 (I136261,I136244,I9110);
nor I_7876 (I136278,I136261,I136162);
and I_7877 (I136295,I136179,I136278);
or I_7878 (I136312,I136012,I136295);
DFFARX1 I_7879  ( .D(I136312), .CLK(I2350), .RSTB(I135933), .Q(I135910) );
not I_7880 (I136343,I136261);
nor I_7881 (I136360,I135950,I136343);
nand I_7882 (I135913,I135995,I136360);
nand I_7883 (I135907,I136131,I136343);
DFFARX1 I_7884  ( .D(I136261), .CLK(I2350), .RSTB(I135933), .Q(I135901) );
DFFARX1 I_7885  ( .D(I9104), .CLK(I2350), .RSTB(I135933), .Q(I136419) );
nand I_7886 (I135919,I136419,I136029);
DFFARX1 I_7887  ( .D(I136419), .CLK(I2350), .RSTB(I135933), .Q(I136450) );
not I_7888 (I135904,I136450);
and I_7889 (I135898,I136419,I136097);
not I_7890 (I136528,I2357);
or I_7891 (I136545,I49196,I49193);
not I_7892 (I136511,I136545);
DFFARX1 I_7893  ( .D(I136545), .CLK(I2350), .RSTB(I136528), .Q(I136490) );
or I_7894 (I136590,I49187,I49196);
nor I_7895 (I136607,I49205,I49178);
nor I_7896 (I136624,I136607,I136545);
not I_7897 (I136641,I49205);
and I_7898 (I136658,I136641,I49199);
nor I_7899 (I136675,I136658,I49193);
DFFARX1 I_7900  ( .D(I136675), .CLK(I2350), .RSTB(I136528), .Q(I136692) );
nor I_7901 (I136709,I49181,I49208);
DFFARX1 I_7902  ( .D(I136709), .CLK(I2350), .RSTB(I136528), .Q(I136726) );
nor I_7903 (I136517,I136726,I136675);
not I_7904 (I136757,I136726);
nor I_7905 (I136774,I49181,I49187);
nand I_7906 (I136791,I136675,I136774);
and I_7907 (I136808,I136590,I136791);
DFFARX1 I_7908  ( .D(I136808), .CLK(I2350), .RSTB(I136528), .Q(I136520) );
DFFARX1 I_7909  ( .D(I49184), .CLK(I2350), .RSTB(I136528), .Q(I136839) );
and I_7910 (I136856,I136839,I49190);
nor I_7911 (I136873,I136856,I136757);
and I_7912 (I136890,I136774,I136873);
or I_7913 (I136907,I136607,I136890);
DFFARX1 I_7914  ( .D(I136907), .CLK(I2350), .RSTB(I136528), .Q(I136505) );
not I_7915 (I136938,I136856);
nor I_7916 (I136955,I136545,I136938);
nand I_7917 (I136508,I136590,I136955);
nand I_7918 (I136502,I136726,I136938);
DFFARX1 I_7919  ( .D(I136856), .CLK(I2350), .RSTB(I136528), .Q(I136496) );
DFFARX1 I_7920  ( .D(I49202), .CLK(I2350), .RSTB(I136528), .Q(I137014) );
nand I_7921 (I136514,I137014,I136624);
DFFARX1 I_7922  ( .D(I137014), .CLK(I2350), .RSTB(I136528), .Q(I137045) );
not I_7923 (I136499,I137045);
and I_7924 (I136493,I137014,I136692);
not I_7925 (I137123,I2357);
or I_7926 (I137140,I88695,I88692);
not I_7927 (I137106,I137140);
DFFARX1 I_7928  ( .D(I137140), .CLK(I2350), .RSTB(I137123), .Q(I137085) );
or I_7929 (I137185,I88710,I88695);
nor I_7930 (I137202,I88701,I88686);
nor I_7931 (I137219,I137202,I137140);
not I_7932 (I137236,I88701);
and I_7933 (I137253,I137236,I88704);
nor I_7934 (I137270,I137253,I88692);
DFFARX1 I_7935  ( .D(I137270), .CLK(I2350), .RSTB(I137123), .Q(I137287) );
nor I_7936 (I137304,I88689,I88698);
DFFARX1 I_7937  ( .D(I137304), .CLK(I2350), .RSTB(I137123), .Q(I137321) );
nor I_7938 (I137112,I137321,I137270);
not I_7939 (I137352,I137321);
nor I_7940 (I137369,I88689,I88710);
nand I_7941 (I137386,I137270,I137369);
and I_7942 (I137403,I137185,I137386);
DFFARX1 I_7943  ( .D(I137403), .CLK(I2350), .RSTB(I137123), .Q(I137115) );
DFFARX1 I_7944  ( .D(I88707), .CLK(I2350), .RSTB(I137123), .Q(I137434) );
and I_7945 (I137451,I137434,I88716);
nor I_7946 (I137468,I137451,I137352);
and I_7947 (I137485,I137369,I137468);
or I_7948 (I137502,I137202,I137485);
DFFARX1 I_7949  ( .D(I137502), .CLK(I2350), .RSTB(I137123), .Q(I137100) );
not I_7950 (I137533,I137451);
nor I_7951 (I137550,I137140,I137533);
nand I_7952 (I137103,I137185,I137550);
nand I_7953 (I137097,I137321,I137533);
DFFARX1 I_7954  ( .D(I137451), .CLK(I2350), .RSTB(I137123), .Q(I137091) );
DFFARX1 I_7955  ( .D(I88713), .CLK(I2350), .RSTB(I137123), .Q(I137609) );
nand I_7956 (I137109,I137609,I137219);
DFFARX1 I_7957  ( .D(I137609), .CLK(I2350), .RSTB(I137123), .Q(I137640) );
not I_7958 (I137094,I137640);
and I_7959 (I137088,I137609,I137287);
not I_7960 (I137718,I2357);
not I_7961 (I137735,I317150);
nor I_7962 (I137752,I317147,I317138);
nand I_7963 (I137769,I137752,I317141);
nor I_7964 (I137786,I137735,I317147);
nand I_7965 (I137803,I137786,I317135);
not I_7966 (I137820,I137803);
not I_7967 (I137837,I317147);
nor I_7968 (I137707,I137803,I137837);
not I_7969 (I137868,I137837);
nand I_7970 (I137692,I137803,I137868);
not I_7971 (I137899,I317156);
nor I_7972 (I137916,I137899,I317159);
and I_7973 (I137933,I137916,I317144);
or I_7974 (I137950,I137933,I317132);
DFFARX1 I_7975  ( .D(I137950), .CLK(I2350), .RSTB(I137718), .Q(I137967) );
nor I_7976 (I137984,I137967,I137820);
DFFARX1 I_7977  ( .D(I137967), .CLK(I2350), .RSTB(I137718), .Q(I138001) );
not I_7978 (I137689,I138001);
nand I_7979 (I138032,I137735,I317156);
and I_7980 (I138049,I138032,I137984);
DFFARX1 I_7981  ( .D(I138032), .CLK(I2350), .RSTB(I137718), .Q(I137686) );
DFFARX1 I_7982  ( .D(I317153), .CLK(I2350), .RSTB(I137718), .Q(I138080) );
nor I_7983 (I138097,I138080,I137803);
nand I_7984 (I137704,I137967,I138097);
nor I_7985 (I138128,I138080,I137868);
not I_7986 (I137701,I138080);
nand I_7987 (I138159,I138080,I137769);
and I_7988 (I138176,I137837,I138159);
DFFARX1 I_7989  ( .D(I138176), .CLK(I2350), .RSTB(I137718), .Q(I137680) );
DFFARX1 I_7990  ( .D(I138080), .CLK(I2350), .RSTB(I137718), .Q(I137683) );
DFFARX1 I_7991  ( .D(I317162), .CLK(I2350), .RSTB(I137718), .Q(I138221) );
not I_7992 (I138238,I138221);
nand I_7993 (I138255,I138238,I137803);
and I_7994 (I138272,I138032,I138255);
DFFARX1 I_7995  ( .D(I138272), .CLK(I2350), .RSTB(I137718), .Q(I137710) );
or I_7996 (I138303,I138238,I138049);
DFFARX1 I_7997  ( .D(I138303), .CLK(I2350), .RSTB(I137718), .Q(I137695) );
nand I_7998 (I137698,I138238,I138128);
not I_7999 (I138381,I2357);
not I_8000 (I138398,I85374);
nor I_8001 (I138415,I85380,I85386);
nand I_8002 (I138432,I138415,I85389);
nor I_8003 (I138449,I138398,I85380);
nand I_8004 (I138466,I138449,I85371);
not I_8005 (I138483,I138466);
not I_8006 (I138500,I85380);
nor I_8007 (I138370,I138466,I138500);
not I_8008 (I138531,I138500);
nand I_8009 (I138355,I138466,I138531);
not I_8010 (I138562,I85383);
nor I_8011 (I138579,I138562,I85377);
and I_8012 (I138596,I138579,I85392);
or I_8013 (I138613,I138596,I85398);
DFFARX1 I_8014  ( .D(I138613), .CLK(I2350), .RSTB(I138381), .Q(I138630) );
nor I_8015 (I138647,I138630,I138483);
DFFARX1 I_8016  ( .D(I138630), .CLK(I2350), .RSTB(I138381), .Q(I138664) );
not I_8017 (I138352,I138664);
nand I_8018 (I138695,I138398,I85383);
and I_8019 (I138712,I138695,I138647);
DFFARX1 I_8020  ( .D(I138695), .CLK(I2350), .RSTB(I138381), .Q(I138349) );
DFFARX1 I_8021  ( .D(I85395), .CLK(I2350), .RSTB(I138381), .Q(I138743) );
nor I_8022 (I138760,I138743,I138466);
nand I_8023 (I138367,I138630,I138760);
nor I_8024 (I138791,I138743,I138531);
not I_8025 (I138364,I138743);
nand I_8026 (I138822,I138743,I138432);
and I_8027 (I138839,I138500,I138822);
DFFARX1 I_8028  ( .D(I138839), .CLK(I2350), .RSTB(I138381), .Q(I138343) );
DFFARX1 I_8029  ( .D(I138743), .CLK(I2350), .RSTB(I138381), .Q(I138346) );
DFFARX1 I_8030  ( .D(I85401), .CLK(I2350), .RSTB(I138381), .Q(I138884) );
not I_8031 (I138901,I138884);
nand I_8032 (I138918,I138901,I138466);
and I_8033 (I138935,I138695,I138918);
DFFARX1 I_8034  ( .D(I138935), .CLK(I2350), .RSTB(I138381), .Q(I138373) );
or I_8035 (I138966,I138901,I138712);
DFFARX1 I_8036  ( .D(I138966), .CLK(I2350), .RSTB(I138381), .Q(I138358) );
nand I_8037 (I138361,I138901,I138791);
not I_8038 (I139044,I2357);
not I_8039 (I139061,I332608);
nor I_8040 (I139078,I332626,I332617);
nand I_8041 (I139095,I139078,I332623);
nor I_8042 (I139112,I139061,I332626);
nand I_8043 (I139129,I139112,I332629);
not I_8044 (I139146,I139129);
not I_8045 (I139163,I332626);
nor I_8046 (I139033,I139129,I139163);
not I_8047 (I139194,I139163);
nand I_8048 (I139018,I139129,I139194);
not I_8049 (I139225,I332605);
nor I_8050 (I139242,I139225,I332620);
and I_8051 (I139259,I139242,I332602);
or I_8052 (I139276,I139259,I332611);
DFFARX1 I_8053  ( .D(I139276), .CLK(I2350), .RSTB(I139044), .Q(I139293) );
nor I_8054 (I139310,I139293,I139146);
DFFARX1 I_8055  ( .D(I139293), .CLK(I2350), .RSTB(I139044), .Q(I139327) );
not I_8056 (I139015,I139327);
nand I_8057 (I139358,I139061,I332605);
and I_8058 (I139375,I139358,I139310);
DFFARX1 I_8059  ( .D(I139358), .CLK(I2350), .RSTB(I139044), .Q(I139012) );
DFFARX1 I_8060  ( .D(I332614), .CLK(I2350), .RSTB(I139044), .Q(I139406) );
nor I_8061 (I139423,I139406,I139129);
nand I_8062 (I139030,I139293,I139423);
nor I_8063 (I139454,I139406,I139194);
not I_8064 (I139027,I139406);
nand I_8065 (I139485,I139406,I139095);
and I_8066 (I139502,I139163,I139485);
DFFARX1 I_8067  ( .D(I139502), .CLK(I2350), .RSTB(I139044), .Q(I139006) );
DFFARX1 I_8068  ( .D(I139406), .CLK(I2350), .RSTB(I139044), .Q(I139009) );
DFFARX1 I_8069  ( .D(I332632), .CLK(I2350), .RSTB(I139044), .Q(I139547) );
not I_8070 (I139564,I139547);
nand I_8071 (I139581,I139564,I139129);
and I_8072 (I139598,I139358,I139581);
DFFARX1 I_8073  ( .D(I139598), .CLK(I2350), .RSTB(I139044), .Q(I139036) );
or I_8074 (I139629,I139564,I139375);
DFFARX1 I_8075  ( .D(I139629), .CLK(I2350), .RSTB(I139044), .Q(I139021) );
nand I_8076 (I139024,I139564,I139454);
not I_8077 (I139707,I2357);
not I_8078 (I139724,I208871);
nor I_8079 (I139741,I208868,I208886);
nand I_8080 (I139758,I139741,I208889);
nor I_8081 (I139775,I139724,I208868);
nand I_8082 (I139792,I139775,I208874);
not I_8083 (I139809,I139792);
not I_8084 (I139826,I208868);
nor I_8085 (I139696,I139792,I139826);
not I_8086 (I139857,I139826);
nand I_8087 (I139681,I139792,I139857);
not I_8088 (I139888,I208883);
nor I_8089 (I139905,I139888,I208865);
and I_8090 (I139922,I139905,I208859);
or I_8091 (I139939,I139922,I208877);
DFFARX1 I_8092  ( .D(I139939), .CLK(I2350), .RSTB(I139707), .Q(I139956) );
nor I_8093 (I139973,I139956,I139809);
DFFARX1 I_8094  ( .D(I139956), .CLK(I2350), .RSTB(I139707), .Q(I139990) );
not I_8095 (I139678,I139990);
nand I_8096 (I140021,I139724,I208883);
and I_8097 (I140038,I140021,I139973);
DFFARX1 I_8098  ( .D(I140021), .CLK(I2350), .RSTB(I139707), .Q(I139675) );
DFFARX1 I_8099  ( .D(I208862), .CLK(I2350), .RSTB(I139707), .Q(I140069) );
nor I_8100 (I140086,I140069,I139792);
nand I_8101 (I139693,I139956,I140086);
nor I_8102 (I140117,I140069,I139857);
not I_8103 (I139690,I140069);
nand I_8104 (I140148,I140069,I139758);
and I_8105 (I140165,I139826,I140148);
DFFARX1 I_8106  ( .D(I140165), .CLK(I2350), .RSTB(I139707), .Q(I139669) );
DFFARX1 I_8107  ( .D(I140069), .CLK(I2350), .RSTB(I139707), .Q(I139672) );
DFFARX1 I_8108  ( .D(I208880), .CLK(I2350), .RSTB(I139707), .Q(I140210) );
not I_8109 (I140227,I140210);
nand I_8110 (I140244,I140227,I139792);
and I_8111 (I140261,I140021,I140244);
DFFARX1 I_8112  ( .D(I140261), .CLK(I2350), .RSTB(I139707), .Q(I139699) );
or I_8113 (I140292,I140227,I140038);
DFFARX1 I_8114  ( .D(I140292), .CLK(I2350), .RSTB(I139707), .Q(I139684) );
nand I_8115 (I139687,I140227,I140117);
not I_8116 (I140370,I2357);
not I_8117 (I140387,I313580);
nor I_8118 (I140404,I313577,I313568);
nand I_8119 (I140421,I140404,I313571);
nor I_8120 (I140438,I140387,I313577);
nand I_8121 (I140455,I140438,I313565);
not I_8122 (I140472,I140455);
not I_8123 (I140489,I313577);
nor I_8124 (I140359,I140455,I140489);
not I_8125 (I140520,I140489);
nand I_8126 (I140344,I140455,I140520);
not I_8127 (I140551,I313586);
nor I_8128 (I140568,I140551,I313589);
and I_8129 (I140585,I140568,I313574);
or I_8130 (I140602,I140585,I313562);
DFFARX1 I_8131  ( .D(I140602), .CLK(I2350), .RSTB(I140370), .Q(I140619) );
nor I_8132 (I140636,I140619,I140472);
DFFARX1 I_8133  ( .D(I140619), .CLK(I2350), .RSTB(I140370), .Q(I140653) );
not I_8134 (I140341,I140653);
nand I_8135 (I140684,I140387,I313586);
and I_8136 (I140701,I140684,I140636);
DFFARX1 I_8137  ( .D(I140684), .CLK(I2350), .RSTB(I140370), .Q(I140338) );
DFFARX1 I_8138  ( .D(I313583), .CLK(I2350), .RSTB(I140370), .Q(I140732) );
nor I_8139 (I140749,I140732,I140455);
nand I_8140 (I140356,I140619,I140749);
nor I_8141 (I140780,I140732,I140520);
not I_8142 (I140353,I140732);
nand I_8143 (I140811,I140732,I140421);
and I_8144 (I140828,I140489,I140811);
DFFARX1 I_8145  ( .D(I140828), .CLK(I2350), .RSTB(I140370), .Q(I140332) );
DFFARX1 I_8146  ( .D(I140732), .CLK(I2350), .RSTB(I140370), .Q(I140335) );
DFFARX1 I_8147  ( .D(I313592), .CLK(I2350), .RSTB(I140370), .Q(I140873) );
not I_8148 (I140890,I140873);
nand I_8149 (I140907,I140890,I140455);
and I_8150 (I140924,I140684,I140907);
DFFARX1 I_8151  ( .D(I140924), .CLK(I2350), .RSTB(I140370), .Q(I140362) );
or I_8152 (I140955,I140890,I140701);
DFFARX1 I_8153  ( .D(I140955), .CLK(I2350), .RSTB(I140370), .Q(I140347) );
nand I_8154 (I140350,I140890,I140780);
not I_8155 (I141033,I2357);
not I_8156 (I141050,I274992);
nor I_8157 (I141067,I275013,I275019);
nand I_8158 (I141084,I141067,I275007);
nor I_8159 (I141101,I141050,I275013);
nand I_8160 (I141118,I141101,I274989);
not I_8161 (I141135,I141118);
not I_8162 (I141152,I275013);
nor I_8163 (I141022,I141118,I141152);
not I_8164 (I141183,I141152);
nand I_8165 (I141007,I141118,I141183);
not I_8166 (I141214,I274995);
nor I_8167 (I141231,I141214,I275016);
and I_8168 (I141248,I141231,I275004);
or I_8169 (I141265,I141248,I275010);
DFFARX1 I_8170  ( .D(I141265), .CLK(I2350), .RSTB(I141033), .Q(I141282) );
nor I_8171 (I141299,I141282,I141135);
DFFARX1 I_8172  ( .D(I141282), .CLK(I2350), .RSTB(I141033), .Q(I141316) );
not I_8173 (I141004,I141316);
nand I_8174 (I141347,I141050,I274995);
and I_8175 (I141364,I141347,I141299);
DFFARX1 I_8176  ( .D(I141347), .CLK(I2350), .RSTB(I141033), .Q(I141001) );
DFFARX1 I_8177  ( .D(I275001), .CLK(I2350), .RSTB(I141033), .Q(I141395) );
nor I_8178 (I141412,I141395,I141118);
nand I_8179 (I141019,I141282,I141412);
nor I_8180 (I141443,I141395,I141183);
not I_8181 (I141016,I141395);
nand I_8182 (I141474,I141395,I141084);
and I_8183 (I141491,I141152,I141474);
DFFARX1 I_8184  ( .D(I141491), .CLK(I2350), .RSTB(I141033), .Q(I140995) );
DFFARX1 I_8185  ( .D(I141395), .CLK(I2350), .RSTB(I141033), .Q(I140998) );
DFFARX1 I_8186  ( .D(I274998), .CLK(I2350), .RSTB(I141033), .Q(I141536) );
not I_8187 (I141553,I141536);
nand I_8188 (I141570,I141553,I141118);
and I_8189 (I141587,I141347,I141570);
DFFARX1 I_8190  ( .D(I141587), .CLK(I2350), .RSTB(I141033), .Q(I141025) );
or I_8191 (I141618,I141553,I141364);
DFFARX1 I_8192  ( .D(I141618), .CLK(I2350), .RSTB(I141033), .Q(I141010) );
nand I_8193 (I141013,I141553,I141443);
not I_8194 (I141696,I2357);
not I_8195 (I141713,I58228);
nor I_8196 (I141730,I58225,I58249);
nand I_8197 (I141747,I141730,I58246);
nor I_8198 (I141764,I141713,I58225);
nand I_8199 (I141781,I141764,I58252);
not I_8200 (I141798,I141781);
not I_8201 (I141815,I58225);
nor I_8202 (I141685,I141781,I141815);
not I_8203 (I141846,I141815);
nand I_8204 (I141670,I141781,I141846);
not I_8205 (I141877,I58243);
nor I_8206 (I141894,I141877,I58234);
and I_8207 (I141911,I141894,I58231);
or I_8208 (I141928,I141911,I58240);
DFFARX1 I_8209  ( .D(I141928), .CLK(I2350), .RSTB(I141696), .Q(I141945) );
nor I_8210 (I141962,I141945,I141798);
DFFARX1 I_8211  ( .D(I141945), .CLK(I2350), .RSTB(I141696), .Q(I141979) );
not I_8212 (I141667,I141979);
nand I_8213 (I142010,I141713,I58243);
and I_8214 (I142027,I142010,I141962);
DFFARX1 I_8215  ( .D(I142010), .CLK(I2350), .RSTB(I141696), .Q(I141664) );
DFFARX1 I_8216  ( .D(I58222), .CLK(I2350), .RSTB(I141696), .Q(I142058) );
nor I_8217 (I142075,I142058,I141781);
nand I_8218 (I141682,I141945,I142075);
nor I_8219 (I142106,I142058,I141846);
not I_8220 (I141679,I142058);
nand I_8221 (I142137,I142058,I141747);
and I_8222 (I142154,I141815,I142137);
DFFARX1 I_8223  ( .D(I142154), .CLK(I2350), .RSTB(I141696), .Q(I141658) );
DFFARX1 I_8224  ( .D(I142058), .CLK(I2350), .RSTB(I141696), .Q(I141661) );
DFFARX1 I_8225  ( .D(I58237), .CLK(I2350), .RSTB(I141696), .Q(I142199) );
not I_8226 (I142216,I142199);
nand I_8227 (I142233,I142216,I141781);
and I_8228 (I142250,I142010,I142233);
DFFARX1 I_8229  ( .D(I142250), .CLK(I2350), .RSTB(I141696), .Q(I141688) );
or I_8230 (I142281,I142216,I142027);
DFFARX1 I_8231  ( .D(I142281), .CLK(I2350), .RSTB(I141696), .Q(I141673) );
nand I_8232 (I141676,I142216,I142106);
not I_8233 (I142359,I2357);
not I_8234 (I142376,I357768);
nor I_8235 (I142393,I357786,I357777);
nand I_8236 (I142410,I142393,I357783);
nor I_8237 (I142427,I142376,I357786);
nand I_8238 (I142444,I142427,I357789);
not I_8239 (I142461,I142444);
not I_8240 (I142478,I357786);
nor I_8241 (I142348,I142444,I142478);
not I_8242 (I142509,I142478);
nand I_8243 (I142333,I142444,I142509);
not I_8244 (I142540,I357765);
nor I_8245 (I142557,I142540,I357780);
and I_8246 (I142574,I142557,I357762);
or I_8247 (I142591,I142574,I357771);
DFFARX1 I_8248  ( .D(I142591), .CLK(I2350), .RSTB(I142359), .Q(I142608) );
nor I_8249 (I142625,I142608,I142461);
DFFARX1 I_8250  ( .D(I142608), .CLK(I2350), .RSTB(I142359), .Q(I142642) );
not I_8251 (I142330,I142642);
nand I_8252 (I142673,I142376,I357765);
and I_8253 (I142690,I142673,I142625);
DFFARX1 I_8254  ( .D(I142673), .CLK(I2350), .RSTB(I142359), .Q(I142327) );
DFFARX1 I_8255  ( .D(I357774), .CLK(I2350), .RSTB(I142359), .Q(I142721) );
nor I_8256 (I142738,I142721,I142444);
nand I_8257 (I142345,I142608,I142738);
nor I_8258 (I142769,I142721,I142509);
not I_8259 (I142342,I142721);
nand I_8260 (I142800,I142721,I142410);
and I_8261 (I142817,I142478,I142800);
DFFARX1 I_8262  ( .D(I142817), .CLK(I2350), .RSTB(I142359), .Q(I142321) );
DFFARX1 I_8263  ( .D(I142721), .CLK(I2350), .RSTB(I142359), .Q(I142324) );
DFFARX1 I_8264  ( .D(I357792), .CLK(I2350), .RSTB(I142359), .Q(I142862) );
not I_8265 (I142879,I142862);
nand I_8266 (I142896,I142879,I142444);
and I_8267 (I142913,I142673,I142896);
DFFARX1 I_8268  ( .D(I142913), .CLK(I2350), .RSTB(I142359), .Q(I142351) );
or I_8269 (I142944,I142879,I142690);
DFFARX1 I_8270  ( .D(I142944), .CLK(I2350), .RSTB(I142359), .Q(I142336) );
nand I_8271 (I142339,I142879,I142769);
not I_8272 (I143022,I2357);
not I_8273 (I143039,I69856);
nor I_8274 (I143056,I69853,I69877);
nand I_8275 (I143073,I143056,I69874);
nor I_8276 (I143090,I143039,I69853);
nand I_8277 (I143107,I143090,I69880);
not I_8278 (I143124,I143107);
not I_8279 (I143141,I69853);
nor I_8280 (I143011,I143107,I143141);
not I_8281 (I143172,I143141);
nand I_8282 (I142996,I143107,I143172);
not I_8283 (I143203,I69871);
nor I_8284 (I143220,I143203,I69862);
and I_8285 (I143237,I143220,I69859);
or I_8286 (I143254,I143237,I69868);
DFFARX1 I_8287  ( .D(I143254), .CLK(I2350), .RSTB(I143022), .Q(I143271) );
nor I_8288 (I143288,I143271,I143124);
DFFARX1 I_8289  ( .D(I143271), .CLK(I2350), .RSTB(I143022), .Q(I143305) );
not I_8290 (I142993,I143305);
nand I_8291 (I143336,I143039,I69871);
and I_8292 (I143353,I143336,I143288);
DFFARX1 I_8293  ( .D(I143336), .CLK(I2350), .RSTB(I143022), .Q(I142990) );
DFFARX1 I_8294  ( .D(I69850), .CLK(I2350), .RSTB(I143022), .Q(I143384) );
nor I_8295 (I143401,I143384,I143107);
nand I_8296 (I143008,I143271,I143401);
nor I_8297 (I143432,I143384,I143172);
not I_8298 (I143005,I143384);
nand I_8299 (I143463,I143384,I143073);
and I_8300 (I143480,I143141,I143463);
DFFARX1 I_8301  ( .D(I143480), .CLK(I2350), .RSTB(I143022), .Q(I142984) );
DFFARX1 I_8302  ( .D(I143384), .CLK(I2350), .RSTB(I143022), .Q(I142987) );
DFFARX1 I_8303  ( .D(I69865), .CLK(I2350), .RSTB(I143022), .Q(I143525) );
not I_8304 (I143542,I143525);
nand I_8305 (I143559,I143542,I143107);
and I_8306 (I143576,I143336,I143559);
DFFARX1 I_8307  ( .D(I143576), .CLK(I2350), .RSTB(I143022), .Q(I143014) );
or I_8308 (I143607,I143542,I143353);
DFFARX1 I_8309  ( .D(I143607), .CLK(I2350), .RSTB(I143022), .Q(I142999) );
nand I_8310 (I143002,I143542,I143432);
not I_8311 (I143685,I2357);
not I_8312 (I143702,I201119);
nor I_8313 (I143719,I201116,I201134);
nand I_8314 (I143736,I143719,I201137);
nor I_8315 (I143753,I143702,I201116);
nand I_8316 (I143770,I143753,I201122);
not I_8317 (I143787,I143770);
not I_8318 (I143804,I201116);
nor I_8319 (I143674,I143770,I143804);
not I_8320 (I143835,I143804);
nand I_8321 (I143659,I143770,I143835);
not I_8322 (I143866,I201131);
nor I_8323 (I143883,I143866,I201113);
and I_8324 (I143900,I143883,I201107);
or I_8325 (I143917,I143900,I201125);
DFFARX1 I_8326  ( .D(I143917), .CLK(I2350), .RSTB(I143685), .Q(I143934) );
nor I_8327 (I143951,I143934,I143787);
DFFARX1 I_8328  ( .D(I143934), .CLK(I2350), .RSTB(I143685), .Q(I143968) );
not I_8329 (I143656,I143968);
nand I_8330 (I143999,I143702,I201131);
and I_8331 (I144016,I143999,I143951);
DFFARX1 I_8332  ( .D(I143999), .CLK(I2350), .RSTB(I143685), .Q(I143653) );
DFFARX1 I_8333  ( .D(I201110), .CLK(I2350), .RSTB(I143685), .Q(I144047) );
nor I_8334 (I144064,I144047,I143770);
nand I_8335 (I143671,I143934,I144064);
nor I_8336 (I144095,I144047,I143835);
not I_8337 (I143668,I144047);
nand I_8338 (I144126,I144047,I143736);
and I_8339 (I144143,I143804,I144126);
DFFARX1 I_8340  ( .D(I144143), .CLK(I2350), .RSTB(I143685), .Q(I143647) );
DFFARX1 I_8341  ( .D(I144047), .CLK(I2350), .RSTB(I143685), .Q(I143650) );
DFFARX1 I_8342  ( .D(I201128), .CLK(I2350), .RSTB(I143685), .Q(I144188) );
not I_8343 (I144205,I144188);
nand I_8344 (I144222,I144205,I143770);
and I_8345 (I144239,I143999,I144222);
DFFARX1 I_8346  ( .D(I144239), .CLK(I2350), .RSTB(I143685), .Q(I143677) );
or I_8347 (I144270,I144205,I144016);
DFFARX1 I_8348  ( .D(I144270), .CLK(I2350), .RSTB(I143685), .Q(I143662) );
nand I_8349 (I143665,I144205,I144095);
not I_8350 (I144348,I2357);
not I_8351 (I144365,I262594);
nor I_8352 (I144382,I262606,I262588);
nand I_8353 (I144399,I144382,I262609);
nor I_8354 (I144416,I144365,I262606);
nand I_8355 (I144433,I144416,I262600);
not I_8356 (I144450,I144433);
not I_8357 (I144467,I262606);
nor I_8358 (I144337,I144433,I144467);
not I_8359 (I144498,I144467);
nand I_8360 (I144322,I144433,I144498);
not I_8361 (I144529,I262591);
nor I_8362 (I144546,I144529,I262585);
and I_8363 (I144563,I144546,I262597);
or I_8364 (I144580,I144563,I262582);
DFFARX1 I_8365  ( .D(I144580), .CLK(I2350), .RSTB(I144348), .Q(I144597) );
nor I_8366 (I144614,I144597,I144450);
DFFARX1 I_8367  ( .D(I144597), .CLK(I2350), .RSTB(I144348), .Q(I144631) );
not I_8368 (I144319,I144631);
nand I_8369 (I144662,I144365,I262591);
and I_8370 (I144679,I144662,I144614);
DFFARX1 I_8371  ( .D(I144662), .CLK(I2350), .RSTB(I144348), .Q(I144316) );
DFFARX1 I_8372  ( .D(I262579), .CLK(I2350), .RSTB(I144348), .Q(I144710) );
nor I_8373 (I144727,I144710,I144433);
nand I_8374 (I144334,I144597,I144727);
nor I_8375 (I144758,I144710,I144498);
not I_8376 (I144331,I144710);
nand I_8377 (I144789,I144710,I144399);
and I_8378 (I144806,I144467,I144789);
DFFARX1 I_8379  ( .D(I144806), .CLK(I2350), .RSTB(I144348), .Q(I144310) );
DFFARX1 I_8380  ( .D(I144710), .CLK(I2350), .RSTB(I144348), .Q(I144313) );
DFFARX1 I_8381  ( .D(I262603), .CLK(I2350), .RSTB(I144348), .Q(I144851) );
not I_8382 (I144868,I144851);
nand I_8383 (I144885,I144868,I144433);
and I_8384 (I144902,I144662,I144885);
DFFARX1 I_8385  ( .D(I144902), .CLK(I2350), .RSTB(I144348), .Q(I144340) );
or I_8386 (I144933,I144868,I144679);
DFFARX1 I_8387  ( .D(I144933), .CLK(I2350), .RSTB(I144348), .Q(I144325) );
nand I_8388 (I144328,I144868,I144758);
not I_8389 (I145011,I2357);
not I_8390 (I145028,I16964);
nor I_8391 (I145045,I16970,I16973);
nand I_8392 (I145062,I145045,I16949);
nor I_8393 (I145079,I145028,I16970);
nand I_8394 (I145096,I145079,I16958);
not I_8395 (I145113,I145096);
not I_8396 (I145130,I16970);
nor I_8397 (I145000,I145096,I145130);
not I_8398 (I145161,I145130);
nand I_8399 (I144985,I145096,I145161);
not I_8400 (I145192,I16952);
nor I_8401 (I145209,I145192,I16976);
and I_8402 (I145226,I145209,I16946);
or I_8403 (I145243,I145226,I16955);
DFFARX1 I_8404  ( .D(I145243), .CLK(I2350), .RSTB(I145011), .Q(I145260) );
nor I_8405 (I145277,I145260,I145113);
DFFARX1 I_8406  ( .D(I145260), .CLK(I2350), .RSTB(I145011), .Q(I145294) );
not I_8407 (I144982,I145294);
nand I_8408 (I145325,I145028,I16952);
and I_8409 (I145342,I145325,I145277);
DFFARX1 I_8410  ( .D(I145325), .CLK(I2350), .RSTB(I145011), .Q(I144979) );
DFFARX1 I_8411  ( .D(I16961), .CLK(I2350), .RSTB(I145011), .Q(I145373) );
nor I_8412 (I145390,I145373,I145096);
nand I_8413 (I144997,I145260,I145390);
nor I_8414 (I145421,I145373,I145161);
not I_8415 (I144994,I145373);
nand I_8416 (I145452,I145373,I145062);
and I_8417 (I145469,I145130,I145452);
DFFARX1 I_8418  ( .D(I145469), .CLK(I2350), .RSTB(I145011), .Q(I144973) );
DFFARX1 I_8419  ( .D(I145373), .CLK(I2350), .RSTB(I145011), .Q(I144976) );
DFFARX1 I_8420  ( .D(I16967), .CLK(I2350), .RSTB(I145011), .Q(I145514) );
not I_8421 (I145531,I145514);
nand I_8422 (I145548,I145531,I145096);
and I_8423 (I145565,I145325,I145548);
DFFARX1 I_8424  ( .D(I145565), .CLK(I2350), .RSTB(I145011), .Q(I145003) );
or I_8425 (I145596,I145531,I145342);
DFFARX1 I_8426  ( .D(I145596), .CLK(I2350), .RSTB(I145011), .Q(I144988) );
nand I_8427 (I144991,I145531,I145421);
not I_8428 (I145674,I2357);
not I_8429 (I145691,I382781);
nor I_8430 (I145708,I382772,I382778);
nand I_8431 (I145725,I145708,I382790);
nor I_8432 (I145742,I145691,I382772);
nand I_8433 (I145759,I145742,I382775);
not I_8434 (I145776,I145759);
not I_8435 (I145793,I382772);
nor I_8436 (I145663,I145759,I145793);
not I_8437 (I145824,I145793);
nand I_8438 (I145648,I145759,I145824);
not I_8439 (I145855,I382799);
nor I_8440 (I145872,I145855,I382793);
and I_8441 (I145889,I145872,I382784);
or I_8442 (I145906,I145889,I382769);
DFFARX1 I_8443  ( .D(I145906), .CLK(I2350), .RSTB(I145674), .Q(I145923) );
nor I_8444 (I145940,I145923,I145776);
DFFARX1 I_8445  ( .D(I145923), .CLK(I2350), .RSTB(I145674), .Q(I145957) );
not I_8446 (I145645,I145957);
nand I_8447 (I145988,I145691,I382799);
and I_8448 (I146005,I145988,I145940);
DFFARX1 I_8449  ( .D(I145988), .CLK(I2350), .RSTB(I145674), .Q(I145642) );
DFFARX1 I_8450  ( .D(I382787), .CLK(I2350), .RSTB(I145674), .Q(I146036) );
nor I_8451 (I146053,I146036,I145759);
nand I_8452 (I145660,I145923,I146053);
nor I_8453 (I146084,I146036,I145824);
not I_8454 (I145657,I146036);
nand I_8455 (I146115,I146036,I145725);
and I_8456 (I146132,I145793,I146115);
DFFARX1 I_8457  ( .D(I146132), .CLK(I2350), .RSTB(I145674), .Q(I145636) );
DFFARX1 I_8458  ( .D(I146036), .CLK(I2350), .RSTB(I145674), .Q(I145639) );
DFFARX1 I_8459  ( .D(I382796), .CLK(I2350), .RSTB(I145674), .Q(I146177) );
not I_8460 (I146194,I146177);
nand I_8461 (I146211,I146194,I145759);
and I_8462 (I146228,I145988,I146211);
DFFARX1 I_8463  ( .D(I146228), .CLK(I2350), .RSTB(I145674), .Q(I145666) );
or I_8464 (I146259,I146194,I146005);
DFFARX1 I_8465  ( .D(I146259), .CLK(I2350), .RSTB(I145674), .Q(I145651) );
nand I_8466 (I145654,I146194,I146084);
not I_8467 (I146337,I2357);
not I_8468 (I146354,I199827);
nor I_8469 (I146371,I199824,I199842);
nand I_8470 (I146388,I146371,I199845);
nor I_8471 (I146405,I146354,I199824);
nand I_8472 (I146422,I146405,I199830);
not I_8473 (I146439,I146422);
not I_8474 (I146456,I199824);
nor I_8475 (I146326,I146422,I146456);
not I_8476 (I146487,I146456);
nand I_8477 (I146311,I146422,I146487);
not I_8478 (I146518,I199839);
nor I_8479 (I146535,I146518,I199821);
and I_8480 (I146552,I146535,I199815);
or I_8481 (I146569,I146552,I199833);
DFFARX1 I_8482  ( .D(I146569), .CLK(I2350), .RSTB(I146337), .Q(I146586) );
nor I_8483 (I146603,I146586,I146439);
DFFARX1 I_8484  ( .D(I146586), .CLK(I2350), .RSTB(I146337), .Q(I146620) );
not I_8485 (I146308,I146620);
nand I_8486 (I146651,I146354,I199839);
and I_8487 (I146668,I146651,I146603);
DFFARX1 I_8488  ( .D(I146651), .CLK(I2350), .RSTB(I146337), .Q(I146305) );
DFFARX1 I_8489  ( .D(I199818), .CLK(I2350), .RSTB(I146337), .Q(I146699) );
nor I_8490 (I146716,I146699,I146422);
nand I_8491 (I146323,I146586,I146716);
nor I_8492 (I146747,I146699,I146487);
not I_8493 (I146320,I146699);
nand I_8494 (I146778,I146699,I146388);
and I_8495 (I146795,I146456,I146778);
DFFARX1 I_8496  ( .D(I146795), .CLK(I2350), .RSTB(I146337), .Q(I146299) );
DFFARX1 I_8497  ( .D(I146699), .CLK(I2350), .RSTB(I146337), .Q(I146302) );
DFFARX1 I_8498  ( .D(I199836), .CLK(I2350), .RSTB(I146337), .Q(I146840) );
not I_8499 (I146857,I146840);
nand I_8500 (I146874,I146857,I146422);
and I_8501 (I146891,I146651,I146874);
DFFARX1 I_8502  ( .D(I146891), .CLK(I2350), .RSTB(I146337), .Q(I146329) );
or I_8503 (I146922,I146857,I146668);
DFFARX1 I_8504  ( .D(I146922), .CLK(I2350), .RSTB(I146337), .Q(I146314) );
nand I_8505 (I146317,I146857,I146747);
not I_8506 (I147000,I2357);
not I_8507 (I147017,I13598);
nor I_8508 (I147034,I13604,I13607);
nand I_8509 (I147051,I147034,I13583);
nor I_8510 (I147068,I147017,I13604);
nand I_8511 (I147085,I147068,I13592);
not I_8512 (I147102,I147085);
not I_8513 (I147119,I13604);
nor I_8514 (I146989,I147085,I147119);
not I_8515 (I147150,I147119);
nand I_8516 (I146974,I147085,I147150);
not I_8517 (I147181,I13586);
nor I_8518 (I147198,I147181,I13610);
and I_8519 (I147215,I147198,I13580);
or I_8520 (I147232,I147215,I13589);
DFFARX1 I_8521  ( .D(I147232), .CLK(I2350), .RSTB(I147000), .Q(I147249) );
nor I_8522 (I147266,I147249,I147102);
DFFARX1 I_8523  ( .D(I147249), .CLK(I2350), .RSTB(I147000), .Q(I147283) );
not I_8524 (I146971,I147283);
nand I_8525 (I147314,I147017,I13586);
and I_8526 (I147331,I147314,I147266);
DFFARX1 I_8527  ( .D(I147314), .CLK(I2350), .RSTB(I147000), .Q(I146968) );
DFFARX1 I_8528  ( .D(I13595), .CLK(I2350), .RSTB(I147000), .Q(I147362) );
nor I_8529 (I147379,I147362,I147085);
nand I_8530 (I146986,I147249,I147379);
nor I_8531 (I147410,I147362,I147150);
not I_8532 (I146983,I147362);
nand I_8533 (I147441,I147362,I147051);
and I_8534 (I147458,I147119,I147441);
DFFARX1 I_8535  ( .D(I147458), .CLK(I2350), .RSTB(I147000), .Q(I146962) );
DFFARX1 I_8536  ( .D(I147362), .CLK(I2350), .RSTB(I147000), .Q(I146965) );
DFFARX1 I_8537  ( .D(I13601), .CLK(I2350), .RSTB(I147000), .Q(I147503) );
not I_8538 (I147520,I147503);
nand I_8539 (I147537,I147520,I147085);
and I_8540 (I147554,I147314,I147537);
DFFARX1 I_8541  ( .D(I147554), .CLK(I2350), .RSTB(I147000), .Q(I146992) );
or I_8542 (I147585,I147520,I147331);
DFFARX1 I_8543  ( .D(I147585), .CLK(I2350), .RSTB(I147000), .Q(I146977) );
nand I_8544 (I146980,I147520,I147410);
not I_8545 (I147663,I2357);
not I_8546 (I147680,I99960);
nor I_8547 (I147697,I99966,I99972);
nand I_8548 (I147714,I147697,I99975);
nor I_8549 (I147731,I147680,I99966);
nand I_8550 (I147748,I147731,I99957);
not I_8551 (I147765,I147748);
not I_8552 (I147782,I99966);
nor I_8553 (I147652,I147748,I147782);
not I_8554 (I147813,I147782);
nand I_8555 (I147637,I147748,I147813);
not I_8556 (I147844,I99969);
nor I_8557 (I147861,I147844,I99963);
and I_8558 (I147878,I147861,I99978);
or I_8559 (I147895,I147878,I99984);
DFFARX1 I_8560  ( .D(I147895), .CLK(I2350), .RSTB(I147663), .Q(I147912) );
nor I_8561 (I147929,I147912,I147765);
DFFARX1 I_8562  ( .D(I147912), .CLK(I2350), .RSTB(I147663), .Q(I147946) );
not I_8563 (I147634,I147946);
nand I_8564 (I147977,I147680,I99969);
and I_8565 (I147994,I147977,I147929);
DFFARX1 I_8566  ( .D(I147977), .CLK(I2350), .RSTB(I147663), .Q(I147631) );
DFFARX1 I_8567  ( .D(I99981), .CLK(I2350), .RSTB(I147663), .Q(I148025) );
nor I_8568 (I148042,I148025,I147748);
nand I_8569 (I147649,I147912,I148042);
nor I_8570 (I148073,I148025,I147813);
not I_8571 (I147646,I148025);
nand I_8572 (I148104,I148025,I147714);
and I_8573 (I148121,I147782,I148104);
DFFARX1 I_8574  ( .D(I148121), .CLK(I2350), .RSTB(I147663), .Q(I147625) );
DFFARX1 I_8575  ( .D(I148025), .CLK(I2350), .RSTB(I147663), .Q(I147628) );
DFFARX1 I_8576  ( .D(I99987), .CLK(I2350), .RSTB(I147663), .Q(I148166) );
not I_8577 (I148183,I148166);
nand I_8578 (I148200,I148183,I147748);
and I_8579 (I148217,I147977,I148200);
DFFARX1 I_8580  ( .D(I148217), .CLK(I2350), .RSTB(I147663), .Q(I147655) );
or I_8581 (I148248,I148183,I147994);
DFFARX1 I_8582  ( .D(I148248), .CLK(I2350), .RSTB(I147663), .Q(I147640) );
nand I_8583 (I147643,I148183,I148073);
not I_8584 (I148326,I2357);
not I_8585 (I148343,I379154);
nor I_8586 (I148360,I379172,I379163);
nand I_8587 (I148377,I148360,I379169);
nor I_8588 (I148394,I148343,I379172);
nand I_8589 (I148411,I148394,I379175);
not I_8590 (I148428,I148411);
not I_8591 (I148445,I379172);
nor I_8592 (I148315,I148411,I148445);
not I_8593 (I148476,I148445);
nand I_8594 (I148300,I148411,I148476);
not I_8595 (I148507,I379151);
nor I_8596 (I148524,I148507,I379166);
and I_8597 (I148541,I148524,I379148);
or I_8598 (I148558,I148541,I379157);
DFFARX1 I_8599  ( .D(I148558), .CLK(I2350), .RSTB(I148326), .Q(I148575) );
nor I_8600 (I148592,I148575,I148428);
DFFARX1 I_8601  ( .D(I148575), .CLK(I2350), .RSTB(I148326), .Q(I148609) );
not I_8602 (I148297,I148609);
nand I_8603 (I148640,I148343,I379151);
and I_8604 (I148657,I148640,I148592);
DFFARX1 I_8605  ( .D(I148640), .CLK(I2350), .RSTB(I148326), .Q(I148294) );
DFFARX1 I_8606  ( .D(I379160), .CLK(I2350), .RSTB(I148326), .Q(I148688) );
nor I_8607 (I148705,I148688,I148411);
nand I_8608 (I148312,I148575,I148705);
nor I_8609 (I148736,I148688,I148476);
not I_8610 (I148309,I148688);
nand I_8611 (I148767,I148688,I148377);
and I_8612 (I148784,I148445,I148767);
DFFARX1 I_8613  ( .D(I148784), .CLK(I2350), .RSTB(I148326), .Q(I148288) );
DFFARX1 I_8614  ( .D(I148688), .CLK(I2350), .RSTB(I148326), .Q(I148291) );
DFFARX1 I_8615  ( .D(I379178), .CLK(I2350), .RSTB(I148326), .Q(I148829) );
not I_8616 (I148846,I148829);
nand I_8617 (I148863,I148846,I148411);
and I_8618 (I148880,I148640,I148863);
DFFARX1 I_8619  ( .D(I148880), .CLK(I2350), .RSTB(I148326), .Q(I148318) );
or I_8620 (I148911,I148846,I148657);
DFFARX1 I_8621  ( .D(I148911), .CLK(I2350), .RSTB(I148326), .Q(I148303) );
nand I_8622 (I148306,I148846,I148736);
not I_8623 (I148989,I2357);
not I_8624 (I149006,I37556);
nor I_8625 (I149023,I37553,I37577);
nand I_8626 (I149040,I149023,I37574);
nor I_8627 (I149057,I149006,I37553);
nand I_8628 (I149074,I149057,I37580);
not I_8629 (I149091,I149074);
not I_8630 (I149108,I37553);
nor I_8631 (I148978,I149074,I149108);
not I_8632 (I149139,I149108);
nand I_8633 (I148963,I149074,I149139);
not I_8634 (I149170,I37571);
nor I_8635 (I149187,I149170,I37562);
and I_8636 (I149204,I149187,I37559);
or I_8637 (I149221,I149204,I37568);
DFFARX1 I_8638  ( .D(I149221), .CLK(I2350), .RSTB(I148989), .Q(I149238) );
nor I_8639 (I149255,I149238,I149091);
DFFARX1 I_8640  ( .D(I149238), .CLK(I2350), .RSTB(I148989), .Q(I149272) );
not I_8641 (I148960,I149272);
nand I_8642 (I149303,I149006,I37571);
and I_8643 (I149320,I149303,I149255);
DFFARX1 I_8644  ( .D(I149303), .CLK(I2350), .RSTB(I148989), .Q(I148957) );
DFFARX1 I_8645  ( .D(I37550), .CLK(I2350), .RSTB(I148989), .Q(I149351) );
nor I_8646 (I149368,I149351,I149074);
nand I_8647 (I148975,I149238,I149368);
nor I_8648 (I149399,I149351,I149139);
not I_8649 (I148972,I149351);
nand I_8650 (I149430,I149351,I149040);
and I_8651 (I149447,I149108,I149430);
DFFARX1 I_8652  ( .D(I149447), .CLK(I2350), .RSTB(I148989), .Q(I148951) );
DFFARX1 I_8653  ( .D(I149351), .CLK(I2350), .RSTB(I148989), .Q(I148954) );
DFFARX1 I_8654  ( .D(I37565), .CLK(I2350), .RSTB(I148989), .Q(I149492) );
not I_8655 (I149509,I149492);
nand I_8656 (I149526,I149509,I149074);
and I_8657 (I149543,I149303,I149526);
DFFARX1 I_8658  ( .D(I149543), .CLK(I2350), .RSTB(I148989), .Q(I148981) );
or I_8659 (I149574,I149509,I149320);
DFFARX1 I_8660  ( .D(I149574), .CLK(I2350), .RSTB(I148989), .Q(I148966) );
nand I_8661 (I148969,I149509,I149399);
not I_8662 (I149652,I2357);
not I_8663 (I149669,I305845);
nor I_8664 (I149686,I305854,I305836);
nand I_8665 (I149703,I149686,I305857);
nor I_8666 (I149720,I149669,I305854);
nand I_8667 (I149737,I149720,I305848);
not I_8668 (I149754,I149737);
not I_8669 (I149771,I305854);
nor I_8670 (I149641,I149737,I149771);
not I_8671 (I149802,I149771);
nand I_8672 (I149626,I149737,I149802);
not I_8673 (I149833,I305842);
nor I_8674 (I149850,I149833,I305833);
and I_8675 (I149867,I149850,I305830);
or I_8676 (I149884,I149867,I305827);
DFFARX1 I_8677  ( .D(I149884), .CLK(I2350), .RSTB(I149652), .Q(I149901) );
nor I_8678 (I149918,I149901,I149754);
DFFARX1 I_8679  ( .D(I149901), .CLK(I2350), .RSTB(I149652), .Q(I149935) );
not I_8680 (I149623,I149935);
nand I_8681 (I149966,I149669,I305842);
and I_8682 (I149983,I149966,I149918);
DFFARX1 I_8683  ( .D(I149966), .CLK(I2350), .RSTB(I149652), .Q(I149620) );
DFFARX1 I_8684  ( .D(I305851), .CLK(I2350), .RSTB(I149652), .Q(I150014) );
nor I_8685 (I150031,I150014,I149737);
nand I_8686 (I149638,I149901,I150031);
nor I_8687 (I150062,I150014,I149802);
not I_8688 (I149635,I150014);
nand I_8689 (I150093,I150014,I149703);
and I_8690 (I150110,I149771,I150093);
DFFARX1 I_8691  ( .D(I150110), .CLK(I2350), .RSTB(I149652), .Q(I149614) );
DFFARX1 I_8692  ( .D(I150014), .CLK(I2350), .RSTB(I149652), .Q(I149617) );
DFFARX1 I_8693  ( .D(I305839), .CLK(I2350), .RSTB(I149652), .Q(I150155) );
not I_8694 (I150172,I150155);
nand I_8695 (I150189,I150172,I149737);
and I_8696 (I150206,I149966,I150189);
DFFARX1 I_8697  ( .D(I150206), .CLK(I2350), .RSTB(I149652), .Q(I149644) );
or I_8698 (I150237,I150172,I149983);
DFFARX1 I_8699  ( .D(I150237), .CLK(I2350), .RSTB(I149652), .Q(I149629) );
nand I_8700 (I149632,I150172,I150062);
not I_8701 (I150315,I2357);
not I_8702 (I150332,I117468);
nor I_8703 (I150349,I117462,I117453);
nand I_8704 (I150366,I150349,I117465);
nor I_8705 (I150383,I150332,I117462);
nand I_8706 (I150400,I150383,I117480);
not I_8707 (I150417,I150400);
not I_8708 (I150434,I117462);
nor I_8709 (I150304,I150400,I150434);
not I_8710 (I150465,I150434);
nand I_8711 (I150289,I150400,I150465);
not I_8712 (I150496,I117456);
nor I_8713 (I150513,I150496,I117450);
and I_8714 (I150530,I150513,I117477);
or I_8715 (I150547,I150530,I117474);
DFFARX1 I_8716  ( .D(I150547), .CLK(I2350), .RSTB(I150315), .Q(I150564) );
nor I_8717 (I150581,I150564,I150417);
DFFARX1 I_8718  ( .D(I150564), .CLK(I2350), .RSTB(I150315), .Q(I150598) );
not I_8719 (I150286,I150598);
nand I_8720 (I150629,I150332,I117456);
and I_8721 (I150646,I150629,I150581);
DFFARX1 I_8722  ( .D(I150629), .CLK(I2350), .RSTB(I150315), .Q(I150283) );
DFFARX1 I_8723  ( .D(I117471), .CLK(I2350), .RSTB(I150315), .Q(I150677) );
nor I_8724 (I150694,I150677,I150400);
nand I_8725 (I150301,I150564,I150694);
nor I_8726 (I150725,I150677,I150465);
not I_8727 (I150298,I150677);
nand I_8728 (I150756,I150677,I150366);
and I_8729 (I150773,I150434,I150756);
DFFARX1 I_8730  ( .D(I150773), .CLK(I2350), .RSTB(I150315), .Q(I150277) );
DFFARX1 I_8731  ( .D(I150677), .CLK(I2350), .RSTB(I150315), .Q(I150280) );
DFFARX1 I_8732  ( .D(I117459), .CLK(I2350), .RSTB(I150315), .Q(I150818) );
not I_8733 (I150835,I150818);
nand I_8734 (I150852,I150835,I150400);
and I_8735 (I150869,I150629,I150852);
DFFARX1 I_8736  ( .D(I150869), .CLK(I2350), .RSTB(I150315), .Q(I150307) );
or I_8737 (I150900,I150835,I150646);
DFFARX1 I_8738  ( .D(I150900), .CLK(I2350), .RSTB(I150315), .Q(I150292) );
nand I_8739 (I150295,I150835,I150725);
not I_8740 (I150978,I2357);
not I_8741 (I150995,I22574);
nor I_8742 (I151012,I22580,I22583);
nand I_8743 (I151029,I151012,I22559);
nor I_8744 (I151046,I150995,I22580);
nand I_8745 (I151063,I151046,I22568);
not I_8746 (I151080,I151063);
not I_8747 (I151097,I22580);
nor I_8748 (I150967,I151063,I151097);
not I_8749 (I151128,I151097);
nand I_8750 (I150952,I151063,I151128);
not I_8751 (I151159,I22562);
nor I_8752 (I151176,I151159,I22586);
and I_8753 (I151193,I151176,I22556);
or I_8754 (I151210,I151193,I22565);
DFFARX1 I_8755  ( .D(I151210), .CLK(I2350), .RSTB(I150978), .Q(I151227) );
nor I_8756 (I151244,I151227,I151080);
DFFARX1 I_8757  ( .D(I151227), .CLK(I2350), .RSTB(I150978), .Q(I151261) );
not I_8758 (I150949,I151261);
nand I_8759 (I151292,I150995,I22562);
and I_8760 (I151309,I151292,I151244);
DFFARX1 I_8761  ( .D(I151292), .CLK(I2350), .RSTB(I150978), .Q(I150946) );
DFFARX1 I_8762  ( .D(I22571), .CLK(I2350), .RSTB(I150978), .Q(I151340) );
nor I_8763 (I151357,I151340,I151063);
nand I_8764 (I150964,I151227,I151357);
nor I_8765 (I151388,I151340,I151128);
not I_8766 (I150961,I151340);
nand I_8767 (I151419,I151340,I151029);
and I_8768 (I151436,I151097,I151419);
DFFARX1 I_8769  ( .D(I151436), .CLK(I2350), .RSTB(I150978), .Q(I150940) );
DFFARX1 I_8770  ( .D(I151340), .CLK(I2350), .RSTB(I150978), .Q(I150943) );
DFFARX1 I_8771  ( .D(I22577), .CLK(I2350), .RSTB(I150978), .Q(I151481) );
not I_8772 (I151498,I151481);
nand I_8773 (I151515,I151498,I151063);
and I_8774 (I151532,I151292,I151515);
DFFARX1 I_8775  ( .D(I151532), .CLK(I2350), .RSTB(I150978), .Q(I150970) );
or I_8776 (I151563,I151498,I151309);
DFFARX1 I_8777  ( .D(I151563), .CLK(I2350), .RSTB(I150978), .Q(I150955) );
nand I_8778 (I150958,I151498,I151388);
not I_8779 (I151641,I2357);
not I_8780 (I151658,I45954);
nor I_8781 (I151675,I45951,I45975);
nand I_8782 (I151692,I151675,I45972);
nor I_8783 (I151709,I151658,I45951);
nand I_8784 (I151726,I151709,I45978);
not I_8785 (I151743,I151726);
not I_8786 (I151760,I45951);
nor I_8787 (I151630,I151726,I151760);
not I_8788 (I151791,I151760);
nand I_8789 (I151615,I151726,I151791);
not I_8790 (I151822,I45969);
nor I_8791 (I151839,I151822,I45960);
and I_8792 (I151856,I151839,I45957);
or I_8793 (I151873,I151856,I45966);
DFFARX1 I_8794  ( .D(I151873), .CLK(I2350), .RSTB(I151641), .Q(I151890) );
nor I_8795 (I151907,I151890,I151743);
DFFARX1 I_8796  ( .D(I151890), .CLK(I2350), .RSTB(I151641), .Q(I151924) );
not I_8797 (I151612,I151924);
nand I_8798 (I151955,I151658,I45969);
and I_8799 (I151972,I151955,I151907);
DFFARX1 I_8800  ( .D(I151955), .CLK(I2350), .RSTB(I151641), .Q(I151609) );
DFFARX1 I_8801  ( .D(I45948), .CLK(I2350), .RSTB(I151641), .Q(I152003) );
nor I_8802 (I152020,I152003,I151726);
nand I_8803 (I151627,I151890,I152020);
nor I_8804 (I152051,I152003,I151791);
not I_8805 (I151624,I152003);
nand I_8806 (I152082,I152003,I151692);
and I_8807 (I152099,I151760,I152082);
DFFARX1 I_8808  ( .D(I152099), .CLK(I2350), .RSTB(I151641), .Q(I151603) );
DFFARX1 I_8809  ( .D(I152003), .CLK(I2350), .RSTB(I151641), .Q(I151606) );
DFFARX1 I_8810  ( .D(I45963), .CLK(I2350), .RSTB(I151641), .Q(I152144) );
not I_8811 (I152161,I152144);
nand I_8812 (I152178,I152161,I151726);
and I_8813 (I152195,I151955,I152178);
DFFARX1 I_8814  ( .D(I152195), .CLK(I2350), .RSTB(I151641), .Q(I151633) );
or I_8815 (I152226,I152161,I151972);
DFFARX1 I_8816  ( .D(I152226), .CLK(I2350), .RSTB(I151641), .Q(I151618) );
nand I_8817 (I151621,I152161,I152051);
not I_8818 (I152304,I2357);
not I_8819 (I152321,I201765);
nor I_8820 (I152338,I201762,I201780);
nand I_8821 (I152355,I152338,I201783);
nor I_8822 (I152372,I152321,I201762);
nand I_8823 (I152389,I152372,I201768);
not I_8824 (I152406,I152389);
not I_8825 (I152423,I201762);
nor I_8826 (I152293,I152389,I152423);
not I_8827 (I152454,I152423);
nand I_8828 (I152278,I152389,I152454);
not I_8829 (I152485,I201777);
nor I_8830 (I152502,I152485,I201759);
and I_8831 (I152519,I152502,I201753);
or I_8832 (I152536,I152519,I201771);
DFFARX1 I_8833  ( .D(I152536), .CLK(I2350), .RSTB(I152304), .Q(I152553) );
nor I_8834 (I152570,I152553,I152406);
DFFARX1 I_8835  ( .D(I152553), .CLK(I2350), .RSTB(I152304), .Q(I152587) );
not I_8836 (I152275,I152587);
nand I_8837 (I152618,I152321,I201777);
and I_8838 (I152635,I152618,I152570);
DFFARX1 I_8839  ( .D(I152618), .CLK(I2350), .RSTB(I152304), .Q(I152272) );
DFFARX1 I_8840  ( .D(I201756), .CLK(I2350), .RSTB(I152304), .Q(I152666) );
nor I_8841 (I152683,I152666,I152389);
nand I_8842 (I152290,I152553,I152683);
nor I_8843 (I152714,I152666,I152454);
not I_8844 (I152287,I152666);
nand I_8845 (I152745,I152666,I152355);
and I_8846 (I152762,I152423,I152745);
DFFARX1 I_8847  ( .D(I152762), .CLK(I2350), .RSTB(I152304), .Q(I152266) );
DFFARX1 I_8848  ( .D(I152666), .CLK(I2350), .RSTB(I152304), .Q(I152269) );
DFFARX1 I_8849  ( .D(I201774), .CLK(I2350), .RSTB(I152304), .Q(I152807) );
not I_8850 (I152824,I152807);
nand I_8851 (I152841,I152824,I152389);
and I_8852 (I152858,I152618,I152841);
DFFARX1 I_8853  ( .D(I152858), .CLK(I2350), .RSTB(I152304), .Q(I152296) );
or I_8854 (I152889,I152824,I152635);
DFFARX1 I_8855  ( .D(I152889), .CLK(I2350), .RSTB(I152304), .Q(I152281) );
nand I_8856 (I152284,I152824,I152714);
not I_8857 (I152967,I2357);
not I_8858 (I152984,I302275);
nor I_8859 (I153001,I302284,I302266);
nand I_8860 (I153018,I153001,I302287);
nor I_8861 (I153035,I152984,I302284);
nand I_8862 (I153052,I153035,I302278);
not I_8863 (I153069,I153052);
not I_8864 (I153086,I302284);
nor I_8865 (I152956,I153052,I153086);
not I_8866 (I153117,I153086);
nand I_8867 (I152941,I153052,I153117);
not I_8868 (I153148,I302272);
nor I_8869 (I153165,I153148,I302263);
and I_8870 (I153182,I153165,I302260);
or I_8871 (I153199,I153182,I302257);
DFFARX1 I_8872  ( .D(I153199), .CLK(I2350), .RSTB(I152967), .Q(I153216) );
nor I_8873 (I153233,I153216,I153069);
DFFARX1 I_8874  ( .D(I153216), .CLK(I2350), .RSTB(I152967), .Q(I153250) );
not I_8875 (I152938,I153250);
nand I_8876 (I153281,I152984,I302272);
and I_8877 (I153298,I153281,I153233);
DFFARX1 I_8878  ( .D(I153281), .CLK(I2350), .RSTB(I152967), .Q(I152935) );
DFFARX1 I_8879  ( .D(I302281), .CLK(I2350), .RSTB(I152967), .Q(I153329) );
nor I_8880 (I153346,I153329,I153052);
nand I_8881 (I152953,I153216,I153346);
nor I_8882 (I153377,I153329,I153117);
not I_8883 (I152950,I153329);
nand I_8884 (I153408,I153329,I153018);
and I_8885 (I153425,I153086,I153408);
DFFARX1 I_8886  ( .D(I153425), .CLK(I2350), .RSTB(I152967), .Q(I152929) );
DFFARX1 I_8887  ( .D(I153329), .CLK(I2350), .RSTB(I152967), .Q(I152932) );
DFFARX1 I_8888  ( .D(I302269), .CLK(I2350), .RSTB(I152967), .Q(I153470) );
not I_8889 (I153487,I153470);
nand I_8890 (I153504,I153487,I153052);
and I_8891 (I153521,I153281,I153504);
DFFARX1 I_8892  ( .D(I153521), .CLK(I2350), .RSTB(I152967), .Q(I152959) );
or I_8893 (I153552,I153487,I153298);
DFFARX1 I_8894  ( .D(I153552), .CLK(I2350), .RSTB(I152967), .Q(I152944) );
nand I_8895 (I152947,I153487,I153377);
not I_8896 (I153630,I2357);
not I_8897 (I153647,I273836);
nor I_8898 (I153664,I273857,I273863);
nand I_8899 (I153681,I153664,I273851);
nor I_8900 (I153698,I153647,I273857);
nand I_8901 (I153715,I153698,I273833);
not I_8902 (I153732,I153715);
not I_8903 (I153749,I273857);
nor I_8904 (I153619,I153715,I153749);
not I_8905 (I153780,I153749);
nand I_8906 (I153604,I153715,I153780);
not I_8907 (I153811,I273839);
nor I_8908 (I153828,I153811,I273860);
and I_8909 (I153845,I153828,I273848);
or I_8910 (I153862,I153845,I273854);
DFFARX1 I_8911  ( .D(I153862), .CLK(I2350), .RSTB(I153630), .Q(I153879) );
nor I_8912 (I153896,I153879,I153732);
DFFARX1 I_8913  ( .D(I153879), .CLK(I2350), .RSTB(I153630), .Q(I153913) );
not I_8914 (I153601,I153913);
nand I_8915 (I153944,I153647,I273839);
and I_8916 (I153961,I153944,I153896);
DFFARX1 I_8917  ( .D(I153944), .CLK(I2350), .RSTB(I153630), .Q(I153598) );
DFFARX1 I_8918  ( .D(I273845), .CLK(I2350), .RSTB(I153630), .Q(I153992) );
nor I_8919 (I154009,I153992,I153715);
nand I_8920 (I153616,I153879,I154009);
nor I_8921 (I154040,I153992,I153780);
not I_8922 (I153613,I153992);
nand I_8923 (I154071,I153992,I153681);
and I_8924 (I154088,I153749,I154071);
DFFARX1 I_8925  ( .D(I154088), .CLK(I2350), .RSTB(I153630), .Q(I153592) );
DFFARX1 I_8926  ( .D(I153992), .CLK(I2350), .RSTB(I153630), .Q(I153595) );
DFFARX1 I_8927  ( .D(I273842), .CLK(I2350), .RSTB(I153630), .Q(I154133) );
not I_8928 (I154150,I154133);
nand I_8929 (I154167,I154150,I153715);
and I_8930 (I154184,I153944,I154167);
DFFARX1 I_8931  ( .D(I154184), .CLK(I2350), .RSTB(I153630), .Q(I153622) );
or I_8932 (I154215,I154150,I153961);
DFFARX1 I_8933  ( .D(I154215), .CLK(I2350), .RSTB(I153630), .Q(I153607) );
nand I_8934 (I153610,I154150,I154040);
not I_8935 (I154293,I2357);
not I_8936 (I154310,I108579);
nor I_8937 (I154327,I108585,I108591);
nand I_8938 (I154344,I154327,I108594);
nor I_8939 (I154361,I154310,I108585);
nand I_8940 (I154378,I154361,I108576);
not I_8941 (I154395,I154378);
not I_8942 (I154412,I108585);
nor I_8943 (I154282,I154378,I154412);
not I_8944 (I154443,I154412);
nand I_8945 (I154267,I154378,I154443);
not I_8946 (I154474,I108588);
nor I_8947 (I154491,I154474,I108582);
and I_8948 (I154508,I154491,I108597);
or I_8949 (I154525,I154508,I108603);
DFFARX1 I_8950  ( .D(I154525), .CLK(I2350), .RSTB(I154293), .Q(I154542) );
nor I_8951 (I154559,I154542,I154395);
DFFARX1 I_8952  ( .D(I154542), .CLK(I2350), .RSTB(I154293), .Q(I154576) );
not I_8953 (I154264,I154576);
nand I_8954 (I154607,I154310,I108588);
and I_8955 (I154624,I154607,I154559);
DFFARX1 I_8956  ( .D(I154607), .CLK(I2350), .RSTB(I154293), .Q(I154261) );
DFFARX1 I_8957  ( .D(I108600), .CLK(I2350), .RSTB(I154293), .Q(I154655) );
nor I_8958 (I154672,I154655,I154378);
nand I_8959 (I154279,I154542,I154672);
nor I_8960 (I154703,I154655,I154443);
not I_8961 (I154276,I154655);
nand I_8962 (I154734,I154655,I154344);
and I_8963 (I154751,I154412,I154734);
DFFARX1 I_8964  ( .D(I154751), .CLK(I2350), .RSTB(I154293), .Q(I154255) );
DFFARX1 I_8965  ( .D(I154655), .CLK(I2350), .RSTB(I154293), .Q(I154258) );
DFFARX1 I_8966  ( .D(I108606), .CLK(I2350), .RSTB(I154293), .Q(I154796) );
not I_8967 (I154813,I154796);
nand I_8968 (I154830,I154813,I154378);
and I_8969 (I154847,I154607,I154830);
DFFARX1 I_8970  ( .D(I154847), .CLK(I2350), .RSTB(I154293), .Q(I154285) );
or I_8971 (I154878,I154813,I154624);
DFFARX1 I_8972  ( .D(I154878), .CLK(I2350), .RSTB(I154293), .Q(I154270) );
nand I_8973 (I154273,I154813,I154703);
not I_8974 (I154956,I2357);
not I_8975 (I154973,I279665);
nor I_8976 (I154990,I279674,I279656);
nand I_8977 (I155007,I154990,I279677);
nor I_8978 (I155024,I154973,I279674);
nand I_8979 (I155041,I155024,I279668);
not I_8980 (I155058,I155041);
not I_8981 (I155075,I279674);
nor I_8982 (I154945,I155041,I155075);
not I_8983 (I155106,I155075);
nand I_8984 (I154930,I155041,I155106);
not I_8985 (I155137,I279662);
nor I_8986 (I155154,I155137,I279653);
and I_8987 (I155171,I155154,I279650);
or I_8988 (I155188,I155171,I279647);
DFFARX1 I_8989  ( .D(I155188), .CLK(I2350), .RSTB(I154956), .Q(I155205) );
nor I_8990 (I155222,I155205,I155058);
DFFARX1 I_8991  ( .D(I155205), .CLK(I2350), .RSTB(I154956), .Q(I155239) );
not I_8992 (I154927,I155239);
nand I_8993 (I155270,I154973,I279662);
and I_8994 (I155287,I155270,I155222);
DFFARX1 I_8995  ( .D(I155270), .CLK(I2350), .RSTB(I154956), .Q(I154924) );
DFFARX1 I_8996  ( .D(I279671), .CLK(I2350), .RSTB(I154956), .Q(I155318) );
nor I_8997 (I155335,I155318,I155041);
nand I_8998 (I154942,I155205,I155335);
nor I_8999 (I155366,I155318,I155106);
not I_9000 (I154939,I155318);
nand I_9001 (I155397,I155318,I155007);
and I_9002 (I155414,I155075,I155397);
DFFARX1 I_9003  ( .D(I155414), .CLK(I2350), .RSTB(I154956), .Q(I154918) );
DFFARX1 I_9004  ( .D(I155318), .CLK(I2350), .RSTB(I154956), .Q(I154921) );
DFFARX1 I_9005  ( .D(I279659), .CLK(I2350), .RSTB(I154956), .Q(I155459) );
not I_9006 (I155476,I155459);
nand I_9007 (I155493,I155476,I155041);
and I_9008 (I155510,I155270,I155493);
DFFARX1 I_9009  ( .D(I155510), .CLK(I2350), .RSTB(I154956), .Q(I154948) );
or I_9010 (I155541,I155476,I155287);
DFFARX1 I_9011  ( .D(I155541), .CLK(I2350), .RSTB(I154956), .Q(I154933) );
nand I_9012 (I154936,I155476,I155366);
not I_9013 (I155619,I2357);
not I_9014 (I155636,I204349);
nor I_9015 (I155653,I204346,I204364);
nand I_9016 (I155670,I155653,I204367);
nor I_9017 (I155687,I155636,I204346);
nand I_9018 (I155704,I155687,I204352);
not I_9019 (I155721,I155704);
not I_9020 (I155738,I204346);
nor I_9021 (I155608,I155704,I155738);
not I_9022 (I155769,I155738);
nand I_9023 (I155593,I155704,I155769);
not I_9024 (I155800,I204361);
nor I_9025 (I155817,I155800,I204343);
and I_9026 (I155834,I155817,I204337);
or I_9027 (I155851,I155834,I204355);
DFFARX1 I_9028  ( .D(I155851), .CLK(I2350), .RSTB(I155619), .Q(I155868) );
nor I_9029 (I155885,I155868,I155721);
DFFARX1 I_9030  ( .D(I155868), .CLK(I2350), .RSTB(I155619), .Q(I155902) );
not I_9031 (I155590,I155902);
nand I_9032 (I155933,I155636,I204361);
and I_9033 (I155950,I155933,I155885);
DFFARX1 I_9034  ( .D(I155933), .CLK(I2350), .RSTB(I155619), .Q(I155587) );
DFFARX1 I_9035  ( .D(I204340), .CLK(I2350), .RSTB(I155619), .Q(I155981) );
nor I_9036 (I155998,I155981,I155704);
nand I_9037 (I155605,I155868,I155998);
nor I_9038 (I156029,I155981,I155769);
not I_9039 (I155602,I155981);
nand I_9040 (I156060,I155981,I155670);
and I_9041 (I156077,I155738,I156060);
DFFARX1 I_9042  ( .D(I156077), .CLK(I2350), .RSTB(I155619), .Q(I155581) );
DFFARX1 I_9043  ( .D(I155981), .CLK(I2350), .RSTB(I155619), .Q(I155584) );
DFFARX1 I_9044  ( .D(I204358), .CLK(I2350), .RSTB(I155619), .Q(I156122) );
not I_9045 (I156139,I156122);
nand I_9046 (I156156,I156139,I155704);
and I_9047 (I156173,I155933,I156156);
DFFARX1 I_9048  ( .D(I156173), .CLK(I2350), .RSTB(I155619), .Q(I155611) );
or I_9049 (I156204,I156139,I155950);
DFFARX1 I_9050  ( .D(I156204), .CLK(I2350), .RSTB(I155619), .Q(I155596) );
nand I_9051 (I155599,I156139,I156029);
not I_9052 (I156282,I2357);
not I_9053 (I156299,I377267);
nor I_9054 (I156316,I377285,I377276);
nand I_9055 (I156333,I156316,I377282);
nor I_9056 (I156350,I156299,I377285);
nand I_9057 (I156367,I156350,I377288);
not I_9058 (I156384,I156367);
not I_9059 (I156401,I377285);
nor I_9060 (I156271,I156367,I156401);
not I_9061 (I156432,I156401);
nand I_9062 (I156256,I156367,I156432);
not I_9063 (I156463,I377264);
nor I_9064 (I156480,I156463,I377279);
and I_9065 (I156497,I156480,I377261);
or I_9066 (I156514,I156497,I377270);
DFFARX1 I_9067  ( .D(I156514), .CLK(I2350), .RSTB(I156282), .Q(I156531) );
nor I_9068 (I156548,I156531,I156384);
DFFARX1 I_9069  ( .D(I156531), .CLK(I2350), .RSTB(I156282), .Q(I156565) );
not I_9070 (I156253,I156565);
nand I_9071 (I156596,I156299,I377264);
and I_9072 (I156613,I156596,I156548);
DFFARX1 I_9073  ( .D(I156596), .CLK(I2350), .RSTB(I156282), .Q(I156250) );
DFFARX1 I_9074  ( .D(I377273), .CLK(I2350), .RSTB(I156282), .Q(I156644) );
nor I_9075 (I156661,I156644,I156367);
nand I_9076 (I156268,I156531,I156661);
nor I_9077 (I156692,I156644,I156432);
not I_9078 (I156265,I156644);
nand I_9079 (I156723,I156644,I156333);
and I_9080 (I156740,I156401,I156723);
DFFARX1 I_9081  ( .D(I156740), .CLK(I2350), .RSTB(I156282), .Q(I156244) );
DFFARX1 I_9082  ( .D(I156644), .CLK(I2350), .RSTB(I156282), .Q(I156247) );
DFFARX1 I_9083  ( .D(I377291), .CLK(I2350), .RSTB(I156282), .Q(I156785) );
not I_9084 (I156802,I156785);
nand I_9085 (I156819,I156802,I156367);
and I_9086 (I156836,I156596,I156819);
DFFARX1 I_9087  ( .D(I156836), .CLK(I2350), .RSTB(I156282), .Q(I156274) );
or I_9088 (I156867,I156802,I156613);
DFFARX1 I_9089  ( .D(I156867), .CLK(I2350), .RSTB(I156282), .Q(I156259) );
nand I_9090 (I156262,I156802,I156692);
not I_9091 (I156945,I2357);
not I_9092 (I156962,I30450);
nor I_9093 (I156979,I30447,I30471);
nand I_9094 (I156996,I156979,I30468);
nor I_9095 (I157013,I156962,I30447);
nand I_9096 (I157030,I157013,I30474);
not I_9097 (I157047,I157030);
not I_9098 (I157064,I30447);
nor I_9099 (I156934,I157030,I157064);
not I_9100 (I157095,I157064);
nand I_9101 (I156919,I157030,I157095);
not I_9102 (I157126,I30465);
nor I_9103 (I157143,I157126,I30456);
and I_9104 (I157160,I157143,I30453);
or I_9105 (I157177,I157160,I30462);
DFFARX1 I_9106  ( .D(I157177), .CLK(I2350), .RSTB(I156945), .Q(I157194) );
nor I_9107 (I157211,I157194,I157047);
DFFARX1 I_9108  ( .D(I157194), .CLK(I2350), .RSTB(I156945), .Q(I157228) );
not I_9109 (I156916,I157228);
nand I_9110 (I157259,I156962,I30465);
and I_9111 (I157276,I157259,I157211);
DFFARX1 I_9112  ( .D(I157259), .CLK(I2350), .RSTB(I156945), .Q(I156913) );
DFFARX1 I_9113  ( .D(I30444), .CLK(I2350), .RSTB(I156945), .Q(I157307) );
nor I_9114 (I157324,I157307,I157030);
nand I_9115 (I156931,I157194,I157324);
nor I_9116 (I157355,I157307,I157095);
not I_9117 (I156928,I157307);
nand I_9118 (I157386,I157307,I156996);
and I_9119 (I157403,I157064,I157386);
DFFARX1 I_9120  ( .D(I157403), .CLK(I2350), .RSTB(I156945), .Q(I156907) );
DFFARX1 I_9121  ( .D(I157307), .CLK(I2350), .RSTB(I156945), .Q(I156910) );
DFFARX1 I_9122  ( .D(I30459), .CLK(I2350), .RSTB(I156945), .Q(I157448) );
not I_9123 (I157465,I157448);
nand I_9124 (I157482,I157465,I157030);
and I_9125 (I157499,I157259,I157482);
DFFARX1 I_9126  ( .D(I157499), .CLK(I2350), .RSTB(I156945), .Q(I156937) );
or I_9127 (I157530,I157465,I157276);
DFFARX1 I_9128  ( .D(I157530), .CLK(I2350), .RSTB(I156945), .Q(I156922) );
nand I_9129 (I156925,I157465,I157355);
not I_9130 (I157608,I2357);
not I_9131 (I157625,I87363);
nor I_9132 (I157642,I87369,I87375);
nand I_9133 (I157659,I157642,I87378);
nor I_9134 (I157676,I157625,I87369);
nand I_9135 (I157693,I157676,I87360);
not I_9136 (I157710,I157693);
not I_9137 (I157727,I87369);
nor I_9138 (I157597,I157693,I157727);
not I_9139 (I157758,I157727);
nand I_9140 (I157582,I157693,I157758);
not I_9141 (I157789,I87372);
nor I_9142 (I157806,I157789,I87366);
and I_9143 (I157823,I157806,I87381);
or I_9144 (I157840,I157823,I87387);
DFFARX1 I_9145  ( .D(I157840), .CLK(I2350), .RSTB(I157608), .Q(I157857) );
nor I_9146 (I157874,I157857,I157710);
DFFARX1 I_9147  ( .D(I157857), .CLK(I2350), .RSTB(I157608), .Q(I157891) );
not I_9148 (I157579,I157891);
nand I_9149 (I157922,I157625,I87372);
and I_9150 (I157939,I157922,I157874);
DFFARX1 I_9151  ( .D(I157922), .CLK(I2350), .RSTB(I157608), .Q(I157576) );
DFFARX1 I_9152  ( .D(I87384), .CLK(I2350), .RSTB(I157608), .Q(I157970) );
nor I_9153 (I157987,I157970,I157693);
nand I_9154 (I157594,I157857,I157987);
nor I_9155 (I158018,I157970,I157758);
not I_9156 (I157591,I157970);
nand I_9157 (I158049,I157970,I157659);
and I_9158 (I158066,I157727,I158049);
DFFARX1 I_9159  ( .D(I158066), .CLK(I2350), .RSTB(I157608), .Q(I157570) );
DFFARX1 I_9160  ( .D(I157970), .CLK(I2350), .RSTB(I157608), .Q(I157573) );
DFFARX1 I_9161  ( .D(I87390), .CLK(I2350), .RSTB(I157608), .Q(I158111) );
not I_9162 (I158128,I158111);
nand I_9163 (I158145,I158128,I157693);
and I_9164 (I158162,I157922,I158145);
DFFARX1 I_9165  ( .D(I158162), .CLK(I2350), .RSTB(I157608), .Q(I157600) );
or I_9166 (I158193,I158128,I157939);
DFFARX1 I_9167  ( .D(I158193), .CLK(I2350), .RSTB(I157608), .Q(I157585) );
nand I_9168 (I157588,I158128,I158018);
not I_9169 (I158271,I2357);
not I_9170 (I158288,I3500);
nor I_9171 (I158305,I3506,I3509);
nand I_9172 (I158322,I158305,I3485);
nor I_9173 (I158339,I158288,I3506);
nand I_9174 (I158356,I158339,I3494);
not I_9175 (I158373,I158356);
not I_9176 (I158390,I3506);
nor I_9177 (I158260,I158356,I158390);
not I_9178 (I158421,I158390);
nand I_9179 (I158245,I158356,I158421);
not I_9180 (I158452,I3488);
nor I_9181 (I158469,I158452,I3512);
and I_9182 (I158486,I158469,I3482);
or I_9183 (I158503,I158486,I3491);
DFFARX1 I_9184  ( .D(I158503), .CLK(I2350), .RSTB(I158271), .Q(I158520) );
nor I_9185 (I158537,I158520,I158373);
DFFARX1 I_9186  ( .D(I158520), .CLK(I2350), .RSTB(I158271), .Q(I158554) );
not I_9187 (I158242,I158554);
nand I_9188 (I158585,I158288,I3488);
and I_9189 (I158602,I158585,I158537);
DFFARX1 I_9190  ( .D(I158585), .CLK(I2350), .RSTB(I158271), .Q(I158239) );
DFFARX1 I_9191  ( .D(I3497), .CLK(I2350), .RSTB(I158271), .Q(I158633) );
nor I_9192 (I158650,I158633,I158356);
nand I_9193 (I158257,I158520,I158650);
nor I_9194 (I158681,I158633,I158421);
not I_9195 (I158254,I158633);
nand I_9196 (I158712,I158633,I158322);
and I_9197 (I158729,I158390,I158712);
DFFARX1 I_9198  ( .D(I158729), .CLK(I2350), .RSTB(I158271), .Q(I158233) );
DFFARX1 I_9199  ( .D(I158633), .CLK(I2350), .RSTB(I158271), .Q(I158236) );
DFFARX1 I_9200  ( .D(I3503), .CLK(I2350), .RSTB(I158271), .Q(I158774) );
not I_9201 (I158791,I158774);
nand I_9202 (I158808,I158791,I158356);
and I_9203 (I158825,I158585,I158808);
DFFARX1 I_9204  ( .D(I158825), .CLK(I2350), .RSTB(I158271), .Q(I158263) );
or I_9205 (I158856,I158791,I158602);
DFFARX1 I_9206  ( .D(I158856), .CLK(I2350), .RSTB(I158271), .Q(I158248) );
nand I_9207 (I158251,I158791,I158681);
not I_9208 (I158934,I2357);
not I_9209 (I158951,I277882);
nor I_9210 (I158968,I277903,I277909);
nand I_9211 (I158985,I158968,I277897);
nor I_9212 (I159002,I158951,I277903);
nand I_9213 (I159019,I159002,I277879);
not I_9214 (I159036,I159019);
not I_9215 (I159053,I277903);
nor I_9216 (I158923,I159019,I159053);
not I_9217 (I159084,I159053);
nand I_9218 (I158908,I159019,I159084);
not I_9219 (I159115,I277885);
nor I_9220 (I159132,I159115,I277906);
and I_9221 (I159149,I159132,I277894);
or I_9222 (I159166,I159149,I277900);
DFFARX1 I_9223  ( .D(I159166), .CLK(I2350), .RSTB(I158934), .Q(I159183) );
nor I_9224 (I159200,I159183,I159036);
DFFARX1 I_9225  ( .D(I159183), .CLK(I2350), .RSTB(I158934), .Q(I159217) );
not I_9226 (I158905,I159217);
nand I_9227 (I159248,I158951,I277885);
and I_9228 (I159265,I159248,I159200);
DFFARX1 I_9229  ( .D(I159248), .CLK(I2350), .RSTB(I158934), .Q(I158902) );
DFFARX1 I_9230  ( .D(I277891), .CLK(I2350), .RSTB(I158934), .Q(I159296) );
nor I_9231 (I159313,I159296,I159019);
nand I_9232 (I158920,I159183,I159313);
nor I_9233 (I159344,I159296,I159084);
not I_9234 (I158917,I159296);
nand I_9235 (I159375,I159296,I158985);
and I_9236 (I159392,I159053,I159375);
DFFARX1 I_9237  ( .D(I159392), .CLK(I2350), .RSTB(I158934), .Q(I158896) );
DFFARX1 I_9238  ( .D(I159296), .CLK(I2350), .RSTB(I158934), .Q(I158899) );
DFFARX1 I_9239  ( .D(I277888), .CLK(I2350), .RSTB(I158934), .Q(I159437) );
not I_9240 (I159454,I159437);
nand I_9241 (I159471,I159454,I159019);
and I_9242 (I159488,I159248,I159471);
DFFARX1 I_9243  ( .D(I159488), .CLK(I2350), .RSTB(I158934), .Q(I158926) );
or I_9244 (I159519,I159454,I159265);
DFFARX1 I_9245  ( .D(I159519), .CLK(I2350), .RSTB(I158934), .Q(I158911) );
nand I_9246 (I158914,I159454,I159344);
not I_9247 (I159597,I2357);
not I_9248 (I159614,I272680);
nor I_9249 (I159631,I272701,I272707);
nand I_9250 (I159648,I159631,I272695);
nor I_9251 (I159665,I159614,I272701);
nand I_9252 (I159682,I159665,I272677);
not I_9253 (I159699,I159682);
not I_9254 (I159716,I272701);
nor I_9255 (I159586,I159682,I159716);
not I_9256 (I159747,I159716);
nand I_9257 (I159571,I159682,I159747);
not I_9258 (I159778,I272683);
nor I_9259 (I159795,I159778,I272704);
and I_9260 (I159812,I159795,I272692);
or I_9261 (I159829,I159812,I272698);
DFFARX1 I_9262  ( .D(I159829), .CLK(I2350), .RSTB(I159597), .Q(I159846) );
nor I_9263 (I159863,I159846,I159699);
DFFARX1 I_9264  ( .D(I159846), .CLK(I2350), .RSTB(I159597), .Q(I159880) );
not I_9265 (I159568,I159880);
nand I_9266 (I159911,I159614,I272683);
and I_9267 (I159928,I159911,I159863);
DFFARX1 I_9268  ( .D(I159911), .CLK(I2350), .RSTB(I159597), .Q(I159565) );
DFFARX1 I_9269  ( .D(I272689), .CLK(I2350), .RSTB(I159597), .Q(I159959) );
nor I_9270 (I159976,I159959,I159682);
nand I_9271 (I159583,I159846,I159976);
nor I_9272 (I160007,I159959,I159747);
not I_9273 (I159580,I159959);
nand I_9274 (I160038,I159959,I159648);
and I_9275 (I160055,I159716,I160038);
DFFARX1 I_9276  ( .D(I160055), .CLK(I2350), .RSTB(I159597), .Q(I159559) );
DFFARX1 I_9277  ( .D(I159959), .CLK(I2350), .RSTB(I159597), .Q(I159562) );
DFFARX1 I_9278  ( .D(I272686), .CLK(I2350), .RSTB(I159597), .Q(I160100) );
not I_9279 (I160117,I160100);
nand I_9280 (I160134,I160117,I159682);
and I_9281 (I160151,I159911,I160134);
DFFARX1 I_9282  ( .D(I160151), .CLK(I2350), .RSTB(I159597), .Q(I159589) );
or I_9283 (I160182,I160117,I159928);
DFFARX1 I_9284  ( .D(I160182), .CLK(I2350), .RSTB(I159597), .Q(I159574) );
nand I_9285 (I159577,I160117,I160007);
not I_9286 (I160260,I2357);
not I_9287 (I160277,I330240);
nor I_9288 (I160294,I330237,I330228);
nand I_9289 (I160311,I160294,I330231);
nor I_9290 (I160328,I160277,I330237);
nand I_9291 (I160345,I160328,I330225);
not I_9292 (I160362,I160345);
not I_9293 (I160379,I330237);
nor I_9294 (I160249,I160345,I160379);
not I_9295 (I160410,I160379);
nand I_9296 (I160234,I160345,I160410);
not I_9297 (I160441,I330246);
nor I_9298 (I160458,I160441,I330249);
and I_9299 (I160475,I160458,I330234);
or I_9300 (I160492,I160475,I330222);
DFFARX1 I_9301  ( .D(I160492), .CLK(I2350), .RSTB(I160260), .Q(I160509) );
nor I_9302 (I160526,I160509,I160362);
DFFARX1 I_9303  ( .D(I160509), .CLK(I2350), .RSTB(I160260), .Q(I160543) );
not I_9304 (I160231,I160543);
nand I_9305 (I160574,I160277,I330246);
and I_9306 (I160591,I160574,I160526);
DFFARX1 I_9307  ( .D(I160574), .CLK(I2350), .RSTB(I160260), .Q(I160228) );
DFFARX1 I_9308  ( .D(I330243), .CLK(I2350), .RSTB(I160260), .Q(I160622) );
nor I_9309 (I160639,I160622,I160345);
nand I_9310 (I160246,I160509,I160639);
nor I_9311 (I160670,I160622,I160410);
not I_9312 (I160243,I160622);
nand I_9313 (I160701,I160622,I160311);
and I_9314 (I160718,I160379,I160701);
DFFARX1 I_9315  ( .D(I160718), .CLK(I2350), .RSTB(I160260), .Q(I160222) );
DFFARX1 I_9316  ( .D(I160622), .CLK(I2350), .RSTB(I160260), .Q(I160225) );
DFFARX1 I_9317  ( .D(I330252), .CLK(I2350), .RSTB(I160260), .Q(I160763) );
not I_9318 (I160780,I160763);
nand I_9319 (I160797,I160780,I160345);
and I_9320 (I160814,I160574,I160797);
DFFARX1 I_9321  ( .D(I160814), .CLK(I2350), .RSTB(I160260), .Q(I160252) );
or I_9322 (I160845,I160780,I160591);
DFFARX1 I_9323  ( .D(I160845), .CLK(I2350), .RSTB(I160260), .Q(I160237) );
nand I_9324 (I160240,I160780,I160670);
not I_9325 (I160923,I2357);
not I_9326 (I160940,I36264);
nor I_9327 (I160957,I36261,I36285);
nand I_9328 (I160974,I160957,I36282);
nor I_9329 (I160991,I160940,I36261);
nand I_9330 (I161008,I160991,I36288);
not I_9331 (I161025,I161008);
not I_9332 (I161042,I36261);
nor I_9333 (I160912,I161008,I161042);
not I_9334 (I161073,I161042);
nand I_9335 (I160897,I161008,I161073);
not I_9336 (I161104,I36279);
nor I_9337 (I161121,I161104,I36270);
and I_9338 (I161138,I161121,I36267);
or I_9339 (I161155,I161138,I36276);
DFFARX1 I_9340  ( .D(I161155), .CLK(I2350), .RSTB(I160923), .Q(I161172) );
nor I_9341 (I161189,I161172,I161025);
DFFARX1 I_9342  ( .D(I161172), .CLK(I2350), .RSTB(I160923), .Q(I161206) );
not I_9343 (I160894,I161206);
nand I_9344 (I161237,I160940,I36279);
and I_9345 (I161254,I161237,I161189);
DFFARX1 I_9346  ( .D(I161237), .CLK(I2350), .RSTB(I160923), .Q(I160891) );
DFFARX1 I_9347  ( .D(I36258), .CLK(I2350), .RSTB(I160923), .Q(I161285) );
nor I_9348 (I161302,I161285,I161008);
nand I_9349 (I160909,I161172,I161302);
nor I_9350 (I161333,I161285,I161073);
not I_9351 (I160906,I161285);
nand I_9352 (I161364,I161285,I160974);
and I_9353 (I161381,I161042,I161364);
DFFARX1 I_9354  ( .D(I161381), .CLK(I2350), .RSTB(I160923), .Q(I160885) );
DFFARX1 I_9355  ( .D(I161285), .CLK(I2350), .RSTB(I160923), .Q(I160888) );
DFFARX1 I_9356  ( .D(I36273), .CLK(I2350), .RSTB(I160923), .Q(I161426) );
not I_9357 (I161443,I161426);
nand I_9358 (I161460,I161443,I161008);
and I_9359 (I161477,I161237,I161460);
DFFARX1 I_9360  ( .D(I161477), .CLK(I2350), .RSTB(I160923), .Q(I160915) );
or I_9361 (I161508,I161443,I161254);
DFFARX1 I_9362  ( .D(I161508), .CLK(I2350), .RSTB(I160923), .Q(I160900) );
nand I_9363 (I160903,I161443,I161333);
not I_9364 (I161586,I2357);
not I_9365 (I161603,I67918);
nor I_9366 (I161620,I67915,I67939);
nand I_9367 (I161637,I161620,I67936);
nor I_9368 (I161654,I161603,I67915);
nand I_9369 (I161671,I161654,I67942);
not I_9370 (I161688,I161671);
not I_9371 (I161705,I67915);
nor I_9372 (I161575,I161671,I161705);
not I_9373 (I161736,I161705);
nand I_9374 (I161560,I161671,I161736);
not I_9375 (I161767,I67933);
nor I_9376 (I161784,I161767,I67924);
and I_9377 (I161801,I161784,I67921);
or I_9378 (I161818,I161801,I67930);
DFFARX1 I_9379  ( .D(I161818), .CLK(I2350), .RSTB(I161586), .Q(I161835) );
nor I_9380 (I161852,I161835,I161688);
DFFARX1 I_9381  ( .D(I161835), .CLK(I2350), .RSTB(I161586), .Q(I161869) );
not I_9382 (I161557,I161869);
nand I_9383 (I161900,I161603,I67933);
and I_9384 (I161917,I161900,I161852);
DFFARX1 I_9385  ( .D(I161900), .CLK(I2350), .RSTB(I161586), .Q(I161554) );
DFFARX1 I_9386  ( .D(I67912), .CLK(I2350), .RSTB(I161586), .Q(I161948) );
nor I_9387 (I161965,I161948,I161671);
nand I_9388 (I161572,I161835,I161965);
nor I_9389 (I161996,I161948,I161736);
not I_9390 (I161569,I161948);
nand I_9391 (I162027,I161948,I161637);
and I_9392 (I162044,I161705,I162027);
DFFARX1 I_9393  ( .D(I162044), .CLK(I2350), .RSTB(I161586), .Q(I161548) );
DFFARX1 I_9394  ( .D(I161948), .CLK(I2350), .RSTB(I161586), .Q(I161551) );
DFFARX1 I_9395  ( .D(I67927), .CLK(I2350), .RSTB(I161586), .Q(I162089) );
not I_9396 (I162106,I162089);
nand I_9397 (I162123,I162106,I161671);
and I_9398 (I162140,I161900,I162123);
DFFARX1 I_9399  ( .D(I162140), .CLK(I2350), .RSTB(I161586), .Q(I161578) );
or I_9400 (I162171,I162106,I161917);
DFFARX1 I_9401  ( .D(I162171), .CLK(I2350), .RSTB(I161586), .Q(I161563) );
nand I_9402 (I161566,I162106,I161996);
not I_9403 (I162249,I2357);
not I_9404 (I162266,I392607);
nor I_9405 (I162283,I392598,I392604);
nand I_9406 (I162300,I162283,I392616);
nor I_9407 (I162317,I162266,I392598);
nand I_9408 (I162334,I162317,I392601);
not I_9409 (I162351,I162334);
not I_9410 (I162368,I392598);
nor I_9411 (I162238,I162334,I162368);
not I_9412 (I162399,I162368);
nand I_9413 (I162223,I162334,I162399);
not I_9414 (I162430,I392625);
nor I_9415 (I162447,I162430,I392619);
and I_9416 (I162464,I162447,I392610);
or I_9417 (I162481,I162464,I392595);
DFFARX1 I_9418  ( .D(I162481), .CLK(I2350), .RSTB(I162249), .Q(I162498) );
nor I_9419 (I162515,I162498,I162351);
DFFARX1 I_9420  ( .D(I162498), .CLK(I2350), .RSTB(I162249), .Q(I162532) );
not I_9421 (I162220,I162532);
nand I_9422 (I162563,I162266,I392625);
and I_9423 (I162580,I162563,I162515);
DFFARX1 I_9424  ( .D(I162563), .CLK(I2350), .RSTB(I162249), .Q(I162217) );
DFFARX1 I_9425  ( .D(I392613), .CLK(I2350), .RSTB(I162249), .Q(I162611) );
nor I_9426 (I162628,I162611,I162334);
nand I_9427 (I162235,I162498,I162628);
nor I_9428 (I162659,I162611,I162399);
not I_9429 (I162232,I162611);
nand I_9430 (I162690,I162611,I162300);
and I_9431 (I162707,I162368,I162690);
DFFARX1 I_9432  ( .D(I162707), .CLK(I2350), .RSTB(I162249), .Q(I162211) );
DFFARX1 I_9433  ( .D(I162611), .CLK(I2350), .RSTB(I162249), .Q(I162214) );
DFFARX1 I_9434  ( .D(I392622), .CLK(I2350), .RSTB(I162249), .Q(I162752) );
not I_9435 (I162769,I162752);
nand I_9436 (I162786,I162769,I162334);
and I_9437 (I162803,I162563,I162786);
DFFARX1 I_9438  ( .D(I162803), .CLK(I2350), .RSTB(I162249), .Q(I162241) );
or I_9439 (I162834,I162769,I162580);
DFFARX1 I_9440  ( .D(I162834), .CLK(I2350), .RSTB(I162249), .Q(I162226) );
nand I_9441 (I162229,I162769,I162659);
not I_9442 (I162912,I2357);
not I_9443 (I162929,I102612);
nor I_9444 (I162946,I102618,I102624);
nand I_9445 (I162963,I162946,I102627);
nor I_9446 (I162980,I162929,I102618);
nand I_9447 (I162997,I162980,I102609);
not I_9448 (I163014,I162997);
not I_9449 (I163031,I102618);
nor I_9450 (I162901,I162997,I163031);
not I_9451 (I163062,I163031);
nand I_9452 (I162886,I162997,I163062);
not I_9453 (I163093,I102621);
nor I_9454 (I163110,I163093,I102615);
and I_9455 (I163127,I163110,I102630);
or I_9456 (I163144,I163127,I102636);
DFFARX1 I_9457  ( .D(I163144), .CLK(I2350), .RSTB(I162912), .Q(I163161) );
nor I_9458 (I163178,I163161,I163014);
DFFARX1 I_9459  ( .D(I163161), .CLK(I2350), .RSTB(I162912), .Q(I163195) );
not I_9460 (I162883,I163195);
nand I_9461 (I163226,I162929,I102621);
and I_9462 (I163243,I163226,I163178);
DFFARX1 I_9463  ( .D(I163226), .CLK(I2350), .RSTB(I162912), .Q(I162880) );
DFFARX1 I_9464  ( .D(I102633), .CLK(I2350), .RSTB(I162912), .Q(I163274) );
nor I_9465 (I163291,I163274,I162997);
nand I_9466 (I162898,I163161,I163291);
nor I_9467 (I163322,I163274,I163062);
not I_9468 (I162895,I163274);
nand I_9469 (I163353,I163274,I162963);
and I_9470 (I163370,I163031,I163353);
DFFARX1 I_9471  ( .D(I163370), .CLK(I2350), .RSTB(I162912), .Q(I162874) );
DFFARX1 I_9472  ( .D(I163274), .CLK(I2350), .RSTB(I162912), .Q(I162877) );
DFFARX1 I_9473  ( .D(I102639), .CLK(I2350), .RSTB(I162912), .Q(I163415) );
not I_9474 (I163432,I163415);
nand I_9475 (I163449,I163432,I162997);
and I_9476 (I163466,I163226,I163449);
DFFARX1 I_9477  ( .D(I163466), .CLK(I2350), .RSTB(I162912), .Q(I162904) );
or I_9478 (I163497,I163432,I163243);
DFFARX1 I_9479  ( .D(I163497), .CLK(I2350), .RSTB(I162912), .Q(I162889) );
nand I_9480 (I162892,I163432,I163322);
not I_9481 (I163575,I2357);
not I_9482 (I163592,I131162);
nor I_9483 (I163609,I131135,I131138);
nand I_9484 (I163626,I163609,I131150);
nor I_9485 (I163643,I163592,I131135);
nand I_9486 (I163660,I163643,I131156);
not I_9487 (I163677,I163660);
not I_9488 (I163694,I131135);
nor I_9489 (I163564,I163660,I163694);
not I_9490 (I163725,I163694);
nand I_9491 (I163549,I163660,I163725);
not I_9492 (I163756,I131159);
nor I_9493 (I163773,I163756,I131141);
and I_9494 (I163790,I163773,I131144);
or I_9495 (I163807,I163790,I131165);
DFFARX1 I_9496  ( .D(I163807), .CLK(I2350), .RSTB(I163575), .Q(I163824) );
nor I_9497 (I163841,I163824,I163677);
DFFARX1 I_9498  ( .D(I163824), .CLK(I2350), .RSTB(I163575), .Q(I163858) );
not I_9499 (I163546,I163858);
nand I_9500 (I163889,I163592,I131159);
and I_9501 (I163906,I163889,I163841);
DFFARX1 I_9502  ( .D(I163889), .CLK(I2350), .RSTB(I163575), .Q(I163543) );
DFFARX1 I_9503  ( .D(I131147), .CLK(I2350), .RSTB(I163575), .Q(I163937) );
nor I_9504 (I163954,I163937,I163660);
nand I_9505 (I163561,I163824,I163954);
nor I_9506 (I163985,I163937,I163725);
not I_9507 (I163558,I163937);
nand I_9508 (I164016,I163937,I163626);
and I_9509 (I164033,I163694,I164016);
DFFARX1 I_9510  ( .D(I164033), .CLK(I2350), .RSTB(I163575), .Q(I163537) );
DFFARX1 I_9511  ( .D(I163937), .CLK(I2350), .RSTB(I163575), .Q(I163540) );
DFFARX1 I_9512  ( .D(I131153), .CLK(I2350), .RSTB(I163575), .Q(I164078) );
not I_9513 (I164095,I164078);
nand I_9514 (I164112,I164095,I163660);
and I_9515 (I164129,I163889,I164112);
DFFARX1 I_9516  ( .D(I164129), .CLK(I2350), .RSTB(I163575), .Q(I163567) );
or I_9517 (I164160,I164095,I163906);
DFFARX1 I_9518  ( .D(I164160), .CLK(I2350), .RSTB(I163575), .Q(I163552) );
nand I_9519 (I163555,I164095,I163985);
not I_9520 (I164238,I2357);
not I_9521 (I164255,I116873);
nor I_9522 (I164272,I116867,I116858);
nand I_9523 (I164289,I164272,I116870);
nor I_9524 (I164306,I164255,I116867);
nand I_9525 (I164323,I164306,I116885);
not I_9526 (I164340,I164323);
not I_9527 (I164357,I116867);
nor I_9528 (I164227,I164323,I164357);
not I_9529 (I164388,I164357);
nand I_9530 (I164212,I164323,I164388);
not I_9531 (I164419,I116861);
nor I_9532 (I164436,I164419,I116855);
and I_9533 (I164453,I164436,I116882);
or I_9534 (I164470,I164453,I116879);
DFFARX1 I_9535  ( .D(I164470), .CLK(I2350), .RSTB(I164238), .Q(I164487) );
nor I_9536 (I164504,I164487,I164340);
DFFARX1 I_9537  ( .D(I164487), .CLK(I2350), .RSTB(I164238), .Q(I164521) );
not I_9538 (I164209,I164521);
nand I_9539 (I164552,I164255,I116861);
and I_9540 (I164569,I164552,I164504);
DFFARX1 I_9541  ( .D(I164552), .CLK(I2350), .RSTB(I164238), .Q(I164206) );
DFFARX1 I_9542  ( .D(I116876), .CLK(I2350), .RSTB(I164238), .Q(I164600) );
nor I_9543 (I164617,I164600,I164323);
nand I_9544 (I164224,I164487,I164617);
nor I_9545 (I164648,I164600,I164388);
not I_9546 (I164221,I164600);
nand I_9547 (I164679,I164600,I164289);
and I_9548 (I164696,I164357,I164679);
DFFARX1 I_9549  ( .D(I164696), .CLK(I2350), .RSTB(I164238), .Q(I164200) );
DFFARX1 I_9550  ( .D(I164600), .CLK(I2350), .RSTB(I164238), .Q(I164203) );
DFFARX1 I_9551  ( .D(I116864), .CLK(I2350), .RSTB(I164238), .Q(I164741) );
not I_9552 (I164758,I164741);
nand I_9553 (I164775,I164758,I164323);
and I_9554 (I164792,I164552,I164775);
DFFARX1 I_9555  ( .D(I164792), .CLK(I2350), .RSTB(I164238), .Q(I164230) );
or I_9556 (I164823,I164758,I164569);
DFFARX1 I_9557  ( .D(I164823), .CLK(I2350), .RSTB(I164238), .Q(I164215) );
nand I_9558 (I164218,I164758,I164648);
not I_9559 (I164901,I2357);
not I_9560 (I164918,I320125);
nor I_9561 (I164935,I320122,I320113);
nand I_9562 (I164952,I164935,I320116);
nor I_9563 (I164969,I164918,I320122);
nand I_9564 (I164986,I164969,I320110);
not I_9565 (I165003,I164986);
not I_9566 (I165020,I320122);
nor I_9567 (I164890,I164986,I165020);
not I_9568 (I165051,I165020);
nand I_9569 (I164875,I164986,I165051);
not I_9570 (I165082,I320131);
nor I_9571 (I165099,I165082,I320134);
and I_9572 (I165116,I165099,I320119);
or I_9573 (I165133,I165116,I320107);
DFFARX1 I_9574  ( .D(I165133), .CLK(I2350), .RSTB(I164901), .Q(I165150) );
nor I_9575 (I165167,I165150,I165003);
DFFARX1 I_9576  ( .D(I165150), .CLK(I2350), .RSTB(I164901), .Q(I165184) );
not I_9577 (I164872,I165184);
nand I_9578 (I165215,I164918,I320131);
and I_9579 (I165232,I165215,I165167);
DFFARX1 I_9580  ( .D(I165215), .CLK(I2350), .RSTB(I164901), .Q(I164869) );
DFFARX1 I_9581  ( .D(I320128), .CLK(I2350), .RSTB(I164901), .Q(I165263) );
nor I_9582 (I165280,I165263,I164986);
nand I_9583 (I164887,I165150,I165280);
nor I_9584 (I165311,I165263,I165051);
not I_9585 (I164884,I165263);
nand I_9586 (I165342,I165263,I164952);
and I_9587 (I165359,I165020,I165342);
DFFARX1 I_9588  ( .D(I165359), .CLK(I2350), .RSTB(I164901), .Q(I164863) );
DFFARX1 I_9589  ( .D(I165263), .CLK(I2350), .RSTB(I164901), .Q(I164866) );
DFFARX1 I_9590  ( .D(I320137), .CLK(I2350), .RSTB(I164901), .Q(I165404) );
not I_9591 (I165421,I165404);
nand I_9592 (I165438,I165421,I164986);
and I_9593 (I165455,I165215,I165438);
DFFARX1 I_9594  ( .D(I165455), .CLK(I2350), .RSTB(I164901), .Q(I164893) );
or I_9595 (I165486,I165421,I165232);
DFFARX1 I_9596  ( .D(I165486), .CLK(I2350), .RSTB(I164901), .Q(I164878) );
nand I_9597 (I164881,I165421,I165311);
not I_9598 (I165564,I2357);
not I_9599 (I165581,I371606);
nor I_9600 (I165598,I371624,I371615);
nand I_9601 (I165615,I165598,I371621);
nor I_9602 (I165632,I165581,I371624);
nand I_9603 (I165649,I165632,I371627);
not I_9604 (I165666,I165649);
not I_9605 (I165683,I371624);
nor I_9606 (I165553,I165649,I165683);
not I_9607 (I165714,I165683);
nand I_9608 (I165538,I165649,I165714);
not I_9609 (I165745,I371603);
nor I_9610 (I165762,I165745,I371618);
and I_9611 (I165779,I165762,I371600);
or I_9612 (I165796,I165779,I371609);
DFFARX1 I_9613  ( .D(I165796), .CLK(I2350), .RSTB(I165564), .Q(I165813) );
nor I_9614 (I165830,I165813,I165666);
DFFARX1 I_9615  ( .D(I165813), .CLK(I2350), .RSTB(I165564), .Q(I165847) );
not I_9616 (I165535,I165847);
nand I_9617 (I165878,I165581,I371603);
and I_9618 (I165895,I165878,I165830);
DFFARX1 I_9619  ( .D(I165878), .CLK(I2350), .RSTB(I165564), .Q(I165532) );
DFFARX1 I_9620  ( .D(I371612), .CLK(I2350), .RSTB(I165564), .Q(I165926) );
nor I_9621 (I165943,I165926,I165649);
nand I_9622 (I165550,I165813,I165943);
nor I_9623 (I165974,I165926,I165714);
not I_9624 (I165547,I165926);
nand I_9625 (I166005,I165926,I165615);
and I_9626 (I166022,I165683,I166005);
DFFARX1 I_9627  ( .D(I166022), .CLK(I2350), .RSTB(I165564), .Q(I165526) );
DFFARX1 I_9628  ( .D(I165926), .CLK(I2350), .RSTB(I165564), .Q(I165529) );
DFFARX1 I_9629  ( .D(I371630), .CLK(I2350), .RSTB(I165564), .Q(I166067) );
not I_9630 (I166084,I166067);
nand I_9631 (I166101,I166084,I165649);
and I_9632 (I166118,I165878,I166101);
DFFARX1 I_9633  ( .D(I166118), .CLK(I2350), .RSTB(I165564), .Q(I165556) );
or I_9634 (I166149,I166084,I165895);
DFFARX1 I_9635  ( .D(I166149), .CLK(I2350), .RSTB(I165564), .Q(I165541) );
nand I_9636 (I165544,I166084,I165974);
not I_9637 (I166227,I2357);
not I_9638 (I166244,I366574);
nor I_9639 (I166261,I366592,I366583);
nand I_9640 (I166278,I166261,I366589);
nor I_9641 (I166295,I166244,I366592);
nand I_9642 (I166312,I166295,I366595);
not I_9643 (I166329,I166312);
not I_9644 (I166346,I366592);
nor I_9645 (I166216,I166312,I166346);
not I_9646 (I166377,I166346);
nand I_9647 (I166201,I166312,I166377);
not I_9648 (I166408,I366571);
nor I_9649 (I166425,I166408,I366586);
and I_9650 (I166442,I166425,I366568);
or I_9651 (I166459,I166442,I366577);
DFFARX1 I_9652  ( .D(I166459), .CLK(I2350), .RSTB(I166227), .Q(I166476) );
nor I_9653 (I166493,I166476,I166329);
DFFARX1 I_9654  ( .D(I166476), .CLK(I2350), .RSTB(I166227), .Q(I166510) );
not I_9655 (I166198,I166510);
nand I_9656 (I166541,I166244,I366571);
and I_9657 (I166558,I166541,I166493);
DFFARX1 I_9658  ( .D(I166541), .CLK(I2350), .RSTB(I166227), .Q(I166195) );
DFFARX1 I_9659  ( .D(I366580), .CLK(I2350), .RSTB(I166227), .Q(I166589) );
nor I_9660 (I166606,I166589,I166312);
nand I_9661 (I166213,I166476,I166606);
nor I_9662 (I166637,I166589,I166377);
not I_9663 (I166210,I166589);
nand I_9664 (I166668,I166589,I166278);
and I_9665 (I166685,I166346,I166668);
DFFARX1 I_9666  ( .D(I166685), .CLK(I2350), .RSTB(I166227), .Q(I166189) );
DFFARX1 I_9667  ( .D(I166589), .CLK(I2350), .RSTB(I166227), .Q(I166192) );
DFFARX1 I_9668  ( .D(I366598), .CLK(I2350), .RSTB(I166227), .Q(I166730) );
not I_9669 (I166747,I166730);
nand I_9670 (I166764,I166747,I166312);
and I_9671 (I166781,I166541,I166764);
DFFARX1 I_9672  ( .D(I166781), .CLK(I2350), .RSTB(I166227), .Q(I166219) );
or I_9673 (I166812,I166747,I166558);
DFFARX1 I_9674  ( .D(I166812), .CLK(I2350), .RSTB(I166227), .Q(I166204) );
nand I_9675 (I166207,I166747,I166637);
not I_9676 (I166890,I2357);
not I_9677 (I166907,I42724);
nor I_9678 (I166924,I42721,I42745);
nand I_9679 (I166941,I166924,I42742);
nor I_9680 (I166958,I166907,I42721);
nand I_9681 (I166975,I166958,I42748);
not I_9682 (I166992,I166975);
not I_9683 (I167009,I42721);
nor I_9684 (I166879,I166975,I167009);
not I_9685 (I167040,I167009);
nand I_9686 (I166864,I166975,I167040);
not I_9687 (I167071,I42739);
nor I_9688 (I167088,I167071,I42730);
and I_9689 (I167105,I167088,I42727);
or I_9690 (I167122,I167105,I42736);
DFFARX1 I_9691  ( .D(I167122), .CLK(I2350), .RSTB(I166890), .Q(I167139) );
nor I_9692 (I167156,I167139,I166992);
DFFARX1 I_9693  ( .D(I167139), .CLK(I2350), .RSTB(I166890), .Q(I167173) );
not I_9694 (I166861,I167173);
nand I_9695 (I167204,I166907,I42739);
and I_9696 (I167221,I167204,I167156);
DFFARX1 I_9697  ( .D(I167204), .CLK(I2350), .RSTB(I166890), .Q(I166858) );
DFFARX1 I_9698  ( .D(I42718), .CLK(I2350), .RSTB(I166890), .Q(I167252) );
nor I_9699 (I167269,I167252,I166975);
nand I_9700 (I166876,I167139,I167269);
nor I_9701 (I167300,I167252,I167040);
not I_9702 (I166873,I167252);
nand I_9703 (I167331,I167252,I166941);
and I_9704 (I167348,I167009,I167331);
DFFARX1 I_9705  ( .D(I167348), .CLK(I2350), .RSTB(I166890), .Q(I166852) );
DFFARX1 I_9706  ( .D(I167252), .CLK(I2350), .RSTB(I166890), .Q(I166855) );
DFFARX1 I_9707  ( .D(I42733), .CLK(I2350), .RSTB(I166890), .Q(I167393) );
not I_9708 (I167410,I167393);
nand I_9709 (I167427,I167410,I166975);
and I_9710 (I167444,I167204,I167427);
DFFARX1 I_9711  ( .D(I167444), .CLK(I2350), .RSTB(I166890), .Q(I166882) );
or I_9712 (I167475,I167410,I167221);
DFFARX1 I_9713  ( .D(I167475), .CLK(I2350), .RSTB(I166890), .Q(I166867) );
nand I_9714 (I166870,I167410,I167300);
not I_9715 (I167553,I2357);
not I_9716 (I167570,I210809);
nor I_9717 (I167587,I210806,I210824);
nand I_9718 (I167604,I167587,I210827);
nor I_9719 (I167621,I167570,I210806);
nand I_9720 (I167638,I167621,I210812);
not I_9721 (I167655,I167638);
not I_9722 (I167672,I210806);
nor I_9723 (I167542,I167638,I167672);
not I_9724 (I167703,I167672);
nand I_9725 (I167527,I167638,I167703);
not I_9726 (I167734,I210821);
nor I_9727 (I167751,I167734,I210803);
and I_9728 (I167768,I167751,I210797);
or I_9729 (I167785,I167768,I210815);
DFFARX1 I_9730  ( .D(I167785), .CLK(I2350), .RSTB(I167553), .Q(I167802) );
nor I_9731 (I167819,I167802,I167655);
DFFARX1 I_9732  ( .D(I167802), .CLK(I2350), .RSTB(I167553), .Q(I167836) );
not I_9733 (I167524,I167836);
nand I_9734 (I167867,I167570,I210821);
and I_9735 (I167884,I167867,I167819);
DFFARX1 I_9736  ( .D(I167867), .CLK(I2350), .RSTB(I167553), .Q(I167521) );
DFFARX1 I_9737  ( .D(I210800), .CLK(I2350), .RSTB(I167553), .Q(I167915) );
nor I_9738 (I167932,I167915,I167638);
nand I_9739 (I167539,I167802,I167932);
nor I_9740 (I167963,I167915,I167703);
not I_9741 (I167536,I167915);
nand I_9742 (I167994,I167915,I167604);
and I_9743 (I168011,I167672,I167994);
DFFARX1 I_9744  ( .D(I168011), .CLK(I2350), .RSTB(I167553), .Q(I167515) );
DFFARX1 I_9745  ( .D(I167915), .CLK(I2350), .RSTB(I167553), .Q(I167518) );
DFFARX1 I_9746  ( .D(I210818), .CLK(I2350), .RSTB(I167553), .Q(I168056) );
not I_9747 (I168073,I168056);
nand I_9748 (I168090,I168073,I167638);
and I_9749 (I168107,I167867,I168090);
DFFARX1 I_9750  ( .D(I168107), .CLK(I2350), .RSTB(I167553), .Q(I167545) );
or I_9751 (I168138,I168073,I167884);
DFFARX1 I_9752  ( .D(I168138), .CLK(I2350), .RSTB(I167553), .Q(I167530) );
nand I_9753 (I167533,I168073,I167963);
not I_9754 (I168216,I2357);
not I_9755 (I168233,I111231);
nor I_9756 (I168250,I111237,I111243);
nand I_9757 (I168267,I168250,I111246);
nor I_9758 (I168284,I168233,I111237);
nand I_9759 (I168301,I168284,I111228);
not I_9760 (I168318,I168301);
not I_9761 (I168335,I111237);
nor I_9762 (I168205,I168301,I168335);
not I_9763 (I168366,I168335);
nand I_9764 (I168190,I168301,I168366);
not I_9765 (I168397,I111240);
nor I_9766 (I168414,I168397,I111234);
and I_9767 (I168431,I168414,I111249);
or I_9768 (I168448,I168431,I111255);
DFFARX1 I_9769  ( .D(I168448), .CLK(I2350), .RSTB(I168216), .Q(I168465) );
nor I_9770 (I168482,I168465,I168318);
DFFARX1 I_9771  ( .D(I168465), .CLK(I2350), .RSTB(I168216), .Q(I168499) );
not I_9772 (I168187,I168499);
nand I_9773 (I168530,I168233,I111240);
and I_9774 (I168547,I168530,I168482);
DFFARX1 I_9775  ( .D(I168530), .CLK(I2350), .RSTB(I168216), .Q(I168184) );
DFFARX1 I_9776  ( .D(I111252), .CLK(I2350), .RSTB(I168216), .Q(I168578) );
nor I_9777 (I168595,I168578,I168301);
nand I_9778 (I168202,I168465,I168595);
nor I_9779 (I168626,I168578,I168366);
not I_9780 (I168199,I168578);
nand I_9781 (I168657,I168578,I168267);
and I_9782 (I168674,I168335,I168657);
DFFARX1 I_9783  ( .D(I168674), .CLK(I2350), .RSTB(I168216), .Q(I168178) );
DFFARX1 I_9784  ( .D(I168578), .CLK(I2350), .RSTB(I168216), .Q(I168181) );
DFFARX1 I_9785  ( .D(I111258), .CLK(I2350), .RSTB(I168216), .Q(I168719) );
not I_9786 (I168736,I168719);
nand I_9787 (I168753,I168736,I168301);
and I_9788 (I168770,I168530,I168753);
DFFARX1 I_9789  ( .D(I168770), .CLK(I2350), .RSTB(I168216), .Q(I168208) );
or I_9790 (I168801,I168736,I168547);
DFFARX1 I_9791  ( .D(I168801), .CLK(I2350), .RSTB(I168216), .Q(I168193) );
nand I_9792 (I168196,I168736,I168626);
not I_9793 (I168879,I2357);
not I_9794 (I168896,I290375);
nor I_9795 (I168913,I290384,I290366);
nand I_9796 (I168930,I168913,I290387);
nor I_9797 (I168947,I168896,I290384);
nand I_9798 (I168964,I168947,I290378);
not I_9799 (I168981,I168964);
not I_9800 (I168998,I290384);
nor I_9801 (I168868,I168964,I168998);
not I_9802 (I169029,I168998);
nand I_9803 (I168853,I168964,I169029);
not I_9804 (I169060,I290372);
nor I_9805 (I169077,I169060,I290363);
and I_9806 (I169094,I169077,I290360);
or I_9807 (I169111,I169094,I290357);
DFFARX1 I_9808  ( .D(I169111), .CLK(I2350), .RSTB(I168879), .Q(I169128) );
nor I_9809 (I169145,I169128,I168981);
DFFARX1 I_9810  ( .D(I169128), .CLK(I2350), .RSTB(I168879), .Q(I169162) );
not I_9811 (I168850,I169162);
nand I_9812 (I169193,I168896,I290372);
and I_9813 (I169210,I169193,I169145);
DFFARX1 I_9814  ( .D(I169193), .CLK(I2350), .RSTB(I168879), .Q(I168847) );
DFFARX1 I_9815  ( .D(I290381), .CLK(I2350), .RSTB(I168879), .Q(I169241) );
nor I_9816 (I169258,I169241,I168964);
nand I_9817 (I168865,I169128,I169258);
nor I_9818 (I169289,I169241,I169029);
not I_9819 (I168862,I169241);
nand I_9820 (I169320,I169241,I168930);
and I_9821 (I169337,I168998,I169320);
DFFARX1 I_9822  ( .D(I169337), .CLK(I2350), .RSTB(I168879), .Q(I168841) );
DFFARX1 I_9823  ( .D(I169241), .CLK(I2350), .RSTB(I168879), .Q(I168844) );
DFFARX1 I_9824  ( .D(I290369), .CLK(I2350), .RSTB(I168879), .Q(I169382) );
not I_9825 (I169399,I169382);
nand I_9826 (I169416,I169399,I168964);
and I_9827 (I169433,I169193,I169416);
DFFARX1 I_9828  ( .D(I169433), .CLK(I2350), .RSTB(I168879), .Q(I168871) );
or I_9829 (I169464,I169399,I169210);
DFFARX1 I_9830  ( .D(I169464), .CLK(I2350), .RSTB(I168879), .Q(I168856) );
nand I_9831 (I168859,I169399,I169289);
not I_9832 (I169542,I2357);
not I_9833 (I169559,I317745);
nor I_9834 (I169576,I317742,I317733);
nand I_9835 (I169593,I169576,I317736);
nor I_9836 (I169610,I169559,I317742);
nand I_9837 (I169627,I169610,I317730);
not I_9838 (I169644,I169627);
not I_9839 (I169661,I317742);
nor I_9840 (I169531,I169627,I169661);
not I_9841 (I169692,I169661);
nand I_9842 (I169516,I169627,I169692);
not I_9843 (I169723,I317751);
nor I_9844 (I169740,I169723,I317754);
and I_9845 (I169757,I169740,I317739);
or I_9846 (I169774,I169757,I317727);
DFFARX1 I_9847  ( .D(I169774), .CLK(I2350), .RSTB(I169542), .Q(I169791) );
nor I_9848 (I169808,I169791,I169644);
DFFARX1 I_9849  ( .D(I169791), .CLK(I2350), .RSTB(I169542), .Q(I169825) );
not I_9850 (I169513,I169825);
nand I_9851 (I169856,I169559,I317751);
and I_9852 (I169873,I169856,I169808);
DFFARX1 I_9853  ( .D(I169856), .CLK(I2350), .RSTB(I169542), .Q(I169510) );
DFFARX1 I_9854  ( .D(I317748), .CLK(I2350), .RSTB(I169542), .Q(I169904) );
nor I_9855 (I169921,I169904,I169627);
nand I_9856 (I169528,I169791,I169921);
nor I_9857 (I169952,I169904,I169692);
not I_9858 (I169525,I169904);
nand I_9859 (I169983,I169904,I169593);
and I_9860 (I170000,I169661,I169983);
DFFARX1 I_9861  ( .D(I170000), .CLK(I2350), .RSTB(I169542), .Q(I169504) );
DFFARX1 I_9862  ( .D(I169904), .CLK(I2350), .RSTB(I169542), .Q(I169507) );
DFFARX1 I_9863  ( .D(I317757), .CLK(I2350), .RSTB(I169542), .Q(I170045) );
not I_9864 (I170062,I170045);
nand I_9865 (I170079,I170062,I169627);
and I_9866 (I170096,I169856,I170079);
DFFARX1 I_9867  ( .D(I170096), .CLK(I2350), .RSTB(I169542), .Q(I169534) );
or I_9868 (I170127,I170062,I169873);
DFFARX1 I_9869  ( .D(I170127), .CLK(I2350), .RSTB(I169542), .Q(I169519) );
nand I_9870 (I169522,I170062,I169952);
not I_9871 (I170205,I2357);
not I_9872 (I170222,I57582);
nor I_9873 (I170239,I57579,I57603);
nand I_9874 (I170256,I170239,I57600);
nor I_9875 (I170273,I170222,I57579);
nand I_9876 (I170290,I170273,I57606);
not I_9877 (I170307,I170290);
not I_9878 (I170324,I57579);
nor I_9879 (I170194,I170290,I170324);
not I_9880 (I170355,I170324);
nand I_9881 (I170179,I170290,I170355);
not I_9882 (I170386,I57597);
nor I_9883 (I170403,I170386,I57588);
and I_9884 (I170420,I170403,I57585);
or I_9885 (I170437,I170420,I57594);
DFFARX1 I_9886  ( .D(I170437), .CLK(I2350), .RSTB(I170205), .Q(I170454) );
nor I_9887 (I170471,I170454,I170307);
DFFARX1 I_9888  ( .D(I170454), .CLK(I2350), .RSTB(I170205), .Q(I170488) );
not I_9889 (I170176,I170488);
nand I_9890 (I170519,I170222,I57597);
and I_9891 (I170536,I170519,I170471);
DFFARX1 I_9892  ( .D(I170519), .CLK(I2350), .RSTB(I170205), .Q(I170173) );
DFFARX1 I_9893  ( .D(I57576), .CLK(I2350), .RSTB(I170205), .Q(I170567) );
nor I_9894 (I170584,I170567,I170290);
nand I_9895 (I170191,I170454,I170584);
nor I_9896 (I170615,I170567,I170355);
not I_9897 (I170188,I170567);
nand I_9898 (I170646,I170567,I170256);
and I_9899 (I170663,I170324,I170646);
DFFARX1 I_9900  ( .D(I170663), .CLK(I2350), .RSTB(I170205), .Q(I170167) );
DFFARX1 I_9901  ( .D(I170567), .CLK(I2350), .RSTB(I170205), .Q(I170170) );
DFFARX1 I_9902  ( .D(I57591), .CLK(I2350), .RSTB(I170205), .Q(I170708) );
not I_9903 (I170725,I170708);
nand I_9904 (I170742,I170725,I170290);
and I_9905 (I170759,I170519,I170742);
DFFARX1 I_9906  ( .D(I170759), .CLK(I2350), .RSTB(I170205), .Q(I170197) );
or I_9907 (I170790,I170725,I170536);
DFFARX1 I_9908  ( .D(I170790), .CLK(I2350), .RSTB(I170205), .Q(I170182) );
nand I_9909 (I170185,I170725,I170615);
not I_9910 (I170868,I2357);
not I_9911 (I170885,I270927);
nor I_9912 (I170902,I270924,I270921);
nand I_9913 (I170919,I170902,I270909);
nor I_9914 (I170936,I170885,I270924);
nand I_9915 (I170953,I170936,I270930);
not I_9916 (I170970,I170953);
not I_9917 (I170987,I270924);
nor I_9918 (I170857,I170953,I170987);
not I_9919 (I171018,I170987);
nand I_9920 (I170842,I170953,I171018);
not I_9921 (I171049,I270912);
nor I_9922 (I171066,I171049,I270918);
and I_9923 (I171083,I171066,I270915);
or I_9924 (I171100,I171083,I270939);
DFFARX1 I_9925  ( .D(I171100), .CLK(I2350), .RSTB(I170868), .Q(I171117) );
nor I_9926 (I171134,I171117,I170970);
DFFARX1 I_9927  ( .D(I171117), .CLK(I2350), .RSTB(I170868), .Q(I171151) );
not I_9928 (I170839,I171151);
nand I_9929 (I171182,I170885,I270912);
and I_9930 (I171199,I171182,I171134);
DFFARX1 I_9931  ( .D(I171182), .CLK(I2350), .RSTB(I170868), .Q(I170836) );
DFFARX1 I_9932  ( .D(I270936), .CLK(I2350), .RSTB(I170868), .Q(I171230) );
nor I_9933 (I171247,I171230,I170953);
nand I_9934 (I170854,I171117,I171247);
nor I_9935 (I171278,I171230,I171018);
not I_9936 (I170851,I171230);
nand I_9937 (I171309,I171230,I170919);
and I_9938 (I171326,I170987,I171309);
DFFARX1 I_9939  ( .D(I171326), .CLK(I2350), .RSTB(I170868), .Q(I170830) );
DFFARX1 I_9940  ( .D(I171230), .CLK(I2350), .RSTB(I170868), .Q(I170833) );
DFFARX1 I_9941  ( .D(I270933), .CLK(I2350), .RSTB(I170868), .Q(I171371) );
not I_9942 (I171388,I171371);
nand I_9943 (I171405,I171388,I170953);
and I_9944 (I171422,I171182,I171405);
DFFARX1 I_9945  ( .D(I171422), .CLK(I2350), .RSTB(I170868), .Q(I170860) );
or I_9946 (I171453,I171388,I171199);
DFFARX1 I_9947  ( .D(I171453), .CLK(I2350), .RSTB(I170868), .Q(I170845) );
nand I_9948 (I170848,I171388,I171278);
not I_9949 (I171531,I2357);
not I_9950 (I171548,I208225);
nor I_9951 (I171565,I208222,I208240);
nand I_9952 (I171582,I171565,I208243);
nor I_9953 (I171599,I171548,I208222);
nand I_9954 (I171616,I171599,I208228);
not I_9955 (I171633,I171616);
not I_9956 (I171650,I208222);
nor I_9957 (I171520,I171616,I171650);
not I_9958 (I171681,I171650);
nand I_9959 (I171505,I171616,I171681);
not I_9960 (I171712,I208237);
nor I_9961 (I171729,I171712,I208219);
and I_9962 (I171746,I171729,I208213);
or I_9963 (I171763,I171746,I208231);
DFFARX1 I_9964  ( .D(I171763), .CLK(I2350), .RSTB(I171531), .Q(I171780) );
nor I_9965 (I171797,I171780,I171633);
DFFARX1 I_9966  ( .D(I171780), .CLK(I2350), .RSTB(I171531), .Q(I171814) );
not I_9967 (I171502,I171814);
nand I_9968 (I171845,I171548,I208237);
and I_9969 (I171862,I171845,I171797);
DFFARX1 I_9970  ( .D(I171845), .CLK(I2350), .RSTB(I171531), .Q(I171499) );
DFFARX1 I_9971  ( .D(I208216), .CLK(I2350), .RSTB(I171531), .Q(I171893) );
nor I_9972 (I171910,I171893,I171616);
nand I_9973 (I171517,I171780,I171910);
nor I_9974 (I171941,I171893,I171681);
not I_9975 (I171514,I171893);
nand I_9976 (I171972,I171893,I171582);
and I_9977 (I171989,I171650,I171972);
DFFARX1 I_9978  ( .D(I171989), .CLK(I2350), .RSTB(I171531), .Q(I171493) );
DFFARX1 I_9979  ( .D(I171893), .CLK(I2350), .RSTB(I171531), .Q(I171496) );
DFFARX1 I_9980  ( .D(I208234), .CLK(I2350), .RSTB(I171531), .Q(I172034) );
not I_9981 (I172051,I172034);
nand I_9982 (I172068,I172051,I171616);
and I_9983 (I172085,I171845,I172068);
DFFARX1 I_9984  ( .D(I172085), .CLK(I2350), .RSTB(I171531), .Q(I171523) );
or I_9985 (I172116,I172051,I171862);
DFFARX1 I_9986  ( .D(I172116), .CLK(I2350), .RSTB(I171531), .Q(I171508) );
nand I_9987 (I171511,I172051,I171941);
not I_9988 (I172194,I2357);
not I_9989 (I172211,I252190);
nor I_9990 (I172228,I252202,I252184);
nand I_9991 (I172245,I172228,I252205);
nor I_9992 (I172262,I172211,I252202);
nand I_9993 (I172279,I172262,I252196);
not I_9994 (I172296,I172279);
not I_9995 (I172313,I252202);
nor I_9996 (I172183,I172279,I172313);
not I_9997 (I172344,I172313);
nand I_9998 (I172168,I172279,I172344);
not I_9999 (I172375,I252187);
nor I_10000 (I172392,I172375,I252181);
and I_10001 (I172409,I172392,I252193);
or I_10002 (I172426,I172409,I252178);
DFFARX1 I_10003  ( .D(I172426), .CLK(I2350), .RSTB(I172194), .Q(I172443) );
nor I_10004 (I172460,I172443,I172296);
DFFARX1 I_10005  ( .D(I172443), .CLK(I2350), .RSTB(I172194), .Q(I172477) );
not I_10006 (I172165,I172477);
nand I_10007 (I172508,I172211,I252187);
and I_10008 (I172525,I172508,I172460);
DFFARX1 I_10009  ( .D(I172508), .CLK(I2350), .RSTB(I172194), .Q(I172162) );
DFFARX1 I_10010  ( .D(I252175), .CLK(I2350), .RSTB(I172194), .Q(I172556) );
nor I_10011 (I172573,I172556,I172279);
nand I_10012 (I172180,I172443,I172573);
nor I_10013 (I172604,I172556,I172344);
not I_10014 (I172177,I172556);
nand I_10015 (I172635,I172556,I172245);
and I_10016 (I172652,I172313,I172635);
DFFARX1 I_10017  ( .D(I172652), .CLK(I2350), .RSTB(I172194), .Q(I172156) );
DFFARX1 I_10018  ( .D(I172556), .CLK(I2350), .RSTB(I172194), .Q(I172159) );
DFFARX1 I_10019  ( .D(I252199), .CLK(I2350), .RSTB(I172194), .Q(I172697) );
not I_10020 (I172714,I172697);
nand I_10021 (I172731,I172714,I172279);
and I_10022 (I172748,I172508,I172731);
DFFARX1 I_10023  ( .D(I172748), .CLK(I2350), .RSTB(I172194), .Q(I172186) );
or I_10024 (I172779,I172714,I172525);
DFFARX1 I_10025  ( .D(I172779), .CLK(I2350), .RSTB(I172194), .Q(I172171) );
nand I_10026 (I172174,I172714,I172604);
not I_10027 (I172857,I2357);
not I_10028 (I172874,I119848);
nor I_10029 (I172891,I119842,I119833);
nand I_10030 (I172908,I172891,I119845);
nor I_10031 (I172925,I172874,I119842);
nand I_10032 (I172942,I172925,I119860);
not I_10033 (I172959,I172942);
not I_10034 (I172976,I119842);
nor I_10035 (I172846,I172942,I172976);
not I_10036 (I173007,I172976);
nand I_10037 (I172831,I172942,I173007);
not I_10038 (I173038,I119836);
nor I_10039 (I173055,I173038,I119830);
and I_10040 (I173072,I173055,I119857);
or I_10041 (I173089,I173072,I119854);
DFFARX1 I_10042  ( .D(I173089), .CLK(I2350), .RSTB(I172857), .Q(I173106) );
nor I_10043 (I173123,I173106,I172959);
DFFARX1 I_10044  ( .D(I173106), .CLK(I2350), .RSTB(I172857), .Q(I173140) );
not I_10045 (I172828,I173140);
nand I_10046 (I173171,I172874,I119836);
and I_10047 (I173188,I173171,I173123);
DFFARX1 I_10048  ( .D(I173171), .CLK(I2350), .RSTB(I172857), .Q(I172825) );
DFFARX1 I_10049  ( .D(I119851), .CLK(I2350), .RSTB(I172857), .Q(I173219) );
nor I_10050 (I173236,I173219,I172942);
nand I_10051 (I172843,I173106,I173236);
nor I_10052 (I173267,I173219,I173007);
not I_10053 (I172840,I173219);
nand I_10054 (I173298,I173219,I172908);
and I_10055 (I173315,I172976,I173298);
DFFARX1 I_10056  ( .D(I173315), .CLK(I2350), .RSTB(I172857), .Q(I172819) );
DFFARX1 I_10057  ( .D(I173219), .CLK(I2350), .RSTB(I172857), .Q(I172822) );
DFFARX1 I_10058  ( .D(I119839), .CLK(I2350), .RSTB(I172857), .Q(I173360) );
not I_10059 (I173377,I173360);
nand I_10060 (I173394,I173377,I172942);
and I_10061 (I173411,I173171,I173394);
DFFARX1 I_10062  ( .D(I173411), .CLK(I2350), .RSTB(I172857), .Q(I172849) );
or I_10063 (I173442,I173377,I173188);
DFFARX1 I_10064  ( .D(I173442), .CLK(I2350), .RSTB(I172857), .Q(I172834) );
nand I_10065 (I172837,I173377,I173267);
not I_10066 (I173520,I2357);
not I_10067 (I173537,I360913);
nor I_10068 (I173554,I360931,I360922);
nand I_10069 (I173571,I173554,I360928);
nor I_10070 (I173588,I173537,I360931);
nand I_10071 (I173605,I173588,I360934);
not I_10072 (I173622,I173605);
not I_10073 (I173639,I360931);
nor I_10074 (I173509,I173605,I173639);
not I_10075 (I173670,I173639);
nand I_10076 (I173494,I173605,I173670);
not I_10077 (I173701,I360910);
nor I_10078 (I173718,I173701,I360925);
and I_10079 (I173735,I173718,I360907);
or I_10080 (I173752,I173735,I360916);
DFFARX1 I_10081  ( .D(I173752), .CLK(I2350), .RSTB(I173520), .Q(I173769) );
nor I_10082 (I173786,I173769,I173622);
DFFARX1 I_10083  ( .D(I173769), .CLK(I2350), .RSTB(I173520), .Q(I173803) );
not I_10084 (I173491,I173803);
nand I_10085 (I173834,I173537,I360910);
and I_10086 (I173851,I173834,I173786);
DFFARX1 I_10087  ( .D(I173834), .CLK(I2350), .RSTB(I173520), .Q(I173488) );
DFFARX1 I_10088  ( .D(I360919), .CLK(I2350), .RSTB(I173520), .Q(I173882) );
nor I_10089 (I173899,I173882,I173605);
nand I_10090 (I173506,I173769,I173899);
nor I_10091 (I173930,I173882,I173670);
not I_10092 (I173503,I173882);
nand I_10093 (I173961,I173882,I173571);
and I_10094 (I173978,I173639,I173961);
DFFARX1 I_10095  ( .D(I173978), .CLK(I2350), .RSTB(I173520), .Q(I173482) );
DFFARX1 I_10096  ( .D(I173882), .CLK(I2350), .RSTB(I173520), .Q(I173485) );
DFFARX1 I_10097  ( .D(I360937), .CLK(I2350), .RSTB(I173520), .Q(I174023) );
not I_10098 (I174040,I174023);
nand I_10099 (I174057,I174040,I173605);
and I_10100 (I174074,I173834,I174057);
DFFARX1 I_10101  ( .D(I174074), .CLK(I2350), .RSTB(I173520), .Q(I173512) );
or I_10102 (I174105,I174040,I173851);
DFFARX1 I_10103  ( .D(I174105), .CLK(I2350), .RSTB(I173520), .Q(I173497) );
nand I_10104 (I173500,I174040,I173930);
not I_10105 (I174183,I2357);
not I_10106 (I174200,I229543);
nor I_10107 (I174217,I229540,I229558);
nand I_10108 (I174234,I174217,I229561);
nor I_10109 (I174251,I174200,I229540);
nand I_10110 (I174268,I174251,I229546);
not I_10111 (I174285,I174268);
not I_10112 (I174302,I229540);
nor I_10113 (I174172,I174268,I174302);
not I_10114 (I174333,I174302);
nand I_10115 (I174157,I174268,I174333);
not I_10116 (I174364,I229555);
nor I_10117 (I174381,I174364,I229537);
and I_10118 (I174398,I174381,I229531);
or I_10119 (I174415,I174398,I229549);
DFFARX1 I_10120  ( .D(I174415), .CLK(I2350), .RSTB(I174183), .Q(I174432) );
nor I_10121 (I174449,I174432,I174285);
DFFARX1 I_10122  ( .D(I174432), .CLK(I2350), .RSTB(I174183), .Q(I174466) );
not I_10123 (I174154,I174466);
nand I_10124 (I174497,I174200,I229555);
and I_10125 (I174514,I174497,I174449);
DFFARX1 I_10126  ( .D(I174497), .CLK(I2350), .RSTB(I174183), .Q(I174151) );
DFFARX1 I_10127  ( .D(I229534), .CLK(I2350), .RSTB(I174183), .Q(I174545) );
nor I_10128 (I174562,I174545,I174268);
nand I_10129 (I174169,I174432,I174562);
nor I_10130 (I174593,I174545,I174333);
not I_10131 (I174166,I174545);
nand I_10132 (I174624,I174545,I174234);
and I_10133 (I174641,I174302,I174624);
DFFARX1 I_10134  ( .D(I174641), .CLK(I2350), .RSTB(I174183), .Q(I174145) );
DFFARX1 I_10135  ( .D(I174545), .CLK(I2350), .RSTB(I174183), .Q(I174148) );
DFFARX1 I_10136  ( .D(I229552), .CLK(I2350), .RSTB(I174183), .Q(I174686) );
not I_10137 (I174703,I174686);
nand I_10138 (I174720,I174703,I174268);
and I_10139 (I174737,I174497,I174720);
DFFARX1 I_10140  ( .D(I174737), .CLK(I2350), .RSTB(I174183), .Q(I174175) );
or I_10141 (I174768,I174703,I174514);
DFFARX1 I_10142  ( .D(I174768), .CLK(I2350), .RSTB(I174183), .Q(I174160) );
nand I_10143 (I174163,I174703,I174593);
not I_10144 (I174846,I2357);
not I_10145 (I174863,I235215);
nor I_10146 (I174880,I235218,I235224);
nand I_10147 (I174897,I174880,I235230);
nor I_10148 (I174914,I174863,I235218);
nand I_10149 (I174931,I174914,I235209);
not I_10150 (I174948,I174931);
not I_10151 (I174965,I235218);
nor I_10152 (I174835,I174931,I174965);
not I_10153 (I174996,I174965);
nand I_10154 (I174820,I174931,I174996);
not I_10155 (I175027,I235221);
nor I_10156 (I175044,I175027,I235236);
and I_10157 (I175061,I175044,I235239);
or I_10158 (I175078,I175061,I235212);
DFFARX1 I_10159  ( .D(I175078), .CLK(I2350), .RSTB(I174846), .Q(I175095) );
nor I_10160 (I175112,I175095,I174948);
DFFARX1 I_10161  ( .D(I175095), .CLK(I2350), .RSTB(I174846), .Q(I175129) );
not I_10162 (I174817,I175129);
nand I_10163 (I175160,I174863,I235221);
and I_10164 (I175177,I175160,I175112);
DFFARX1 I_10165  ( .D(I175160), .CLK(I2350), .RSTB(I174846), .Q(I174814) );
DFFARX1 I_10166  ( .D(I235233), .CLK(I2350), .RSTB(I174846), .Q(I175208) );
nor I_10167 (I175225,I175208,I174931);
nand I_10168 (I174832,I175095,I175225);
nor I_10169 (I175256,I175208,I174996);
not I_10170 (I174829,I175208);
nand I_10171 (I175287,I175208,I174897);
and I_10172 (I175304,I174965,I175287);
DFFARX1 I_10173  ( .D(I175304), .CLK(I2350), .RSTB(I174846), .Q(I174808) );
DFFARX1 I_10174  ( .D(I175208), .CLK(I2350), .RSTB(I174846), .Q(I174811) );
DFFARX1 I_10175  ( .D(I235227), .CLK(I2350), .RSTB(I174846), .Q(I175349) );
not I_10176 (I175366,I175349);
nand I_10177 (I175383,I175366,I174931);
and I_10178 (I175400,I175160,I175383);
DFFARX1 I_10179  ( .D(I175400), .CLK(I2350), .RSTB(I174846), .Q(I174838) );
or I_10180 (I175431,I175366,I175177);
DFFARX1 I_10181  ( .D(I175431), .CLK(I2350), .RSTB(I174846), .Q(I174823) );
nand I_10182 (I174826,I175366,I175256);
not I_10183 (I175509,I2357);
not I_10184 (I175526,I372235);
nor I_10185 (I175543,I372253,I372244);
nand I_10186 (I175560,I175543,I372250);
nor I_10187 (I175577,I175526,I372253);
nand I_10188 (I175594,I175577,I372256);
not I_10189 (I175611,I175594);
not I_10190 (I175628,I372253);
nor I_10191 (I175498,I175594,I175628);
not I_10192 (I175659,I175628);
nand I_10193 (I175483,I175594,I175659);
not I_10194 (I175690,I372232);
nor I_10195 (I175707,I175690,I372247);
and I_10196 (I175724,I175707,I372229);
or I_10197 (I175741,I175724,I372238);
DFFARX1 I_10198  ( .D(I175741), .CLK(I2350), .RSTB(I175509), .Q(I175758) );
nor I_10199 (I175775,I175758,I175611);
DFFARX1 I_10200  ( .D(I175758), .CLK(I2350), .RSTB(I175509), .Q(I175792) );
not I_10201 (I175480,I175792);
nand I_10202 (I175823,I175526,I372232);
and I_10203 (I175840,I175823,I175775);
DFFARX1 I_10204  ( .D(I175823), .CLK(I2350), .RSTB(I175509), .Q(I175477) );
DFFARX1 I_10205  ( .D(I372241), .CLK(I2350), .RSTB(I175509), .Q(I175871) );
nor I_10206 (I175888,I175871,I175594);
nand I_10207 (I175495,I175758,I175888);
nor I_10208 (I175919,I175871,I175659);
not I_10209 (I175492,I175871);
nand I_10210 (I175950,I175871,I175560);
and I_10211 (I175967,I175628,I175950);
DFFARX1 I_10212  ( .D(I175967), .CLK(I2350), .RSTB(I175509), .Q(I175471) );
DFFARX1 I_10213  ( .D(I175871), .CLK(I2350), .RSTB(I175509), .Q(I175474) );
DFFARX1 I_10214  ( .D(I372259), .CLK(I2350), .RSTB(I175509), .Q(I176012) );
not I_10215 (I176029,I176012);
nand I_10216 (I176046,I176029,I175594);
and I_10217 (I176063,I175823,I176046);
DFFARX1 I_10218  ( .D(I176063), .CLK(I2350), .RSTB(I175509), .Q(I175501) );
or I_10219 (I176094,I176029,I175840);
DFFARX1 I_10220  ( .D(I176094), .CLK(I2350), .RSTB(I175509), .Q(I175486) );
nand I_10221 (I175489,I176029,I175919);
not I_10222 (I176172,I2357);
not I_10223 (I176189,I365945);
nor I_10224 (I176206,I365963,I365954);
nand I_10225 (I176223,I176206,I365960);
nor I_10226 (I176240,I176189,I365963);
nand I_10227 (I176257,I176240,I365966);
not I_10228 (I176274,I176257);
not I_10229 (I176291,I365963);
nor I_10230 (I176161,I176257,I176291);
not I_10231 (I176322,I176291);
nand I_10232 (I176146,I176257,I176322);
not I_10233 (I176353,I365942);
nor I_10234 (I176370,I176353,I365957);
and I_10235 (I176387,I176370,I365939);
or I_10236 (I176404,I176387,I365948);
DFFARX1 I_10237  ( .D(I176404), .CLK(I2350), .RSTB(I176172), .Q(I176421) );
nor I_10238 (I176438,I176421,I176274);
DFFARX1 I_10239  ( .D(I176421), .CLK(I2350), .RSTB(I176172), .Q(I176455) );
not I_10240 (I176143,I176455);
nand I_10241 (I176486,I176189,I365942);
and I_10242 (I176503,I176486,I176438);
DFFARX1 I_10243  ( .D(I176486), .CLK(I2350), .RSTB(I176172), .Q(I176140) );
DFFARX1 I_10244  ( .D(I365951), .CLK(I2350), .RSTB(I176172), .Q(I176534) );
nor I_10245 (I176551,I176534,I176257);
nand I_10246 (I176158,I176421,I176551);
nor I_10247 (I176582,I176534,I176322);
not I_10248 (I176155,I176534);
nand I_10249 (I176613,I176534,I176223);
and I_10250 (I176630,I176291,I176613);
DFFARX1 I_10251  ( .D(I176630), .CLK(I2350), .RSTB(I176172), .Q(I176134) );
DFFARX1 I_10252  ( .D(I176534), .CLK(I2350), .RSTB(I176172), .Q(I176137) );
DFFARX1 I_10253  ( .D(I365969), .CLK(I2350), .RSTB(I176172), .Q(I176675) );
not I_10254 (I176692,I176675);
nand I_10255 (I176709,I176692,I176257);
and I_10256 (I176726,I176486,I176709);
DFFARX1 I_10257  ( .D(I176726), .CLK(I2350), .RSTB(I176172), .Q(I176164) );
or I_10258 (I176757,I176692,I176503);
DFFARX1 I_10259  ( .D(I176757), .CLK(I2350), .RSTB(I176172), .Q(I176149) );
nand I_10260 (I176152,I176692,I176582);
not I_10261 (I176835,I2357);
not I_10262 (I176852,I277304);
nor I_10263 (I176869,I277325,I277331);
nand I_10264 (I176886,I176869,I277319);
nor I_10265 (I176903,I176852,I277325);
nand I_10266 (I176920,I176903,I277301);
not I_10267 (I176937,I176920);
not I_10268 (I176954,I277325);
nor I_10269 (I176824,I176920,I176954);
not I_10270 (I176985,I176954);
nand I_10271 (I176809,I176920,I176985);
not I_10272 (I177016,I277307);
nor I_10273 (I177033,I177016,I277328);
and I_10274 (I177050,I177033,I277316);
or I_10275 (I177067,I177050,I277322);
DFFARX1 I_10276  ( .D(I177067), .CLK(I2350), .RSTB(I176835), .Q(I177084) );
nor I_10277 (I177101,I177084,I176937);
DFFARX1 I_10278  ( .D(I177084), .CLK(I2350), .RSTB(I176835), .Q(I177118) );
not I_10279 (I176806,I177118);
nand I_10280 (I177149,I176852,I277307);
and I_10281 (I177166,I177149,I177101);
DFFARX1 I_10282  ( .D(I177149), .CLK(I2350), .RSTB(I176835), .Q(I176803) );
DFFARX1 I_10283  ( .D(I277313), .CLK(I2350), .RSTB(I176835), .Q(I177197) );
nor I_10284 (I177214,I177197,I176920);
nand I_10285 (I176821,I177084,I177214);
nor I_10286 (I177245,I177197,I176985);
not I_10287 (I176818,I177197);
nand I_10288 (I177276,I177197,I176886);
and I_10289 (I177293,I176954,I177276);
DFFARX1 I_10290  ( .D(I177293), .CLK(I2350), .RSTB(I176835), .Q(I176797) );
DFFARX1 I_10291  ( .D(I177197), .CLK(I2350), .RSTB(I176835), .Q(I176800) );
DFFARX1 I_10292  ( .D(I277310), .CLK(I2350), .RSTB(I176835), .Q(I177338) );
not I_10293 (I177355,I177338);
nand I_10294 (I177372,I177355,I176920);
and I_10295 (I177389,I177149,I177372);
DFFARX1 I_10296  ( .D(I177389), .CLK(I2350), .RSTB(I176835), .Q(I176827) );
or I_10297 (I177420,I177355,I177166);
DFFARX1 I_10298  ( .D(I177420), .CLK(I2350), .RSTB(I176835), .Q(I176812) );
nand I_10299 (I176815,I177355,I177245);
not I_10300 (I177498,I2357);
not I_10301 (I177515,I362171);
nor I_10302 (I177532,I362189,I362180);
nand I_10303 (I177549,I177532,I362186);
nor I_10304 (I177566,I177515,I362189);
nand I_10305 (I177583,I177566,I362192);
not I_10306 (I177600,I177583);
not I_10307 (I177617,I362189);
nor I_10308 (I177487,I177583,I177617);
not I_10309 (I177648,I177617);
nand I_10310 (I177472,I177583,I177648);
not I_10311 (I177679,I362168);
nor I_10312 (I177696,I177679,I362183);
and I_10313 (I177713,I177696,I362165);
or I_10314 (I177730,I177713,I362174);
DFFARX1 I_10315  ( .D(I177730), .CLK(I2350), .RSTB(I177498), .Q(I177747) );
nor I_10316 (I177764,I177747,I177600);
DFFARX1 I_10317  ( .D(I177747), .CLK(I2350), .RSTB(I177498), .Q(I177781) );
not I_10318 (I177469,I177781);
nand I_10319 (I177812,I177515,I362168);
and I_10320 (I177829,I177812,I177764);
DFFARX1 I_10321  ( .D(I177812), .CLK(I2350), .RSTB(I177498), .Q(I177466) );
DFFARX1 I_10322  ( .D(I362177), .CLK(I2350), .RSTB(I177498), .Q(I177860) );
nor I_10323 (I177877,I177860,I177583);
nand I_10324 (I177484,I177747,I177877);
nor I_10325 (I177908,I177860,I177648);
not I_10326 (I177481,I177860);
nand I_10327 (I177939,I177860,I177549);
and I_10328 (I177956,I177617,I177939);
DFFARX1 I_10329  ( .D(I177956), .CLK(I2350), .RSTB(I177498), .Q(I177460) );
DFFARX1 I_10330  ( .D(I177860), .CLK(I2350), .RSTB(I177498), .Q(I177463) );
DFFARX1 I_10331  ( .D(I362195), .CLK(I2350), .RSTB(I177498), .Q(I178001) );
not I_10332 (I178018,I178001);
nand I_10333 (I178035,I178018,I177583);
and I_10334 (I178052,I177812,I178035);
DFFARX1 I_10335  ( .D(I178052), .CLK(I2350), .RSTB(I177498), .Q(I177490) );
or I_10336 (I178083,I178018,I177829);
DFFARX1 I_10337  ( .D(I178083), .CLK(I2350), .RSTB(I177498), .Q(I177475) );
nand I_10338 (I177478,I178018,I177908);
not I_10339 (I178161,I2357);
not I_10340 (I178178,I132947);
nor I_10341 (I178195,I132920,I132923);
nand I_10342 (I178212,I178195,I132935);
nor I_10343 (I178229,I178178,I132920);
nand I_10344 (I178246,I178229,I132941);
not I_10345 (I178263,I178246);
not I_10346 (I178280,I132920);
nor I_10347 (I178150,I178246,I178280);
not I_10348 (I178311,I178280);
nand I_10349 (I178135,I178246,I178311);
not I_10350 (I178342,I132944);
nor I_10351 (I178359,I178342,I132926);
and I_10352 (I178376,I178359,I132929);
or I_10353 (I178393,I178376,I132950);
DFFARX1 I_10354  ( .D(I178393), .CLK(I2350), .RSTB(I178161), .Q(I178410) );
nor I_10355 (I178427,I178410,I178263);
DFFARX1 I_10356  ( .D(I178410), .CLK(I2350), .RSTB(I178161), .Q(I178444) );
not I_10357 (I178132,I178444);
nand I_10358 (I178475,I178178,I132944);
and I_10359 (I178492,I178475,I178427);
DFFARX1 I_10360  ( .D(I178475), .CLK(I2350), .RSTB(I178161), .Q(I178129) );
DFFARX1 I_10361  ( .D(I132932), .CLK(I2350), .RSTB(I178161), .Q(I178523) );
nor I_10362 (I178540,I178523,I178246);
nand I_10363 (I178147,I178410,I178540);
nor I_10364 (I178571,I178523,I178311);
not I_10365 (I178144,I178523);
nand I_10366 (I178602,I178523,I178212);
and I_10367 (I178619,I178280,I178602);
DFFARX1 I_10368  ( .D(I178619), .CLK(I2350), .RSTB(I178161), .Q(I178123) );
DFFARX1 I_10369  ( .D(I178523), .CLK(I2350), .RSTB(I178161), .Q(I178126) );
DFFARX1 I_10370  ( .D(I132938), .CLK(I2350), .RSTB(I178161), .Q(I178664) );
not I_10371 (I178681,I178664);
nand I_10372 (I178698,I178681,I178246);
and I_10373 (I178715,I178475,I178698);
DFFARX1 I_10374  ( .D(I178715), .CLK(I2350), .RSTB(I178161), .Q(I178153) );
or I_10375 (I178746,I178681,I178492);
DFFARX1 I_10376  ( .D(I178746), .CLK(I2350), .RSTB(I178161), .Q(I178138) );
nand I_10377 (I178141,I178681,I178571);
not I_10378 (I178824,I2357);
not I_10379 (I178841,I121038);
nor I_10380 (I178858,I121032,I121023);
nand I_10381 (I178875,I178858,I121035);
nor I_10382 (I178892,I178841,I121032);
nand I_10383 (I178909,I178892,I121050);
not I_10384 (I178926,I178909);
not I_10385 (I178943,I121032);
nor I_10386 (I178813,I178909,I178943);
not I_10387 (I178974,I178943);
nand I_10388 (I178798,I178909,I178974);
not I_10389 (I179005,I121026);
nor I_10390 (I179022,I179005,I121020);
and I_10391 (I179039,I179022,I121047);
or I_10392 (I179056,I179039,I121044);
DFFARX1 I_10393  ( .D(I179056), .CLK(I2350), .RSTB(I178824), .Q(I179073) );
nor I_10394 (I179090,I179073,I178926);
DFFARX1 I_10395  ( .D(I179073), .CLK(I2350), .RSTB(I178824), .Q(I179107) );
not I_10396 (I178795,I179107);
nand I_10397 (I179138,I178841,I121026);
and I_10398 (I179155,I179138,I179090);
DFFARX1 I_10399  ( .D(I179138), .CLK(I2350), .RSTB(I178824), .Q(I178792) );
DFFARX1 I_10400  ( .D(I121041), .CLK(I2350), .RSTB(I178824), .Q(I179186) );
nor I_10401 (I179203,I179186,I178909);
nand I_10402 (I178810,I179073,I179203);
nor I_10403 (I179234,I179186,I178974);
not I_10404 (I178807,I179186);
nand I_10405 (I179265,I179186,I178875);
and I_10406 (I179282,I178943,I179265);
DFFARX1 I_10407  ( .D(I179282), .CLK(I2350), .RSTB(I178824), .Q(I178786) );
DFFARX1 I_10408  ( .D(I179186), .CLK(I2350), .RSTB(I178824), .Q(I178789) );
DFFARX1 I_10409  ( .D(I121029), .CLK(I2350), .RSTB(I178824), .Q(I179327) );
not I_10410 (I179344,I179327);
nand I_10411 (I179361,I179344,I178909);
and I_10412 (I179378,I179138,I179361);
DFFARX1 I_10413  ( .D(I179378), .CLK(I2350), .RSTB(I178824), .Q(I178816) );
or I_10414 (I179409,I179344,I179155);
DFFARX1 I_10415  ( .D(I179409), .CLK(I2350), .RSTB(I178824), .Q(I178801) );
nand I_10416 (I178804,I179344,I179234);
not I_10417 (I179487,I2357);
not I_10418 (I179504,I374122);
nor I_10419 (I179521,I374140,I374131);
nand I_10420 (I179538,I179521,I374137);
nor I_10421 (I179555,I179504,I374140);
nand I_10422 (I179572,I179555,I374143);
not I_10423 (I179589,I179572);
not I_10424 (I179606,I374140);
nor I_10425 (I179476,I179572,I179606);
not I_10426 (I179637,I179606);
nand I_10427 (I179461,I179572,I179637);
not I_10428 (I179668,I374119);
nor I_10429 (I179685,I179668,I374134);
and I_10430 (I179702,I179685,I374116);
or I_10431 (I179719,I179702,I374125);
DFFARX1 I_10432  ( .D(I179719), .CLK(I2350), .RSTB(I179487), .Q(I179736) );
nor I_10433 (I179753,I179736,I179589);
DFFARX1 I_10434  ( .D(I179736), .CLK(I2350), .RSTB(I179487), .Q(I179770) );
not I_10435 (I179458,I179770);
nand I_10436 (I179801,I179504,I374119);
and I_10437 (I179818,I179801,I179753);
DFFARX1 I_10438  ( .D(I179801), .CLK(I2350), .RSTB(I179487), .Q(I179455) );
DFFARX1 I_10439  ( .D(I374128), .CLK(I2350), .RSTB(I179487), .Q(I179849) );
nor I_10440 (I179866,I179849,I179572);
nand I_10441 (I179473,I179736,I179866);
nor I_10442 (I179897,I179849,I179637);
not I_10443 (I179470,I179849);
nand I_10444 (I179928,I179849,I179538);
and I_10445 (I179945,I179606,I179928);
DFFARX1 I_10446  ( .D(I179945), .CLK(I2350), .RSTB(I179487), .Q(I179449) );
DFFARX1 I_10447  ( .D(I179849), .CLK(I2350), .RSTB(I179487), .Q(I179452) );
DFFARX1 I_10448  ( .D(I374146), .CLK(I2350), .RSTB(I179487), .Q(I179990) );
not I_10449 (I180007,I179990);
nand I_10450 (I180024,I180007,I179572);
and I_10451 (I180041,I179801,I180024);
DFFARX1 I_10452  ( .D(I180041), .CLK(I2350), .RSTB(I179487), .Q(I179479) );
or I_10453 (I180072,I180007,I179818);
DFFARX1 I_10454  ( .D(I180072), .CLK(I2350), .RSTB(I179487), .Q(I179464) );
nand I_10455 (I179467,I180007,I179897);
not I_10456 (I180150,I2357);
not I_10457 (I180167,I367203);
nor I_10458 (I180184,I367221,I367212);
nand I_10459 (I180201,I180184,I367218);
nor I_10460 (I180218,I180167,I367221);
nand I_10461 (I180235,I180218,I367224);
not I_10462 (I180252,I180235);
not I_10463 (I180269,I367221);
nor I_10464 (I180139,I180235,I180269);
not I_10465 (I180300,I180269);
nand I_10466 (I180124,I180235,I180300);
not I_10467 (I180331,I367200);
nor I_10468 (I180348,I180331,I367215);
and I_10469 (I180365,I180348,I367197);
or I_10470 (I180382,I180365,I367206);
DFFARX1 I_10471  ( .D(I180382), .CLK(I2350), .RSTB(I180150), .Q(I180399) );
nor I_10472 (I180416,I180399,I180252);
DFFARX1 I_10473  ( .D(I180399), .CLK(I2350), .RSTB(I180150), .Q(I180433) );
not I_10474 (I180121,I180433);
nand I_10475 (I180464,I180167,I367200);
and I_10476 (I180481,I180464,I180416);
DFFARX1 I_10477  ( .D(I180464), .CLK(I2350), .RSTB(I180150), .Q(I180118) );
DFFARX1 I_10478  ( .D(I367209), .CLK(I2350), .RSTB(I180150), .Q(I180512) );
nor I_10479 (I180529,I180512,I180235);
nand I_10480 (I180136,I180399,I180529);
nor I_10481 (I180560,I180512,I180300);
not I_10482 (I180133,I180512);
nand I_10483 (I180591,I180512,I180201);
and I_10484 (I180608,I180269,I180591);
DFFARX1 I_10485  ( .D(I180608), .CLK(I2350), .RSTB(I180150), .Q(I180112) );
DFFARX1 I_10486  ( .D(I180512), .CLK(I2350), .RSTB(I180150), .Q(I180115) );
DFFARX1 I_10487  ( .D(I367227), .CLK(I2350), .RSTB(I180150), .Q(I180653) );
not I_10488 (I180670,I180653);
nand I_10489 (I180687,I180670,I180235);
and I_10490 (I180704,I180464,I180687);
DFFARX1 I_10491  ( .D(I180704), .CLK(I2350), .RSTB(I180150), .Q(I180142) );
or I_10492 (I180735,I180670,I180481);
DFFARX1 I_10493  ( .D(I180735), .CLK(I2350), .RSTB(I180150), .Q(I180127) );
nand I_10494 (I180130,I180670,I180560);
not I_10495 (I180813,I2357);
not I_10496 (I180830,I249878);
nor I_10497 (I180847,I249890,I249872);
nand I_10498 (I180864,I180847,I249893);
nor I_10499 (I180881,I180830,I249890);
nand I_10500 (I180898,I180881,I249884);
not I_10501 (I180915,I180898);
not I_10502 (I180932,I249890);
nor I_10503 (I180802,I180898,I180932);
not I_10504 (I180963,I180932);
nand I_10505 (I180787,I180898,I180963);
not I_10506 (I180994,I249875);
nor I_10507 (I181011,I180994,I249869);
and I_10508 (I181028,I181011,I249881);
or I_10509 (I181045,I181028,I249866);
DFFARX1 I_10510  ( .D(I181045), .CLK(I2350), .RSTB(I180813), .Q(I181062) );
nor I_10511 (I181079,I181062,I180915);
DFFARX1 I_10512  ( .D(I181062), .CLK(I2350), .RSTB(I180813), .Q(I181096) );
not I_10513 (I180784,I181096);
nand I_10514 (I181127,I180830,I249875);
and I_10515 (I181144,I181127,I181079);
DFFARX1 I_10516  ( .D(I181127), .CLK(I2350), .RSTB(I180813), .Q(I180781) );
DFFARX1 I_10517  ( .D(I249863), .CLK(I2350), .RSTB(I180813), .Q(I181175) );
nor I_10518 (I181192,I181175,I180898);
nand I_10519 (I180799,I181062,I181192);
nor I_10520 (I181223,I181175,I180963);
not I_10521 (I180796,I181175);
nand I_10522 (I181254,I181175,I180864);
and I_10523 (I181271,I180932,I181254);
DFFARX1 I_10524  ( .D(I181271), .CLK(I2350), .RSTB(I180813), .Q(I180775) );
DFFARX1 I_10525  ( .D(I181175), .CLK(I2350), .RSTB(I180813), .Q(I180778) );
DFFARX1 I_10526  ( .D(I249887), .CLK(I2350), .RSTB(I180813), .Q(I181316) );
not I_10527 (I181333,I181316);
nand I_10528 (I181350,I181333,I180898);
and I_10529 (I181367,I181127,I181350);
DFFARX1 I_10530  ( .D(I181367), .CLK(I2350), .RSTB(I180813), .Q(I180805) );
or I_10531 (I181398,I181333,I181144);
DFFARX1 I_10532  ( .D(I181398), .CLK(I2350), .RSTB(I180813), .Q(I180790) );
nand I_10533 (I180793,I181333,I181223);
not I_10534 (I181476,I2357);
not I_10535 (I181493,I264328);
nor I_10536 (I181510,I264340,I264322);
nand I_10537 (I181527,I181510,I264343);
nor I_10538 (I181544,I181493,I264340);
nand I_10539 (I181561,I181544,I264334);
not I_10540 (I181578,I181561);
not I_10541 (I181595,I264340);
nor I_10542 (I181465,I181561,I181595);
not I_10543 (I181626,I181595);
nand I_10544 (I181450,I181561,I181626);
not I_10545 (I181657,I264325);
nor I_10546 (I181674,I181657,I264319);
and I_10547 (I181691,I181674,I264331);
or I_10548 (I181708,I181691,I264316);
DFFARX1 I_10549  ( .D(I181708), .CLK(I2350), .RSTB(I181476), .Q(I181725) );
nor I_10550 (I181742,I181725,I181578);
DFFARX1 I_10551  ( .D(I181725), .CLK(I2350), .RSTB(I181476), .Q(I181759) );
not I_10552 (I181447,I181759);
nand I_10553 (I181790,I181493,I264325);
and I_10554 (I181807,I181790,I181742);
DFFARX1 I_10555  ( .D(I181790), .CLK(I2350), .RSTB(I181476), .Q(I181444) );
DFFARX1 I_10556  ( .D(I264313), .CLK(I2350), .RSTB(I181476), .Q(I181838) );
nor I_10557 (I181855,I181838,I181561);
nand I_10558 (I181462,I181725,I181855);
nor I_10559 (I181886,I181838,I181626);
not I_10560 (I181459,I181838);
nand I_10561 (I181917,I181838,I181527);
and I_10562 (I181934,I181595,I181917);
DFFARX1 I_10563  ( .D(I181934), .CLK(I2350), .RSTB(I181476), .Q(I181438) );
DFFARX1 I_10564  ( .D(I181838), .CLK(I2350), .RSTB(I181476), .Q(I181441) );
DFFARX1 I_10565  ( .D(I264337), .CLK(I2350), .RSTB(I181476), .Q(I181979) );
not I_10566 (I181996,I181979);
nand I_10567 (I182013,I181996,I181561);
and I_10568 (I182030,I181790,I182013);
DFFARX1 I_10569  ( .D(I182030), .CLK(I2350), .RSTB(I181476), .Q(I181468) );
or I_10570 (I182061,I181996,I181807);
DFFARX1 I_10571  ( .D(I182061), .CLK(I2350), .RSTB(I181476), .Q(I181453) );
nand I_10572 (I181456,I181996,I181886);
not I_10573 (I182139,I2357);
not I_10574 (I182156,I92004);
nor I_10575 (I182173,I92010,I92016);
nand I_10576 (I182190,I182173,I92019);
nor I_10577 (I182207,I182156,I92010);
nand I_10578 (I182224,I182207,I92001);
not I_10579 (I182241,I182224);
not I_10580 (I182258,I92010);
nor I_10581 (I182128,I182224,I182258);
not I_10582 (I182289,I182258);
nand I_10583 (I182113,I182224,I182289);
not I_10584 (I182320,I92013);
nor I_10585 (I182337,I182320,I92007);
and I_10586 (I182354,I182337,I92022);
or I_10587 (I182371,I182354,I92028);
DFFARX1 I_10588  ( .D(I182371), .CLK(I2350), .RSTB(I182139), .Q(I182388) );
nor I_10589 (I182405,I182388,I182241);
DFFARX1 I_10590  ( .D(I182388), .CLK(I2350), .RSTB(I182139), .Q(I182422) );
not I_10591 (I182110,I182422);
nand I_10592 (I182453,I182156,I92013);
and I_10593 (I182470,I182453,I182405);
DFFARX1 I_10594  ( .D(I182453), .CLK(I2350), .RSTB(I182139), .Q(I182107) );
DFFARX1 I_10595  ( .D(I92025), .CLK(I2350), .RSTB(I182139), .Q(I182501) );
nor I_10596 (I182518,I182501,I182224);
nand I_10597 (I182125,I182388,I182518);
nor I_10598 (I182549,I182501,I182289);
not I_10599 (I182122,I182501);
nand I_10600 (I182580,I182501,I182190);
and I_10601 (I182597,I182258,I182580);
DFFARX1 I_10602  ( .D(I182597), .CLK(I2350), .RSTB(I182139), .Q(I182101) );
DFFARX1 I_10603  ( .D(I182501), .CLK(I2350), .RSTB(I182139), .Q(I182104) );
DFFARX1 I_10604  ( .D(I92031), .CLK(I2350), .RSTB(I182139), .Q(I182642) );
not I_10605 (I182659,I182642);
nand I_10606 (I182676,I182659,I182224);
and I_10607 (I182693,I182453,I182676);
DFFARX1 I_10608  ( .D(I182693), .CLK(I2350), .RSTB(I182139), .Q(I182131) );
or I_10609 (I182724,I182659,I182470);
DFFARX1 I_10610  ( .D(I182724), .CLK(I2350), .RSTB(I182139), .Q(I182116) );
nand I_10611 (I182119,I182659,I182549);
not I_10612 (I182802,I2357);
not I_10613 (I182819,I365316);
nor I_10614 (I182836,I365334,I365325);
nand I_10615 (I182853,I182836,I365331);
nor I_10616 (I182870,I182819,I365334);
nand I_10617 (I182887,I182870,I365337);
not I_10618 (I182904,I182887);
not I_10619 (I182921,I365334);
nor I_10620 (I182791,I182887,I182921);
not I_10621 (I182952,I182921);
nand I_10622 (I182776,I182887,I182952);
not I_10623 (I182983,I365313);
nor I_10624 (I183000,I182983,I365328);
and I_10625 (I183017,I183000,I365310);
or I_10626 (I183034,I183017,I365319);
DFFARX1 I_10627  ( .D(I183034), .CLK(I2350), .RSTB(I182802), .Q(I183051) );
nor I_10628 (I183068,I183051,I182904);
DFFARX1 I_10629  ( .D(I183051), .CLK(I2350), .RSTB(I182802), .Q(I183085) );
not I_10630 (I182773,I183085);
nand I_10631 (I183116,I182819,I365313);
and I_10632 (I183133,I183116,I183068);
DFFARX1 I_10633  ( .D(I183116), .CLK(I2350), .RSTB(I182802), .Q(I182770) );
DFFARX1 I_10634  ( .D(I365322), .CLK(I2350), .RSTB(I182802), .Q(I183164) );
nor I_10635 (I183181,I183164,I182887);
nand I_10636 (I182788,I183051,I183181);
nor I_10637 (I183212,I183164,I182952);
not I_10638 (I182785,I183164);
nand I_10639 (I183243,I183164,I182853);
and I_10640 (I183260,I182921,I183243);
DFFARX1 I_10641  ( .D(I183260), .CLK(I2350), .RSTB(I182802), .Q(I182764) );
DFFARX1 I_10642  ( .D(I183164), .CLK(I2350), .RSTB(I182802), .Q(I182767) );
DFFARX1 I_10643  ( .D(I365340), .CLK(I2350), .RSTB(I182802), .Q(I183305) );
not I_10644 (I183322,I183305);
nand I_10645 (I183339,I183322,I182887);
and I_10646 (I183356,I183116,I183339);
DFFARX1 I_10647  ( .D(I183356), .CLK(I2350), .RSTB(I182802), .Q(I182794) );
or I_10648 (I183387,I183322,I183133);
DFFARX1 I_10649  ( .D(I183387), .CLK(I2350), .RSTB(I182802), .Q(I182779) );
nand I_10650 (I182782,I183322,I183212);
not I_10651 (I183465,I2357);
not I_10652 (I183482,I289780);
nor I_10653 (I183499,I289789,I289771);
nand I_10654 (I183516,I183499,I289792);
nor I_10655 (I183533,I183482,I289789);
nand I_10656 (I183550,I183533,I289783);
not I_10657 (I183567,I183550);
not I_10658 (I183584,I289789);
nor I_10659 (I183454,I183550,I183584);
not I_10660 (I183615,I183584);
nand I_10661 (I183439,I183550,I183615);
not I_10662 (I183646,I289777);
nor I_10663 (I183663,I183646,I289768);
and I_10664 (I183680,I183663,I289765);
or I_10665 (I183697,I183680,I289762);
DFFARX1 I_10666  ( .D(I183697), .CLK(I2350), .RSTB(I183465), .Q(I183714) );
nor I_10667 (I183731,I183714,I183567);
DFFARX1 I_10668  ( .D(I183714), .CLK(I2350), .RSTB(I183465), .Q(I183748) );
not I_10669 (I183436,I183748);
nand I_10670 (I183779,I183482,I289777);
and I_10671 (I183796,I183779,I183731);
DFFARX1 I_10672  ( .D(I183779), .CLK(I2350), .RSTB(I183465), .Q(I183433) );
DFFARX1 I_10673  ( .D(I289786), .CLK(I2350), .RSTB(I183465), .Q(I183827) );
nor I_10674 (I183844,I183827,I183550);
nand I_10675 (I183451,I183714,I183844);
nor I_10676 (I183875,I183827,I183615);
not I_10677 (I183448,I183827);
nand I_10678 (I183906,I183827,I183516);
and I_10679 (I183923,I183584,I183906);
DFFARX1 I_10680  ( .D(I183923), .CLK(I2350), .RSTB(I183465), .Q(I183427) );
DFFARX1 I_10681  ( .D(I183827), .CLK(I2350), .RSTB(I183465), .Q(I183430) );
DFFARX1 I_10682  ( .D(I289774), .CLK(I2350), .RSTB(I183465), .Q(I183968) );
not I_10683 (I183985,I183968);
nand I_10684 (I184002,I183985,I183550);
and I_10685 (I184019,I183779,I184002);
DFFARX1 I_10686  ( .D(I184019), .CLK(I2350), .RSTB(I183465), .Q(I183457) );
or I_10687 (I184050,I183985,I183796);
DFFARX1 I_10688  ( .D(I184050), .CLK(I2350), .RSTB(I183465), .Q(I183442) );
nand I_10689 (I183445,I183985,I183875);
not I_10690 (I184128,I2357);
not I_10691 (I184145,I77608);
nor I_10692 (I184162,I77605,I77629);
nand I_10693 (I184179,I184162,I77626);
nor I_10694 (I184196,I184145,I77605);
nand I_10695 (I184213,I184196,I77632);
not I_10696 (I184230,I184213);
not I_10697 (I184247,I77605);
nor I_10698 (I184117,I184213,I184247);
not I_10699 (I184278,I184247);
nand I_10700 (I184102,I184213,I184278);
not I_10701 (I184309,I77623);
nor I_10702 (I184326,I184309,I77614);
and I_10703 (I184343,I184326,I77611);
or I_10704 (I184360,I184343,I77620);
DFFARX1 I_10705  ( .D(I184360), .CLK(I2350), .RSTB(I184128), .Q(I184377) );
nor I_10706 (I184394,I184377,I184230);
DFFARX1 I_10707  ( .D(I184377), .CLK(I2350), .RSTB(I184128), .Q(I184411) );
not I_10708 (I184099,I184411);
nand I_10709 (I184442,I184145,I77623);
and I_10710 (I184459,I184442,I184394);
DFFARX1 I_10711  ( .D(I184442), .CLK(I2350), .RSTB(I184128), .Q(I184096) );
DFFARX1 I_10712  ( .D(I77602), .CLK(I2350), .RSTB(I184128), .Q(I184490) );
nor I_10713 (I184507,I184490,I184213);
nand I_10714 (I184114,I184377,I184507);
nor I_10715 (I184538,I184490,I184278);
not I_10716 (I184111,I184490);
nand I_10717 (I184569,I184490,I184179);
and I_10718 (I184586,I184247,I184569);
DFFARX1 I_10719  ( .D(I184586), .CLK(I2350), .RSTB(I184128), .Q(I184090) );
DFFARX1 I_10720  ( .D(I184490), .CLK(I2350), .RSTB(I184128), .Q(I184093) );
DFFARX1 I_10721  ( .D(I77617), .CLK(I2350), .RSTB(I184128), .Q(I184631) );
not I_10722 (I184648,I184631);
nand I_10723 (I184665,I184648,I184213);
and I_10724 (I184682,I184442,I184665);
DFFARX1 I_10725  ( .D(I184682), .CLK(I2350), .RSTB(I184128), .Q(I184120) );
or I_10726 (I184713,I184648,I184459);
DFFARX1 I_10727  ( .D(I184713), .CLK(I2350), .RSTB(I184128), .Q(I184105) );
nand I_10728 (I184108,I184648,I184538);
not I_10729 (I184791,I2357);
not I_10730 (I184808,I255658);
nor I_10731 (I184825,I255670,I255652);
nand I_10732 (I184842,I184825,I255673);
nor I_10733 (I184859,I184808,I255670);
nand I_10734 (I184876,I184859,I255664);
not I_10735 (I184893,I184876);
not I_10736 (I184910,I255670);
nor I_10737 (I184780,I184876,I184910);
not I_10738 (I184941,I184910);
nand I_10739 (I184765,I184876,I184941);
not I_10740 (I184972,I255655);
nor I_10741 (I184989,I184972,I255649);
and I_10742 (I185006,I184989,I255661);
or I_10743 (I185023,I185006,I255646);
DFFARX1 I_10744  ( .D(I185023), .CLK(I2350), .RSTB(I184791), .Q(I185040) );
nor I_10745 (I185057,I185040,I184893);
DFFARX1 I_10746  ( .D(I185040), .CLK(I2350), .RSTB(I184791), .Q(I185074) );
not I_10747 (I184762,I185074);
nand I_10748 (I185105,I184808,I255655);
and I_10749 (I185122,I185105,I185057);
DFFARX1 I_10750  ( .D(I185105), .CLK(I2350), .RSTB(I184791), .Q(I184759) );
DFFARX1 I_10751  ( .D(I255643), .CLK(I2350), .RSTB(I184791), .Q(I185153) );
nor I_10752 (I185170,I185153,I184876);
nand I_10753 (I184777,I185040,I185170);
nor I_10754 (I185201,I185153,I184941);
not I_10755 (I184774,I185153);
nand I_10756 (I185232,I185153,I184842);
and I_10757 (I185249,I184910,I185232);
DFFARX1 I_10758  ( .D(I185249), .CLK(I2350), .RSTB(I184791), .Q(I184753) );
DFFARX1 I_10759  ( .D(I185153), .CLK(I2350), .RSTB(I184791), .Q(I184756) );
DFFARX1 I_10760  ( .D(I255667), .CLK(I2350), .RSTB(I184791), .Q(I185294) );
not I_10761 (I185311,I185294);
nand I_10762 (I185328,I185311,I184876);
and I_10763 (I185345,I185105,I185328);
DFFARX1 I_10764  ( .D(I185345), .CLK(I2350), .RSTB(I184791), .Q(I184783) );
or I_10765 (I185376,I185311,I185122);
DFFARX1 I_10766  ( .D(I185376), .CLK(I2350), .RSTB(I184791), .Q(I184768) );
nand I_10767 (I184771,I185311,I185201);
not I_10768 (I185454,I2357);
not I_10769 (I185471,I358397);
nor I_10770 (I185488,I358415,I358406);
nand I_10771 (I185505,I185488,I358412);
nor I_10772 (I185522,I185471,I358415);
nand I_10773 (I185539,I185522,I358418);
not I_10774 (I185556,I185539);
not I_10775 (I185573,I358415);
nor I_10776 (I185443,I185539,I185573);
not I_10777 (I185604,I185573);
nand I_10778 (I185428,I185539,I185604);
not I_10779 (I185635,I358394);
nor I_10780 (I185652,I185635,I358409);
and I_10781 (I185669,I185652,I358391);
or I_10782 (I185686,I185669,I358400);
DFFARX1 I_10783  ( .D(I185686), .CLK(I2350), .RSTB(I185454), .Q(I185703) );
nor I_10784 (I185720,I185703,I185556);
DFFARX1 I_10785  ( .D(I185703), .CLK(I2350), .RSTB(I185454), .Q(I185737) );
not I_10786 (I185425,I185737);
nand I_10787 (I185768,I185471,I358394);
and I_10788 (I185785,I185768,I185720);
DFFARX1 I_10789  ( .D(I185768), .CLK(I2350), .RSTB(I185454), .Q(I185422) );
DFFARX1 I_10790  ( .D(I358403), .CLK(I2350), .RSTB(I185454), .Q(I185816) );
nor I_10791 (I185833,I185816,I185539);
nand I_10792 (I185440,I185703,I185833);
nor I_10793 (I185864,I185816,I185604);
not I_10794 (I185437,I185816);
nand I_10795 (I185895,I185816,I185505);
and I_10796 (I185912,I185573,I185895);
DFFARX1 I_10797  ( .D(I185912), .CLK(I2350), .RSTB(I185454), .Q(I185416) );
DFFARX1 I_10798  ( .D(I185816), .CLK(I2350), .RSTB(I185454), .Q(I185419) );
DFFARX1 I_10799  ( .D(I358421), .CLK(I2350), .RSTB(I185454), .Q(I185957) );
not I_10800 (I185974,I185957);
nand I_10801 (I185991,I185974,I185539);
and I_10802 (I186008,I185768,I185991);
DFFARX1 I_10803  ( .D(I186008), .CLK(I2350), .RSTB(I185454), .Q(I185446) );
or I_10804 (I186039,I185974,I185785);
DFFARX1 I_10805  ( .D(I186039), .CLK(I2350), .RSTB(I185454), .Q(I185431) );
nand I_10806 (I185434,I185974,I185864);
not I_10807 (I186117,I2357);
not I_10808 (I186134,I245254);
nor I_10809 (I186151,I245266,I245248);
nand I_10810 (I186168,I186151,I245269);
nor I_10811 (I186185,I186134,I245266);
nand I_10812 (I186202,I186185,I245260);
not I_10813 (I186219,I186202);
not I_10814 (I186236,I245266);
nor I_10815 (I186106,I186202,I186236);
not I_10816 (I186267,I186236);
nand I_10817 (I186091,I186202,I186267);
not I_10818 (I186298,I245251);
nor I_10819 (I186315,I186298,I245245);
and I_10820 (I186332,I186315,I245257);
or I_10821 (I186349,I186332,I245242);
DFFARX1 I_10822  ( .D(I186349), .CLK(I2350), .RSTB(I186117), .Q(I186366) );
nor I_10823 (I186383,I186366,I186219);
DFFARX1 I_10824  ( .D(I186366), .CLK(I2350), .RSTB(I186117), .Q(I186400) );
not I_10825 (I186088,I186400);
nand I_10826 (I186431,I186134,I245251);
and I_10827 (I186448,I186431,I186383);
DFFARX1 I_10828  ( .D(I186431), .CLK(I2350), .RSTB(I186117), .Q(I186085) );
DFFARX1 I_10829  ( .D(I245239), .CLK(I2350), .RSTB(I186117), .Q(I186479) );
nor I_10830 (I186496,I186479,I186202);
nand I_10831 (I186103,I186366,I186496);
nor I_10832 (I186527,I186479,I186267);
not I_10833 (I186100,I186479);
nand I_10834 (I186558,I186479,I186168);
and I_10835 (I186575,I186236,I186558);
DFFARX1 I_10836  ( .D(I186575), .CLK(I2350), .RSTB(I186117), .Q(I186079) );
DFFARX1 I_10837  ( .D(I186479), .CLK(I2350), .RSTB(I186117), .Q(I186082) );
DFFARX1 I_10838  ( .D(I245263), .CLK(I2350), .RSTB(I186117), .Q(I186620) );
not I_10839 (I186637,I186620);
nand I_10840 (I186654,I186637,I186202);
and I_10841 (I186671,I186431,I186654);
DFFARX1 I_10842  ( .D(I186671), .CLK(I2350), .RSTB(I186117), .Q(I186109) );
or I_10843 (I186702,I186637,I186448);
DFFARX1 I_10844  ( .D(I186702), .CLK(I2350), .RSTB(I186117), .Q(I186094) );
nand I_10845 (I186097,I186637,I186527);
not I_10846 (I186780,I2357);
not I_10847 (I186797,I308225);
nor I_10848 (I186814,I308234,I308216);
nand I_10849 (I186831,I186814,I308237);
nor I_10850 (I186848,I186797,I308234);
nand I_10851 (I186865,I186848,I308228);
not I_10852 (I186882,I186865);
not I_10853 (I186899,I308234);
nor I_10854 (I186769,I186865,I186899);
not I_10855 (I186930,I186899);
nand I_10856 (I186754,I186865,I186930);
not I_10857 (I186961,I308222);
nor I_10858 (I186978,I186961,I308213);
and I_10859 (I186995,I186978,I308210);
or I_10860 (I187012,I186995,I308207);
DFFARX1 I_10861  ( .D(I187012), .CLK(I2350), .RSTB(I186780), .Q(I187029) );
nor I_10862 (I187046,I187029,I186882);
DFFARX1 I_10863  ( .D(I187029), .CLK(I2350), .RSTB(I186780), .Q(I187063) );
not I_10864 (I186751,I187063);
nand I_10865 (I187094,I186797,I308222);
and I_10866 (I187111,I187094,I187046);
DFFARX1 I_10867  ( .D(I187094), .CLK(I2350), .RSTB(I186780), .Q(I186748) );
DFFARX1 I_10868  ( .D(I308231), .CLK(I2350), .RSTB(I186780), .Q(I187142) );
nor I_10869 (I187159,I187142,I186865);
nand I_10870 (I186766,I187029,I187159);
nor I_10871 (I187190,I187142,I186930);
not I_10872 (I186763,I187142);
nand I_10873 (I187221,I187142,I186831);
and I_10874 (I187238,I186899,I187221);
DFFARX1 I_10875  ( .D(I187238), .CLK(I2350), .RSTB(I186780), .Q(I186742) );
DFFARX1 I_10876  ( .D(I187142), .CLK(I2350), .RSTB(I186780), .Q(I186745) );
DFFARX1 I_10877  ( .D(I308219), .CLK(I2350), .RSTB(I186780), .Q(I187283) );
not I_10878 (I187300,I187283);
nand I_10879 (I187317,I187300,I186865);
and I_10880 (I187334,I187094,I187317);
DFFARX1 I_10881  ( .D(I187334), .CLK(I2350), .RSTB(I186780), .Q(I186772) );
or I_10882 (I187365,I187300,I187111);
DFFARX1 I_10883  ( .D(I187365), .CLK(I2350), .RSTB(I186780), .Q(I186757) );
nand I_10884 (I186760,I187300,I187190);
not I_10885 (I187443,I2357);
not I_10886 (I187460,I285615);
nor I_10887 (I187477,I285624,I285606);
nand I_10888 (I187494,I187477,I285627);
nor I_10889 (I187511,I187460,I285624);
nand I_10890 (I187528,I187511,I285618);
not I_10891 (I187545,I187528);
not I_10892 (I187562,I285624);
nor I_10893 (I187432,I187528,I187562);
not I_10894 (I187593,I187562);
nand I_10895 (I187417,I187528,I187593);
not I_10896 (I187624,I285612);
nor I_10897 (I187641,I187624,I285603);
and I_10898 (I187658,I187641,I285600);
or I_10899 (I187675,I187658,I285597);
DFFARX1 I_10900  ( .D(I187675), .CLK(I2350), .RSTB(I187443), .Q(I187692) );
nor I_10901 (I187709,I187692,I187545);
DFFARX1 I_10902  ( .D(I187692), .CLK(I2350), .RSTB(I187443), .Q(I187726) );
not I_10903 (I187414,I187726);
nand I_10904 (I187757,I187460,I285612);
and I_10905 (I187774,I187757,I187709);
DFFARX1 I_10906  ( .D(I187757), .CLK(I2350), .RSTB(I187443), .Q(I187411) );
DFFARX1 I_10907  ( .D(I285621), .CLK(I2350), .RSTB(I187443), .Q(I187805) );
nor I_10908 (I187822,I187805,I187528);
nand I_10909 (I187429,I187692,I187822);
nor I_10910 (I187853,I187805,I187593);
not I_10911 (I187426,I187805);
nand I_10912 (I187884,I187805,I187494);
and I_10913 (I187901,I187562,I187884);
DFFARX1 I_10914  ( .D(I187901), .CLK(I2350), .RSTB(I187443), .Q(I187405) );
DFFARX1 I_10915  ( .D(I187805), .CLK(I2350), .RSTB(I187443), .Q(I187408) );
DFFARX1 I_10916  ( .D(I285609), .CLK(I2350), .RSTB(I187443), .Q(I187946) );
not I_10917 (I187963,I187946);
nand I_10918 (I187980,I187963,I187528);
and I_10919 (I187997,I187757,I187980);
DFFARX1 I_10920  ( .D(I187997), .CLK(I2350), .RSTB(I187443), .Q(I187435) );
or I_10921 (I188028,I187963,I187774);
DFFARX1 I_10922  ( .D(I188028), .CLK(I2350), .RSTB(I187443), .Q(I187420) );
nand I_10923 (I187423,I187963,I187853);
not I_10924 (I188106,I2357);
not I_10925 (I188123,I38848);
nor I_10926 (I188140,I38845,I38869);
nand I_10927 (I188157,I188140,I38866);
nor I_10928 (I188174,I188123,I38845);
nand I_10929 (I188191,I188174,I38872);
not I_10930 (I188208,I188191);
not I_10931 (I188225,I38845);
nor I_10932 (I188095,I188191,I188225);
not I_10933 (I188256,I188225);
nand I_10934 (I188080,I188191,I188256);
not I_10935 (I188287,I38863);
nor I_10936 (I188304,I188287,I38854);
and I_10937 (I188321,I188304,I38851);
or I_10938 (I188338,I188321,I38860);
DFFARX1 I_10939  ( .D(I188338), .CLK(I2350), .RSTB(I188106), .Q(I188355) );
nor I_10940 (I188372,I188355,I188208);
DFFARX1 I_10941  ( .D(I188355), .CLK(I2350), .RSTB(I188106), .Q(I188389) );
not I_10942 (I188077,I188389);
nand I_10943 (I188420,I188123,I38863);
and I_10944 (I188437,I188420,I188372);
DFFARX1 I_10945  ( .D(I188420), .CLK(I2350), .RSTB(I188106), .Q(I188074) );
DFFARX1 I_10946  ( .D(I38842), .CLK(I2350), .RSTB(I188106), .Q(I188468) );
nor I_10947 (I188485,I188468,I188191);
nand I_10948 (I188092,I188355,I188485);
nor I_10949 (I188516,I188468,I188256);
not I_10950 (I188089,I188468);
nand I_10951 (I188547,I188468,I188157);
and I_10952 (I188564,I188225,I188547);
DFFARX1 I_10953  ( .D(I188564), .CLK(I2350), .RSTB(I188106), .Q(I188068) );
DFFARX1 I_10954  ( .D(I188468), .CLK(I2350), .RSTB(I188106), .Q(I188071) );
DFFARX1 I_10955  ( .D(I38857), .CLK(I2350), .RSTB(I188106), .Q(I188609) );
not I_10956 (I188626,I188609);
nand I_10957 (I188643,I188626,I188191);
and I_10958 (I188660,I188420,I188643);
DFFARX1 I_10959  ( .D(I188660), .CLK(I2350), .RSTB(I188106), .Q(I188098) );
or I_10960 (I188691,I188626,I188437);
DFFARX1 I_10961  ( .D(I188691), .CLK(I2350), .RSTB(I188106), .Q(I188083) );
nand I_10962 (I188086,I188626,I188516);
not I_10963 (I188769,I2357);
not I_10964 (I188786,I134732);
nor I_10965 (I188803,I134705,I134708);
nand I_10966 (I188820,I188803,I134720);
nor I_10967 (I188837,I188786,I134705);
nand I_10968 (I188854,I188837,I134726);
not I_10969 (I188871,I188854);
not I_10970 (I188888,I134705);
nor I_10971 (I188758,I188854,I188888);
not I_10972 (I188919,I188888);
nand I_10973 (I188743,I188854,I188919);
not I_10974 (I188950,I134729);
nor I_10975 (I188967,I188950,I134711);
and I_10976 (I188984,I188967,I134714);
or I_10977 (I189001,I188984,I134735);
DFFARX1 I_10978  ( .D(I189001), .CLK(I2350), .RSTB(I188769), .Q(I189018) );
nor I_10979 (I189035,I189018,I188871);
DFFARX1 I_10980  ( .D(I189018), .CLK(I2350), .RSTB(I188769), .Q(I189052) );
not I_10981 (I188740,I189052);
nand I_10982 (I189083,I188786,I134729);
and I_10983 (I189100,I189083,I189035);
DFFARX1 I_10984  ( .D(I189083), .CLK(I2350), .RSTB(I188769), .Q(I188737) );
DFFARX1 I_10985  ( .D(I134717), .CLK(I2350), .RSTB(I188769), .Q(I189131) );
nor I_10986 (I189148,I189131,I188854);
nand I_10987 (I188755,I189018,I189148);
nor I_10988 (I189179,I189131,I188919);
not I_10989 (I188752,I189131);
nand I_10990 (I189210,I189131,I188820);
and I_10991 (I189227,I188888,I189210);
DFFARX1 I_10992  ( .D(I189227), .CLK(I2350), .RSTB(I188769), .Q(I188731) );
DFFARX1 I_10993  ( .D(I189131), .CLK(I2350), .RSTB(I188769), .Q(I188734) );
DFFARX1 I_10994  ( .D(I134723), .CLK(I2350), .RSTB(I188769), .Q(I189272) );
not I_10995 (I189289,I189272);
nand I_10996 (I189306,I189289,I188854);
and I_10997 (I189323,I189083,I189306);
DFFARX1 I_10998  ( .D(I189323), .CLK(I2350), .RSTB(I188769), .Q(I188761) );
or I_10999 (I189354,I189289,I189100);
DFFARX1 I_11000  ( .D(I189354), .CLK(I2350), .RSTB(I188769), .Q(I188746) );
nand I_11001 (I188749,I189289,I189179);
not I_11002 (I189432,I2357);
not I_11003 (I189449,I227605);
nor I_11004 (I189466,I227602,I227620);
nand I_11005 (I189483,I189466,I227623);
nor I_11006 (I189500,I189449,I227602);
nand I_11007 (I189517,I189500,I227608);
not I_11008 (I189534,I189517);
not I_11009 (I189551,I227602);
nor I_11010 (I189421,I189517,I189551);
not I_11011 (I189582,I189551);
nand I_11012 (I189406,I189517,I189582);
not I_11013 (I189613,I227617);
nor I_11014 (I189630,I189613,I227599);
and I_11015 (I189647,I189630,I227593);
or I_11016 (I189664,I189647,I227611);
DFFARX1 I_11017  ( .D(I189664), .CLK(I2350), .RSTB(I189432), .Q(I189681) );
nor I_11018 (I189698,I189681,I189534);
DFFARX1 I_11019  ( .D(I189681), .CLK(I2350), .RSTB(I189432), .Q(I189715) );
not I_11020 (I189403,I189715);
nand I_11021 (I189746,I189449,I227617);
and I_11022 (I189763,I189746,I189698);
DFFARX1 I_11023  ( .D(I189746), .CLK(I2350), .RSTB(I189432), .Q(I189400) );
DFFARX1 I_11024  ( .D(I227596), .CLK(I2350), .RSTB(I189432), .Q(I189794) );
nor I_11025 (I189811,I189794,I189517);
nand I_11026 (I189418,I189681,I189811);
nor I_11027 (I189842,I189794,I189582);
not I_11028 (I189415,I189794);
nand I_11029 (I189873,I189794,I189483);
and I_11030 (I189890,I189551,I189873);
DFFARX1 I_11031  ( .D(I189890), .CLK(I2350), .RSTB(I189432), .Q(I189394) );
DFFARX1 I_11032  ( .D(I189794), .CLK(I2350), .RSTB(I189432), .Q(I189397) );
DFFARX1 I_11033  ( .D(I227614), .CLK(I2350), .RSTB(I189432), .Q(I189935) );
not I_11034 (I189952,I189935);
nand I_11035 (I189969,I189952,I189517);
and I_11036 (I189986,I189746,I189969);
DFFARX1 I_11037  ( .D(I189986), .CLK(I2350), .RSTB(I189432), .Q(I189424) );
or I_11038 (I190017,I189952,I189763);
DFFARX1 I_11039  ( .D(I190017), .CLK(I2350), .RSTB(I189432), .Q(I189409) );
nand I_11040 (I189412,I189952,I189842);
not I_11041 (I190095,I2357);
not I_11042 (I190112,I355881);
nor I_11043 (I190129,I355899,I355890);
nand I_11044 (I190146,I190129,I355896);
nor I_11045 (I190163,I190112,I355899);
nand I_11046 (I190180,I190163,I355902);
not I_11047 (I190197,I190180);
not I_11048 (I190214,I355899);
nor I_11049 (I190084,I190180,I190214);
not I_11050 (I190245,I190214);
nand I_11051 (I190069,I190180,I190245);
not I_11052 (I190276,I355878);
nor I_11053 (I190293,I190276,I355893);
and I_11054 (I190310,I190293,I355875);
or I_11055 (I190327,I190310,I355884);
DFFARX1 I_11056  ( .D(I190327), .CLK(I2350), .RSTB(I190095), .Q(I190344) );
nor I_11057 (I190361,I190344,I190197);
DFFARX1 I_11058  ( .D(I190344), .CLK(I2350), .RSTB(I190095), .Q(I190378) );
not I_11059 (I190066,I190378);
nand I_11060 (I190409,I190112,I355878);
and I_11061 (I190426,I190409,I190361);
DFFARX1 I_11062  ( .D(I190409), .CLK(I2350), .RSTB(I190095), .Q(I190063) );
DFFARX1 I_11063  ( .D(I355887), .CLK(I2350), .RSTB(I190095), .Q(I190457) );
nor I_11064 (I190474,I190457,I190180);
nand I_11065 (I190081,I190344,I190474);
nor I_11066 (I190505,I190457,I190245);
not I_11067 (I190078,I190457);
nand I_11068 (I190536,I190457,I190146);
and I_11069 (I190553,I190214,I190536);
DFFARX1 I_11070  ( .D(I190553), .CLK(I2350), .RSTB(I190095), .Q(I190057) );
DFFARX1 I_11071  ( .D(I190457), .CLK(I2350), .RSTB(I190095), .Q(I190060) );
DFFARX1 I_11072  ( .D(I355905), .CLK(I2350), .RSTB(I190095), .Q(I190598) );
not I_11073 (I190615,I190598);
nand I_11074 (I190632,I190615,I190180);
and I_11075 (I190649,I190409,I190632);
DFFARX1 I_11076  ( .D(I190649), .CLK(I2350), .RSTB(I190095), .Q(I190087) );
or I_11077 (I190680,I190615,I190426);
DFFARX1 I_11078  ( .D(I190680), .CLK(I2350), .RSTB(I190095), .Q(I190072) );
nand I_11079 (I190075,I190615,I190505);
not I_11080 (I190758,I2357);
not I_11081 (I190775,I10793);
nor I_11082 (I190792,I10799,I10802);
nand I_11083 (I190809,I190792,I10778);
nor I_11084 (I190826,I190775,I10799);
nand I_11085 (I190843,I190826,I10787);
not I_11086 (I190860,I190843);
not I_11087 (I190877,I10799);
nor I_11088 (I190747,I190843,I190877);
not I_11089 (I190908,I190877);
nand I_11090 (I190732,I190843,I190908);
not I_11091 (I190939,I10781);
nor I_11092 (I190956,I190939,I10805);
and I_11093 (I190973,I190956,I10775);
or I_11094 (I190990,I190973,I10784);
DFFARX1 I_11095  ( .D(I190990), .CLK(I2350), .RSTB(I190758), .Q(I191007) );
nor I_11096 (I191024,I191007,I190860);
DFFARX1 I_11097  ( .D(I191007), .CLK(I2350), .RSTB(I190758), .Q(I191041) );
not I_11098 (I190729,I191041);
nand I_11099 (I191072,I190775,I10781);
and I_11100 (I191089,I191072,I191024);
DFFARX1 I_11101  ( .D(I191072), .CLK(I2350), .RSTB(I190758), .Q(I190726) );
DFFARX1 I_11102  ( .D(I10790), .CLK(I2350), .RSTB(I190758), .Q(I191120) );
nor I_11103 (I191137,I191120,I190843);
nand I_11104 (I190744,I191007,I191137);
nor I_11105 (I191168,I191120,I190908);
not I_11106 (I190741,I191120);
nand I_11107 (I191199,I191120,I190809);
and I_11108 (I191216,I190877,I191199);
DFFARX1 I_11109  ( .D(I191216), .CLK(I2350), .RSTB(I190758), .Q(I190720) );
DFFARX1 I_11110  ( .D(I191120), .CLK(I2350), .RSTB(I190758), .Q(I190723) );
DFFARX1 I_11111  ( .D(I10796), .CLK(I2350), .RSTB(I190758), .Q(I191261) );
not I_11112 (I191278,I191261);
nand I_11113 (I191295,I191278,I190843);
and I_11114 (I191312,I191072,I191295);
DFFARX1 I_11115  ( .D(I191312), .CLK(I2350), .RSTB(I190758), .Q(I190750) );
or I_11116 (I191343,I191278,I191089);
DFFARX1 I_11117  ( .D(I191343), .CLK(I2350), .RSTB(I190758), .Q(I190735) );
nand I_11118 (I190738,I191278,I191168);
not I_11119 (I191421,I2357);
not I_11120 (I191438,I390295);
nor I_11121 (I191455,I390286,I390292);
nand I_11122 (I191472,I191455,I390304);
nor I_11123 (I191489,I191438,I390286);
nand I_11124 (I191506,I191489,I390289);
not I_11125 (I191523,I191506);
not I_11126 (I191540,I390286);
nor I_11127 (I191410,I191506,I191540);
not I_11128 (I191571,I191540);
nand I_11129 (I191395,I191506,I191571);
not I_11130 (I191602,I390313);
nor I_11131 (I191619,I191602,I390307);
and I_11132 (I191636,I191619,I390298);
or I_11133 (I191653,I191636,I390283);
DFFARX1 I_11134  ( .D(I191653), .CLK(I2350), .RSTB(I191421), .Q(I191670) );
nor I_11135 (I191687,I191670,I191523);
DFFARX1 I_11136  ( .D(I191670), .CLK(I2350), .RSTB(I191421), .Q(I191704) );
not I_11137 (I191392,I191704);
nand I_11138 (I191735,I191438,I390313);
and I_11139 (I191752,I191735,I191687);
DFFARX1 I_11140  ( .D(I191735), .CLK(I2350), .RSTB(I191421), .Q(I191389) );
DFFARX1 I_11141  ( .D(I390301), .CLK(I2350), .RSTB(I191421), .Q(I191783) );
nor I_11142 (I191800,I191783,I191506);
nand I_11143 (I191407,I191670,I191800);
nor I_11144 (I191831,I191783,I191571);
not I_11145 (I191404,I191783);
nand I_11146 (I191862,I191783,I191472);
and I_11147 (I191879,I191540,I191862);
DFFARX1 I_11148  ( .D(I191879), .CLK(I2350), .RSTB(I191421), .Q(I191383) );
DFFARX1 I_11149  ( .D(I191783), .CLK(I2350), .RSTB(I191421), .Q(I191386) );
DFFARX1 I_11150  ( .D(I390310), .CLK(I2350), .RSTB(I191421), .Q(I191924) );
not I_11151 (I191941,I191924);
nand I_11152 (I191958,I191941,I191506);
and I_11153 (I191975,I191735,I191958);
DFFARX1 I_11154  ( .D(I191975), .CLK(I2350), .RSTB(I191421), .Q(I191413) );
or I_11155 (I192006,I191941,I191752);
DFFARX1 I_11156  ( .D(I192006), .CLK(I2350), .RSTB(I191421), .Q(I191398) );
nand I_11157 (I191401,I191941,I191831);
not I_11158 (I192084,I2357);
not I_11159 (I192101,I34326);
nor I_11160 (I192118,I34323,I34347);
nand I_11161 (I192135,I192118,I34344);
nor I_11162 (I192152,I192101,I34323);
nand I_11163 (I192169,I192152,I34350);
not I_11164 (I192186,I192169);
not I_11165 (I192203,I34323);
nor I_11166 (I192073,I192169,I192203);
not I_11167 (I192234,I192203);
nand I_11168 (I192058,I192169,I192234);
not I_11169 (I192265,I34341);
nor I_11170 (I192282,I192265,I34332);
and I_11171 (I192299,I192282,I34329);
or I_11172 (I192316,I192299,I34338);
DFFARX1 I_11173  ( .D(I192316), .CLK(I2350), .RSTB(I192084), .Q(I192333) );
nor I_11174 (I192350,I192333,I192186);
DFFARX1 I_11175  ( .D(I192333), .CLK(I2350), .RSTB(I192084), .Q(I192367) );
not I_11176 (I192055,I192367);
nand I_11177 (I192398,I192101,I34341);
and I_11178 (I192415,I192398,I192350);
DFFARX1 I_11179  ( .D(I192398), .CLK(I2350), .RSTB(I192084), .Q(I192052) );
DFFARX1 I_11180  ( .D(I34320), .CLK(I2350), .RSTB(I192084), .Q(I192446) );
nor I_11181 (I192463,I192446,I192169);
nand I_11182 (I192070,I192333,I192463);
nor I_11183 (I192494,I192446,I192234);
not I_11184 (I192067,I192446);
nand I_11185 (I192525,I192446,I192135);
and I_11186 (I192542,I192203,I192525);
DFFARX1 I_11187  ( .D(I192542), .CLK(I2350), .RSTB(I192084), .Q(I192046) );
DFFARX1 I_11188  ( .D(I192446), .CLK(I2350), .RSTB(I192084), .Q(I192049) );
DFFARX1 I_11189  ( .D(I34335), .CLK(I2350), .RSTB(I192084), .Q(I192587) );
not I_11190 (I192604,I192587);
nand I_11191 (I192621,I192604,I192169);
and I_11192 (I192638,I192398,I192621);
DFFARX1 I_11193  ( .D(I192638), .CLK(I2350), .RSTB(I192084), .Q(I192076) );
or I_11194 (I192669,I192604,I192415);
DFFARX1 I_11195  ( .D(I192669), .CLK(I2350), .RSTB(I192084), .Q(I192061) );
nand I_11196 (I192064,I192604,I192494);
not I_11197 (I192747,I2357);
not I_11198 (I192764,I4052);
nor I_11199 (I192781,I4067,I4061);
nand I_11200 (I192798,I192781,I4070);
nor I_11201 (I192815,I192764,I4067);
nand I_11202 (I192832,I192815,I4046);
DFFARX1 I_11203  ( .D(I192832), .CLK(I2350), .RSTB(I192747), .Q(I192849) );
not I_11204 (I192718,I192849);
not I_11205 (I192880,I4067);
not I_11206 (I192897,I192880);
not I_11207 (I192914,I4043);
nor I_11208 (I192931,I192914,I4058);
and I_11209 (I192948,I192931,I4064);
or I_11210 (I192965,I192948,I4073);
DFFARX1 I_11211  ( .D(I192965), .CLK(I2350), .RSTB(I192747), .Q(I192982) );
DFFARX1 I_11212  ( .D(I192982), .CLK(I2350), .RSTB(I192747), .Q(I192715) );
DFFARX1 I_11213  ( .D(I192982), .CLK(I2350), .RSTB(I192747), .Q(I193013) );
DFFARX1 I_11214  ( .D(I192982), .CLK(I2350), .RSTB(I192747), .Q(I192709) );
nand I_11215 (I193044,I192764,I4043);
nand I_11216 (I193061,I193044,I192798);
and I_11217 (I193078,I192880,I193061);
DFFARX1 I_11218  ( .D(I193078), .CLK(I2350), .RSTB(I192747), .Q(I192739) );
and I_11219 (I192712,I193044,I193013);
DFFARX1 I_11220  ( .D(I4055), .CLK(I2350), .RSTB(I192747), .Q(I193123) );
nor I_11221 (I192736,I193123,I193044);
nor I_11222 (I193154,I193123,I192798);
nand I_11223 (I192733,I192832,I193154);
not I_11224 (I192730,I193123);
DFFARX1 I_11225  ( .D(I4049), .CLK(I2350), .RSTB(I192747), .Q(I193199) );
not I_11226 (I193216,I193199);
nor I_11227 (I193233,I193216,I192897);
and I_11228 (I193250,I193123,I193233);
or I_11229 (I193267,I193044,I193250);
DFFARX1 I_11230  ( .D(I193267), .CLK(I2350), .RSTB(I192747), .Q(I192724) );
not I_11231 (I193298,I193216);
nor I_11232 (I193315,I193123,I193298);
nand I_11233 (I192727,I193216,I193315);
nand I_11234 (I192721,I192880,I193298);
not I_11235 (I193393,I2357);
not I_11236 (I193410,I159583);
nor I_11237 (I193427,I159562,I159574);
nand I_11238 (I193444,I193427,I159577);
nor I_11239 (I193461,I193410,I159562);
nand I_11240 (I193478,I193461,I159559);
DFFARX1 I_11241  ( .D(I193478), .CLK(I2350), .RSTB(I193393), .Q(I193495) );
not I_11242 (I193364,I193495);
not I_11243 (I193526,I159562);
not I_11244 (I193543,I193526);
not I_11245 (I193560,I159580);
nor I_11246 (I193577,I193560,I159571);
and I_11247 (I193594,I193577,I159565);
or I_11248 (I193611,I193594,I159589);
DFFARX1 I_11249  ( .D(I193611), .CLK(I2350), .RSTB(I193393), .Q(I193628) );
DFFARX1 I_11250  ( .D(I193628), .CLK(I2350), .RSTB(I193393), .Q(I193361) );
DFFARX1 I_11251  ( .D(I193628), .CLK(I2350), .RSTB(I193393), .Q(I193659) );
DFFARX1 I_11252  ( .D(I193628), .CLK(I2350), .RSTB(I193393), .Q(I193355) );
nand I_11253 (I193690,I193410,I159580);
nand I_11254 (I193707,I193690,I193444);
and I_11255 (I193724,I193526,I193707);
DFFARX1 I_11256  ( .D(I193724), .CLK(I2350), .RSTB(I193393), .Q(I193385) );
and I_11257 (I193358,I193690,I193659);
DFFARX1 I_11258  ( .D(I159586), .CLK(I2350), .RSTB(I193393), .Q(I193769) );
nor I_11259 (I193382,I193769,I193690);
nor I_11260 (I193800,I193769,I193444);
nand I_11261 (I193379,I193478,I193800);
not I_11262 (I193376,I193769);
DFFARX1 I_11263  ( .D(I159568), .CLK(I2350), .RSTB(I193393), .Q(I193845) );
not I_11264 (I193862,I193845);
nor I_11265 (I193879,I193862,I193543);
and I_11266 (I193896,I193769,I193879);
or I_11267 (I193913,I193690,I193896);
DFFARX1 I_11268  ( .D(I193913), .CLK(I2350), .RSTB(I193393), .Q(I193370) );
not I_11269 (I193944,I193862);
nor I_11270 (I193961,I193769,I193944);
nand I_11271 (I193373,I193862,I193961);
nand I_11272 (I193367,I193526,I193944);
not I_11273 (I194039,I2357);
not I_11274 (I194056,I321315);
nor I_11275 (I194073,I321303,I321312);
nand I_11276 (I194090,I194073,I321327);
nor I_11277 (I194107,I194056,I321303);
nand I_11278 (I194124,I194107,I321309);
DFFARX1 I_11279  ( .D(I194124), .CLK(I2350), .RSTB(I194039), .Q(I194141) );
not I_11280 (I194010,I194141);
not I_11281 (I194172,I321303);
not I_11282 (I194189,I194172);
not I_11283 (I194206,I321297);
nor I_11284 (I194223,I194206,I321318);
and I_11285 (I194240,I194223,I321300);
or I_11286 (I194257,I194240,I321306);
DFFARX1 I_11287  ( .D(I194257), .CLK(I2350), .RSTB(I194039), .Q(I194274) );
DFFARX1 I_11288  ( .D(I194274), .CLK(I2350), .RSTB(I194039), .Q(I194007) );
DFFARX1 I_11289  ( .D(I194274), .CLK(I2350), .RSTB(I194039), .Q(I194305) );
DFFARX1 I_11290  ( .D(I194274), .CLK(I2350), .RSTB(I194039), .Q(I194001) );
nand I_11291 (I194336,I194056,I321297);
nand I_11292 (I194353,I194336,I194090);
and I_11293 (I194370,I194172,I194353);
DFFARX1 I_11294  ( .D(I194370), .CLK(I2350), .RSTB(I194039), .Q(I194031) );
and I_11295 (I194004,I194336,I194305);
DFFARX1 I_11296  ( .D(I321324), .CLK(I2350), .RSTB(I194039), .Q(I194415) );
nor I_11297 (I194028,I194415,I194336);
nor I_11298 (I194446,I194415,I194090);
nand I_11299 (I194025,I194124,I194446);
not I_11300 (I194022,I194415);
DFFARX1 I_11301  ( .D(I321321), .CLK(I2350), .RSTB(I194039), .Q(I194491) );
not I_11302 (I194508,I194491);
nor I_11303 (I194525,I194508,I194189);
and I_11304 (I194542,I194415,I194525);
or I_11305 (I194559,I194336,I194542);
DFFARX1 I_11306  ( .D(I194559), .CLK(I2350), .RSTB(I194039), .Q(I194016) );
not I_11307 (I194590,I194508);
nor I_11308 (I194607,I194415,I194590);
nand I_11309 (I194019,I194508,I194607);
nand I_11310 (I194013,I194172,I194590);
not I_11311 (I194685,I2357);
not I_11312 (I194702,I20882);
nor I_11313 (I194719,I20897,I20891);
nand I_11314 (I194736,I194719,I20900);
nor I_11315 (I194753,I194702,I20897);
nand I_11316 (I194770,I194753,I20876);
DFFARX1 I_11317  ( .D(I194770), .CLK(I2350), .RSTB(I194685), .Q(I194787) );
not I_11318 (I194656,I194787);
not I_11319 (I194818,I20897);
not I_11320 (I194835,I194818);
not I_11321 (I194852,I20873);
nor I_11322 (I194869,I194852,I20888);
and I_11323 (I194886,I194869,I20894);
or I_11324 (I194903,I194886,I20903);
DFFARX1 I_11325  ( .D(I194903), .CLK(I2350), .RSTB(I194685), .Q(I194920) );
DFFARX1 I_11326  ( .D(I194920), .CLK(I2350), .RSTB(I194685), .Q(I194653) );
DFFARX1 I_11327  ( .D(I194920), .CLK(I2350), .RSTB(I194685), .Q(I194951) );
DFFARX1 I_11328  ( .D(I194920), .CLK(I2350), .RSTB(I194685), .Q(I194647) );
nand I_11329 (I194982,I194702,I20873);
nand I_11330 (I194999,I194982,I194736);
and I_11331 (I195016,I194818,I194999);
DFFARX1 I_11332  ( .D(I195016), .CLK(I2350), .RSTB(I194685), .Q(I194677) );
and I_11333 (I194650,I194982,I194951);
DFFARX1 I_11334  ( .D(I20885), .CLK(I2350), .RSTB(I194685), .Q(I195061) );
nor I_11335 (I194674,I195061,I194982);
nor I_11336 (I195092,I195061,I194736);
nand I_11337 (I194671,I194770,I195092);
not I_11338 (I194668,I195061);
DFFARX1 I_11339  ( .D(I20879), .CLK(I2350), .RSTB(I194685), .Q(I195137) );
not I_11340 (I195154,I195137);
nor I_11341 (I195171,I195154,I194835);
and I_11342 (I195188,I195061,I195171);
or I_11343 (I195205,I194982,I195188);
DFFARX1 I_11344  ( .D(I195205), .CLK(I2350), .RSTB(I194685), .Q(I194662) );
not I_11345 (I195236,I195154);
nor I_11346 (I195253,I195061,I195236);
nand I_11347 (I194665,I195154,I195253);
nand I_11348 (I194659,I194818,I195236);
not I_11349 (I195331,I2357);
not I_11350 (I195348,I304646);
nor I_11351 (I195365,I304658,I304652);
nand I_11352 (I195382,I195365,I304637);
nor I_11353 (I195399,I195348,I304658);
nand I_11354 (I195416,I195399,I304664);
DFFARX1 I_11355  ( .D(I195416), .CLK(I2350), .RSTB(I195331), .Q(I195433) );
not I_11356 (I195302,I195433);
not I_11357 (I195464,I304658);
not I_11358 (I195481,I195464);
not I_11359 (I195498,I304661);
nor I_11360 (I195515,I195498,I304643);
and I_11361 (I195532,I195515,I304640);
or I_11362 (I195549,I195532,I304667);
DFFARX1 I_11363  ( .D(I195549), .CLK(I2350), .RSTB(I195331), .Q(I195566) );
DFFARX1 I_11364  ( .D(I195566), .CLK(I2350), .RSTB(I195331), .Q(I195299) );
DFFARX1 I_11365  ( .D(I195566), .CLK(I2350), .RSTB(I195331), .Q(I195597) );
DFFARX1 I_11366  ( .D(I195566), .CLK(I2350), .RSTB(I195331), .Q(I195293) );
nand I_11367 (I195628,I195348,I304661);
nand I_11368 (I195645,I195628,I195382);
and I_11369 (I195662,I195464,I195645);
DFFARX1 I_11370  ( .D(I195662), .CLK(I2350), .RSTB(I195331), .Q(I195323) );
and I_11371 (I195296,I195628,I195597);
DFFARX1 I_11372  ( .D(I304655), .CLK(I2350), .RSTB(I195331), .Q(I195707) );
nor I_11373 (I195320,I195707,I195628);
nor I_11374 (I195738,I195707,I195382);
nand I_11375 (I195317,I195416,I195738);
not I_11376 (I195314,I195707);
DFFARX1 I_11377  ( .D(I304649), .CLK(I2350), .RSTB(I195331), .Q(I195783) );
not I_11378 (I195800,I195783);
nor I_11379 (I195817,I195800,I195481);
and I_11380 (I195834,I195707,I195817);
or I_11381 (I195851,I195628,I195834);
DFFARX1 I_11382  ( .D(I195851), .CLK(I2350), .RSTB(I195331), .Q(I195308) );
not I_11383 (I195882,I195800);
nor I_11384 (I195899,I195707,I195882);
nand I_11385 (I195311,I195800,I195899);
nand I_11386 (I195305,I195464,I195882);
not I_11387 (I195977,I2357);
not I_11388 (I195994,I76977);
nor I_11389 (I196011,I76968,I76959);
nand I_11390 (I196028,I196011,I76974);
nor I_11391 (I196045,I195994,I76968);
nand I_11392 (I196062,I196045,I76971);
DFFARX1 I_11393  ( .D(I196062), .CLK(I2350), .RSTB(I195977), .Q(I196079) );
not I_11394 (I195948,I196079);
not I_11395 (I196110,I76968);
not I_11396 (I196127,I196110);
not I_11397 (I196144,I76980);
nor I_11398 (I196161,I196144,I76965);
and I_11399 (I196178,I196161,I76983);
or I_11400 (I196195,I196178,I76956);
DFFARX1 I_11401  ( .D(I196195), .CLK(I2350), .RSTB(I195977), .Q(I196212) );
DFFARX1 I_11402  ( .D(I196212), .CLK(I2350), .RSTB(I195977), .Q(I195945) );
DFFARX1 I_11403  ( .D(I196212), .CLK(I2350), .RSTB(I195977), .Q(I196243) );
DFFARX1 I_11404  ( .D(I196212), .CLK(I2350), .RSTB(I195977), .Q(I195939) );
nand I_11405 (I196274,I195994,I76980);
nand I_11406 (I196291,I196274,I196028);
and I_11407 (I196308,I196110,I196291);
DFFARX1 I_11408  ( .D(I196308), .CLK(I2350), .RSTB(I195977), .Q(I195969) );
and I_11409 (I195942,I196274,I196243);
DFFARX1 I_11410  ( .D(I76986), .CLK(I2350), .RSTB(I195977), .Q(I196353) );
nor I_11411 (I195966,I196353,I196274);
nor I_11412 (I196384,I196353,I196028);
nand I_11413 (I195963,I196062,I196384);
not I_11414 (I195960,I196353);
DFFARX1 I_11415  ( .D(I76962), .CLK(I2350), .RSTB(I195977), .Q(I196429) );
not I_11416 (I196446,I196429);
nor I_11417 (I196463,I196446,I196127);
and I_11418 (I196480,I196353,I196463);
or I_11419 (I196497,I196274,I196480);
DFFARX1 I_11420  ( .D(I196497), .CLK(I2350), .RSTB(I195977), .Q(I195954) );
not I_11421 (I196528,I196446);
nor I_11422 (I196545,I196353,I196528);
nand I_11423 (I195957,I196446,I196545);
nand I_11424 (I195951,I196110,I196528);
not I_11425 (I196623,I2357);
not I_11426 (I196640,I112557);
nor I_11427 (I196657,I112578,I112560);
nand I_11428 (I196674,I196657,I112584);
nor I_11429 (I196691,I196640,I112578);
nand I_11430 (I196708,I196691,I112581);
DFFARX1 I_11431  ( .D(I196708), .CLK(I2350), .RSTB(I196623), .Q(I196725) );
not I_11432 (I196594,I196725);
not I_11433 (I196756,I112578);
not I_11434 (I196773,I196756);
not I_11435 (I196790,I112575);
nor I_11436 (I196807,I196790,I112554);
and I_11437 (I196824,I196807,I112566);
or I_11438 (I196841,I196824,I112563);
DFFARX1 I_11439  ( .D(I196841), .CLK(I2350), .RSTB(I196623), .Q(I196858) );
DFFARX1 I_11440  ( .D(I196858), .CLK(I2350), .RSTB(I196623), .Q(I196591) );
DFFARX1 I_11441  ( .D(I196858), .CLK(I2350), .RSTB(I196623), .Q(I196889) );
DFFARX1 I_11442  ( .D(I196858), .CLK(I2350), .RSTB(I196623), .Q(I196585) );
nand I_11443 (I196920,I196640,I112575);
nand I_11444 (I196937,I196920,I196674);
and I_11445 (I196954,I196756,I196937);
DFFARX1 I_11446  ( .D(I196954), .CLK(I2350), .RSTB(I196623), .Q(I196615) );
and I_11447 (I196588,I196920,I196889);
DFFARX1 I_11448  ( .D(I112569), .CLK(I2350), .RSTB(I196623), .Q(I196999) );
nor I_11449 (I196612,I196999,I196920);
nor I_11450 (I197030,I196999,I196674);
nand I_11451 (I196609,I196708,I197030);
not I_11452 (I196606,I196999);
DFFARX1 I_11453  ( .D(I112572), .CLK(I2350), .RSTB(I196623), .Q(I197075) );
not I_11454 (I197092,I197075);
nor I_11455 (I197109,I197092,I196773);
and I_11456 (I197126,I196999,I197109);
or I_11457 (I197143,I196920,I197126);
DFFARX1 I_11458  ( .D(I197143), .CLK(I2350), .RSTB(I196623), .Q(I196600) );
not I_11459 (I197174,I197092);
nor I_11460 (I197191,I196999,I197174);
nand I_11461 (I196603,I197092,I197191);
nand I_11462 (I196597,I196756,I197174);
not I_11463 (I197269,I2357);
not I_11464 (I197286,I261438);
nor I_11465 (I197303,I261441,I261423);
nand I_11466 (I197320,I197303,I261450);
nor I_11467 (I197337,I197286,I261441);
nand I_11468 (I197354,I197337,I261429);
DFFARX1 I_11469  ( .D(I197354), .CLK(I2350), .RSTB(I197269), .Q(I197371) );
not I_11470 (I197240,I197371);
not I_11471 (I197402,I261441);
not I_11472 (I197419,I197402);
not I_11473 (I197436,I261435);
nor I_11474 (I197453,I197436,I261447);
and I_11475 (I197470,I197453,I261453);
or I_11476 (I197487,I197470,I261432);
DFFARX1 I_11477  ( .D(I197487), .CLK(I2350), .RSTB(I197269), .Q(I197504) );
DFFARX1 I_11478  ( .D(I197504), .CLK(I2350), .RSTB(I197269), .Q(I197237) );
DFFARX1 I_11479  ( .D(I197504), .CLK(I2350), .RSTB(I197269), .Q(I197535) );
DFFARX1 I_11480  ( .D(I197504), .CLK(I2350), .RSTB(I197269), .Q(I197231) );
nand I_11481 (I197566,I197286,I261435);
nand I_11482 (I197583,I197566,I197320);
and I_11483 (I197600,I197402,I197583);
DFFARX1 I_11484  ( .D(I197600), .CLK(I2350), .RSTB(I197269), .Q(I197261) );
and I_11485 (I197234,I197566,I197535);
DFFARX1 I_11486  ( .D(I261444), .CLK(I2350), .RSTB(I197269), .Q(I197645) );
nor I_11487 (I197258,I197645,I197566);
nor I_11488 (I197676,I197645,I197320);
nand I_11489 (I197255,I197354,I197676);
not I_11490 (I197252,I197645);
DFFARX1 I_11491  ( .D(I261426), .CLK(I2350), .RSTB(I197269), .Q(I197721) );
not I_11492 (I197738,I197721);
nor I_11493 (I197755,I197738,I197419);
and I_11494 (I197772,I197645,I197755);
or I_11495 (I197789,I197566,I197772);
DFFARX1 I_11496  ( .D(I197789), .CLK(I2350), .RSTB(I197269), .Q(I197246) );
not I_11497 (I197820,I197738);
nor I_11498 (I197837,I197645,I197820);
nand I_11499 (I197249,I197738,I197837);
nand I_11500 (I197243,I197402,I197820);
not I_11501 (I197915,I2357);
not I_11502 (I197932,I15272);
nor I_11503 (I197949,I15287,I15281);
nand I_11504 (I197966,I197949,I15290);
nor I_11505 (I197983,I197932,I15287);
nand I_11506 (I198000,I197983,I15266);
DFFARX1 I_11507  ( .D(I198000), .CLK(I2350), .RSTB(I197915), .Q(I198017) );
not I_11508 (I197886,I198017);
not I_11509 (I198048,I15287);
not I_11510 (I198065,I198048);
not I_11511 (I198082,I15263);
nor I_11512 (I198099,I198082,I15278);
and I_11513 (I198116,I198099,I15284);
or I_11514 (I198133,I198116,I15293);
DFFARX1 I_11515  ( .D(I198133), .CLK(I2350), .RSTB(I197915), .Q(I198150) );
DFFARX1 I_11516  ( .D(I198150), .CLK(I2350), .RSTB(I197915), .Q(I197883) );
DFFARX1 I_11517  ( .D(I198150), .CLK(I2350), .RSTB(I197915), .Q(I198181) );
DFFARX1 I_11518  ( .D(I198150), .CLK(I2350), .RSTB(I197915), .Q(I197877) );
nand I_11519 (I198212,I197932,I15263);
nand I_11520 (I198229,I198212,I197966);
and I_11521 (I198246,I198048,I198229);
DFFARX1 I_11522  ( .D(I198246), .CLK(I2350), .RSTB(I197915), .Q(I197907) );
and I_11523 (I197880,I198212,I198181);
DFFARX1 I_11524  ( .D(I15275), .CLK(I2350), .RSTB(I197915), .Q(I198291) );
nor I_11525 (I197904,I198291,I198212);
nor I_11526 (I198322,I198291,I197966);
nand I_11527 (I197901,I198000,I198322);
not I_11528 (I197898,I198291);
DFFARX1 I_11529  ( .D(I15269), .CLK(I2350), .RSTB(I197915), .Q(I198367) );
not I_11530 (I198384,I198367);
nor I_11531 (I198401,I198384,I198065);
and I_11532 (I198418,I198291,I198401);
or I_11533 (I198435,I198212,I198418);
DFFARX1 I_11534  ( .D(I198435), .CLK(I2350), .RSTB(I197915), .Q(I197892) );
not I_11535 (I198466,I198384);
nor I_11536 (I198483,I198291,I198466);
nand I_11537 (I197895,I198384,I198483);
nand I_11538 (I197889,I198048,I198466);
not I_11539 (I198561,I2357);
not I_11540 (I198578,I369105);
nor I_11541 (I198595,I369102,I369087);
nand I_11542 (I198612,I198595,I369096);
nor I_11543 (I198629,I198578,I369102);
nand I_11544 (I198646,I198629,I369111);
DFFARX1 I_11545  ( .D(I198646), .CLK(I2350), .RSTB(I198561), .Q(I198663) );
not I_11546 (I198532,I198663);
not I_11547 (I198694,I369102);
not I_11548 (I198711,I198694);
not I_11549 (I198728,I369084);
nor I_11550 (I198745,I198728,I369090);
and I_11551 (I198762,I198745,I369114);
or I_11552 (I198779,I198762,I369108);
DFFARX1 I_11553  ( .D(I198779), .CLK(I2350), .RSTB(I198561), .Q(I198796) );
DFFARX1 I_11554  ( .D(I198796), .CLK(I2350), .RSTB(I198561), .Q(I198529) );
DFFARX1 I_11555  ( .D(I198796), .CLK(I2350), .RSTB(I198561), .Q(I198827) );
DFFARX1 I_11556  ( .D(I198796), .CLK(I2350), .RSTB(I198561), .Q(I198523) );
nand I_11557 (I198858,I198578,I369084);
nand I_11558 (I198875,I198858,I198612);
and I_11559 (I198892,I198694,I198875);
DFFARX1 I_11560  ( .D(I198892), .CLK(I2350), .RSTB(I198561), .Q(I198553) );
and I_11561 (I198526,I198858,I198827);
DFFARX1 I_11562  ( .D(I369093), .CLK(I2350), .RSTB(I198561), .Q(I198937) );
nor I_11563 (I198550,I198937,I198858);
nor I_11564 (I198968,I198937,I198612);
nand I_11565 (I198547,I198646,I198968);
not I_11566 (I198544,I198937);
DFFARX1 I_11567  ( .D(I369099), .CLK(I2350), .RSTB(I198561), .Q(I199013) );
not I_11568 (I199030,I199013);
nor I_11569 (I199047,I199030,I198711);
and I_11570 (I199064,I198937,I199047);
or I_11571 (I199081,I198858,I199064);
DFFARX1 I_11572  ( .D(I199081), .CLK(I2350), .RSTB(I198561), .Q(I198538) );
not I_11573 (I199112,I199030);
nor I_11574 (I199129,I198937,I199112);
nand I_11575 (I198541,I199030,I199129);
nand I_11576 (I198535,I198694,I199112);
not I_11577 (I199207,I2357);
not I_11578 (I199224,I124001);
nor I_11579 (I199241,I124007,I124004);
nand I_11580 (I199258,I199241,I123998);
nor I_11581 (I199275,I199224,I124007);
nand I_11582 (I199292,I199275,I124022);
DFFARX1 I_11583  ( .D(I199292), .CLK(I2350), .RSTB(I199207), .Q(I199309) );
not I_11584 (I199178,I199309);
not I_11585 (I199340,I124007);
not I_11586 (I199357,I199340);
not I_11587 (I199374,I124019);
nor I_11588 (I199391,I199374,I124010);
and I_11589 (I199408,I199391,I123995);
or I_11590 (I199425,I199408,I124016);
DFFARX1 I_11591  ( .D(I199425), .CLK(I2350), .RSTB(I199207), .Q(I199442) );
DFFARX1 I_11592  ( .D(I199442), .CLK(I2350), .RSTB(I199207), .Q(I199175) );
DFFARX1 I_11593  ( .D(I199442), .CLK(I2350), .RSTB(I199207), .Q(I199473) );
DFFARX1 I_11594  ( .D(I199442), .CLK(I2350), .RSTB(I199207), .Q(I199169) );
nand I_11595 (I199504,I199224,I124019);
nand I_11596 (I199521,I199504,I199258);
and I_11597 (I199538,I199340,I199521);
DFFARX1 I_11598  ( .D(I199538), .CLK(I2350), .RSTB(I199207), .Q(I199199) );
and I_11599 (I199172,I199504,I199473);
DFFARX1 I_11600  ( .D(I124013), .CLK(I2350), .RSTB(I199207), .Q(I199583) );
nor I_11601 (I199196,I199583,I199504);
nor I_11602 (I199614,I199583,I199258);
nand I_11603 (I199193,I199292,I199614);
not I_11604 (I199190,I199583);
DFFARX1 I_11605  ( .D(I124025), .CLK(I2350), .RSTB(I199207), .Q(I199659) );
not I_11606 (I199676,I199659);
nor I_11607 (I199693,I199676,I199357);
and I_11608 (I199710,I199583,I199693);
or I_11609 (I199727,I199504,I199710);
DFFARX1 I_11610  ( .D(I199727), .CLK(I2350), .RSTB(I199207), .Q(I199184) );
not I_11611 (I199758,I199676);
nor I_11612 (I199775,I199583,I199758);
nand I_11613 (I199187,I199676,I199775);
nand I_11614 (I199181,I199340,I199758);
not I_11615 (I199853,I2357);
not I_11616 (I199870,I324885);
nor I_11617 (I199887,I324873,I324882);
nand I_11618 (I199904,I199887,I324897);
nor I_11619 (I199921,I199870,I324873);
nand I_11620 (I199938,I199921,I324879);
DFFARX1 I_11621  ( .D(I199938), .CLK(I2350), .RSTB(I199853), .Q(I199955) );
not I_11622 (I199824,I199955);
not I_11623 (I199986,I324873);
not I_11624 (I200003,I199986);
not I_11625 (I200020,I324867);
nor I_11626 (I200037,I200020,I324888);
and I_11627 (I200054,I200037,I324870);
or I_11628 (I200071,I200054,I324876);
DFFARX1 I_11629  ( .D(I200071), .CLK(I2350), .RSTB(I199853), .Q(I200088) );
DFFARX1 I_11630  ( .D(I200088), .CLK(I2350), .RSTB(I199853), .Q(I199821) );
DFFARX1 I_11631  ( .D(I200088), .CLK(I2350), .RSTB(I199853), .Q(I200119) );
DFFARX1 I_11632  ( .D(I200088), .CLK(I2350), .RSTB(I199853), .Q(I199815) );
nand I_11633 (I200150,I199870,I324867);
nand I_11634 (I200167,I200150,I199904);
and I_11635 (I200184,I199986,I200167);
DFFARX1 I_11636  ( .D(I200184), .CLK(I2350), .RSTB(I199853), .Q(I199845) );
and I_11637 (I199818,I200150,I200119);
DFFARX1 I_11638  ( .D(I324894), .CLK(I2350), .RSTB(I199853), .Q(I200229) );
nor I_11639 (I199842,I200229,I200150);
nor I_11640 (I200260,I200229,I199904);
nand I_11641 (I199839,I199938,I200260);
not I_11642 (I199836,I200229);
DFFARX1 I_11643  ( .D(I324891), .CLK(I2350), .RSTB(I199853), .Q(I200305) );
not I_11644 (I200322,I200305);
nor I_11645 (I200339,I200322,I200003);
and I_11646 (I200356,I200229,I200339);
or I_11647 (I200373,I200150,I200356);
DFFARX1 I_11648  ( .D(I200373), .CLK(I2350), .RSTB(I199853), .Q(I199830) );
not I_11649 (I200404,I200322);
nor I_11650 (I200421,I200229,I200404);
nand I_11651 (I199833,I200322,I200421);
nand I_11652 (I199827,I199986,I200404);
not I_11653 (I200499,I2357);
not I_11654 (I200516,I91341);
nor I_11655 (I200533,I91362,I91344);
nand I_11656 (I200550,I200533,I91368);
nor I_11657 (I200567,I200516,I91362);
nand I_11658 (I200584,I200567,I91365);
DFFARX1 I_11659  ( .D(I200584), .CLK(I2350), .RSTB(I200499), .Q(I200601) );
not I_11660 (I200470,I200601);
not I_11661 (I200632,I91362);
not I_11662 (I200649,I200632);
not I_11663 (I200666,I91359);
nor I_11664 (I200683,I200666,I91338);
and I_11665 (I200700,I200683,I91350);
or I_11666 (I200717,I200700,I91347);
DFFARX1 I_11667  ( .D(I200717), .CLK(I2350), .RSTB(I200499), .Q(I200734) );
DFFARX1 I_11668  ( .D(I200734), .CLK(I2350), .RSTB(I200499), .Q(I200467) );
DFFARX1 I_11669  ( .D(I200734), .CLK(I2350), .RSTB(I200499), .Q(I200765) );
DFFARX1 I_11670  ( .D(I200734), .CLK(I2350), .RSTB(I200499), .Q(I200461) );
nand I_11671 (I200796,I200516,I91359);
nand I_11672 (I200813,I200796,I200550);
and I_11673 (I200830,I200632,I200813);
DFFARX1 I_11674  ( .D(I200830), .CLK(I2350), .RSTB(I200499), .Q(I200491) );
and I_11675 (I200464,I200796,I200765);
DFFARX1 I_11676  ( .D(I91353), .CLK(I2350), .RSTB(I200499), .Q(I200875) );
nor I_11677 (I200488,I200875,I200796);
nor I_11678 (I200906,I200875,I200550);
nand I_11679 (I200485,I200584,I200906);
not I_11680 (I200482,I200875);
DFFARX1 I_11681  ( .D(I91356), .CLK(I2350), .RSTB(I200499), .Q(I200951) );
not I_11682 (I200968,I200951);
nor I_11683 (I200985,I200968,I200649);
and I_11684 (I201002,I200875,I200985);
or I_11685 (I201019,I200796,I201002);
DFFARX1 I_11686  ( .D(I201019), .CLK(I2350), .RSTB(I200499), .Q(I200476) );
not I_11687 (I201050,I200968);
nor I_11688 (I201067,I200875,I201050);
nand I_11689 (I200479,I200968,I201067);
nand I_11690 (I200473,I200632,I201050);
not I_11691 (I201145,I2357);
not I_11692 (I201162,I2335);
nor I_11693 (I201179,I1359,I1319);
nand I_11694 (I201196,I201179,I2263);
nor I_11695 (I201213,I201162,I1359);
nand I_11696 (I201230,I201213,I1855);
DFFARX1 I_11697  ( .D(I201230), .CLK(I2350), .RSTB(I201145), .Q(I201247) );
not I_11698 (I201116,I201247);
not I_11699 (I201278,I1359);
not I_11700 (I201295,I201278);
not I_11701 (I201312,I1751);
nor I_11702 (I201329,I201312,I1695);
and I_11703 (I201346,I201329,I1847);
or I_11704 (I201363,I201346,I1215);
DFFARX1 I_11705  ( .D(I201363), .CLK(I2350), .RSTB(I201145), .Q(I201380) );
DFFARX1 I_11706  ( .D(I201380), .CLK(I2350), .RSTB(I201145), .Q(I201113) );
DFFARX1 I_11707  ( .D(I201380), .CLK(I2350), .RSTB(I201145), .Q(I201411) );
DFFARX1 I_11708  ( .D(I201380), .CLK(I2350), .RSTB(I201145), .Q(I201107) );
nand I_11709 (I201442,I201162,I1751);
nand I_11710 (I201459,I201442,I201196);
and I_11711 (I201476,I201278,I201459);
DFFARX1 I_11712  ( .D(I201476), .CLK(I2350), .RSTB(I201145), .Q(I201137) );
and I_11713 (I201110,I201442,I201411);
DFFARX1 I_11714  ( .D(I1519), .CLK(I2350), .RSTB(I201145), .Q(I201521) );
nor I_11715 (I201134,I201521,I201442);
nor I_11716 (I201552,I201521,I201196);
nand I_11717 (I201131,I201230,I201552);
not I_11718 (I201128,I201521);
DFFARX1 I_11719  ( .D(I1463), .CLK(I2350), .RSTB(I201145), .Q(I201597) );
not I_11720 (I201614,I201597);
nor I_11721 (I201631,I201614,I201295);
and I_11722 (I201648,I201521,I201631);
or I_11723 (I201665,I201442,I201648);
DFFARX1 I_11724  ( .D(I201665), .CLK(I2350), .RSTB(I201145), .Q(I201122) );
not I_11725 (I201696,I201614);
nor I_11726 (I201713,I201521,I201696);
nand I_11727 (I201125,I201614,I201713);
nand I_11728 (I201119,I201278,I201696);
not I_11729 (I201791,I2357);
not I_11730 (I201808,I373508);
nor I_11731 (I201825,I373505,I373490);
nand I_11732 (I201842,I201825,I373499);
nor I_11733 (I201859,I201808,I373505);
nand I_11734 (I201876,I201859,I373514);
DFFARX1 I_11735  ( .D(I201876), .CLK(I2350), .RSTB(I201791), .Q(I201893) );
not I_11736 (I201762,I201893);
not I_11737 (I201924,I373505);
not I_11738 (I201941,I201924);
not I_11739 (I201958,I373487);
nor I_11740 (I201975,I201958,I373493);
and I_11741 (I201992,I201975,I373517);
or I_11742 (I202009,I201992,I373511);
DFFARX1 I_11743  ( .D(I202009), .CLK(I2350), .RSTB(I201791), .Q(I202026) );
DFFARX1 I_11744  ( .D(I202026), .CLK(I2350), .RSTB(I201791), .Q(I201759) );
DFFARX1 I_11745  ( .D(I202026), .CLK(I2350), .RSTB(I201791), .Q(I202057) );
DFFARX1 I_11746  ( .D(I202026), .CLK(I2350), .RSTB(I201791), .Q(I201753) );
nand I_11747 (I202088,I201808,I373487);
nand I_11748 (I202105,I202088,I201842);
and I_11749 (I202122,I201924,I202105);
DFFARX1 I_11750  ( .D(I202122), .CLK(I2350), .RSTB(I201791), .Q(I201783) );
and I_11751 (I201756,I202088,I202057);
DFFARX1 I_11752  ( .D(I373496), .CLK(I2350), .RSTB(I201791), .Q(I202167) );
nor I_11753 (I201780,I202167,I202088);
nor I_11754 (I202198,I202167,I201842);
nand I_11755 (I201777,I201876,I202198);
not I_11756 (I201774,I202167);
DFFARX1 I_11757  ( .D(I373502), .CLK(I2350), .RSTB(I201791), .Q(I202243) );
not I_11758 (I202260,I202243);
nor I_11759 (I202277,I202260,I201941);
and I_11760 (I202294,I202167,I202277);
or I_11761 (I202311,I202088,I202294);
DFFARX1 I_11762  ( .D(I202311), .CLK(I2350), .RSTB(I201791), .Q(I201768) );
not I_11763 (I202342,I202260);
nor I_11764 (I202359,I202167,I202342);
nand I_11765 (I201771,I202260,I202359);
nand I_11766 (I201765,I201924,I202342);
not I_11767 (I202437,I2357);
not I_11768 (I202454,I42093);
nor I_11769 (I202471,I42084,I42075);
nand I_11770 (I202488,I202471,I42090);
nor I_11771 (I202505,I202454,I42084);
nand I_11772 (I202522,I202505,I42087);
DFFARX1 I_11773  ( .D(I202522), .CLK(I2350), .RSTB(I202437), .Q(I202539) );
not I_11774 (I202408,I202539);
not I_11775 (I202570,I42084);
not I_11776 (I202587,I202570);
not I_11777 (I202604,I42096);
nor I_11778 (I202621,I202604,I42081);
and I_11779 (I202638,I202621,I42099);
or I_11780 (I202655,I202638,I42072);
DFFARX1 I_11781  ( .D(I202655), .CLK(I2350), .RSTB(I202437), .Q(I202672) );
DFFARX1 I_11782  ( .D(I202672), .CLK(I2350), .RSTB(I202437), .Q(I202405) );
DFFARX1 I_11783  ( .D(I202672), .CLK(I2350), .RSTB(I202437), .Q(I202703) );
DFFARX1 I_11784  ( .D(I202672), .CLK(I2350), .RSTB(I202437), .Q(I202399) );
nand I_11785 (I202734,I202454,I42096);
nand I_11786 (I202751,I202734,I202488);
and I_11787 (I202768,I202570,I202751);
DFFARX1 I_11788  ( .D(I202768), .CLK(I2350), .RSTB(I202437), .Q(I202429) );
and I_11789 (I202402,I202734,I202703);
DFFARX1 I_11790  ( .D(I42102), .CLK(I2350), .RSTB(I202437), .Q(I202813) );
nor I_11791 (I202426,I202813,I202734);
nor I_11792 (I202844,I202813,I202488);
nand I_11793 (I202423,I202522,I202844);
not I_11794 (I202420,I202813);
DFFARX1 I_11795  ( .D(I42078), .CLK(I2350), .RSTB(I202437), .Q(I202889) );
not I_11796 (I202906,I202889);
nor I_11797 (I202923,I202906,I202587);
and I_11798 (I202940,I202813,I202923);
or I_11799 (I202957,I202734,I202940);
DFFARX1 I_11800  ( .D(I202957), .CLK(I2350), .RSTB(I202437), .Q(I202414) );
not I_11801 (I202988,I202906);
nor I_11802 (I203005,I202813,I202988);
nand I_11803 (I202417,I202906,I203005);
nand I_11804 (I202411,I202570,I202988);
not I_11805 (I203083,I2357);
not I_11806 (I203100,I2183);
nor I_11807 (I203117,I2071,I1575);
nand I_11808 (I203134,I203117,I2223);
nor I_11809 (I203151,I203100,I2071);
nand I_11810 (I203168,I203151,I2199);
DFFARX1 I_11811  ( .D(I203168), .CLK(I2350), .RSTB(I203083), .Q(I203185) );
not I_11812 (I203054,I203185);
not I_11813 (I203216,I2071);
not I_11814 (I203233,I203216);
not I_11815 (I203250,I2231);
nor I_11816 (I203267,I203250,I1343);
and I_11817 (I203284,I203267,I1263);
or I_11818 (I203301,I203284,I1975);
DFFARX1 I_11819  ( .D(I203301), .CLK(I2350), .RSTB(I203083), .Q(I203318) );
DFFARX1 I_11820  ( .D(I203318), .CLK(I2350), .RSTB(I203083), .Q(I203051) );
DFFARX1 I_11821  ( .D(I203318), .CLK(I2350), .RSTB(I203083), .Q(I203349) );
DFFARX1 I_11822  ( .D(I203318), .CLK(I2350), .RSTB(I203083), .Q(I203045) );
nand I_11823 (I203380,I203100,I2231);
nand I_11824 (I203397,I203380,I203134);
and I_11825 (I203414,I203216,I203397);
DFFARX1 I_11826  ( .D(I203414), .CLK(I2350), .RSTB(I203083), .Q(I203075) );
and I_11827 (I203048,I203380,I203349);
DFFARX1 I_11828  ( .D(I1679), .CLK(I2350), .RSTB(I203083), .Q(I203459) );
nor I_11829 (I203072,I203459,I203380);
nor I_11830 (I203490,I203459,I203134);
nand I_11831 (I203069,I203168,I203490);
not I_11832 (I203066,I203459);
DFFARX1 I_11833  ( .D(I1831), .CLK(I2350), .RSTB(I203083), .Q(I203535) );
not I_11834 (I203552,I203535);
nor I_11835 (I203569,I203552,I203233);
and I_11836 (I203586,I203459,I203569);
or I_11837 (I203603,I203380,I203586);
DFFARX1 I_11838  ( .D(I203603), .CLK(I2350), .RSTB(I203083), .Q(I203060) );
not I_11839 (I203634,I203552);
nor I_11840 (I203651,I203459,I203634);
nand I_11841 (I203063,I203552,I203651);
nand I_11842 (I203057,I203216,I203634);
not I_11843 (I203729,I2357);
not I_11844 (I203746,I61473);
nor I_11845 (I203763,I61464,I61455);
nand I_11846 (I203780,I203763,I61470);
nor I_11847 (I203797,I203746,I61464);
nand I_11848 (I203814,I203797,I61467);
DFFARX1 I_11849  ( .D(I203814), .CLK(I2350), .RSTB(I203729), .Q(I203831) );
not I_11850 (I203700,I203831);
not I_11851 (I203862,I61464);
not I_11852 (I203879,I203862);
not I_11853 (I203896,I61476);
nor I_11854 (I203913,I203896,I61461);
and I_11855 (I203930,I203913,I61479);
or I_11856 (I203947,I203930,I61452);
DFFARX1 I_11857  ( .D(I203947), .CLK(I2350), .RSTB(I203729), .Q(I203964) );
DFFARX1 I_11858  ( .D(I203964), .CLK(I2350), .RSTB(I203729), .Q(I203697) );
DFFARX1 I_11859  ( .D(I203964), .CLK(I2350), .RSTB(I203729), .Q(I203995) );
DFFARX1 I_11860  ( .D(I203964), .CLK(I2350), .RSTB(I203729), .Q(I203691) );
nand I_11861 (I204026,I203746,I61476);
nand I_11862 (I204043,I204026,I203780);
and I_11863 (I204060,I203862,I204043);
DFFARX1 I_11864  ( .D(I204060), .CLK(I2350), .RSTB(I203729), .Q(I203721) );
and I_11865 (I203694,I204026,I203995);
DFFARX1 I_11866  ( .D(I61482), .CLK(I2350), .RSTB(I203729), .Q(I204105) );
nor I_11867 (I203718,I204105,I204026);
nor I_11868 (I204136,I204105,I203780);
nand I_11869 (I203715,I203814,I204136);
not I_11870 (I203712,I204105);
DFFARX1 I_11871  ( .D(I61458), .CLK(I2350), .RSTB(I203729), .Q(I204181) );
not I_11872 (I204198,I204181);
nor I_11873 (I204215,I204198,I203879);
and I_11874 (I204232,I204105,I204215);
or I_11875 (I204249,I204026,I204232);
DFFARX1 I_11876  ( .D(I204249), .CLK(I2350), .RSTB(I203729), .Q(I203706) );
not I_11877 (I204280,I204198);
nor I_11878 (I204297,I204105,I204280);
nand I_11879 (I203709,I204198,I204297);
nand I_11880 (I203703,I203862,I204280);
not I_11881 (I204375,I2357);
not I_11882 (I204392,I246988);
nor I_11883 (I204409,I246991,I246973);
nand I_11884 (I204426,I204409,I247000);
nor I_11885 (I204443,I204392,I246991);
nand I_11886 (I204460,I204443,I246979);
DFFARX1 I_11887  ( .D(I204460), .CLK(I2350), .RSTB(I204375), .Q(I204477) );
not I_11888 (I204346,I204477);
not I_11889 (I204508,I246991);
not I_11890 (I204525,I204508);
not I_11891 (I204542,I246985);
nor I_11892 (I204559,I204542,I246997);
and I_11893 (I204576,I204559,I247003);
or I_11894 (I204593,I204576,I246982);
DFFARX1 I_11895  ( .D(I204593), .CLK(I2350), .RSTB(I204375), .Q(I204610) );
DFFARX1 I_11896  ( .D(I204610), .CLK(I2350), .RSTB(I204375), .Q(I204343) );
DFFARX1 I_11897  ( .D(I204610), .CLK(I2350), .RSTB(I204375), .Q(I204641) );
DFFARX1 I_11898  ( .D(I204610), .CLK(I2350), .RSTB(I204375), .Q(I204337) );
nand I_11899 (I204672,I204392,I246985);
nand I_11900 (I204689,I204672,I204426);
and I_11901 (I204706,I204508,I204689);
DFFARX1 I_11902  ( .D(I204706), .CLK(I2350), .RSTB(I204375), .Q(I204367) );
and I_11903 (I204340,I204672,I204641);
DFFARX1 I_11904  ( .D(I246994), .CLK(I2350), .RSTB(I204375), .Q(I204751) );
nor I_11905 (I204364,I204751,I204672);
nor I_11906 (I204782,I204751,I204426);
nand I_11907 (I204361,I204460,I204782);
not I_11908 (I204358,I204751);
DFFARX1 I_11909  ( .D(I246976), .CLK(I2350), .RSTB(I204375), .Q(I204827) );
not I_11910 (I204844,I204827);
nor I_11911 (I204861,I204844,I204525);
and I_11912 (I204878,I204751,I204861);
or I_11913 (I204895,I204672,I204878);
DFFARX1 I_11914  ( .D(I204895), .CLK(I2350), .RSTB(I204375), .Q(I204352) );
not I_11915 (I204926,I204844);
nor I_11916 (I204943,I204751,I204926);
nand I_11917 (I204355,I204844,I204943);
nand I_11918 (I204349,I204508,I204926);
not I_11919 (I205021,I2357);
not I_11920 (I205038,I276741);
nor I_11921 (I205055,I276747,I276732);
nand I_11922 (I205072,I205055,I276726);
nor I_11923 (I205089,I205038,I276747);
nand I_11924 (I205106,I205089,I276753);
DFFARX1 I_11925  ( .D(I205106), .CLK(I2350), .RSTB(I205021), .Q(I205123) );
not I_11926 (I204992,I205123);
not I_11927 (I205154,I276747);
not I_11928 (I205171,I205154);
not I_11929 (I205188,I276738);
nor I_11930 (I205205,I205188,I276744);
and I_11931 (I205222,I205205,I276750);
or I_11932 (I205239,I205222,I276723);
DFFARX1 I_11933  ( .D(I205239), .CLK(I2350), .RSTB(I205021), .Q(I205256) );
DFFARX1 I_11934  ( .D(I205256), .CLK(I2350), .RSTB(I205021), .Q(I204989) );
DFFARX1 I_11935  ( .D(I205256), .CLK(I2350), .RSTB(I205021), .Q(I205287) );
DFFARX1 I_11936  ( .D(I205256), .CLK(I2350), .RSTB(I205021), .Q(I204983) );
nand I_11937 (I205318,I205038,I276738);
nand I_11938 (I205335,I205318,I205072);
and I_11939 (I205352,I205154,I205335);
DFFARX1 I_11940  ( .D(I205352), .CLK(I2350), .RSTB(I205021), .Q(I205013) );
and I_11941 (I204986,I205318,I205287);
DFFARX1 I_11942  ( .D(I276729), .CLK(I2350), .RSTB(I205021), .Q(I205397) );
nor I_11943 (I205010,I205397,I205318);
nor I_11944 (I205428,I205397,I205072);
nand I_11945 (I205007,I205106,I205428);
not I_11946 (I205004,I205397);
DFFARX1 I_11947  ( .D(I276735), .CLK(I2350), .RSTB(I205021), .Q(I205473) );
not I_11948 (I205490,I205473);
nor I_11949 (I205507,I205490,I205171);
and I_11950 (I205524,I205397,I205507);
or I_11951 (I205541,I205318,I205524);
DFFARX1 I_11952  ( .D(I205541), .CLK(I2350), .RSTB(I205021), .Q(I204998) );
not I_11953 (I205572,I205490);
nor I_11954 (I205589,I205397,I205572);
nand I_11955 (I205001,I205490,I205589);
nand I_11956 (I204995,I205154,I205572);
not I_11957 (I205667,I2357);
not I_11958 (I205684,I29819);
nor I_11959 (I205701,I29810,I29801);
nand I_11960 (I205718,I205701,I29816);
nor I_11961 (I205735,I205684,I29810);
nand I_11962 (I205752,I205735,I29813);
DFFARX1 I_11963  ( .D(I205752), .CLK(I2350), .RSTB(I205667), .Q(I205769) );
not I_11964 (I205638,I205769);
not I_11965 (I205800,I29810);
not I_11966 (I205817,I205800);
not I_11967 (I205834,I29822);
nor I_11968 (I205851,I205834,I29807);
and I_11969 (I205868,I205851,I29825);
or I_11970 (I205885,I205868,I29798);
DFFARX1 I_11971  ( .D(I205885), .CLK(I2350), .RSTB(I205667), .Q(I205902) );
DFFARX1 I_11972  ( .D(I205902), .CLK(I2350), .RSTB(I205667), .Q(I205635) );
DFFARX1 I_11973  ( .D(I205902), .CLK(I2350), .RSTB(I205667), .Q(I205933) );
DFFARX1 I_11974  ( .D(I205902), .CLK(I2350), .RSTB(I205667), .Q(I205629) );
nand I_11975 (I205964,I205684,I29822);
nand I_11976 (I205981,I205964,I205718);
and I_11977 (I205998,I205800,I205981);
DFFARX1 I_11978  ( .D(I205998), .CLK(I2350), .RSTB(I205667), .Q(I205659) );
and I_11979 (I205632,I205964,I205933);
DFFARX1 I_11980  ( .D(I29828), .CLK(I2350), .RSTB(I205667), .Q(I206043) );
nor I_11981 (I205656,I206043,I205964);
nor I_11982 (I206074,I206043,I205718);
nand I_11983 (I205653,I205752,I206074);
not I_11984 (I205650,I206043);
DFFARX1 I_11985  ( .D(I29804), .CLK(I2350), .RSTB(I205667), .Q(I206119) );
not I_11986 (I206136,I206119);
nor I_11987 (I206153,I206136,I205817);
and I_11988 (I206170,I206043,I206153);
or I_11989 (I206187,I205964,I206170);
DFFARX1 I_11990  ( .D(I206187), .CLK(I2350), .RSTB(I205667), .Q(I205644) );
not I_11991 (I206218,I206136);
nor I_11992 (I206235,I206043,I206218);
nand I_11993 (I205647,I206136,I206235);
nand I_11994 (I205641,I205800,I206218);
not I_11995 (I206313,I2357);
not I_11996 (I206330,I31111);
nor I_11997 (I206347,I31102,I31093);
nand I_11998 (I206364,I206347,I31108);
nor I_11999 (I206381,I206330,I31102);
nand I_12000 (I206398,I206381,I31105);
DFFARX1 I_12001  ( .D(I206398), .CLK(I2350), .RSTB(I206313), .Q(I206415) );
not I_12002 (I206284,I206415);
not I_12003 (I206446,I31102);
not I_12004 (I206463,I206446);
not I_12005 (I206480,I31114);
nor I_12006 (I206497,I206480,I31099);
and I_12007 (I206514,I206497,I31117);
or I_12008 (I206531,I206514,I31090);
DFFARX1 I_12009  ( .D(I206531), .CLK(I2350), .RSTB(I206313), .Q(I206548) );
DFFARX1 I_12010  ( .D(I206548), .CLK(I2350), .RSTB(I206313), .Q(I206281) );
DFFARX1 I_12011  ( .D(I206548), .CLK(I2350), .RSTB(I206313), .Q(I206579) );
DFFARX1 I_12012  ( .D(I206548), .CLK(I2350), .RSTB(I206313), .Q(I206275) );
nand I_12013 (I206610,I206330,I31114);
nand I_12014 (I206627,I206610,I206364);
and I_12015 (I206644,I206446,I206627);
DFFARX1 I_12016  ( .D(I206644), .CLK(I2350), .RSTB(I206313), .Q(I206305) );
and I_12017 (I206278,I206610,I206579);
DFFARX1 I_12018  ( .D(I31120), .CLK(I2350), .RSTB(I206313), .Q(I206689) );
nor I_12019 (I206302,I206689,I206610);
nor I_12020 (I206720,I206689,I206364);
nand I_12021 (I206299,I206398,I206720);
not I_12022 (I206296,I206689);
DFFARX1 I_12023  ( .D(I31096), .CLK(I2350), .RSTB(I206313), .Q(I206765) );
not I_12024 (I206782,I206765);
nor I_12025 (I206799,I206782,I206463);
and I_12026 (I206816,I206689,I206799);
or I_12027 (I206833,I206610,I206816);
DFFARX1 I_12028  ( .D(I206833), .CLK(I2350), .RSTB(I206313), .Q(I206290) );
not I_12029 (I206864,I206782);
nor I_12030 (I206881,I206689,I206864);
nand I_12031 (I206293,I206782,I206881);
nand I_12032 (I206287,I206446,I206864);
not I_12033 (I206959,I2357);
not I_12034 (I206976,I81499);
nor I_12035 (I206993,I81490,I81481);
nand I_12036 (I207010,I206993,I81496);
nor I_12037 (I207027,I206976,I81490);
nand I_12038 (I207044,I207027,I81493);
DFFARX1 I_12039  ( .D(I207044), .CLK(I2350), .RSTB(I206959), .Q(I207061) );
not I_12040 (I206930,I207061);
not I_12041 (I207092,I81490);
not I_12042 (I207109,I207092);
not I_12043 (I207126,I81502);
nor I_12044 (I207143,I207126,I81487);
and I_12045 (I207160,I207143,I81505);
or I_12046 (I207177,I207160,I81478);
DFFARX1 I_12047  ( .D(I207177), .CLK(I2350), .RSTB(I206959), .Q(I207194) );
DFFARX1 I_12048  ( .D(I207194), .CLK(I2350), .RSTB(I206959), .Q(I206927) );
DFFARX1 I_12049  ( .D(I207194), .CLK(I2350), .RSTB(I206959), .Q(I207225) );
DFFARX1 I_12050  ( .D(I207194), .CLK(I2350), .RSTB(I206959), .Q(I206921) );
nand I_12051 (I207256,I206976,I81502);
nand I_12052 (I207273,I207256,I207010);
and I_12053 (I207290,I207092,I207273);
DFFARX1 I_12054  ( .D(I207290), .CLK(I2350), .RSTB(I206959), .Q(I206951) );
and I_12055 (I206924,I207256,I207225);
DFFARX1 I_12056  ( .D(I81508), .CLK(I2350), .RSTB(I206959), .Q(I207335) );
nor I_12057 (I206948,I207335,I207256);
nor I_12058 (I207366,I207335,I207010);
nand I_12059 (I206945,I207044,I207366);
not I_12060 (I206942,I207335);
DFFARX1 I_12061  ( .D(I81484), .CLK(I2350), .RSTB(I206959), .Q(I207411) );
not I_12062 (I207428,I207411);
nor I_12063 (I207445,I207428,I207109);
and I_12064 (I207462,I207335,I207445);
or I_12065 (I207479,I207256,I207462);
DFFARX1 I_12066  ( .D(I207479), .CLK(I2350), .RSTB(I206959), .Q(I206936) );
not I_12067 (I207510,I207428);
nor I_12068 (I207527,I207335,I207510);
nand I_12069 (I206939,I207428,I207527);
nand I_12070 (I206933,I207092,I207510);
not I_12071 (I207605,I2357);
not I_12072 (I207622,I188092);
nor I_12073 (I207639,I188071,I188083);
nand I_12074 (I207656,I207639,I188086);
nor I_12075 (I207673,I207622,I188071);
nand I_12076 (I207690,I207673,I188068);
DFFARX1 I_12077  ( .D(I207690), .CLK(I2350), .RSTB(I207605), .Q(I207707) );
not I_12078 (I207576,I207707);
not I_12079 (I207738,I188071);
not I_12080 (I207755,I207738);
not I_12081 (I207772,I188089);
nor I_12082 (I207789,I207772,I188080);
and I_12083 (I207806,I207789,I188074);
or I_12084 (I207823,I207806,I188098);
DFFARX1 I_12085  ( .D(I207823), .CLK(I2350), .RSTB(I207605), .Q(I207840) );
DFFARX1 I_12086  ( .D(I207840), .CLK(I2350), .RSTB(I207605), .Q(I207573) );
DFFARX1 I_12087  ( .D(I207840), .CLK(I2350), .RSTB(I207605), .Q(I207871) );
DFFARX1 I_12088  ( .D(I207840), .CLK(I2350), .RSTB(I207605), .Q(I207567) );
nand I_12089 (I207902,I207622,I188089);
nand I_12090 (I207919,I207902,I207656);
and I_12091 (I207936,I207738,I207919);
DFFARX1 I_12092  ( .D(I207936), .CLK(I2350), .RSTB(I207605), .Q(I207597) );
and I_12093 (I207570,I207902,I207871);
DFFARX1 I_12094  ( .D(I188095), .CLK(I2350), .RSTB(I207605), .Q(I207981) );
nor I_12095 (I207594,I207981,I207902);
nor I_12096 (I208012,I207981,I207656);
nand I_12097 (I207591,I207690,I208012);
not I_12098 (I207588,I207981);
DFFARX1 I_12099  ( .D(I188077), .CLK(I2350), .RSTB(I207605), .Q(I208057) );
not I_12100 (I208074,I208057);
nor I_12101 (I208091,I208074,I207755);
and I_12102 (I208108,I207981,I208091);
or I_12103 (I208125,I207902,I208108);
DFFARX1 I_12104  ( .D(I208125), .CLK(I2350), .RSTB(I207605), .Q(I207582) );
not I_12105 (I208156,I208074);
nor I_12106 (I208173,I207981,I208156);
nand I_12107 (I207585,I208074,I208173);
nand I_12108 (I207579,I207738,I208156);
not I_12109 (I208251,I2357);
not I_12110 (I208268,I342687);
nor I_12111 (I208285,I342684,I342669);
nand I_12112 (I208302,I208285,I342678);
nor I_12113 (I208319,I208268,I342684);
nand I_12114 (I208336,I208319,I342693);
DFFARX1 I_12115  ( .D(I208336), .CLK(I2350), .RSTB(I208251), .Q(I208353) );
not I_12116 (I208222,I208353);
not I_12117 (I208384,I342684);
not I_12118 (I208401,I208384);
not I_12119 (I208418,I342666);
nor I_12120 (I208435,I208418,I342672);
and I_12121 (I208452,I208435,I342696);
or I_12122 (I208469,I208452,I342690);
DFFARX1 I_12123  ( .D(I208469), .CLK(I2350), .RSTB(I208251), .Q(I208486) );
DFFARX1 I_12124  ( .D(I208486), .CLK(I2350), .RSTB(I208251), .Q(I208219) );
DFFARX1 I_12125  ( .D(I208486), .CLK(I2350), .RSTB(I208251), .Q(I208517) );
DFFARX1 I_12126  ( .D(I208486), .CLK(I2350), .RSTB(I208251), .Q(I208213) );
nand I_12127 (I208548,I208268,I342666);
nand I_12128 (I208565,I208548,I208302);
and I_12129 (I208582,I208384,I208565);
DFFARX1 I_12130  ( .D(I208582), .CLK(I2350), .RSTB(I208251), .Q(I208243) );
and I_12131 (I208216,I208548,I208517);
DFFARX1 I_12132  ( .D(I342675), .CLK(I2350), .RSTB(I208251), .Q(I208627) );
nor I_12133 (I208240,I208627,I208548);
nor I_12134 (I208658,I208627,I208302);
nand I_12135 (I208237,I208336,I208658);
not I_12136 (I208234,I208627);
DFFARX1 I_12137  ( .D(I342681), .CLK(I2350), .RSTB(I208251), .Q(I208703) );
not I_12138 (I208720,I208703);
nor I_12139 (I208737,I208720,I208401);
and I_12140 (I208754,I208627,I208737);
or I_12141 (I208771,I208548,I208754);
DFFARX1 I_12142  ( .D(I208771), .CLK(I2350), .RSTB(I208251), .Q(I208228) );
not I_12143 (I208802,I208720);
nor I_12144 (I208819,I208627,I208802);
nand I_12145 (I208231,I208720,I208819);
nand I_12146 (I208225,I208384,I208802);
not I_12147 (I208897,I2357);
not I_12148 (I208914,I361557);
nor I_12149 (I208931,I361554,I361539);
nand I_12150 (I208948,I208931,I361548);
nor I_12151 (I208965,I208914,I361554);
nand I_12152 (I208982,I208965,I361563);
DFFARX1 I_12153  ( .D(I208982), .CLK(I2350), .RSTB(I208897), .Q(I208999) );
not I_12154 (I208868,I208999);
not I_12155 (I209030,I361554);
not I_12156 (I209047,I209030);
not I_12157 (I209064,I361536);
nor I_12158 (I209081,I209064,I361542);
and I_12159 (I209098,I209081,I361566);
or I_12160 (I209115,I209098,I361560);
DFFARX1 I_12161  ( .D(I209115), .CLK(I2350), .RSTB(I208897), .Q(I209132) );
DFFARX1 I_12162  ( .D(I209132), .CLK(I2350), .RSTB(I208897), .Q(I208865) );
DFFARX1 I_12163  ( .D(I209132), .CLK(I2350), .RSTB(I208897), .Q(I209163) );
DFFARX1 I_12164  ( .D(I209132), .CLK(I2350), .RSTB(I208897), .Q(I208859) );
nand I_12165 (I209194,I208914,I361536);
nand I_12166 (I209211,I209194,I208948);
and I_12167 (I209228,I209030,I209211);
DFFARX1 I_12168  ( .D(I209228), .CLK(I2350), .RSTB(I208897), .Q(I208889) );
and I_12169 (I208862,I209194,I209163);
DFFARX1 I_12170  ( .D(I361545), .CLK(I2350), .RSTB(I208897), .Q(I209273) );
nor I_12171 (I208886,I209273,I209194);
nor I_12172 (I209304,I209273,I208948);
nand I_12173 (I208883,I208982,I209304);
not I_12174 (I208880,I209273);
DFFARX1 I_12175  ( .D(I361551), .CLK(I2350), .RSTB(I208897), .Q(I209349) );
not I_12176 (I209366,I209349);
nor I_12177 (I209383,I209366,I209047);
and I_12178 (I209400,I209273,I209383);
or I_12179 (I209417,I209194,I209400);
DFFARX1 I_12180  ( .D(I209417), .CLK(I2350), .RSTB(I208897), .Q(I208874) );
not I_12181 (I209448,I209366);
nor I_12182 (I209465,I209273,I209448);
nand I_12183 (I208877,I209366,I209465);
nand I_12184 (I208871,I209030,I209448);
not I_12185 (I209543,I2357);
not I_12186 (I209560,I376653);
nor I_12187 (I209577,I376650,I376635);
nand I_12188 (I209594,I209577,I376644);
nor I_12189 (I209611,I209560,I376650);
nand I_12190 (I209628,I209611,I376659);
DFFARX1 I_12191  ( .D(I209628), .CLK(I2350), .RSTB(I209543), .Q(I209645) );
not I_12192 (I209514,I209645);
not I_12193 (I209676,I376650);
not I_12194 (I209693,I209676);
not I_12195 (I209710,I376632);
nor I_12196 (I209727,I209710,I376638);
and I_12197 (I209744,I209727,I376662);
or I_12198 (I209761,I209744,I376656);
DFFARX1 I_12199  ( .D(I209761), .CLK(I2350), .RSTB(I209543), .Q(I209778) );
DFFARX1 I_12200  ( .D(I209778), .CLK(I2350), .RSTB(I209543), .Q(I209511) );
DFFARX1 I_12201  ( .D(I209778), .CLK(I2350), .RSTB(I209543), .Q(I209809) );
DFFARX1 I_12202  ( .D(I209778), .CLK(I2350), .RSTB(I209543), .Q(I209505) );
nand I_12203 (I209840,I209560,I376632);
nand I_12204 (I209857,I209840,I209594);
and I_12205 (I209874,I209676,I209857);
DFFARX1 I_12206  ( .D(I209874), .CLK(I2350), .RSTB(I209543), .Q(I209535) );
and I_12207 (I209508,I209840,I209809);
DFFARX1 I_12208  ( .D(I376641), .CLK(I2350), .RSTB(I209543), .Q(I209919) );
nor I_12209 (I209532,I209919,I209840);
nor I_12210 (I209950,I209919,I209594);
nand I_12211 (I209529,I209628,I209950);
not I_12212 (I209526,I209919);
DFFARX1 I_12213  ( .D(I376647), .CLK(I2350), .RSTB(I209543), .Q(I209995) );
not I_12214 (I210012,I209995);
nor I_12215 (I210029,I210012,I209693);
and I_12216 (I210046,I209919,I210029);
or I_12217 (I210063,I209840,I210046);
DFFARX1 I_12218  ( .D(I210063), .CLK(I2350), .RSTB(I209543), .Q(I209520) );
not I_12219 (I210094,I210012);
nor I_12220 (I210111,I209919,I210094);
nand I_12221 (I209523,I210012,I210111);
nand I_12222 (I209517,I209676,I210094);
not I_12223 (I210189,I2357);
not I_12224 (I210206,I393769);
nor I_12225 (I210223,I393754,I393760);
nand I_12226 (I210240,I210223,I393757);
nor I_12227 (I210257,I210206,I393754);
nand I_12228 (I210274,I210257,I393766);
DFFARX1 I_12229  ( .D(I210274), .CLK(I2350), .RSTB(I210189), .Q(I210291) );
not I_12230 (I210160,I210291);
not I_12231 (I210322,I393754);
not I_12232 (I210339,I210322);
not I_12233 (I210356,I393781);
nor I_12234 (I210373,I210356,I393775);
and I_12235 (I210390,I210373,I393772);
or I_12236 (I210407,I210390,I393751);
DFFARX1 I_12237  ( .D(I210407), .CLK(I2350), .RSTB(I210189), .Q(I210424) );
DFFARX1 I_12238  ( .D(I210424), .CLK(I2350), .RSTB(I210189), .Q(I210157) );
DFFARX1 I_12239  ( .D(I210424), .CLK(I2350), .RSTB(I210189), .Q(I210455) );
DFFARX1 I_12240  ( .D(I210424), .CLK(I2350), .RSTB(I210189), .Q(I210151) );
nand I_12241 (I210486,I210206,I393781);
nand I_12242 (I210503,I210486,I210240);
and I_12243 (I210520,I210322,I210503);
DFFARX1 I_12244  ( .D(I210520), .CLK(I2350), .RSTB(I210189), .Q(I210181) );
and I_12245 (I210154,I210486,I210455);
DFFARX1 I_12246  ( .D(I393778), .CLK(I2350), .RSTB(I210189), .Q(I210565) );
nor I_12247 (I210178,I210565,I210486);
nor I_12248 (I210596,I210565,I210240);
nand I_12249 (I210175,I210274,I210596);
not I_12250 (I210172,I210565);
DFFARX1 I_12251  ( .D(I393763), .CLK(I2350), .RSTB(I210189), .Q(I210641) );
not I_12252 (I210658,I210641);
nor I_12253 (I210675,I210658,I210339);
and I_12254 (I210692,I210565,I210675);
or I_12255 (I210709,I210486,I210692);
DFFARX1 I_12256  ( .D(I210709), .CLK(I2350), .RSTB(I210189), .Q(I210166) );
not I_12257 (I210740,I210658);
nor I_12258 (I210757,I210565,I210740);
nand I_12259 (I210169,I210658,I210757);
nand I_12260 (I210163,I210322,I210740);
not I_12261 (I210835,I2357);
not I_12262 (I210852,I291556);
nor I_12263 (I210869,I291568,I291562);
nand I_12264 (I210886,I210869,I291547);
nor I_12265 (I210903,I210852,I291568);
nand I_12266 (I210920,I210903,I291574);
DFFARX1 I_12267  ( .D(I210920), .CLK(I2350), .RSTB(I210835), .Q(I210937) );
not I_12268 (I210806,I210937);
not I_12269 (I210968,I291568);
not I_12270 (I210985,I210968);
not I_12271 (I211002,I291571);
nor I_12272 (I211019,I211002,I291553);
and I_12273 (I211036,I211019,I291550);
or I_12274 (I211053,I211036,I291577);
DFFARX1 I_12275  ( .D(I211053), .CLK(I2350), .RSTB(I210835), .Q(I211070) );
DFFARX1 I_12276  ( .D(I211070), .CLK(I2350), .RSTB(I210835), .Q(I210803) );
DFFARX1 I_12277  ( .D(I211070), .CLK(I2350), .RSTB(I210835), .Q(I211101) );
DFFARX1 I_12278  ( .D(I211070), .CLK(I2350), .RSTB(I210835), .Q(I210797) );
nand I_12279 (I211132,I210852,I291571);
nand I_12280 (I211149,I211132,I210886);
and I_12281 (I211166,I210968,I211149);
DFFARX1 I_12282  ( .D(I211166), .CLK(I2350), .RSTB(I210835), .Q(I210827) );
and I_12283 (I210800,I211132,I211101);
DFFARX1 I_12284  ( .D(I291565), .CLK(I2350), .RSTB(I210835), .Q(I211211) );
nor I_12285 (I210824,I211211,I211132);
nor I_12286 (I211242,I211211,I210886);
nand I_12287 (I210821,I210920,I211242);
not I_12288 (I210818,I211211);
DFFARX1 I_12289  ( .D(I291559), .CLK(I2350), .RSTB(I210835), .Q(I211287) );
not I_12290 (I211304,I211287);
nor I_12291 (I211321,I211304,I210985);
and I_12292 (I211338,I211211,I211321);
or I_12293 (I211355,I211132,I211338);
DFFARX1 I_12294  ( .D(I211355), .CLK(I2350), .RSTB(I210835), .Q(I210812) );
not I_12295 (I211386,I211304);
nor I_12296 (I211403,I211211,I211386);
nand I_12297 (I210815,I211304,I211403);
nand I_12298 (I210809,I210968,I211386);
not I_12299 (I211481,I2357);
not I_12300 (I211498,I174832);
nor I_12301 (I211515,I174811,I174823);
nand I_12302 (I211532,I211515,I174826);
nor I_12303 (I211549,I211498,I174811);
nand I_12304 (I211566,I211549,I174808);
DFFARX1 I_12305  ( .D(I211566), .CLK(I2350), .RSTB(I211481), .Q(I211583) );
not I_12306 (I211452,I211583);
not I_12307 (I211614,I174811);
not I_12308 (I211631,I211614);
not I_12309 (I211648,I174829);
nor I_12310 (I211665,I211648,I174820);
and I_12311 (I211682,I211665,I174814);
or I_12312 (I211699,I211682,I174838);
DFFARX1 I_12313  ( .D(I211699), .CLK(I2350), .RSTB(I211481), .Q(I211716) );
DFFARX1 I_12314  ( .D(I211716), .CLK(I2350), .RSTB(I211481), .Q(I211449) );
DFFARX1 I_12315  ( .D(I211716), .CLK(I2350), .RSTB(I211481), .Q(I211747) );
DFFARX1 I_12316  ( .D(I211716), .CLK(I2350), .RSTB(I211481), .Q(I211443) );
nand I_12317 (I211778,I211498,I174829);
nand I_12318 (I211795,I211778,I211532);
and I_12319 (I211812,I211614,I211795);
DFFARX1 I_12320  ( .D(I211812), .CLK(I2350), .RSTB(I211481), .Q(I211473) );
and I_12321 (I211446,I211778,I211747);
DFFARX1 I_12322  ( .D(I174835), .CLK(I2350), .RSTB(I211481), .Q(I211857) );
nor I_12323 (I211470,I211857,I211778);
nor I_12324 (I211888,I211857,I211532);
nand I_12325 (I211467,I211566,I211888);
not I_12326 (I211464,I211857);
DFFARX1 I_12327  ( .D(I174817), .CLK(I2350), .RSTB(I211481), .Q(I211933) );
not I_12328 (I211950,I211933);
nor I_12329 (I211967,I211950,I211631);
and I_12330 (I211984,I211857,I211967);
or I_12331 (I212001,I211778,I211984);
DFFARX1 I_12332  ( .D(I212001), .CLK(I2350), .RSTB(I211481), .Q(I211458) );
not I_12333 (I212032,I211950);
nor I_12334 (I212049,I211857,I212032);
nand I_12335 (I211461,I211950,I212049);
nand I_12336 (I211455,I211614,I212032);
not I_12337 (I212127,I2357);
not I_12338 (I212144,I321910);
nor I_12339 (I212161,I321898,I321907);
nand I_12340 (I212178,I212161,I321922);
nor I_12341 (I212195,I212144,I321898);
nand I_12342 (I212212,I212195,I321904);
DFFARX1 I_12343  ( .D(I212212), .CLK(I2350), .RSTB(I212127), .Q(I212229) );
not I_12344 (I212098,I212229);
not I_12345 (I212260,I321898);
not I_12346 (I212277,I212260);
not I_12347 (I212294,I321892);
nor I_12348 (I212311,I212294,I321913);
and I_12349 (I212328,I212311,I321895);
or I_12350 (I212345,I212328,I321901);
DFFARX1 I_12351  ( .D(I212345), .CLK(I2350), .RSTB(I212127), .Q(I212362) );
DFFARX1 I_12352  ( .D(I212362), .CLK(I2350), .RSTB(I212127), .Q(I212095) );
DFFARX1 I_12353  ( .D(I212362), .CLK(I2350), .RSTB(I212127), .Q(I212393) );
DFFARX1 I_12354  ( .D(I212362), .CLK(I2350), .RSTB(I212127), .Q(I212089) );
nand I_12355 (I212424,I212144,I321892);
nand I_12356 (I212441,I212424,I212178);
and I_12357 (I212458,I212260,I212441);
DFFARX1 I_12358  ( .D(I212458), .CLK(I2350), .RSTB(I212127), .Q(I212119) );
and I_12359 (I212092,I212424,I212393);
DFFARX1 I_12360  ( .D(I321919), .CLK(I2350), .RSTB(I212127), .Q(I212503) );
nor I_12361 (I212116,I212503,I212424);
nor I_12362 (I212534,I212503,I212178);
nand I_12363 (I212113,I212212,I212534);
not I_12364 (I212110,I212503);
DFFARX1 I_12365  ( .D(I321916), .CLK(I2350), .RSTB(I212127), .Q(I212579) );
not I_12366 (I212596,I212579);
nor I_12367 (I212613,I212596,I212277);
and I_12368 (I212630,I212503,I212613);
or I_12369 (I212647,I212424,I212630);
DFFARX1 I_12370  ( .D(I212647), .CLK(I2350), .RSTB(I212127), .Q(I212104) );
not I_12371 (I212678,I212596);
nor I_12372 (I212695,I212503,I212678);
nand I_12373 (I212107,I212596,I212695);
nand I_12374 (I212101,I212260,I212678);
not I_12375 (I212773,I2357);
not I_12376 (I212790,I4613);
nor I_12377 (I212807,I4628,I4622);
nand I_12378 (I212824,I212807,I4631);
nor I_12379 (I212841,I212790,I4628);
nand I_12380 (I212858,I212841,I4607);
DFFARX1 I_12381  ( .D(I212858), .CLK(I2350), .RSTB(I212773), .Q(I212875) );
not I_12382 (I212744,I212875);
not I_12383 (I212906,I4628);
not I_12384 (I212923,I212906);
not I_12385 (I212940,I4604);
nor I_12386 (I212957,I212940,I4619);
and I_12387 (I212974,I212957,I4625);
or I_12388 (I212991,I212974,I4634);
DFFARX1 I_12389  ( .D(I212991), .CLK(I2350), .RSTB(I212773), .Q(I213008) );
DFFARX1 I_12390  ( .D(I213008), .CLK(I2350), .RSTB(I212773), .Q(I212741) );
DFFARX1 I_12391  ( .D(I213008), .CLK(I2350), .RSTB(I212773), .Q(I213039) );
DFFARX1 I_12392  ( .D(I213008), .CLK(I2350), .RSTB(I212773), .Q(I212735) );
nand I_12393 (I213070,I212790,I4604);
nand I_12394 (I213087,I213070,I212824);
and I_12395 (I213104,I212906,I213087);
DFFARX1 I_12396  ( .D(I213104), .CLK(I2350), .RSTB(I212773), .Q(I212765) );
and I_12397 (I212738,I213070,I213039);
DFFARX1 I_12398  ( .D(I4616), .CLK(I2350), .RSTB(I212773), .Q(I213149) );
nor I_12399 (I212762,I213149,I213070);
nor I_12400 (I213180,I213149,I212824);
nand I_12401 (I212759,I212858,I213180);
not I_12402 (I212756,I213149);
DFFARX1 I_12403  ( .D(I4610), .CLK(I2350), .RSTB(I212773), .Q(I213225) );
not I_12404 (I213242,I213225);
nor I_12405 (I213259,I213242,I212923);
and I_12406 (I213276,I213149,I213259);
or I_12407 (I213293,I213070,I213276);
DFFARX1 I_12408  ( .D(I213293), .CLK(I2350), .RSTB(I212773), .Q(I212750) );
not I_12409 (I213324,I213242);
nor I_12410 (I213341,I213149,I213324);
nand I_12411 (I212753,I213242,I213341);
nand I_12412 (I212747,I212906,I213324);
not I_12413 (I213419,I2357);
not I_12414 (I213436,I348977);
nor I_12415 (I213453,I348974,I348959);
nand I_12416 (I213470,I213453,I348968);
nor I_12417 (I213487,I213436,I348974);
nand I_12418 (I213504,I213487,I348983);
DFFARX1 I_12419  ( .D(I213504), .CLK(I2350), .RSTB(I213419), .Q(I213521) );
not I_12420 (I213390,I213521);
not I_12421 (I213552,I348974);
not I_12422 (I213569,I213552);
not I_12423 (I213586,I348956);
nor I_12424 (I213603,I213586,I348962);
and I_12425 (I213620,I213603,I348986);
or I_12426 (I213637,I213620,I348980);
DFFARX1 I_12427  ( .D(I213637), .CLK(I2350), .RSTB(I213419), .Q(I213654) );
DFFARX1 I_12428  ( .D(I213654), .CLK(I2350), .RSTB(I213419), .Q(I213387) );
DFFARX1 I_12429  ( .D(I213654), .CLK(I2350), .RSTB(I213419), .Q(I213685) );
DFFARX1 I_12430  ( .D(I213654), .CLK(I2350), .RSTB(I213419), .Q(I213381) );
nand I_12431 (I213716,I213436,I348956);
nand I_12432 (I213733,I213716,I213470);
and I_12433 (I213750,I213552,I213733);
DFFARX1 I_12434  ( .D(I213750), .CLK(I2350), .RSTB(I213419), .Q(I213411) );
and I_12435 (I213384,I213716,I213685);
DFFARX1 I_12436  ( .D(I348965), .CLK(I2350), .RSTB(I213419), .Q(I213795) );
nor I_12437 (I213408,I213795,I213716);
nor I_12438 (I213826,I213795,I213470);
nand I_12439 (I213405,I213504,I213826);
not I_12440 (I213402,I213795);
DFFARX1 I_12441  ( .D(I348971), .CLK(I2350), .RSTB(I213419), .Q(I213871) );
not I_12442 (I213888,I213871);
nor I_12443 (I213905,I213888,I213569);
and I_12444 (I213922,I213795,I213905);
or I_12445 (I213939,I213716,I213922);
DFFARX1 I_12446  ( .D(I213939), .CLK(I2350), .RSTB(I213419), .Q(I213396) );
not I_12447 (I213970,I213888);
nor I_12448 (I213987,I213795,I213970);
nand I_12449 (I213399,I213888,I213987);
nand I_12450 (I213393,I213552,I213970);
not I_12451 (I214065,I2357);
not I_12452 (I214082,I80207);
nor I_12453 (I214099,I80198,I80189);
nand I_12454 (I214116,I214099,I80204);
nor I_12455 (I214133,I214082,I80198);
nand I_12456 (I214150,I214133,I80201);
DFFARX1 I_12457  ( .D(I214150), .CLK(I2350), .RSTB(I214065), .Q(I214167) );
not I_12458 (I214036,I214167);
not I_12459 (I214198,I80198);
not I_12460 (I214215,I214198);
not I_12461 (I214232,I80210);
nor I_12462 (I214249,I214232,I80195);
and I_12463 (I214266,I214249,I80213);
or I_12464 (I214283,I214266,I80186);
DFFARX1 I_12465  ( .D(I214283), .CLK(I2350), .RSTB(I214065), .Q(I214300) );
DFFARX1 I_12466  ( .D(I214300), .CLK(I2350), .RSTB(I214065), .Q(I214033) );
DFFARX1 I_12467  ( .D(I214300), .CLK(I2350), .RSTB(I214065), .Q(I214331) );
DFFARX1 I_12468  ( .D(I214300), .CLK(I2350), .RSTB(I214065), .Q(I214027) );
nand I_12469 (I214362,I214082,I80210);
nand I_12470 (I214379,I214362,I214116);
and I_12471 (I214396,I214198,I214379);
DFFARX1 I_12472  ( .D(I214396), .CLK(I2350), .RSTB(I214065), .Q(I214057) );
and I_12473 (I214030,I214362,I214331);
DFFARX1 I_12474  ( .D(I80216), .CLK(I2350), .RSTB(I214065), .Q(I214441) );
nor I_12475 (I214054,I214441,I214362);
nor I_12476 (I214472,I214441,I214116);
nand I_12477 (I214051,I214150,I214472);
not I_12478 (I214048,I214441);
DFFARX1 I_12479  ( .D(I80192), .CLK(I2350), .RSTB(I214065), .Q(I214517) );
not I_12480 (I214534,I214517);
nor I_12481 (I214551,I214534,I214215);
and I_12482 (I214568,I214441,I214551);
or I_12483 (I214585,I214362,I214568);
DFFARX1 I_12484  ( .D(I214585), .CLK(I2350), .RSTB(I214065), .Q(I214042) );
not I_12485 (I214616,I214534);
nor I_12486 (I214633,I214441,I214616);
nand I_12487 (I214045,I214534,I214633);
nand I_12488 (I214039,I214198,I214616);
not I_12489 (I214711,I2357);
not I_12490 (I214728,I23126);
nor I_12491 (I214745,I23141,I23135);
nand I_12492 (I214762,I214745,I23144);
nor I_12493 (I214779,I214728,I23141);
nand I_12494 (I214796,I214779,I23120);
DFFARX1 I_12495  ( .D(I214796), .CLK(I2350), .RSTB(I214711), .Q(I214813) );
not I_12496 (I214682,I214813);
not I_12497 (I214844,I23141);
not I_12498 (I214861,I214844);
not I_12499 (I214878,I23117);
nor I_12500 (I214895,I214878,I23132);
and I_12501 (I214912,I214895,I23138);
or I_12502 (I214929,I214912,I23147);
DFFARX1 I_12503  ( .D(I214929), .CLK(I2350), .RSTB(I214711), .Q(I214946) );
DFFARX1 I_12504  ( .D(I214946), .CLK(I2350), .RSTB(I214711), .Q(I214679) );
DFFARX1 I_12505  ( .D(I214946), .CLK(I2350), .RSTB(I214711), .Q(I214977) );
DFFARX1 I_12506  ( .D(I214946), .CLK(I2350), .RSTB(I214711), .Q(I214673) );
nand I_12507 (I215008,I214728,I23117);
nand I_12508 (I215025,I215008,I214762);
and I_12509 (I215042,I214844,I215025);
DFFARX1 I_12510  ( .D(I215042), .CLK(I2350), .RSTB(I214711), .Q(I214703) );
and I_12511 (I214676,I215008,I214977);
DFFARX1 I_12512  ( .D(I23129), .CLK(I2350), .RSTB(I214711), .Q(I215087) );
nor I_12513 (I214700,I215087,I215008);
nor I_12514 (I215118,I215087,I214762);
nand I_12515 (I214697,I214796,I215118);
not I_12516 (I214694,I215087);
DFFARX1 I_12517  ( .D(I23123), .CLK(I2350), .RSTB(I214711), .Q(I215163) );
not I_12518 (I215180,I215163);
nor I_12519 (I215197,I215180,I214861);
and I_12520 (I215214,I215087,I215197);
or I_12521 (I215231,I215008,I215214);
DFFARX1 I_12522  ( .D(I215231), .CLK(I2350), .RSTB(I214711), .Q(I214688) );
not I_12523 (I215262,I215180);
nor I_12524 (I215279,I215087,I215262);
nand I_12525 (I214691,I215180,I215279);
nand I_12526 (I214685,I214844,I215262);
not I_12527 (I215357,I2357);
not I_12528 (I215374,I360299);
nor I_12529 (I215391,I360296,I360281);
nand I_12530 (I215408,I215391,I360290);
nor I_12531 (I215425,I215374,I360296);
nand I_12532 (I215442,I215425,I360305);
DFFARX1 I_12533  ( .D(I215442), .CLK(I2350), .RSTB(I215357), .Q(I215459) );
not I_12534 (I215328,I215459);
not I_12535 (I215490,I360296);
not I_12536 (I215507,I215490);
not I_12537 (I215524,I360278);
nor I_12538 (I215541,I215524,I360284);
and I_12539 (I215558,I215541,I360308);
or I_12540 (I215575,I215558,I360302);
DFFARX1 I_12541  ( .D(I215575), .CLK(I2350), .RSTB(I215357), .Q(I215592) );
DFFARX1 I_12542  ( .D(I215592), .CLK(I2350), .RSTB(I215357), .Q(I215325) );
DFFARX1 I_12543  ( .D(I215592), .CLK(I2350), .RSTB(I215357), .Q(I215623) );
DFFARX1 I_12544  ( .D(I215592), .CLK(I2350), .RSTB(I215357), .Q(I215319) );
nand I_12545 (I215654,I215374,I360278);
nand I_12546 (I215671,I215654,I215408);
and I_12547 (I215688,I215490,I215671);
DFFARX1 I_12548  ( .D(I215688), .CLK(I2350), .RSTB(I215357), .Q(I215349) );
and I_12549 (I215322,I215654,I215623);
DFFARX1 I_12550  ( .D(I360287), .CLK(I2350), .RSTB(I215357), .Q(I215733) );
nor I_12551 (I215346,I215733,I215654);
nor I_12552 (I215764,I215733,I215408);
nand I_12553 (I215343,I215442,I215764);
not I_12554 (I215340,I215733);
DFFARX1 I_12555  ( .D(I360293), .CLK(I2350), .RSTB(I215357), .Q(I215809) );
not I_12556 (I215826,I215809);
nor I_12557 (I215843,I215826,I215507);
and I_12558 (I215860,I215733,I215843);
or I_12559 (I215877,I215654,I215860);
DFFARX1 I_12560  ( .D(I215877), .CLK(I2350), .RSTB(I215357), .Q(I215334) );
not I_12561 (I215908,I215826);
nor I_12562 (I215925,I215733,I215908);
nand I_12563 (I215337,I215826,I215925);
nand I_12564 (I215331,I215490,I215908);
not I_12565 (I216003,I2357);
not I_12566 (I216020,I364702);
nor I_12567 (I216037,I364699,I364684);
nand I_12568 (I216054,I216037,I364693);
nor I_12569 (I216071,I216020,I364699);
nand I_12570 (I216088,I216071,I364708);
DFFARX1 I_12571  ( .D(I216088), .CLK(I2350), .RSTB(I216003), .Q(I216105) );
not I_12572 (I215974,I216105);
not I_12573 (I216136,I364699);
not I_12574 (I216153,I216136);
not I_12575 (I216170,I364681);
nor I_12576 (I216187,I216170,I364687);
and I_12577 (I216204,I216187,I364711);
or I_12578 (I216221,I216204,I364705);
DFFARX1 I_12579  ( .D(I216221), .CLK(I2350), .RSTB(I216003), .Q(I216238) );
DFFARX1 I_12580  ( .D(I216238), .CLK(I2350), .RSTB(I216003), .Q(I215971) );
DFFARX1 I_12581  ( .D(I216238), .CLK(I2350), .RSTB(I216003), .Q(I216269) );
DFFARX1 I_12582  ( .D(I216238), .CLK(I2350), .RSTB(I216003), .Q(I215965) );
nand I_12583 (I216300,I216020,I364681);
nand I_12584 (I216317,I216300,I216054);
and I_12585 (I216334,I216136,I216317);
DFFARX1 I_12586  ( .D(I216334), .CLK(I2350), .RSTB(I216003), .Q(I215995) );
and I_12587 (I215968,I216300,I216269);
DFFARX1 I_12588  ( .D(I364690), .CLK(I2350), .RSTB(I216003), .Q(I216379) );
nor I_12589 (I215992,I216379,I216300);
nor I_12590 (I216410,I216379,I216054);
nand I_12591 (I215989,I216088,I216410);
not I_12592 (I215986,I216379);
DFFARX1 I_12593  ( .D(I364696), .CLK(I2350), .RSTB(I216003), .Q(I216455) );
not I_12594 (I216472,I216455);
nor I_12595 (I216489,I216472,I216153);
and I_12596 (I216506,I216379,I216489);
or I_12597 (I216523,I216300,I216506);
DFFARX1 I_12598  ( .D(I216523), .CLK(I2350), .RSTB(I216003), .Q(I215980) );
not I_12599 (I216554,I216472);
nor I_12600 (I216571,I216379,I216554);
nand I_12601 (I215983,I216472,I216571);
nand I_12602 (I215977,I216136,I216554);
not I_12603 (I216649,I2357);
not I_12604 (I216666,I295126);
nor I_12605 (I216683,I295138,I295132);
nand I_12606 (I216700,I216683,I295117);
nor I_12607 (I216717,I216666,I295138);
nand I_12608 (I216734,I216717,I295144);
DFFARX1 I_12609  ( .D(I216734), .CLK(I2350), .RSTB(I216649), .Q(I216751) );
not I_12610 (I216620,I216751);
not I_12611 (I216782,I295138);
not I_12612 (I216799,I216782);
not I_12613 (I216816,I295141);
nor I_12614 (I216833,I216816,I295123);
and I_12615 (I216850,I216833,I295120);
or I_12616 (I216867,I216850,I295147);
DFFARX1 I_12617  ( .D(I216867), .CLK(I2350), .RSTB(I216649), .Q(I216884) );
DFFARX1 I_12618  ( .D(I216884), .CLK(I2350), .RSTB(I216649), .Q(I216617) );
DFFARX1 I_12619  ( .D(I216884), .CLK(I2350), .RSTB(I216649), .Q(I216915) );
DFFARX1 I_12620  ( .D(I216884), .CLK(I2350), .RSTB(I216649), .Q(I216611) );
nand I_12621 (I216946,I216666,I295141);
nand I_12622 (I216963,I216946,I216700);
and I_12623 (I216980,I216782,I216963);
DFFARX1 I_12624  ( .D(I216980), .CLK(I2350), .RSTB(I216649), .Q(I216641) );
and I_12625 (I216614,I216946,I216915);
DFFARX1 I_12626  ( .D(I295135), .CLK(I2350), .RSTB(I216649), .Q(I217025) );
nor I_12627 (I216638,I217025,I216946);
nor I_12628 (I217056,I217025,I216700);
nand I_12629 (I216635,I216734,I217056);
not I_12630 (I216632,I217025);
DFFARX1 I_12631  ( .D(I295129), .CLK(I2350), .RSTB(I216649), .Q(I217101) );
not I_12632 (I217118,I217101);
nor I_12633 (I217135,I217118,I216799);
and I_12634 (I217152,I217025,I217135);
or I_12635 (I217169,I216946,I217152);
DFFARX1 I_12636  ( .D(I217169), .CLK(I2350), .RSTB(I216649), .Q(I216626) );
not I_12637 (I217200,I217118);
nor I_12638 (I217217,I217025,I217200);
nand I_12639 (I216629,I217118,I217217);
nand I_12640 (I216623,I216782,I217200);
not I_12641 (I217295,I2357);
not I_12642 (I217312,I105264);
nor I_12643 (I217329,I105285,I105267);
nand I_12644 (I217346,I217329,I105291);
nor I_12645 (I217363,I217312,I105285);
nand I_12646 (I217380,I217363,I105288);
DFFARX1 I_12647  ( .D(I217380), .CLK(I2350), .RSTB(I217295), .Q(I217397) );
not I_12648 (I217266,I217397);
not I_12649 (I217428,I105285);
not I_12650 (I217445,I217428);
not I_12651 (I217462,I105282);
nor I_12652 (I217479,I217462,I105261);
and I_12653 (I217496,I217479,I105273);
or I_12654 (I217513,I217496,I105270);
DFFARX1 I_12655  ( .D(I217513), .CLK(I2350), .RSTB(I217295), .Q(I217530) );
DFFARX1 I_12656  ( .D(I217530), .CLK(I2350), .RSTB(I217295), .Q(I217263) );
DFFARX1 I_12657  ( .D(I217530), .CLK(I2350), .RSTB(I217295), .Q(I217561) );
DFFARX1 I_12658  ( .D(I217530), .CLK(I2350), .RSTB(I217295), .Q(I217257) );
nand I_12659 (I217592,I217312,I105282);
nand I_12660 (I217609,I217592,I217346);
and I_12661 (I217626,I217428,I217609);
DFFARX1 I_12662  ( .D(I217626), .CLK(I2350), .RSTB(I217295), .Q(I217287) );
and I_12663 (I217260,I217592,I217561);
DFFARX1 I_12664  ( .D(I105276), .CLK(I2350), .RSTB(I217295), .Q(I217671) );
nor I_12665 (I217284,I217671,I217592);
nor I_12666 (I217702,I217671,I217346);
nand I_12667 (I217281,I217380,I217702);
not I_12668 (I217278,I217671);
DFFARX1 I_12669  ( .D(I105279), .CLK(I2350), .RSTB(I217295), .Q(I217747) );
not I_12670 (I217764,I217747);
nor I_12671 (I217781,I217764,I217445);
and I_12672 (I217798,I217671,I217781);
or I_12673 (I217815,I217592,I217798);
DFFARX1 I_12674  ( .D(I217815), .CLK(I2350), .RSTB(I217295), .Q(I217272) );
not I_12675 (I217846,I217764);
nor I_12676 (I217863,I217671,I217846);
nand I_12677 (I217275,I217764,I217863);
nand I_12678 (I217269,I217428,I217846);
not I_12679 (I217941,I2357);
not I_12680 (I217958,I389145);
nor I_12681 (I217975,I389130,I389136);
nand I_12682 (I217992,I217975,I389133);
nor I_12683 (I218009,I217958,I389130);
nand I_12684 (I218026,I218009,I389142);
DFFARX1 I_12685  ( .D(I218026), .CLK(I2350), .RSTB(I217941), .Q(I218043) );
not I_12686 (I217912,I218043);
not I_12687 (I218074,I389130);
not I_12688 (I218091,I218074);
not I_12689 (I218108,I389157);
nor I_12690 (I218125,I218108,I389151);
and I_12691 (I218142,I218125,I389148);
or I_12692 (I218159,I218142,I389127);
DFFARX1 I_12693  ( .D(I218159), .CLK(I2350), .RSTB(I217941), .Q(I218176) );
DFFARX1 I_12694  ( .D(I218176), .CLK(I2350), .RSTB(I217941), .Q(I217909) );
DFFARX1 I_12695  ( .D(I218176), .CLK(I2350), .RSTB(I217941), .Q(I218207) );
DFFARX1 I_12696  ( .D(I218176), .CLK(I2350), .RSTB(I217941), .Q(I217903) );
nand I_12697 (I218238,I217958,I389157);
nand I_12698 (I218255,I218238,I217992);
and I_12699 (I218272,I218074,I218255);
DFFARX1 I_12700  ( .D(I218272), .CLK(I2350), .RSTB(I217941), .Q(I217933) );
and I_12701 (I217906,I218238,I218207);
DFFARX1 I_12702  ( .D(I389154), .CLK(I2350), .RSTB(I217941), .Q(I218317) );
nor I_12703 (I217930,I218317,I218238);
nor I_12704 (I218348,I218317,I217992);
nand I_12705 (I217927,I218026,I218348);
not I_12706 (I217924,I218317);
DFFARX1 I_12707  ( .D(I389139), .CLK(I2350), .RSTB(I217941), .Q(I218393) );
not I_12708 (I218410,I218393);
nor I_12709 (I218427,I218410,I218091);
and I_12710 (I218444,I218317,I218427);
or I_12711 (I218461,I218238,I218444);
DFFARX1 I_12712  ( .D(I218461), .CLK(I2350), .RSTB(I217941), .Q(I217918) );
not I_12713 (I218492,I218410);
nor I_12714 (I218509,I218317,I218492);
nand I_12715 (I217921,I218410,I218509);
nand I_12716 (I217915,I218074,I218492);
not I_12717 (I218587,I2357);
not I_12718 (I218604,I60827);
nor I_12719 (I218621,I60818,I60809);
nand I_12720 (I218638,I218621,I60824);
nor I_12721 (I218655,I218604,I60818);
nand I_12722 (I218672,I218655,I60821);
DFFARX1 I_12723  ( .D(I218672), .CLK(I2350), .RSTB(I218587), .Q(I218689) );
not I_12724 (I218558,I218689);
not I_12725 (I218720,I60818);
not I_12726 (I218737,I218720);
not I_12727 (I218754,I60830);
nor I_12728 (I218771,I218754,I60815);
and I_12729 (I218788,I218771,I60833);
or I_12730 (I218805,I218788,I60806);
DFFARX1 I_12731  ( .D(I218805), .CLK(I2350), .RSTB(I218587), .Q(I218822) );
DFFARX1 I_12732  ( .D(I218822), .CLK(I2350), .RSTB(I218587), .Q(I218555) );
DFFARX1 I_12733  ( .D(I218822), .CLK(I2350), .RSTB(I218587), .Q(I218853) );
DFFARX1 I_12734  ( .D(I218822), .CLK(I2350), .RSTB(I218587), .Q(I218549) );
nand I_12735 (I218884,I218604,I60830);
nand I_12736 (I218901,I218884,I218638);
and I_12737 (I218918,I218720,I218901);
DFFARX1 I_12738  ( .D(I218918), .CLK(I2350), .RSTB(I218587), .Q(I218579) );
and I_12739 (I218552,I218884,I218853);
DFFARX1 I_12740  ( .D(I60836), .CLK(I2350), .RSTB(I218587), .Q(I218963) );
nor I_12741 (I218576,I218963,I218884);
nor I_12742 (I218994,I218963,I218638);
nand I_12743 (I218573,I218672,I218994);
not I_12744 (I218570,I218963);
DFFARX1 I_12745  ( .D(I60812), .CLK(I2350), .RSTB(I218587), .Q(I219039) );
not I_12746 (I219056,I219039);
nor I_12747 (I219073,I219056,I218737);
and I_12748 (I219090,I218963,I219073);
or I_12749 (I219107,I218884,I219090);
DFFARX1 I_12750  ( .D(I219107), .CLK(I2350), .RSTB(I218587), .Q(I218564) );
not I_12751 (I219138,I219056);
nor I_12752 (I219155,I218963,I219138);
nand I_12753 (I218567,I219056,I219155);
nand I_12754 (I218561,I218720,I219138);
not I_12755 (I219233,I2357);
not I_12756 (I219250,I95319);
nor I_12757 (I219267,I95340,I95322);
nand I_12758 (I219284,I219267,I95346);
nor I_12759 (I219301,I219250,I95340);
nand I_12760 (I219318,I219301,I95343);
DFFARX1 I_12761  ( .D(I219318), .CLK(I2350), .RSTB(I219233), .Q(I219335) );
not I_12762 (I219204,I219335);
not I_12763 (I219366,I95340);
not I_12764 (I219383,I219366);
not I_12765 (I219400,I95337);
nor I_12766 (I219417,I219400,I95316);
and I_12767 (I219434,I219417,I95328);
or I_12768 (I219451,I219434,I95325);
DFFARX1 I_12769  ( .D(I219451), .CLK(I2350), .RSTB(I219233), .Q(I219468) );
DFFARX1 I_12770  ( .D(I219468), .CLK(I2350), .RSTB(I219233), .Q(I219201) );
DFFARX1 I_12771  ( .D(I219468), .CLK(I2350), .RSTB(I219233), .Q(I219499) );
DFFARX1 I_12772  ( .D(I219468), .CLK(I2350), .RSTB(I219233), .Q(I219195) );
nand I_12773 (I219530,I219250,I95337);
nand I_12774 (I219547,I219530,I219284);
and I_12775 (I219564,I219366,I219547);
DFFARX1 I_12776  ( .D(I219564), .CLK(I2350), .RSTB(I219233), .Q(I219225) );
and I_12777 (I219198,I219530,I219499);
DFFARX1 I_12778  ( .D(I95331), .CLK(I2350), .RSTB(I219233), .Q(I219609) );
nor I_12779 (I219222,I219609,I219530);
nor I_12780 (I219640,I219609,I219284);
nand I_12781 (I219219,I219318,I219640);
not I_12782 (I219216,I219609);
DFFARX1 I_12783  ( .D(I95334), .CLK(I2350), .RSTB(I219233), .Q(I219685) );
not I_12784 (I219702,I219685);
nor I_12785 (I219719,I219702,I219383);
and I_12786 (I219736,I219609,I219719);
or I_12787 (I219753,I219530,I219736);
DFFARX1 I_12788  ( .D(I219753), .CLK(I2350), .RSTB(I219233), .Q(I219210) );
not I_12789 (I219784,I219702);
nor I_12790 (I219801,I219609,I219784);
nand I_12791 (I219213,I219702,I219801);
nand I_12792 (I219207,I219366,I219784);
not I_12793 (I219879,I2357);
not I_12794 (I219896,I342058);
nor I_12795 (I219913,I342055,I342040);
nand I_12796 (I219930,I219913,I342049);
nor I_12797 (I219947,I219896,I342055);
nand I_12798 (I219964,I219947,I342064);
DFFARX1 I_12799  ( .D(I219964), .CLK(I2350), .RSTB(I219879), .Q(I219981) );
not I_12800 (I219850,I219981);
not I_12801 (I220012,I342055);
not I_12802 (I220029,I220012);
not I_12803 (I220046,I342037);
nor I_12804 (I220063,I220046,I342043);
and I_12805 (I220080,I220063,I342067);
or I_12806 (I220097,I220080,I342061);
DFFARX1 I_12807  ( .D(I220097), .CLK(I2350), .RSTB(I219879), .Q(I220114) );
DFFARX1 I_12808  ( .D(I220114), .CLK(I2350), .RSTB(I219879), .Q(I219847) );
DFFARX1 I_12809  ( .D(I220114), .CLK(I2350), .RSTB(I219879), .Q(I220145) );
DFFARX1 I_12810  ( .D(I220114), .CLK(I2350), .RSTB(I219879), .Q(I219841) );
nand I_12811 (I220176,I219896,I342037);
nand I_12812 (I220193,I220176,I219930);
and I_12813 (I220210,I220012,I220193);
DFFARX1 I_12814  ( .D(I220210), .CLK(I2350), .RSTB(I219879), .Q(I219871) );
and I_12815 (I219844,I220176,I220145);
DFFARX1 I_12816  ( .D(I342046), .CLK(I2350), .RSTB(I219879), .Q(I220255) );
nor I_12817 (I219868,I220255,I220176);
nor I_12818 (I220286,I220255,I219930);
nand I_12819 (I219865,I219964,I220286);
not I_12820 (I219862,I220255);
DFFARX1 I_12821  ( .D(I342052), .CLK(I2350), .RSTB(I219879), .Q(I220331) );
not I_12822 (I220348,I220331);
nor I_12823 (I220365,I220348,I220029);
and I_12824 (I220382,I220255,I220365);
or I_12825 (I220399,I220176,I220382);
DFFARX1 I_12826  ( .D(I220399), .CLK(I2350), .RSTB(I219879), .Q(I219856) );
not I_12827 (I220430,I220348);
nor I_12828 (I220447,I220255,I220430);
nand I_12829 (I219859,I220348,I220447);
nand I_12830 (I219853,I220012,I220430);
not I_12831 (I220525,I2357);
not I_12832 (I220542,I25943);
nor I_12833 (I220559,I25934,I25925);
nand I_12834 (I220576,I220559,I25940);
nor I_12835 (I220593,I220542,I25934);
nand I_12836 (I220610,I220593,I25937);
DFFARX1 I_12837  ( .D(I220610), .CLK(I2350), .RSTB(I220525), .Q(I220627) );
not I_12838 (I220496,I220627);
not I_12839 (I220658,I25934);
not I_12840 (I220675,I220658);
not I_12841 (I220692,I25946);
nor I_12842 (I220709,I220692,I25931);
and I_12843 (I220726,I220709,I25949);
or I_12844 (I220743,I220726,I25922);
DFFARX1 I_12845  ( .D(I220743), .CLK(I2350), .RSTB(I220525), .Q(I220760) );
DFFARX1 I_12846  ( .D(I220760), .CLK(I2350), .RSTB(I220525), .Q(I220493) );
DFFARX1 I_12847  ( .D(I220760), .CLK(I2350), .RSTB(I220525), .Q(I220791) );
DFFARX1 I_12848  ( .D(I220760), .CLK(I2350), .RSTB(I220525), .Q(I220487) );
nand I_12849 (I220822,I220542,I25946);
nand I_12850 (I220839,I220822,I220576);
and I_12851 (I220856,I220658,I220839);
DFFARX1 I_12852  ( .D(I220856), .CLK(I2350), .RSTB(I220525), .Q(I220517) );
and I_12853 (I220490,I220822,I220791);
DFFARX1 I_12854  ( .D(I25952), .CLK(I2350), .RSTB(I220525), .Q(I220901) );
nor I_12855 (I220514,I220901,I220822);
nor I_12856 (I220932,I220901,I220576);
nand I_12857 (I220511,I220610,I220932);
not I_12858 (I220508,I220901);
DFFARX1 I_12859  ( .D(I25928), .CLK(I2350), .RSTB(I220525), .Q(I220977) );
not I_12860 (I220994,I220977);
nor I_12861 (I221011,I220994,I220675);
and I_12862 (I221028,I220901,I221011);
or I_12863 (I221045,I220822,I221028);
DFFARX1 I_12864  ( .D(I221045), .CLK(I2350), .RSTB(I220525), .Q(I220502) );
not I_12865 (I221076,I220994);
nor I_12866 (I221093,I220901,I221076);
nand I_12867 (I220505,I220994,I221093);
nand I_12868 (I220499,I220658,I221076);
not I_12869 (I221171,I2357);
not I_12870 (I221188,I167539);
nor I_12871 (I221205,I167518,I167530);
nand I_12872 (I221222,I221205,I167533);
nor I_12873 (I221239,I221188,I167518);
nand I_12874 (I221256,I221239,I167515);
DFFARX1 I_12875  ( .D(I221256), .CLK(I2350), .RSTB(I221171), .Q(I221273) );
not I_12876 (I221142,I221273);
not I_12877 (I221304,I167518);
not I_12878 (I221321,I221304);
not I_12879 (I221338,I167536);
nor I_12880 (I221355,I221338,I167527);
and I_12881 (I221372,I221355,I167521);
or I_12882 (I221389,I221372,I167545);
DFFARX1 I_12883  ( .D(I221389), .CLK(I2350), .RSTB(I221171), .Q(I221406) );
DFFARX1 I_12884  ( .D(I221406), .CLK(I2350), .RSTB(I221171), .Q(I221139) );
DFFARX1 I_12885  ( .D(I221406), .CLK(I2350), .RSTB(I221171), .Q(I221437) );
DFFARX1 I_12886  ( .D(I221406), .CLK(I2350), .RSTB(I221171), .Q(I221133) );
nand I_12887 (I221468,I221188,I167536);
nand I_12888 (I221485,I221468,I221222);
and I_12889 (I221502,I221304,I221485);
DFFARX1 I_12890  ( .D(I221502), .CLK(I2350), .RSTB(I221171), .Q(I221163) );
and I_12891 (I221136,I221468,I221437);
DFFARX1 I_12892  ( .D(I167542), .CLK(I2350), .RSTB(I221171), .Q(I221547) );
nor I_12893 (I221160,I221547,I221468);
nor I_12894 (I221578,I221547,I221222);
nand I_12895 (I221157,I221256,I221578);
not I_12896 (I221154,I221547);
DFFARX1 I_12897  ( .D(I167524), .CLK(I2350), .RSTB(I221171), .Q(I221623) );
not I_12898 (I221640,I221623);
nor I_12899 (I221657,I221640,I221321);
and I_12900 (I221674,I221547,I221657);
or I_12901 (I221691,I221468,I221674);
DFFARX1 I_12902  ( .D(I221691), .CLK(I2350), .RSTB(I221171), .Q(I221148) );
not I_12903 (I221722,I221640);
nor I_12904 (I221739,I221547,I221722);
nand I_12905 (I221151,I221640,I221739);
nand I_12906 (I221145,I221304,I221722);
not I_12907 (I221817,I2357);
not I_12908 (I221834,I95982);
nor I_12909 (I221851,I96003,I95985);
nand I_12910 (I221868,I221851,I96009);
nor I_12911 (I221885,I221834,I96003);
nand I_12912 (I221902,I221885,I96006);
DFFARX1 I_12913  ( .D(I221902), .CLK(I2350), .RSTB(I221817), .Q(I221919) );
not I_12914 (I221788,I221919);
not I_12915 (I221950,I96003);
not I_12916 (I221967,I221950);
not I_12917 (I221984,I96000);
nor I_12918 (I222001,I221984,I95979);
and I_12919 (I222018,I222001,I95991);
or I_12920 (I222035,I222018,I95988);
DFFARX1 I_12921  ( .D(I222035), .CLK(I2350), .RSTB(I221817), .Q(I222052) );
DFFARX1 I_12922  ( .D(I222052), .CLK(I2350), .RSTB(I221817), .Q(I221785) );
DFFARX1 I_12923  ( .D(I222052), .CLK(I2350), .RSTB(I221817), .Q(I222083) );
DFFARX1 I_12924  ( .D(I222052), .CLK(I2350), .RSTB(I221817), .Q(I221779) );
nand I_12925 (I222114,I221834,I96000);
nand I_12926 (I222131,I222114,I221868);
and I_12927 (I222148,I221950,I222131);
DFFARX1 I_12928  ( .D(I222148), .CLK(I2350), .RSTB(I221817), .Q(I221809) );
and I_12929 (I221782,I222114,I222083);
DFFARX1 I_12930  ( .D(I95994), .CLK(I2350), .RSTB(I221817), .Q(I222193) );
nor I_12931 (I221806,I222193,I222114);
nor I_12932 (I222224,I222193,I221868);
nand I_12933 (I221803,I221902,I222224);
not I_12934 (I221800,I222193);
DFFARX1 I_12935  ( .D(I95997), .CLK(I2350), .RSTB(I221817), .Q(I222269) );
not I_12936 (I222286,I222269);
nor I_12937 (I222303,I222286,I221967);
and I_12938 (I222320,I222193,I222303);
or I_12939 (I222337,I222114,I222320);
DFFARX1 I_12940  ( .D(I222337), .CLK(I2350), .RSTB(I221817), .Q(I221794) );
not I_12941 (I222368,I222286);
nor I_12942 (I222385,I222193,I222368);
nand I_12943 (I221797,I222286,I222385);
nand I_12944 (I221791,I221950,I222368);
not I_12945 (I222463,I2357);
not I_12946 (I222480,I170191);
nor I_12947 (I222497,I170170,I170182);
nand I_12948 (I222514,I222497,I170185);
nor I_12949 (I222531,I222480,I170170);
nand I_12950 (I222548,I222531,I170167);
DFFARX1 I_12951  ( .D(I222548), .CLK(I2350), .RSTB(I222463), .Q(I222565) );
not I_12952 (I222434,I222565);
not I_12953 (I222596,I170170);
not I_12954 (I222613,I222596);
not I_12955 (I222630,I170188);
nor I_12956 (I222647,I222630,I170179);
and I_12957 (I222664,I222647,I170173);
or I_12958 (I222681,I222664,I170197);
DFFARX1 I_12959  ( .D(I222681), .CLK(I2350), .RSTB(I222463), .Q(I222698) );
DFFARX1 I_12960  ( .D(I222698), .CLK(I2350), .RSTB(I222463), .Q(I222431) );
DFFARX1 I_12961  ( .D(I222698), .CLK(I2350), .RSTB(I222463), .Q(I222729) );
DFFARX1 I_12962  ( .D(I222698), .CLK(I2350), .RSTB(I222463), .Q(I222425) );
nand I_12963 (I222760,I222480,I170188);
nand I_12964 (I222777,I222760,I222514);
and I_12965 (I222794,I222596,I222777);
DFFARX1 I_12966  ( .D(I222794), .CLK(I2350), .RSTB(I222463), .Q(I222455) );
and I_12967 (I222428,I222760,I222729);
DFFARX1 I_12968  ( .D(I170194), .CLK(I2350), .RSTB(I222463), .Q(I222839) );
nor I_12969 (I222452,I222839,I222760);
nor I_12970 (I222870,I222839,I222514);
nand I_12971 (I222449,I222548,I222870);
not I_12972 (I222446,I222839);
DFFARX1 I_12973  ( .D(I170176), .CLK(I2350), .RSTB(I222463), .Q(I222915) );
not I_12974 (I222932,I222915);
nor I_12975 (I222949,I222932,I222613);
and I_12976 (I222966,I222839,I222949);
or I_12977 (I222983,I222760,I222966);
DFFARX1 I_12978  ( .D(I222983), .CLK(I2350), .RSTB(I222463), .Q(I222440) );
not I_12979 (I223014,I222932);
nor I_12980 (I223031,I222839,I223014);
nand I_12981 (I222443,I222932,I223031);
nand I_12982 (I222437,I222596,I223014);
not I_12983 (I223109,I2357);
not I_12984 (I223126,I346461);
nor I_12985 (I223143,I346458,I346443);
nand I_12986 (I223160,I223143,I346452);
nor I_12987 (I223177,I223126,I346458);
nand I_12988 (I223194,I223177,I346467);
DFFARX1 I_12989  ( .D(I223194), .CLK(I2350), .RSTB(I223109), .Q(I223211) );
not I_12990 (I223080,I223211);
not I_12991 (I223242,I346458);
not I_12992 (I223259,I223242);
not I_12993 (I223276,I346440);
nor I_12994 (I223293,I223276,I346446);
and I_12995 (I223310,I223293,I346470);
or I_12996 (I223327,I223310,I346464);
DFFARX1 I_12997  ( .D(I223327), .CLK(I2350), .RSTB(I223109), .Q(I223344) );
DFFARX1 I_12998  ( .D(I223344), .CLK(I2350), .RSTB(I223109), .Q(I223077) );
DFFARX1 I_12999  ( .D(I223344), .CLK(I2350), .RSTB(I223109), .Q(I223375) );
DFFARX1 I_13000  ( .D(I223344), .CLK(I2350), .RSTB(I223109), .Q(I223071) );
nand I_13001 (I223406,I223126,I346440);
nand I_13002 (I223423,I223406,I223160);
and I_13003 (I223440,I223242,I223423);
DFFARX1 I_13004  ( .D(I223440), .CLK(I2350), .RSTB(I223109), .Q(I223101) );
and I_13005 (I223074,I223406,I223375);
DFFARX1 I_13006  ( .D(I346449), .CLK(I2350), .RSTB(I223109), .Q(I223485) );
nor I_13007 (I223098,I223485,I223406);
nor I_13008 (I223516,I223485,I223160);
nand I_13009 (I223095,I223194,I223516);
not I_13010 (I223092,I223485);
DFFARX1 I_13011  ( .D(I346455), .CLK(I2350), .RSTB(I223109), .Q(I223561) );
not I_13012 (I223578,I223561);
nor I_13013 (I223595,I223578,I223259);
and I_13014 (I223612,I223485,I223595);
or I_13015 (I223629,I223406,I223612);
DFFARX1 I_13016  ( .D(I223629), .CLK(I2350), .RSTB(I223109), .Q(I223086) );
not I_13017 (I223660,I223578);
nor I_13018 (I223677,I223485,I223660);
nand I_13019 (I223089,I223578,I223677);
nand I_13020 (I223083,I223242,I223660);
not I_13021 (I223755,I2357);
not I_13022 (I223772,I154279);
nor I_13023 (I223789,I154258,I154270);
nand I_13024 (I223806,I223789,I154273);
nor I_13025 (I223823,I223772,I154258);
nand I_13026 (I223840,I223823,I154255);
DFFARX1 I_13027  ( .D(I223840), .CLK(I2350), .RSTB(I223755), .Q(I223857) );
not I_13028 (I223726,I223857);
not I_13029 (I223888,I154258);
not I_13030 (I223905,I223888);
not I_13031 (I223922,I154276);
nor I_13032 (I223939,I223922,I154267);
and I_13033 (I223956,I223939,I154261);
or I_13034 (I223973,I223956,I154285);
DFFARX1 I_13035  ( .D(I223973), .CLK(I2350), .RSTB(I223755), .Q(I223990) );
DFFARX1 I_13036  ( .D(I223990), .CLK(I2350), .RSTB(I223755), .Q(I223723) );
DFFARX1 I_13037  ( .D(I223990), .CLK(I2350), .RSTB(I223755), .Q(I224021) );
DFFARX1 I_13038  ( .D(I223990), .CLK(I2350), .RSTB(I223755), .Q(I223717) );
nand I_13039 (I224052,I223772,I154276);
nand I_13040 (I224069,I224052,I223806);
and I_13041 (I224086,I223888,I224069);
DFFARX1 I_13042  ( .D(I224086), .CLK(I2350), .RSTB(I223755), .Q(I223747) );
and I_13043 (I223720,I224052,I224021);
DFFARX1 I_13044  ( .D(I154282), .CLK(I2350), .RSTB(I223755), .Q(I224131) );
nor I_13045 (I223744,I224131,I224052);
nor I_13046 (I224162,I224131,I223806);
nand I_13047 (I223741,I223840,I224162);
not I_13048 (I223738,I224131);
DFFARX1 I_13049  ( .D(I154264), .CLK(I2350), .RSTB(I223755), .Q(I224207) );
not I_13050 (I224224,I224207);
nor I_13051 (I224241,I224224,I223905);
and I_13052 (I224258,I224131,I224241);
or I_13053 (I224275,I224052,I224258);
DFFARX1 I_13054  ( .D(I224275), .CLK(I2350), .RSTB(I223755), .Q(I223732) );
not I_13055 (I224306,I224224);
nor I_13056 (I224323,I224131,I224306);
nand I_13057 (I223735,I224224,I224323);
nand I_13058 (I223729,I223888,I224306);
not I_13059 (I224401,I2357);
not I_13060 (I224418,I234615);
nor I_13061 (I224435,I234624,I234609);
nand I_13062 (I224452,I224435,I234597);
nor I_13063 (I224469,I224418,I234624);
nand I_13064 (I224486,I224469,I234600);
DFFARX1 I_13065  ( .D(I224486), .CLK(I2350), .RSTB(I224401), .Q(I224503) );
not I_13066 (I224372,I224503);
not I_13067 (I224534,I234624);
not I_13068 (I224551,I224534);
not I_13069 (I224568,I234612);
nor I_13070 (I224585,I224568,I234606);
and I_13071 (I224602,I224585,I234603);
or I_13072 (I224619,I224602,I234618);
DFFARX1 I_13073  ( .D(I224619), .CLK(I2350), .RSTB(I224401), .Q(I224636) );
DFFARX1 I_13074  ( .D(I224636), .CLK(I2350), .RSTB(I224401), .Q(I224369) );
DFFARX1 I_13075  ( .D(I224636), .CLK(I2350), .RSTB(I224401), .Q(I224667) );
DFFARX1 I_13076  ( .D(I224636), .CLK(I2350), .RSTB(I224401), .Q(I224363) );
nand I_13077 (I224698,I224418,I234612);
nand I_13078 (I224715,I224698,I224452);
and I_13079 (I224732,I224534,I224715);
DFFARX1 I_13080  ( .D(I224732), .CLK(I2350), .RSTB(I224401), .Q(I224393) );
and I_13081 (I224366,I224698,I224667);
DFFARX1 I_13082  ( .D(I234627), .CLK(I2350), .RSTB(I224401), .Q(I224777) );
nor I_13083 (I224390,I224777,I224698);
nor I_13084 (I224808,I224777,I224452);
nand I_13085 (I224387,I224486,I224808);
not I_13086 (I224384,I224777);
DFFARX1 I_13087  ( .D(I234621), .CLK(I2350), .RSTB(I224401), .Q(I224853) );
not I_13088 (I224870,I224853);
nor I_13089 (I224887,I224870,I224551);
and I_13090 (I224904,I224777,I224887);
or I_13091 (I224921,I224698,I224904);
DFFARX1 I_13092  ( .D(I224921), .CLK(I2350), .RSTB(I224401), .Q(I224378) );
not I_13093 (I224952,I224870);
nor I_13094 (I224969,I224777,I224952);
nand I_13095 (I224381,I224870,I224969);
nand I_13096 (I224375,I224534,I224952);
not I_13097 (I225047,I2357);
not I_13098 (I225064,I13028);
nor I_13099 (I225081,I13043,I13037);
nand I_13100 (I225098,I225081,I13046);
nor I_13101 (I225115,I225064,I13043);
nand I_13102 (I225132,I225115,I13022);
DFFARX1 I_13103  ( .D(I225132), .CLK(I2350), .RSTB(I225047), .Q(I225149) );
not I_13104 (I225018,I225149);
not I_13105 (I225180,I13043);
not I_13106 (I225197,I225180);
not I_13107 (I225214,I13019);
nor I_13108 (I225231,I225214,I13034);
and I_13109 (I225248,I225231,I13040);
or I_13110 (I225265,I225248,I13049);
DFFARX1 I_13111  ( .D(I225265), .CLK(I2350), .RSTB(I225047), .Q(I225282) );
DFFARX1 I_13112  ( .D(I225282), .CLK(I2350), .RSTB(I225047), .Q(I225015) );
DFFARX1 I_13113  ( .D(I225282), .CLK(I2350), .RSTB(I225047), .Q(I225313) );
DFFARX1 I_13114  ( .D(I225282), .CLK(I2350), .RSTB(I225047), .Q(I225009) );
nand I_13115 (I225344,I225064,I13019);
nand I_13116 (I225361,I225344,I225098);
and I_13117 (I225378,I225180,I225361);
DFFARX1 I_13118  ( .D(I225378), .CLK(I2350), .RSTB(I225047), .Q(I225039) );
and I_13119 (I225012,I225344,I225313);
DFFARX1 I_13120  ( .D(I13031), .CLK(I2350), .RSTB(I225047), .Q(I225423) );
nor I_13121 (I225036,I225423,I225344);
nor I_13122 (I225454,I225423,I225098);
nand I_13123 (I225033,I225132,I225454);
not I_13124 (I225030,I225423);
DFFARX1 I_13125  ( .D(I13025), .CLK(I2350), .RSTB(I225047), .Q(I225499) );
not I_13126 (I225516,I225499);
nor I_13127 (I225533,I225516,I225197);
and I_13128 (I225550,I225423,I225533);
or I_13129 (I225567,I225344,I225550);
DFFARX1 I_13130  ( .D(I225567), .CLK(I2350), .RSTB(I225047), .Q(I225024) );
not I_13131 (I225598,I225516);
nor I_13132 (I225615,I225423,I225598);
nand I_13133 (I225027,I225516,I225615);
nand I_13134 (I225021,I225180,I225598);
not I_13135 (I225693,I2357);
not I_13136 (I225710,I121621);
nor I_13137 (I225727,I121627,I121624);
nand I_13138 (I225744,I225727,I121618);
nor I_13139 (I225761,I225710,I121627);
nand I_13140 (I225778,I225761,I121642);
DFFARX1 I_13141  ( .D(I225778), .CLK(I2350), .RSTB(I225693), .Q(I225795) );
not I_13142 (I225664,I225795);
not I_13143 (I225826,I121627);
not I_13144 (I225843,I225826);
not I_13145 (I225860,I121639);
nor I_13146 (I225877,I225860,I121630);
and I_13147 (I225894,I225877,I121615);
or I_13148 (I225911,I225894,I121636);
DFFARX1 I_13149  ( .D(I225911), .CLK(I2350), .RSTB(I225693), .Q(I225928) );
DFFARX1 I_13150  ( .D(I225928), .CLK(I2350), .RSTB(I225693), .Q(I225661) );
DFFARX1 I_13151  ( .D(I225928), .CLK(I2350), .RSTB(I225693), .Q(I225959) );
DFFARX1 I_13152  ( .D(I225928), .CLK(I2350), .RSTB(I225693), .Q(I225655) );
nand I_13153 (I225990,I225710,I121639);
nand I_13154 (I226007,I225990,I225744);
and I_13155 (I226024,I225826,I226007);
DFFARX1 I_13156  ( .D(I226024), .CLK(I2350), .RSTB(I225693), .Q(I225685) );
and I_13157 (I225658,I225990,I225959);
DFFARX1 I_13158  ( .D(I121633), .CLK(I2350), .RSTB(I225693), .Q(I226069) );
nor I_13159 (I225682,I226069,I225990);
nor I_13160 (I226100,I226069,I225744);
nand I_13161 (I225679,I225778,I226100);
not I_13162 (I225676,I226069);
DFFARX1 I_13163  ( .D(I121645), .CLK(I2350), .RSTB(I225693), .Q(I226145) );
not I_13164 (I226162,I226145);
nor I_13165 (I226179,I226162,I225843);
and I_13166 (I226196,I226069,I226179);
or I_13167 (I226213,I225990,I226196);
DFFARX1 I_13168  ( .D(I226213), .CLK(I2350), .RSTB(I225693), .Q(I225670) );
not I_13169 (I226244,I226162);
nor I_13170 (I226261,I226069,I226244);
nand I_13171 (I225673,I226162,I226261);
nand I_13172 (I225667,I225826,I226244);
not I_13173 (I226339,I2357);
not I_13174 (I226356,I174169);
nor I_13175 (I226373,I174148,I174160);
nand I_13176 (I226390,I226373,I174163);
nor I_13177 (I226407,I226356,I174148);
nand I_13178 (I226424,I226407,I174145);
DFFARX1 I_13179  ( .D(I226424), .CLK(I2350), .RSTB(I226339), .Q(I226441) );
not I_13180 (I226310,I226441);
not I_13181 (I226472,I174148);
not I_13182 (I226489,I226472);
not I_13183 (I226506,I174166);
nor I_13184 (I226523,I226506,I174157);
and I_13185 (I226540,I226523,I174151);
or I_13186 (I226557,I226540,I174175);
DFFARX1 I_13187  ( .D(I226557), .CLK(I2350), .RSTB(I226339), .Q(I226574) );
DFFARX1 I_13188  ( .D(I226574), .CLK(I2350), .RSTB(I226339), .Q(I226307) );
DFFARX1 I_13189  ( .D(I226574), .CLK(I2350), .RSTB(I226339), .Q(I226605) );
DFFARX1 I_13190  ( .D(I226574), .CLK(I2350), .RSTB(I226339), .Q(I226301) );
nand I_13191 (I226636,I226356,I174166);
nand I_13192 (I226653,I226636,I226390);
and I_13193 (I226670,I226472,I226653);
DFFARX1 I_13194  ( .D(I226670), .CLK(I2350), .RSTB(I226339), .Q(I226331) );
and I_13195 (I226304,I226636,I226605);
DFFARX1 I_13196  ( .D(I174172), .CLK(I2350), .RSTB(I226339), .Q(I226715) );
nor I_13197 (I226328,I226715,I226636);
nor I_13198 (I226746,I226715,I226390);
nand I_13199 (I226325,I226424,I226746);
not I_13200 (I226322,I226715);
DFFARX1 I_13201  ( .D(I174154), .CLK(I2350), .RSTB(I226339), .Q(I226791) );
not I_13202 (I226808,I226791);
nor I_13203 (I226825,I226808,I226489);
and I_13204 (I226842,I226715,I226825);
or I_13205 (I226859,I226636,I226842);
DFFARX1 I_13206  ( .D(I226859), .CLK(I2350), .RSTB(I226339), .Q(I226316) );
not I_13207 (I226890,I226808);
nor I_13208 (I226907,I226715,I226890);
nand I_13209 (I226319,I226808,I226907);
nand I_13210 (I226313,I226472,I226890);
not I_13211 (I226985,I2357);
not I_13212 (I227002,I172180);
nor I_13213 (I227019,I172159,I172171);
nand I_13214 (I227036,I227019,I172174);
nor I_13215 (I227053,I227002,I172159);
nand I_13216 (I227070,I227053,I172156);
DFFARX1 I_13217  ( .D(I227070), .CLK(I2350), .RSTB(I226985), .Q(I227087) );
not I_13218 (I226956,I227087);
not I_13219 (I227118,I172159);
not I_13220 (I227135,I227118);
not I_13221 (I227152,I172177);
nor I_13222 (I227169,I227152,I172168);
and I_13223 (I227186,I227169,I172162);
or I_13224 (I227203,I227186,I172186);
DFFARX1 I_13225  ( .D(I227203), .CLK(I2350), .RSTB(I226985), .Q(I227220) );
DFFARX1 I_13226  ( .D(I227220), .CLK(I2350), .RSTB(I226985), .Q(I226953) );
DFFARX1 I_13227  ( .D(I227220), .CLK(I2350), .RSTB(I226985), .Q(I227251) );
DFFARX1 I_13228  ( .D(I227220), .CLK(I2350), .RSTB(I226985), .Q(I226947) );
nand I_13229 (I227282,I227002,I172177);
nand I_13230 (I227299,I227282,I227036);
and I_13231 (I227316,I227118,I227299);
DFFARX1 I_13232  ( .D(I227316), .CLK(I2350), .RSTB(I226985), .Q(I226977) );
and I_13233 (I226950,I227282,I227251);
DFFARX1 I_13234  ( .D(I172183), .CLK(I2350), .RSTB(I226985), .Q(I227361) );
nor I_13235 (I226974,I227361,I227282);
nor I_13236 (I227392,I227361,I227036);
nand I_13237 (I226971,I227070,I227392);
not I_13238 (I226968,I227361);
DFFARX1 I_13239  ( .D(I172165), .CLK(I2350), .RSTB(I226985), .Q(I227437) );
not I_13240 (I227454,I227437);
nor I_13241 (I227471,I227454,I227135);
and I_13242 (I227488,I227361,I227471);
or I_13243 (I227505,I227282,I227488);
DFFARX1 I_13244  ( .D(I227505), .CLK(I2350), .RSTB(I226985), .Q(I226962) );
not I_13245 (I227536,I227454);
nor I_13246 (I227553,I227361,I227536);
nand I_13247 (I226965,I227454,I227553);
nand I_13248 (I226959,I227118,I227536);
not I_13249 (I227631,I2357);
not I_13250 (I227648,I376024);
nor I_13251 (I227665,I376021,I376006);
nand I_13252 (I227682,I227665,I376015);
nor I_13253 (I227699,I227648,I376021);
nand I_13254 (I227716,I227699,I376030);
DFFARX1 I_13255  ( .D(I227716), .CLK(I2350), .RSTB(I227631), .Q(I227733) );
not I_13256 (I227602,I227733);
not I_13257 (I227764,I376021);
not I_13258 (I227781,I227764);
not I_13259 (I227798,I376003);
nor I_13260 (I227815,I227798,I376009);
and I_13261 (I227832,I227815,I376033);
or I_13262 (I227849,I227832,I376027);
DFFARX1 I_13263  ( .D(I227849), .CLK(I2350), .RSTB(I227631), .Q(I227866) );
DFFARX1 I_13264  ( .D(I227866), .CLK(I2350), .RSTB(I227631), .Q(I227599) );
DFFARX1 I_13265  ( .D(I227866), .CLK(I2350), .RSTB(I227631), .Q(I227897) );
DFFARX1 I_13266  ( .D(I227866), .CLK(I2350), .RSTB(I227631), .Q(I227593) );
nand I_13267 (I227928,I227648,I376003);
nand I_13268 (I227945,I227928,I227682);
and I_13269 (I227962,I227764,I227945);
DFFARX1 I_13270  ( .D(I227962), .CLK(I2350), .RSTB(I227631), .Q(I227623) );
and I_13271 (I227596,I227928,I227897);
DFFARX1 I_13272  ( .D(I376012), .CLK(I2350), .RSTB(I227631), .Q(I228007) );
nor I_13273 (I227620,I228007,I227928);
nor I_13274 (I228038,I228007,I227682);
nand I_13275 (I227617,I227716,I228038);
not I_13276 (I227614,I228007);
DFFARX1 I_13277  ( .D(I376018), .CLK(I2350), .RSTB(I227631), .Q(I228083) );
not I_13278 (I228100,I228083);
nor I_13279 (I228117,I228100,I227781);
and I_13280 (I228134,I228007,I228117);
or I_13281 (I228151,I227928,I228134);
DFFARX1 I_13282  ( .D(I228151), .CLK(I2350), .RSTB(I227631), .Q(I227608) );
not I_13283 (I228182,I228100);
nor I_13284 (I228199,I228007,I228182);
nand I_13285 (I227611,I228100,I228199);
nand I_13286 (I227605,I227764,I228182);
not I_13287 (I228277,I2357);
not I_13288 (I228294,I343316);
nor I_13289 (I228311,I343313,I343298);
nand I_13290 (I228328,I228311,I343307);
nor I_13291 (I228345,I228294,I343313);
nand I_13292 (I228362,I228345,I343322);
DFFARX1 I_13293  ( .D(I228362), .CLK(I2350), .RSTB(I228277), .Q(I228379) );
not I_13294 (I228248,I228379);
not I_13295 (I228410,I343313);
not I_13296 (I228427,I228410);
not I_13297 (I228444,I343295);
nor I_13298 (I228461,I228444,I343301);
and I_13299 (I228478,I228461,I343325);
or I_13300 (I228495,I228478,I343319);
DFFARX1 I_13301  ( .D(I228495), .CLK(I2350), .RSTB(I228277), .Q(I228512) );
DFFARX1 I_13302  ( .D(I228512), .CLK(I2350), .RSTB(I228277), .Q(I228245) );
DFFARX1 I_13303  ( .D(I228512), .CLK(I2350), .RSTB(I228277), .Q(I228543) );
DFFARX1 I_13304  ( .D(I228512), .CLK(I2350), .RSTB(I228277), .Q(I228239) );
nand I_13305 (I228574,I228294,I343295);
nand I_13306 (I228591,I228574,I228328);
and I_13307 (I228608,I228410,I228591);
DFFARX1 I_13308  ( .D(I228608), .CLK(I2350), .RSTB(I228277), .Q(I228269) );
and I_13309 (I228242,I228574,I228543);
DFFARX1 I_13310  ( .D(I343304), .CLK(I2350), .RSTB(I228277), .Q(I228653) );
nor I_13311 (I228266,I228653,I228574);
nor I_13312 (I228684,I228653,I228328);
nand I_13313 (I228263,I228362,I228684);
not I_13314 (I228260,I228653);
DFFARX1 I_13315  ( .D(I343310), .CLK(I2350), .RSTB(I228277), .Q(I228729) );
not I_13316 (I228746,I228729);
nor I_13317 (I228763,I228746,I228427);
and I_13318 (I228780,I228653,I228763);
or I_13319 (I228797,I228574,I228780);
DFFARX1 I_13320  ( .D(I228797), .CLK(I2350), .RSTB(I228277), .Q(I228254) );
not I_13321 (I228828,I228746);
nor I_13322 (I228845,I228653,I228828);
nand I_13323 (I228257,I228746,I228845);
nand I_13324 (I228251,I228410,I228828);
not I_13325 (I228923,I2357);
not I_13326 (I228940,I134125);
nor I_13327 (I228957,I134113,I134116);
nand I_13328 (I228974,I228957,I134140);
nor I_13329 (I228991,I228940,I134113);
nand I_13330 (I229008,I228991,I134122);
DFFARX1 I_13331  ( .D(I229008), .CLK(I2350), .RSTB(I228923), .Q(I229025) );
not I_13332 (I228894,I229025);
not I_13333 (I229056,I134113);
not I_13334 (I229073,I229056);
not I_13335 (I229090,I134119);
nor I_13336 (I229107,I229090,I134134);
and I_13337 (I229124,I229107,I134110);
or I_13338 (I229141,I229124,I134137);
DFFARX1 I_13339  ( .D(I229141), .CLK(I2350), .RSTB(I228923), .Q(I229158) );
DFFARX1 I_13340  ( .D(I229158), .CLK(I2350), .RSTB(I228923), .Q(I228891) );
DFFARX1 I_13341  ( .D(I229158), .CLK(I2350), .RSTB(I228923), .Q(I229189) );
DFFARX1 I_13342  ( .D(I229158), .CLK(I2350), .RSTB(I228923), .Q(I228885) );
nand I_13343 (I229220,I228940,I134119);
nand I_13344 (I229237,I229220,I228974);
and I_13345 (I229254,I229056,I229237);
DFFARX1 I_13346  ( .D(I229254), .CLK(I2350), .RSTB(I228923), .Q(I228915) );
and I_13347 (I228888,I229220,I229189);
DFFARX1 I_13348  ( .D(I134128), .CLK(I2350), .RSTB(I228923), .Q(I229299) );
nor I_13349 (I228912,I229299,I229220);
nor I_13350 (I229330,I229299,I228974);
nand I_13351 (I228909,I229008,I229330);
not I_13352 (I228906,I229299);
DFFARX1 I_13353  ( .D(I134131), .CLK(I2350), .RSTB(I228923), .Q(I229375) );
not I_13354 (I229392,I229375);
nor I_13355 (I229409,I229392,I229073);
and I_13356 (I229426,I229299,I229409);
or I_13357 (I229443,I229220,I229426);
DFFARX1 I_13358  ( .D(I229443), .CLK(I2350), .RSTB(I228923), .Q(I228900) );
not I_13359 (I229474,I229392);
nor I_13360 (I229491,I229299,I229474);
nand I_13361 (I228903,I229392,I229491);
nand I_13362 (I228897,I229056,I229474);
not I_13363 (I229569,I2357);
not I_13364 (I229586,I264906);
nor I_13365 (I229603,I264909,I264891);
nand I_13366 (I229620,I229603,I264918);
nor I_13367 (I229637,I229586,I264909);
nand I_13368 (I229654,I229637,I264897);
DFFARX1 I_13369  ( .D(I229654), .CLK(I2350), .RSTB(I229569), .Q(I229671) );
not I_13370 (I229540,I229671);
not I_13371 (I229702,I264909);
not I_13372 (I229719,I229702);
not I_13373 (I229736,I264903);
nor I_13374 (I229753,I229736,I264915);
and I_13375 (I229770,I229753,I264921);
or I_13376 (I229787,I229770,I264900);
DFFARX1 I_13377  ( .D(I229787), .CLK(I2350), .RSTB(I229569), .Q(I229804) );
DFFARX1 I_13378  ( .D(I229804), .CLK(I2350), .RSTB(I229569), .Q(I229537) );
DFFARX1 I_13379  ( .D(I229804), .CLK(I2350), .RSTB(I229569), .Q(I229835) );
DFFARX1 I_13380  ( .D(I229804), .CLK(I2350), .RSTB(I229569), .Q(I229531) );
nand I_13381 (I229866,I229586,I264903);
nand I_13382 (I229883,I229866,I229620);
and I_13383 (I229900,I229702,I229883);
DFFARX1 I_13384  ( .D(I229900), .CLK(I2350), .RSTB(I229569), .Q(I229561) );
and I_13385 (I229534,I229866,I229835);
DFFARX1 I_13386  ( .D(I264912), .CLK(I2350), .RSTB(I229569), .Q(I229945) );
nor I_13387 (I229558,I229945,I229866);
nor I_13388 (I229976,I229945,I229620);
nand I_13389 (I229555,I229654,I229976);
not I_13390 (I229552,I229945);
DFFARX1 I_13391  ( .D(I264894), .CLK(I2350), .RSTB(I229569), .Q(I230021) );
not I_13392 (I230038,I230021);
nor I_13393 (I230055,I230038,I229719);
and I_13394 (I230072,I229945,I230055);
or I_13395 (I230089,I229866,I230072);
DFFARX1 I_13396  ( .D(I230089), .CLK(I2350), .RSTB(I229569), .Q(I229546) );
not I_13397 (I230120,I230038);
nor I_13398 (I230137,I229945,I230120);
nand I_13399 (I229549,I230038,I230137);
nand I_13400 (I229543,I229702,I230120);
not I_13401 (I230215,I2357);
not I_13402 (I230232,I232779);
nor I_13403 (I230249,I232788,I232773);
nand I_13404 (I230266,I230249,I232761);
nor I_13405 (I230283,I230232,I232788);
nand I_13406 (I230300,I230283,I232764);
DFFARX1 I_13407  ( .D(I230300), .CLK(I2350), .RSTB(I230215), .Q(I230317) );
not I_13408 (I230186,I230317);
not I_13409 (I230348,I232788);
not I_13410 (I230365,I230348);
not I_13411 (I230382,I232776);
nor I_13412 (I230399,I230382,I232770);
and I_13413 (I230416,I230399,I232767);
or I_13414 (I230433,I230416,I232782);
DFFARX1 I_13415  ( .D(I230433), .CLK(I2350), .RSTB(I230215), .Q(I230450) );
DFFARX1 I_13416  ( .D(I230450), .CLK(I2350), .RSTB(I230215), .Q(I230183) );
DFFARX1 I_13417  ( .D(I230450), .CLK(I2350), .RSTB(I230215), .Q(I230481) );
DFFARX1 I_13418  ( .D(I230450), .CLK(I2350), .RSTB(I230215), .Q(I230177) );
nand I_13419 (I230512,I230232,I232776);
nand I_13420 (I230529,I230512,I230266);
and I_13421 (I230546,I230348,I230529);
DFFARX1 I_13422  ( .D(I230546), .CLK(I2350), .RSTB(I230215), .Q(I230207) );
and I_13423 (I230180,I230512,I230481);
DFFARX1 I_13424  ( .D(I232791), .CLK(I2350), .RSTB(I230215), .Q(I230591) );
nor I_13425 (I230204,I230591,I230512);
nor I_13426 (I230622,I230591,I230266);
nand I_13427 (I230201,I230300,I230622);
not I_13428 (I230198,I230591);
DFFARX1 I_13429  ( .D(I232785), .CLK(I2350), .RSTB(I230215), .Q(I230667) );
not I_13430 (I230684,I230667);
nor I_13431 (I230701,I230684,I230365);
and I_13432 (I230718,I230591,I230701);
or I_13433 (I230735,I230512,I230718);
DFFARX1 I_13434  ( .D(I230735), .CLK(I2350), .RSTB(I230215), .Q(I230192) );
not I_13435 (I230766,I230684);
nor I_13436 (I230783,I230591,I230766);
nand I_13437 (I230195,I230684,I230783);
nand I_13438 (I230189,I230348,I230766);
not I_13439 (I230861,I2357);
not I_13440 (I230878,I237675);
nor I_13441 (I230895,I237684,I237669);
nand I_13442 (I230912,I230895,I237657);
nor I_13443 (I230929,I230878,I237684);
nand I_13444 (I230946,I230929,I237660);
DFFARX1 I_13445  ( .D(I230946), .CLK(I2350), .RSTB(I230861), .Q(I230963) );
not I_13446 (I230832,I230963);
not I_13447 (I230994,I237684);
not I_13448 (I231011,I230994);
not I_13449 (I231028,I237672);
nor I_13450 (I231045,I231028,I237666);
and I_13451 (I231062,I231045,I237663);
or I_13452 (I231079,I231062,I237678);
DFFARX1 I_13453  ( .D(I231079), .CLK(I2350), .RSTB(I230861), .Q(I231096) );
DFFARX1 I_13454  ( .D(I231096), .CLK(I2350), .RSTB(I230861), .Q(I230829) );
DFFARX1 I_13455  ( .D(I231096), .CLK(I2350), .RSTB(I230861), .Q(I231127) );
DFFARX1 I_13456  ( .D(I231096), .CLK(I2350), .RSTB(I230861), .Q(I230823) );
nand I_13457 (I231158,I230878,I237672);
nand I_13458 (I231175,I231158,I230912);
and I_13459 (I231192,I230994,I231175);
DFFARX1 I_13460  ( .D(I231192), .CLK(I2350), .RSTB(I230861), .Q(I230853) );
and I_13461 (I230826,I231158,I231127);
DFFARX1 I_13462  ( .D(I237687), .CLK(I2350), .RSTB(I230861), .Q(I231237) );
nor I_13463 (I230850,I231237,I231158);
nor I_13464 (I231268,I231237,I230912);
nand I_13465 (I230847,I230946,I231268);
not I_13466 (I230844,I231237);
DFFARX1 I_13467  ( .D(I237681), .CLK(I2350), .RSTB(I230861), .Q(I231313) );
not I_13468 (I231330,I231313);
nor I_13469 (I231347,I231330,I231011);
and I_13470 (I231364,I231237,I231347);
or I_13471 (I231381,I231158,I231364);
DFFARX1 I_13472  ( .D(I231381), .CLK(I2350), .RSTB(I230861), .Q(I230838) );
not I_13473 (I231412,I231330);
nor I_13474 (I231429,I231237,I231412);
nand I_13475 (I230841,I231330,I231429);
nand I_13476 (I230835,I230994,I231412);
not I_13477 (I231507,I2357);
not I_13478 (I231524,I147649);
nor I_13479 (I231541,I147628,I147640);
nand I_13480 (I231558,I231541,I147643);
nor I_13481 (I231575,I231524,I147628);
nand I_13482 (I231592,I231575,I147625);
DFFARX1 I_13483  ( .D(I231592), .CLK(I2350), .RSTB(I231507), .Q(I231609) );
not I_13484 (I231478,I231609);
not I_13485 (I231640,I147628);
not I_13486 (I231657,I231640);
not I_13487 (I231674,I147646);
nor I_13488 (I231691,I231674,I147637);
and I_13489 (I231708,I231691,I147631);
or I_13490 (I231725,I231708,I147655);
DFFARX1 I_13491  ( .D(I231725), .CLK(I2350), .RSTB(I231507), .Q(I231742) );
DFFARX1 I_13492  ( .D(I231742), .CLK(I2350), .RSTB(I231507), .Q(I231475) );
DFFARX1 I_13493  ( .D(I231742), .CLK(I2350), .RSTB(I231507), .Q(I231773) );
DFFARX1 I_13494  ( .D(I231742), .CLK(I2350), .RSTB(I231507), .Q(I231469) );
nand I_13495 (I231804,I231524,I147646);
nand I_13496 (I231821,I231804,I231558);
and I_13497 (I231838,I231640,I231821);
DFFARX1 I_13498  ( .D(I231838), .CLK(I2350), .RSTB(I231507), .Q(I231499) );
and I_13499 (I231472,I231804,I231773);
DFFARX1 I_13500  ( .D(I147652), .CLK(I2350), .RSTB(I231507), .Q(I231883) );
nor I_13501 (I231496,I231883,I231804);
nor I_13502 (I231914,I231883,I231558);
nand I_13503 (I231493,I231592,I231914);
not I_13504 (I231490,I231883);
DFFARX1 I_13505  ( .D(I147634), .CLK(I2350), .RSTB(I231507), .Q(I231959) );
not I_13506 (I231976,I231959);
nor I_13507 (I231993,I231976,I231657);
and I_13508 (I232010,I231883,I231993);
or I_13509 (I232027,I231804,I232010);
DFFARX1 I_13510  ( .D(I232027), .CLK(I2350), .RSTB(I231507), .Q(I231484) );
not I_13511 (I232058,I231976);
nor I_13512 (I232075,I231883,I232058);
nand I_13513 (I231487,I231976,I232075);
nand I_13514 (I231481,I231640,I232058);
not I_13515 (I232153,I2357);
not I_13516 (I232170,I68579);
nor I_13517 (I232187,I68570,I68561);
nand I_13518 (I232204,I232187,I68576);
nor I_13519 (I232221,I232170,I68570);
nand I_13520 (I232238,I232221,I68573);
DFFARX1 I_13521  ( .D(I232238), .CLK(I2350), .RSTB(I232153), .Q(I232255) );
not I_13522 (I232124,I232255);
not I_13523 (I232286,I68570);
not I_13524 (I232303,I232286);
not I_13525 (I232320,I68582);
nor I_13526 (I232337,I232320,I68567);
and I_13527 (I232354,I232337,I68585);
or I_13528 (I232371,I232354,I68558);
DFFARX1 I_13529  ( .D(I232371), .CLK(I2350), .RSTB(I232153), .Q(I232388) );
DFFARX1 I_13530  ( .D(I232388), .CLK(I2350), .RSTB(I232153), .Q(I232121) );
DFFARX1 I_13531  ( .D(I232388), .CLK(I2350), .RSTB(I232153), .Q(I232419) );
DFFARX1 I_13532  ( .D(I232388), .CLK(I2350), .RSTB(I232153), .Q(I232115) );
nand I_13533 (I232450,I232170,I68582);
nand I_13534 (I232467,I232450,I232204);
and I_13535 (I232484,I232286,I232467);
DFFARX1 I_13536  ( .D(I232484), .CLK(I2350), .RSTB(I232153), .Q(I232145) );
and I_13537 (I232118,I232450,I232419);
DFFARX1 I_13538  ( .D(I68588), .CLK(I2350), .RSTB(I232153), .Q(I232529) );
nor I_13539 (I232142,I232529,I232450);
nor I_13540 (I232560,I232529,I232204);
nand I_13541 (I232139,I232238,I232560);
not I_13542 (I232136,I232529);
DFFARX1 I_13543  ( .D(I68564), .CLK(I2350), .RSTB(I232153), .Q(I232605) );
not I_13544 (I232622,I232605);
nor I_13545 (I232639,I232622,I232303);
and I_13546 (I232656,I232529,I232639);
or I_13547 (I232673,I232450,I232656);
DFFARX1 I_13548  ( .D(I232673), .CLK(I2350), .RSTB(I232153), .Q(I232130) );
not I_13549 (I232704,I232622);
nor I_13550 (I232721,I232529,I232704);
nand I_13551 (I232133,I232622,I232721);
nand I_13552 (I232127,I232286,I232704);
not I_13553 (I232799,I2357);
or I_13554 (I232816,I66620,I66647);
or I_13555 (I232833,I66635,I66620);
nor I_13556 (I232850,I66644,I66623);
DFFARX1 I_13557  ( .D(I232850), .CLK(I2350), .RSTB(I232799), .Q(I232867) );
DFFARX1 I_13558  ( .D(I232850), .CLK(I2350), .RSTB(I232799), .Q(I232761) );
not I_13559 (I232898,I66644);
and I_13560 (I232915,I232898,I66641);
nor I_13561 (I232932,I232915,I66647);
nor I_13562 (I232949,I66638,I66626);
DFFARX1 I_13563  ( .D(I232949), .CLK(I2350), .RSTB(I232799), .Q(I232966) );
not I_13564 (I232983,I232966);
DFFARX1 I_13565  ( .D(I232966), .CLK(I2350), .RSTB(I232799), .Q(I232770) );
nor I_13566 (I233014,I66638,I66635);
and I_13567 (I232764,I233014,I232867);
DFFARX1 I_13568  ( .D(I66650), .CLK(I2350), .RSTB(I232799), .Q(I233045) );
and I_13569 (I233062,I233045,I66632);
nand I_13570 (I233079,I233062,I232833);
and I_13571 (I233096,I232966,I233079);
DFFARX1 I_13572  ( .D(I233096), .CLK(I2350), .RSTB(I232799), .Q(I232791) );
nor I_13573 (I232788,I233062,I232932);
not I_13574 (I233141,I233062);
nor I_13575 (I233158,I232816,I233141);
nor I_13576 (I233175,I233062,I233014);
nand I_13577 (I232785,I232833,I233175);
nor I_13578 (I233206,I233062,I232983);
not I_13579 (I232782,I233062);
nand I_13580 (I232773,I233062,I232983);
DFFARX1 I_13581  ( .D(I66629), .CLK(I2350), .RSTB(I232799), .Q(I233251) );
and I_13582 (I233268,I233251,I233158);
or I_13583 (I233285,I232816,I233268);
DFFARX1 I_13584  ( .D(I233285), .CLK(I2350), .RSTB(I232799), .Q(I232776) );
nand I_13585 (I232779,I233251,I233206);
nand I_13586 (I233330,I233251,I232932);
and I_13587 (I233347,I232850,I233330);
DFFARX1 I_13588  ( .D(I233347), .CLK(I2350), .RSTB(I232799), .Q(I232767) );
not I_13589 (I233411,I2357);
or I_13590 (I233428,I7997,I7982);
or I_13591 (I233445,I7970,I7997);
nor I_13592 (I233462,I7976,I8000);
DFFARX1 I_13593  ( .D(I233462), .CLK(I2350), .RSTB(I233411), .Q(I233479) );
DFFARX1 I_13594  ( .D(I233462), .CLK(I2350), .RSTB(I233411), .Q(I233373) );
not I_13595 (I233510,I7976);
and I_13596 (I233527,I233510,I7973);
nor I_13597 (I233544,I233527,I7982);
nor I_13598 (I233561,I7988,I7985);
DFFARX1 I_13599  ( .D(I233561), .CLK(I2350), .RSTB(I233411), .Q(I233578) );
not I_13600 (I233595,I233578);
DFFARX1 I_13601  ( .D(I233578), .CLK(I2350), .RSTB(I233411), .Q(I233382) );
nor I_13602 (I233626,I7988,I7970);
and I_13603 (I233376,I233626,I233479);
DFFARX1 I_13604  ( .D(I7979), .CLK(I2350), .RSTB(I233411), .Q(I233657) );
and I_13605 (I233674,I233657,I7994);
nand I_13606 (I233691,I233674,I233445);
and I_13607 (I233708,I233578,I233691);
DFFARX1 I_13608  ( .D(I233708), .CLK(I2350), .RSTB(I233411), .Q(I233403) );
nor I_13609 (I233400,I233674,I233544);
not I_13610 (I233753,I233674);
nor I_13611 (I233770,I233428,I233753);
nor I_13612 (I233787,I233674,I233626);
nand I_13613 (I233397,I233445,I233787);
nor I_13614 (I233818,I233674,I233595);
not I_13615 (I233394,I233674);
nand I_13616 (I233385,I233674,I233595);
DFFARX1 I_13617  ( .D(I7991), .CLK(I2350), .RSTB(I233411), .Q(I233863) );
and I_13618 (I233880,I233863,I233770);
or I_13619 (I233897,I233428,I233880);
DFFARX1 I_13620  ( .D(I233897), .CLK(I2350), .RSTB(I233411), .Q(I233388) );
nand I_13621 (I233391,I233863,I233818);
nand I_13622 (I233942,I233863,I233544);
and I_13623 (I233959,I233462,I233942);
DFFARX1 I_13624  ( .D(I233959), .CLK(I2350), .RSTB(I233411), .Q(I233379) );
not I_13625 (I234023,I2357);
or I_13626 (I234040,I344574,I344577);
or I_13627 (I234057,I344583,I344574);
nor I_13628 (I234074,I344580,I344556);
DFFARX1 I_13629  ( .D(I234074), .CLK(I2350), .RSTB(I234023), .Q(I234091) );
DFFARX1 I_13630  ( .D(I234074), .CLK(I2350), .RSTB(I234023), .Q(I233985) );
not I_13631 (I234122,I344580);
and I_13632 (I234139,I234122,I344559);
nor I_13633 (I234156,I234139,I344577);
nor I_13634 (I234173,I344568,I344553);
DFFARX1 I_13635  ( .D(I234173), .CLK(I2350), .RSTB(I234023), .Q(I234190) );
not I_13636 (I234207,I234190);
DFFARX1 I_13637  ( .D(I234190), .CLK(I2350), .RSTB(I234023), .Q(I233994) );
nor I_13638 (I234238,I344568,I344583);
and I_13639 (I233988,I234238,I234091);
DFFARX1 I_13640  ( .D(I344571), .CLK(I2350), .RSTB(I234023), .Q(I234269) );
and I_13641 (I234286,I234269,I344565);
nand I_13642 (I234303,I234286,I234057);
and I_13643 (I234320,I234190,I234303);
DFFARX1 I_13644  ( .D(I234320), .CLK(I2350), .RSTB(I234023), .Q(I234015) );
nor I_13645 (I234012,I234286,I234156);
not I_13646 (I234365,I234286);
nor I_13647 (I234382,I234040,I234365);
nor I_13648 (I234399,I234286,I234238);
nand I_13649 (I234009,I234057,I234399);
nor I_13650 (I234430,I234286,I234207);
not I_13651 (I234006,I234286);
nand I_13652 (I233997,I234286,I234207);
DFFARX1 I_13653  ( .D(I344562), .CLK(I2350), .RSTB(I234023), .Q(I234475) );
and I_13654 (I234492,I234475,I234382);
or I_13655 (I234509,I234040,I234492);
DFFARX1 I_13656  ( .D(I234509), .CLK(I2350), .RSTB(I234023), .Q(I234000) );
nand I_13657 (I234003,I234475,I234430);
nand I_13658 (I234554,I234475,I234156);
and I_13659 (I234571,I234074,I234554);
DFFARX1 I_13660  ( .D(I234571), .CLK(I2350), .RSTB(I234023), .Q(I233991) );
not I_13661 (I234635,I2357);
or I_13662 (I234652,I230838,I230850);
or I_13663 (I234669,I230832,I230838);
nor I_13664 (I234686,I230853,I230829);
DFFARX1 I_13665  ( .D(I234686), .CLK(I2350), .RSTB(I234635), .Q(I234703) );
DFFARX1 I_13666  ( .D(I234686), .CLK(I2350), .RSTB(I234635), .Q(I234597) );
not I_13667 (I234734,I230853);
and I_13668 (I234751,I234734,I230844);
nor I_13669 (I234768,I234751,I230850);
nor I_13670 (I234785,I230823,I230841);
DFFARX1 I_13671  ( .D(I234785), .CLK(I2350), .RSTB(I234635), .Q(I234802) );
not I_13672 (I234819,I234802);
DFFARX1 I_13673  ( .D(I234802), .CLK(I2350), .RSTB(I234635), .Q(I234606) );
nor I_13674 (I234850,I230823,I230832);
and I_13675 (I234600,I234850,I234703);
DFFARX1 I_13676  ( .D(I230847), .CLK(I2350), .RSTB(I234635), .Q(I234881) );
and I_13677 (I234898,I234881,I230826);
nand I_13678 (I234915,I234898,I234669);
and I_13679 (I234932,I234802,I234915);
DFFARX1 I_13680  ( .D(I234932), .CLK(I2350), .RSTB(I234635), .Q(I234627) );
nor I_13681 (I234624,I234898,I234768);
not I_13682 (I234977,I234898);
nor I_13683 (I234994,I234652,I234977);
nor I_13684 (I235011,I234898,I234850);
nand I_13685 (I234621,I234669,I235011);
nor I_13686 (I235042,I234898,I234819);
not I_13687 (I234618,I234898);
nand I_13688 (I234609,I234898,I234819);
DFFARX1 I_13689  ( .D(I230835), .CLK(I2350), .RSTB(I234635), .Q(I235087) );
and I_13690 (I235104,I235087,I234994);
or I_13691 (I235121,I234652,I235104);
DFFARX1 I_13692  ( .D(I235121), .CLK(I2350), .RSTB(I234635), .Q(I234612) );
nand I_13693 (I234615,I235087,I235042);
nand I_13694 (I235166,I235087,I234768);
and I_13695 (I235183,I234686,I235166);
DFFARX1 I_13696  ( .D(I235183), .CLK(I2350), .RSTB(I234635), .Q(I234603) );
not I_13697 (I235247,I2357);
or I_13698 (I235264,I158908,I158896);
or I_13699 (I235281,I158905,I158908);
nor I_13700 (I235298,I158899,I158920);
DFFARX1 I_13701  ( .D(I235298), .CLK(I2350), .RSTB(I235247), .Q(I235315) );
DFFARX1 I_13702  ( .D(I235298), .CLK(I2350), .RSTB(I235247), .Q(I235209) );
not I_13703 (I235346,I158899);
and I_13704 (I235363,I235346,I158914);
nor I_13705 (I235380,I235363,I158896);
nor I_13706 (I235397,I158911,I158926);
DFFARX1 I_13707  ( .D(I235397), .CLK(I2350), .RSTB(I235247), .Q(I235414) );
not I_13708 (I235431,I235414);
DFFARX1 I_13709  ( .D(I235414), .CLK(I2350), .RSTB(I235247), .Q(I235218) );
nor I_13710 (I235462,I158911,I158905);
and I_13711 (I235212,I235462,I235315);
DFFARX1 I_13712  ( .D(I158923), .CLK(I2350), .RSTB(I235247), .Q(I235493) );
and I_13713 (I235510,I235493,I158902);
nand I_13714 (I235527,I235510,I235281);
and I_13715 (I235544,I235414,I235527);
DFFARX1 I_13716  ( .D(I235544), .CLK(I2350), .RSTB(I235247), .Q(I235239) );
nor I_13717 (I235236,I235510,I235380);
not I_13718 (I235589,I235510);
nor I_13719 (I235606,I235264,I235589);
nor I_13720 (I235623,I235510,I235462);
nand I_13721 (I235233,I235281,I235623);
nor I_13722 (I235654,I235510,I235431);
not I_13723 (I235230,I235510);
nand I_13724 (I235221,I235510,I235431);
DFFARX1 I_13725  ( .D(I158917), .CLK(I2350), .RSTB(I235247), .Q(I235699) );
and I_13726 (I235716,I235699,I235606);
or I_13727 (I235733,I235264,I235716);
DFFARX1 I_13728  ( .D(I235733), .CLK(I2350), .RSTB(I235247), .Q(I235224) );
nand I_13729 (I235227,I235699,I235654);
nand I_13730 (I235778,I235699,I235380);
and I_13731 (I235795,I235298,I235778);
DFFARX1 I_13732  ( .D(I235795), .CLK(I2350), .RSTB(I235247), .Q(I235215) );
not I_13733 (I235859,I2357);
or I_13734 (I235876,I94659,I94680);
or I_13735 (I235893,I94677,I94659);
nor I_13736 (I235910,I94668,I94665);
DFFARX1 I_13737  ( .D(I235910), .CLK(I2350), .RSTB(I235859), .Q(I235927) );
DFFARX1 I_13738  ( .D(I235910), .CLK(I2350), .RSTB(I235859), .Q(I235821) );
not I_13739 (I235958,I94668);
and I_13740 (I235975,I235958,I94674);
nor I_13741 (I235992,I235975,I94680);
nor I_13742 (I236009,I94662,I94653);
DFFARX1 I_13743  ( .D(I236009), .CLK(I2350), .RSTB(I235859), .Q(I236026) );
not I_13744 (I236043,I236026);
DFFARX1 I_13745  ( .D(I236026), .CLK(I2350), .RSTB(I235859), .Q(I235830) );
nor I_13746 (I236074,I94662,I94677);
and I_13747 (I235824,I236074,I235927);
DFFARX1 I_13748  ( .D(I94656), .CLK(I2350), .RSTB(I235859), .Q(I236105) );
and I_13749 (I236122,I236105,I94671);
nand I_13750 (I236139,I236122,I235893);
and I_13751 (I236156,I236026,I236139);
DFFARX1 I_13752  ( .D(I236156), .CLK(I2350), .RSTB(I235859), .Q(I235851) );
nor I_13753 (I235848,I236122,I235992);
not I_13754 (I236201,I236122);
nor I_13755 (I236218,I235876,I236201);
nor I_13756 (I236235,I236122,I236074);
nand I_13757 (I235845,I235893,I236235);
nor I_13758 (I236266,I236122,I236043);
not I_13759 (I235842,I236122);
nand I_13760 (I235833,I236122,I236043);
DFFARX1 I_13761  ( .D(I94683), .CLK(I2350), .RSTB(I235859), .Q(I236311) );
and I_13762 (I236328,I236311,I236218);
or I_13763 (I236345,I235876,I236328);
DFFARX1 I_13764  ( .D(I236345), .CLK(I2350), .RSTB(I235859), .Q(I235836) );
nand I_13765 (I235839,I236311,I236266);
nand I_13766 (I236390,I236311,I235992);
and I_13767 (I236407,I235910,I236390);
DFFARX1 I_13768  ( .D(I236407), .CLK(I2350), .RSTB(I235859), .Q(I235827) );
not I_13769 (I236471,I2357);
or I_13770 (I236488,I135916,I135925);
or I_13771 (I236505,I135910,I135916);
nor I_13772 (I236522,I135904,I135898);
DFFARX1 I_13773  ( .D(I236522), .CLK(I2350), .RSTB(I236471), .Q(I236539) );
DFFARX1 I_13774  ( .D(I236522), .CLK(I2350), .RSTB(I236471), .Q(I236433) );
not I_13775 (I236570,I135904);
and I_13776 (I236587,I236570,I135895);
nor I_13777 (I236604,I236587,I135925);
nor I_13778 (I236621,I135922,I135919);
DFFARX1 I_13779  ( .D(I236621), .CLK(I2350), .RSTB(I236471), .Q(I236638) );
not I_13780 (I236655,I236638);
DFFARX1 I_13781  ( .D(I236638), .CLK(I2350), .RSTB(I236471), .Q(I236442) );
nor I_13782 (I236686,I135922,I135910);
and I_13783 (I236436,I236686,I236539);
DFFARX1 I_13784  ( .D(I135901), .CLK(I2350), .RSTB(I236471), .Q(I236717) );
and I_13785 (I236734,I236717,I135907);
nand I_13786 (I236751,I236734,I236505);
and I_13787 (I236768,I236638,I236751);
DFFARX1 I_13788  ( .D(I236768), .CLK(I2350), .RSTB(I236471), .Q(I236463) );
nor I_13789 (I236460,I236734,I236604);
not I_13790 (I236813,I236734);
nor I_13791 (I236830,I236488,I236813);
nor I_13792 (I236847,I236734,I236686);
nand I_13793 (I236457,I236505,I236847);
nor I_13794 (I236878,I236734,I236655);
not I_13795 (I236454,I236734);
nand I_13796 (I236445,I236734,I236655);
DFFARX1 I_13797  ( .D(I135913), .CLK(I2350), .RSTB(I236471), .Q(I236923) );
and I_13798 (I236940,I236923,I236830);
or I_13799 (I236957,I236488,I236940);
DFFARX1 I_13800  ( .D(I236957), .CLK(I2350), .RSTB(I236471), .Q(I236448) );
nand I_13801 (I236451,I236923,I236878);
nand I_13802 (I237002,I236923,I236604);
and I_13803 (I237019,I236522,I237002);
DFFARX1 I_13804  ( .D(I237019), .CLK(I2350), .RSTB(I236471), .Q(I236439) );
not I_13805 (I237083,I2357);
or I_13806 (I237100,I141007,I140995);
or I_13807 (I237117,I141004,I141007);
nor I_13808 (I237134,I140998,I141019);
DFFARX1 I_13809  ( .D(I237134), .CLK(I2350), .RSTB(I237083), .Q(I237151) );
DFFARX1 I_13810  ( .D(I237134), .CLK(I2350), .RSTB(I237083), .Q(I237045) );
not I_13811 (I237182,I140998);
and I_13812 (I237199,I237182,I141013);
nor I_13813 (I237216,I237199,I140995);
nor I_13814 (I237233,I141010,I141025);
DFFARX1 I_13815  ( .D(I237233), .CLK(I2350), .RSTB(I237083), .Q(I237250) );
not I_13816 (I237267,I237250);
DFFARX1 I_13817  ( .D(I237250), .CLK(I2350), .RSTB(I237083), .Q(I237054) );
nor I_13818 (I237298,I141010,I141004);
and I_13819 (I237048,I237298,I237151);
DFFARX1 I_13820  ( .D(I141022), .CLK(I2350), .RSTB(I237083), .Q(I237329) );
and I_13821 (I237346,I237329,I141001);
nand I_13822 (I237363,I237346,I237117);
and I_13823 (I237380,I237250,I237363);
DFFARX1 I_13824  ( .D(I237380), .CLK(I2350), .RSTB(I237083), .Q(I237075) );
nor I_13825 (I237072,I237346,I237216);
not I_13826 (I237425,I237346);
nor I_13827 (I237442,I237100,I237425);
nor I_13828 (I237459,I237346,I237298);
nand I_13829 (I237069,I237117,I237459);
nor I_13830 (I237490,I237346,I237267);
not I_13831 (I237066,I237346);
nand I_13832 (I237057,I237346,I237267);
DFFARX1 I_13833  ( .D(I141016), .CLK(I2350), .RSTB(I237083), .Q(I237535) );
and I_13834 (I237552,I237535,I237442);
or I_13835 (I237569,I237100,I237552);
DFFARX1 I_13836  ( .D(I237569), .CLK(I2350), .RSTB(I237083), .Q(I237060) );
nand I_13837 (I237063,I237535,I237490);
nand I_13838 (I237614,I237535,I237216);
and I_13839 (I237631,I237134,I237614);
DFFARX1 I_13840  ( .D(I237631), .CLK(I2350), .RSTB(I237083), .Q(I237051) );
not I_13841 (I237695,I2357);
or I_13842 (I237712,I173494,I173482);
or I_13843 (I237729,I173491,I173494);
nor I_13844 (I237746,I173485,I173506);
DFFARX1 I_13845  ( .D(I237746), .CLK(I2350), .RSTB(I237695), .Q(I237763) );
DFFARX1 I_13846  ( .D(I237746), .CLK(I2350), .RSTB(I237695), .Q(I237657) );
not I_13847 (I237794,I173485);
and I_13848 (I237811,I237794,I173500);
nor I_13849 (I237828,I237811,I173482);
nor I_13850 (I237845,I173497,I173512);
DFFARX1 I_13851  ( .D(I237845), .CLK(I2350), .RSTB(I237695), .Q(I237862) );
not I_13852 (I237879,I237862);
DFFARX1 I_13853  ( .D(I237862), .CLK(I2350), .RSTB(I237695), .Q(I237666) );
nor I_13854 (I237910,I173497,I173491);
and I_13855 (I237660,I237910,I237763);
DFFARX1 I_13856  ( .D(I173509), .CLK(I2350), .RSTB(I237695), .Q(I237941) );
and I_13857 (I237958,I237941,I173488);
nand I_13858 (I237975,I237958,I237729);
and I_13859 (I237992,I237862,I237975);
DFFARX1 I_13860  ( .D(I237992), .CLK(I2350), .RSTB(I237695), .Q(I237687) );
nor I_13861 (I237684,I237958,I237828);
not I_13862 (I238037,I237958);
nor I_13863 (I238054,I237712,I238037);
nor I_13864 (I238071,I237958,I237910);
nand I_13865 (I237681,I237729,I238071);
nor I_13866 (I238102,I237958,I237879);
not I_13867 (I237678,I237958);
nand I_13868 (I237669,I237958,I237879);
DFFARX1 I_13869  ( .D(I173503), .CLK(I2350), .RSTB(I237695), .Q(I238147) );
and I_13870 (I238164,I238147,I238054);
or I_13871 (I238181,I237712,I238164);
DFFARX1 I_13872  ( .D(I238181), .CLK(I2350), .RSTB(I237695), .Q(I237672) );
nand I_13873 (I237675,I238147,I238102);
nand I_13874 (I238226,I238147,I237828);
and I_13875 (I238243,I237746,I238226);
DFFARX1 I_13876  ( .D(I238243), .CLK(I2350), .RSTB(I237695), .Q(I237663) );
not I_13877 (I238307,I2357);
or I_13878 (I238324,I164875,I164863);
or I_13879 (I238341,I164872,I164875);
nor I_13880 (I238358,I164866,I164887);
DFFARX1 I_13881  ( .D(I238358), .CLK(I2350), .RSTB(I238307), .Q(I238375) );
DFFARX1 I_13882  ( .D(I238358), .CLK(I2350), .RSTB(I238307), .Q(I238269) );
not I_13883 (I238406,I164866);
and I_13884 (I238423,I238406,I164881);
nor I_13885 (I238440,I238423,I164863);
nor I_13886 (I238457,I164878,I164893);
DFFARX1 I_13887  ( .D(I238457), .CLK(I2350), .RSTB(I238307), .Q(I238474) );
not I_13888 (I238491,I238474);
DFFARX1 I_13889  ( .D(I238474), .CLK(I2350), .RSTB(I238307), .Q(I238278) );
nor I_13890 (I238522,I164878,I164872);
and I_13891 (I238272,I238522,I238375);
DFFARX1 I_13892  ( .D(I164890), .CLK(I2350), .RSTB(I238307), .Q(I238553) );
and I_13893 (I238570,I238553,I164869);
nand I_13894 (I238587,I238570,I238341);
and I_13895 (I238604,I238474,I238587);
DFFARX1 I_13896  ( .D(I238604), .CLK(I2350), .RSTB(I238307), .Q(I238299) );
nor I_13897 (I238296,I238570,I238440);
not I_13898 (I238649,I238570);
nor I_13899 (I238666,I238324,I238649);
nor I_13900 (I238683,I238570,I238522);
nand I_13901 (I238293,I238341,I238683);
nor I_13902 (I238714,I238570,I238491);
not I_13903 (I238290,I238570);
nand I_13904 (I238281,I238570,I238491);
DFFARX1 I_13905  ( .D(I164884), .CLK(I2350), .RSTB(I238307), .Q(I238759) );
and I_13906 (I238776,I238759,I238666);
or I_13907 (I238793,I238324,I238776);
DFFARX1 I_13908  ( .D(I238793), .CLK(I2350), .RSTB(I238307), .Q(I238284) );
nand I_13909 (I238287,I238759,I238714);
nand I_13910 (I238838,I238759,I238440);
and I_13911 (I238855,I238358,I238838);
DFFARX1 I_13912  ( .D(I238855), .CLK(I2350), .RSTB(I238307), .Q(I238275) );
not I_13913 (I238919,I2357);
nand I_13914 (I238936,I103962,I103941);
and I_13915 (I238953,I238936,I103938);
DFFARX1 I_13916  ( .D(I238953), .CLK(I2350), .RSTB(I238919), .Q(I238970) );
not I_13917 (I238987,I238970);
DFFARX1 I_13918  ( .D(I238970), .CLK(I2350), .RSTB(I238919), .Q(I238887) );
nor I_13919 (I239018,I103947,I103941);
DFFARX1 I_13920  ( .D(I103935), .CLK(I2350), .RSTB(I238919), .Q(I239035) );
DFFARX1 I_13921  ( .D(I239035), .CLK(I2350), .RSTB(I238919), .Q(I239052) );
not I_13922 (I238890,I239052);
DFFARX1 I_13923  ( .D(I239035), .CLK(I2350), .RSTB(I238919), .Q(I239083) );
and I_13924 (I238884,I238970,I239083);
nand I_13925 (I239114,I103965,I103956);
and I_13926 (I239131,I239114,I103953);
DFFARX1 I_13927  ( .D(I239131), .CLK(I2350), .RSTB(I238919), .Q(I239148) );
nor I_13928 (I239165,I239148,I238987);
not I_13929 (I239182,I239148);
nand I_13930 (I238893,I238970,I239182);
DFFARX1 I_13931  ( .D(I103950), .CLK(I2350), .RSTB(I238919), .Q(I239213) );
and I_13932 (I239230,I239213,I103959);
nor I_13933 (I239247,I239230,I239148);
nor I_13934 (I239264,I239230,I239182);
nand I_13935 (I238899,I239018,I239264);
not I_13936 (I238902,I239230);
DFFARX1 I_13937  ( .D(I239230), .CLK(I2350), .RSTB(I238919), .Q(I238881) );
DFFARX1 I_13938  ( .D(I103944), .CLK(I2350), .RSTB(I238919), .Q(I239323) );
nand I_13939 (I239340,I239323,I239035);
and I_13940 (I239357,I239018,I239340);
DFFARX1 I_13941  ( .D(I239357), .CLK(I2350), .RSTB(I238919), .Q(I238911) );
nor I_13942 (I238908,I239323,I239230);
and I_13943 (I239402,I239323,I239165);
or I_13944 (I239419,I239018,I239402);
DFFARX1 I_13945  ( .D(I239419), .CLK(I2350), .RSTB(I238919), .Q(I238896) );
nand I_13946 (I238905,I239323,I239247);
not I_13947 (I239497,I2357);
nand I_13948 (I239514,I354006,I354009);
and I_13949 (I239531,I239514,I354015);
DFFARX1 I_13950  ( .D(I239531), .CLK(I2350), .RSTB(I239497), .Q(I239548) );
not I_13951 (I239565,I239548);
DFFARX1 I_13952  ( .D(I239548), .CLK(I2350), .RSTB(I239497), .Q(I239465) );
nor I_13953 (I239596,I354012,I354009);
DFFARX1 I_13954  ( .D(I353991), .CLK(I2350), .RSTB(I239497), .Q(I239613) );
DFFARX1 I_13955  ( .D(I239613), .CLK(I2350), .RSTB(I239497), .Q(I239630) );
not I_13956 (I239468,I239630);
DFFARX1 I_13957  ( .D(I239613), .CLK(I2350), .RSTB(I239497), .Q(I239661) );
and I_13958 (I239462,I239548,I239661);
nand I_13959 (I239692,I353988,I354003);
and I_13960 (I239709,I239692,I354000);
DFFARX1 I_13961  ( .D(I239709), .CLK(I2350), .RSTB(I239497), .Q(I239726) );
nor I_13962 (I239743,I239726,I239565);
not I_13963 (I239760,I239726);
nand I_13964 (I239471,I239548,I239760);
DFFARX1 I_13965  ( .D(I354018), .CLK(I2350), .RSTB(I239497), .Q(I239791) );
and I_13966 (I239808,I239791,I353997);
nor I_13967 (I239825,I239808,I239726);
nor I_13968 (I239842,I239808,I239760);
nand I_13969 (I239477,I239596,I239842);
not I_13970 (I239480,I239808);
DFFARX1 I_13971  ( .D(I239808), .CLK(I2350), .RSTB(I239497), .Q(I239459) );
DFFARX1 I_13972  ( .D(I353994), .CLK(I2350), .RSTB(I239497), .Q(I239901) );
nand I_13973 (I239918,I239901,I239613);
and I_13974 (I239935,I239596,I239918);
DFFARX1 I_13975  ( .D(I239935), .CLK(I2350), .RSTB(I239497), .Q(I239489) );
nor I_13976 (I239486,I239901,I239808);
and I_13977 (I239980,I239901,I239743);
or I_13978 (I239997,I239596,I239980);
DFFARX1 I_13979  ( .D(I239997), .CLK(I2350), .RSTB(I239497), .Q(I239474) );
nand I_13980 (I239483,I239901,I239825);
not I_13981 (I240075,I2357);
nand I_13982 (I240092,I141661,I141688);
and I_13983 (I240109,I240092,I141676);
DFFARX1 I_13984  ( .D(I240109), .CLK(I2350), .RSTB(I240075), .Q(I240126) );
not I_13985 (I240143,I240126);
DFFARX1 I_13986  ( .D(I240126), .CLK(I2350), .RSTB(I240075), .Q(I240043) );
nor I_13987 (I240174,I141664,I141688);
DFFARX1 I_13988  ( .D(I141679), .CLK(I2350), .RSTB(I240075), .Q(I240191) );
DFFARX1 I_13989  ( .D(I240191), .CLK(I2350), .RSTB(I240075), .Q(I240208) );
not I_13990 (I240046,I240208);
DFFARX1 I_13991  ( .D(I240191), .CLK(I2350), .RSTB(I240075), .Q(I240239) );
and I_13992 (I240040,I240126,I240239);
nand I_13993 (I240270,I141673,I141670);
and I_13994 (I240287,I240270,I141667);
DFFARX1 I_13995  ( .D(I240287), .CLK(I2350), .RSTB(I240075), .Q(I240304) );
nor I_13996 (I240321,I240304,I240143);
not I_13997 (I240338,I240304);
nand I_13998 (I240049,I240126,I240338);
DFFARX1 I_13999  ( .D(I141682), .CLK(I2350), .RSTB(I240075), .Q(I240369) );
and I_14000 (I240386,I240369,I141658);
nor I_14001 (I240403,I240386,I240304);
nor I_14002 (I240420,I240386,I240338);
nand I_14003 (I240055,I240174,I240420);
not I_14004 (I240058,I240386);
DFFARX1 I_14005  ( .D(I240386), .CLK(I2350), .RSTB(I240075), .Q(I240037) );
DFFARX1 I_14006  ( .D(I141685), .CLK(I2350), .RSTB(I240075), .Q(I240479) );
nand I_14007 (I240496,I240479,I240191);
and I_14008 (I240513,I240174,I240496);
DFFARX1 I_14009  ( .D(I240513), .CLK(I2350), .RSTB(I240075), .Q(I240067) );
nor I_14010 (I240064,I240479,I240386);
and I_14011 (I240558,I240479,I240321);
or I_14012 (I240575,I240174,I240558);
DFFARX1 I_14013  ( .D(I240575), .CLK(I2350), .RSTB(I240075), .Q(I240052) );
nand I_14014 (I240061,I240479,I240403);
not I_14015 (I240653,I2357);
nand I_14016 (I240670,I359038,I359041);
and I_14017 (I240687,I240670,I359047);
DFFARX1 I_14018  ( .D(I240687), .CLK(I2350), .RSTB(I240653), .Q(I240704) );
not I_14019 (I240721,I240704);
DFFARX1 I_14020  ( .D(I240704), .CLK(I2350), .RSTB(I240653), .Q(I240621) );
nor I_14021 (I240752,I359044,I359041);
DFFARX1 I_14022  ( .D(I359023), .CLK(I2350), .RSTB(I240653), .Q(I240769) );
DFFARX1 I_14023  ( .D(I240769), .CLK(I2350), .RSTB(I240653), .Q(I240786) );
not I_14024 (I240624,I240786);
DFFARX1 I_14025  ( .D(I240769), .CLK(I2350), .RSTB(I240653), .Q(I240817) );
and I_14026 (I240618,I240704,I240817);
nand I_14027 (I240848,I359020,I359035);
and I_14028 (I240865,I240848,I359032);
DFFARX1 I_14029  ( .D(I240865), .CLK(I2350), .RSTB(I240653), .Q(I240882) );
nor I_14030 (I240899,I240882,I240721);
not I_14031 (I240916,I240882);
nand I_14032 (I240627,I240704,I240916);
DFFARX1 I_14033  ( .D(I359050), .CLK(I2350), .RSTB(I240653), .Q(I240947) );
and I_14034 (I240964,I240947,I359029);
nor I_14035 (I240981,I240964,I240882);
nor I_14036 (I240998,I240964,I240916);
nand I_14037 (I240633,I240752,I240998);
not I_14038 (I240636,I240964);
DFFARX1 I_14039  ( .D(I240964), .CLK(I2350), .RSTB(I240653), .Q(I240615) );
DFFARX1 I_14040  ( .D(I359026), .CLK(I2350), .RSTB(I240653), .Q(I241057) );
nand I_14041 (I241074,I241057,I240769);
and I_14042 (I241091,I240752,I241074);
DFFARX1 I_14043  ( .D(I241091), .CLK(I2350), .RSTB(I240653), .Q(I240645) );
nor I_14044 (I240642,I241057,I240964);
and I_14045 (I241136,I241057,I240899);
or I_14046 (I241153,I240752,I241136);
DFFARX1 I_14047  ( .D(I241153), .CLK(I2350), .RSTB(I240653), .Q(I240630) );
nand I_14048 (I240639,I241057,I240981);
not I_14049 (I241231,I2357);
nand I_14050 (I241248,I205644,I205641);
and I_14051 (I241265,I241248,I205653);
DFFARX1 I_14052  ( .D(I241265), .CLK(I2350), .RSTB(I241231), .Q(I241282) );
not I_14053 (I241299,I241282);
DFFARX1 I_14054  ( .D(I241282), .CLK(I2350), .RSTB(I241231), .Q(I241199) );
nor I_14055 (I241330,I205650,I205641);
DFFARX1 I_14056  ( .D(I205656), .CLK(I2350), .RSTB(I241231), .Q(I241347) );
DFFARX1 I_14057  ( .D(I241347), .CLK(I2350), .RSTB(I241231), .Q(I241364) );
not I_14058 (I241202,I241364);
DFFARX1 I_14059  ( .D(I241347), .CLK(I2350), .RSTB(I241231), .Q(I241395) );
and I_14060 (I241196,I241282,I241395);
nand I_14061 (I241426,I205632,I205635);
and I_14062 (I241443,I241426,I205659);
DFFARX1 I_14063  ( .D(I241443), .CLK(I2350), .RSTB(I241231), .Q(I241460) );
nor I_14064 (I241477,I241460,I241299);
not I_14065 (I241494,I241460);
nand I_14066 (I241205,I241282,I241494);
DFFARX1 I_14067  ( .D(I205638), .CLK(I2350), .RSTB(I241231), .Q(I241525) );
and I_14068 (I241542,I241525,I205629);
nor I_14069 (I241559,I241542,I241460);
nor I_14070 (I241576,I241542,I241494);
nand I_14071 (I241211,I241330,I241576);
not I_14072 (I241214,I241542);
DFFARX1 I_14073  ( .D(I241542), .CLK(I2350), .RSTB(I241231), .Q(I241193) );
DFFARX1 I_14074  ( .D(I205647), .CLK(I2350), .RSTB(I241231), .Q(I241635) );
nand I_14075 (I241652,I241635,I241347);
and I_14076 (I241669,I241330,I241652);
DFFARX1 I_14077  ( .D(I241669), .CLK(I2350), .RSTB(I241231), .Q(I241223) );
nor I_14078 (I241220,I241635,I241542);
and I_14079 (I241714,I241635,I241477);
or I_14080 (I241731,I241330,I241714);
DFFARX1 I_14081  ( .D(I241731), .CLK(I2350), .RSTB(I241231), .Q(I241208) );
nand I_14082 (I241217,I241635,I241559);
not I_14083 (I241809,I2357);
nand I_14084 (I241826,I302879,I302867);
and I_14085 (I241843,I241826,I302861);
DFFARX1 I_14086  ( .D(I241843), .CLK(I2350), .RSTB(I241809), .Q(I241860) );
not I_14087 (I241877,I241860);
DFFARX1 I_14088  ( .D(I241860), .CLK(I2350), .RSTB(I241809), .Q(I241777) );
nor I_14089 (I241908,I302858,I302867);
DFFARX1 I_14090  ( .D(I302852), .CLK(I2350), .RSTB(I241809), .Q(I241925) );
DFFARX1 I_14091  ( .D(I241925), .CLK(I2350), .RSTB(I241809), .Q(I241942) );
not I_14092 (I241780,I241942);
DFFARX1 I_14093  ( .D(I241925), .CLK(I2350), .RSTB(I241809), .Q(I241973) );
and I_14094 (I241774,I241860,I241973);
nand I_14095 (I242004,I302855,I302870);
and I_14096 (I242021,I242004,I302882);
DFFARX1 I_14097  ( .D(I242021), .CLK(I2350), .RSTB(I241809), .Q(I242038) );
nor I_14098 (I242055,I242038,I241877);
not I_14099 (I242072,I242038);
nand I_14100 (I241783,I241860,I242072);
DFFARX1 I_14101  ( .D(I302873), .CLK(I2350), .RSTB(I241809), .Q(I242103) );
and I_14102 (I242120,I242103,I302864);
nor I_14103 (I242137,I242120,I242038);
nor I_14104 (I242154,I242120,I242072);
nand I_14105 (I241789,I241908,I242154);
not I_14106 (I241792,I242120);
DFFARX1 I_14107  ( .D(I242120), .CLK(I2350), .RSTB(I241809), .Q(I241771) );
DFFARX1 I_14108  ( .D(I302876), .CLK(I2350), .RSTB(I241809), .Q(I242213) );
nand I_14109 (I242230,I242213,I241925);
and I_14110 (I242247,I241908,I242230);
DFFARX1 I_14111  ( .D(I242247), .CLK(I2350), .RSTB(I241809), .Q(I241801) );
nor I_14112 (I241798,I242213,I242120);
and I_14113 (I242292,I242213,I242055);
or I_14114 (I242309,I241908,I242292);
DFFARX1 I_14115  ( .D(I242309), .CLK(I2350), .RSTB(I241809), .Q(I241786) );
nand I_14116 (I241795,I242213,I242137);
not I_14117 (I242387,I2357);
nand I_14118 (I242404,I48553,I48535);
and I_14119 (I242421,I242404,I48547);
DFFARX1 I_14120  ( .D(I242421), .CLK(I2350), .RSTB(I242387), .Q(I242438) );
not I_14121 (I242455,I242438);
DFFARX1 I_14122  ( .D(I242438), .CLK(I2350), .RSTB(I242387), .Q(I242355) );
nor I_14123 (I242486,I48550,I48535);
DFFARX1 I_14124  ( .D(I48559), .CLK(I2350), .RSTB(I242387), .Q(I242503) );
DFFARX1 I_14125  ( .D(I242503), .CLK(I2350), .RSTB(I242387), .Q(I242520) );
not I_14126 (I242358,I242520);
DFFARX1 I_14127  ( .D(I242503), .CLK(I2350), .RSTB(I242387), .Q(I242551) );
and I_14128 (I242352,I242438,I242551);
nand I_14129 (I242582,I48538,I48562);
and I_14130 (I242599,I242582,I48541);
DFFARX1 I_14131  ( .D(I242599), .CLK(I2350), .RSTB(I242387), .Q(I242616) );
nor I_14132 (I242633,I242616,I242455);
not I_14133 (I242650,I242616);
nand I_14134 (I242361,I242438,I242650);
DFFARX1 I_14135  ( .D(I48544), .CLK(I2350), .RSTB(I242387), .Q(I242681) );
and I_14136 (I242698,I242681,I48556);
nor I_14137 (I242715,I242698,I242616);
nor I_14138 (I242732,I242698,I242650);
nand I_14139 (I242367,I242486,I242732);
not I_14140 (I242370,I242698);
DFFARX1 I_14141  ( .D(I242698), .CLK(I2350), .RSTB(I242387), .Q(I242349) );
DFFARX1 I_14142  ( .D(I48532), .CLK(I2350), .RSTB(I242387), .Q(I242791) );
nand I_14143 (I242808,I242791,I242503);
and I_14144 (I242825,I242486,I242808);
DFFARX1 I_14145  ( .D(I242825), .CLK(I2350), .RSTB(I242387), .Q(I242379) );
nor I_14146 (I242376,I242791,I242698);
and I_14147 (I242870,I242791,I242633);
or I_14148 (I242887,I242486,I242870);
DFFARX1 I_14149  ( .D(I242887), .CLK(I2350), .RSTB(I242387), .Q(I242364) );
nand I_14150 (I242373,I242791,I242715);
not I_14151 (I242965,I2357);
nand I_14152 (I242982,I195308,I195305);
and I_14153 (I242999,I242982,I195317);
DFFARX1 I_14154  ( .D(I242999), .CLK(I2350), .RSTB(I242965), .Q(I243016) );
not I_14155 (I243033,I243016);
DFFARX1 I_14156  ( .D(I243016), .CLK(I2350), .RSTB(I242965), .Q(I242933) );
nor I_14157 (I243064,I195314,I195305);
DFFARX1 I_14158  ( .D(I195320), .CLK(I2350), .RSTB(I242965), .Q(I243081) );
DFFARX1 I_14159  ( .D(I243081), .CLK(I2350), .RSTB(I242965), .Q(I243098) );
not I_14160 (I242936,I243098);
DFFARX1 I_14161  ( .D(I243081), .CLK(I2350), .RSTB(I242965), .Q(I243129) );
and I_14162 (I242930,I243016,I243129);
nand I_14163 (I243160,I195296,I195299);
and I_14164 (I243177,I243160,I195323);
DFFARX1 I_14165  ( .D(I243177), .CLK(I2350), .RSTB(I242965), .Q(I243194) );
nor I_14166 (I243211,I243194,I243033);
not I_14167 (I243228,I243194);
nand I_14168 (I242939,I243016,I243228);
DFFARX1 I_14169  ( .D(I195302), .CLK(I2350), .RSTB(I242965), .Q(I243259) );
and I_14170 (I243276,I243259,I195293);
nor I_14171 (I243293,I243276,I243194);
nor I_14172 (I243310,I243276,I243228);
nand I_14173 (I242945,I243064,I243310);
not I_14174 (I242948,I243276);
DFFARX1 I_14175  ( .D(I243276), .CLK(I2350), .RSTB(I242965), .Q(I242927) );
DFFARX1 I_14176  ( .D(I195311), .CLK(I2350), .RSTB(I242965), .Q(I243369) );
nand I_14177 (I243386,I243369,I243081);
and I_14178 (I243403,I243064,I243386);
DFFARX1 I_14179  ( .D(I243403), .CLK(I2350), .RSTB(I242965), .Q(I242957) );
nor I_14180 (I242954,I243369,I243276);
and I_14181 (I243448,I243369,I243211);
or I_14182 (I243465,I243064,I243448);
DFFARX1 I_14183  ( .D(I243465), .CLK(I2350), .RSTB(I242965), .Q(I242942) );
nand I_14184 (I242951,I243369,I243293);
not I_14185 (I243543,I2357);
nand I_14186 (I243560,I327256,I327253);
and I_14187 (I243577,I243560,I327247);
DFFARX1 I_14188  ( .D(I243577), .CLK(I2350), .RSTB(I243543), .Q(I243594) );
not I_14189 (I243611,I243594);
DFFARX1 I_14190  ( .D(I243594), .CLK(I2350), .RSTB(I243543), .Q(I243511) );
nor I_14191 (I243642,I327268,I327253);
DFFARX1 I_14192  ( .D(I327271), .CLK(I2350), .RSTB(I243543), .Q(I243659) );
DFFARX1 I_14193  ( .D(I243659), .CLK(I2350), .RSTB(I243543), .Q(I243676) );
not I_14194 (I243514,I243676);
DFFARX1 I_14195  ( .D(I243659), .CLK(I2350), .RSTB(I243543), .Q(I243707) );
and I_14196 (I243508,I243594,I243707);
nand I_14197 (I243738,I327274,I327265);
and I_14198 (I243755,I243738,I327277);
DFFARX1 I_14199  ( .D(I243755), .CLK(I2350), .RSTB(I243543), .Q(I243772) );
nor I_14200 (I243789,I243772,I243611);
not I_14201 (I243806,I243772);
nand I_14202 (I243517,I243594,I243806);
DFFARX1 I_14203  ( .D(I327250), .CLK(I2350), .RSTB(I243543), .Q(I243837) );
and I_14204 (I243854,I243837,I327259);
nor I_14205 (I243871,I243854,I243772);
nor I_14206 (I243888,I243854,I243806);
nand I_14207 (I243523,I243642,I243888);
not I_14208 (I243526,I243854);
DFFARX1 I_14209  ( .D(I243854), .CLK(I2350), .RSTB(I243543), .Q(I243505) );
DFFARX1 I_14210  ( .D(I327262), .CLK(I2350), .RSTB(I243543), .Q(I243947) );
nand I_14211 (I243964,I243947,I243659);
and I_14212 (I243981,I243642,I243964);
DFFARX1 I_14213  ( .D(I243981), .CLK(I2350), .RSTB(I243543), .Q(I243535) );
nor I_14214 (I243532,I243947,I243854);
and I_14215 (I244026,I243947,I243789);
or I_14216 (I244043,I243642,I244026);
DFFARX1 I_14217  ( .D(I244043), .CLK(I2350), .RSTB(I243543), .Q(I243520) );
nand I_14218 (I243529,I243947,I243871);
not I_14219 (I244121,I2357);
nand I_14220 (I244138,I52429,I52411);
and I_14221 (I244155,I244138,I52423);
DFFARX1 I_14222  ( .D(I244155), .CLK(I2350), .RSTB(I244121), .Q(I244172) );
not I_14223 (I244189,I244172);
DFFARX1 I_14224  ( .D(I244172), .CLK(I2350), .RSTB(I244121), .Q(I244089) );
nor I_14225 (I244220,I52426,I52411);
DFFARX1 I_14226  ( .D(I52435), .CLK(I2350), .RSTB(I244121), .Q(I244237) );
DFFARX1 I_14227  ( .D(I244237), .CLK(I2350), .RSTB(I244121), .Q(I244254) );
not I_14228 (I244092,I244254);
DFFARX1 I_14229  ( .D(I244237), .CLK(I2350), .RSTB(I244121), .Q(I244285) );
and I_14230 (I244086,I244172,I244285);
nand I_14231 (I244316,I52414,I52438);
and I_14232 (I244333,I244316,I52417);
DFFARX1 I_14233  ( .D(I244333), .CLK(I2350), .RSTB(I244121), .Q(I244350) );
nor I_14234 (I244367,I244350,I244189);
not I_14235 (I244384,I244350);
nand I_14236 (I244095,I244172,I244384);
DFFARX1 I_14237  ( .D(I52420), .CLK(I2350), .RSTB(I244121), .Q(I244415) );
and I_14238 (I244432,I244415,I52432);
nor I_14239 (I244449,I244432,I244350);
nor I_14240 (I244466,I244432,I244384);
nand I_14241 (I244101,I244220,I244466);
not I_14242 (I244104,I244432);
DFFARX1 I_14243  ( .D(I244432), .CLK(I2350), .RSTB(I244121), .Q(I244083) );
DFFARX1 I_14244  ( .D(I52408), .CLK(I2350), .RSTB(I244121), .Q(I244525) );
nand I_14245 (I244542,I244525,I244237);
and I_14246 (I244559,I244220,I244542);
DFFARX1 I_14247  ( .D(I244559), .CLK(I2350), .RSTB(I244121), .Q(I244113) );
nor I_14248 (I244110,I244525,I244432);
and I_14249 (I244604,I244525,I244367);
or I_14250 (I244621,I244220,I244604);
DFFARX1 I_14251  ( .D(I244621), .CLK(I2350), .RSTB(I244121), .Q(I244098) );
nand I_14252 (I244107,I244525,I244449);
not I_14253 (I244699,I2357);
nand I_14254 (I244716,I280864,I280852);
and I_14255 (I244733,I244716,I280846);
DFFARX1 I_14256  ( .D(I244733), .CLK(I2350), .RSTB(I244699), .Q(I244750) );
not I_14257 (I244767,I244750);
DFFARX1 I_14258  ( .D(I244750), .CLK(I2350), .RSTB(I244699), .Q(I244667) );
nor I_14259 (I244798,I280843,I280852);
DFFARX1 I_14260  ( .D(I280837), .CLK(I2350), .RSTB(I244699), .Q(I244815) );
DFFARX1 I_14261  ( .D(I244815), .CLK(I2350), .RSTB(I244699), .Q(I244832) );
not I_14262 (I244670,I244832);
DFFARX1 I_14263  ( .D(I244815), .CLK(I2350), .RSTB(I244699), .Q(I244863) );
and I_14264 (I244664,I244750,I244863);
nand I_14265 (I244894,I280840,I280855);
and I_14266 (I244911,I244894,I280867);
DFFARX1 I_14267  ( .D(I244911), .CLK(I2350), .RSTB(I244699), .Q(I244928) );
nor I_14268 (I244945,I244928,I244767);
not I_14269 (I244962,I244928);
nand I_14270 (I244673,I244750,I244962);
DFFARX1 I_14271  ( .D(I280858), .CLK(I2350), .RSTB(I244699), .Q(I244993) );
and I_14272 (I245010,I244993,I280849);
nor I_14273 (I245027,I245010,I244928);
nor I_14274 (I245044,I245010,I244962);
nand I_14275 (I244679,I244798,I245044);
not I_14276 (I244682,I245010);
DFFARX1 I_14277  ( .D(I245010), .CLK(I2350), .RSTB(I244699), .Q(I244661) );
DFFARX1 I_14278  ( .D(I280861), .CLK(I2350), .RSTB(I244699), .Q(I245103) );
nand I_14279 (I245120,I245103,I244815);
and I_14280 (I245137,I244798,I245120);
DFFARX1 I_14281  ( .D(I245137), .CLK(I2350), .RSTB(I244699), .Q(I244691) );
nor I_14282 (I244688,I245103,I245010);
and I_14283 (I245182,I245103,I244945);
or I_14284 (I245199,I244798,I245182);
DFFARX1 I_14285  ( .D(I245199), .CLK(I2350), .RSTB(I244699), .Q(I244676) );
nand I_14286 (I244685,I245103,I245027);
not I_14287 (I245277,I2357);
nand I_14288 (I245294,I136490,I136493);
and I_14289 (I245311,I245294,I136499);
DFFARX1 I_14290  ( .D(I245311), .CLK(I2350), .RSTB(I245277), .Q(I245328) );
not I_14291 (I245345,I245328);
DFFARX1 I_14292  ( .D(I245328), .CLK(I2350), .RSTB(I245277), .Q(I245245) );
nor I_14293 (I245376,I136511,I136493);
DFFARX1 I_14294  ( .D(I136502), .CLK(I2350), .RSTB(I245277), .Q(I245393) );
DFFARX1 I_14295  ( .D(I245393), .CLK(I2350), .RSTB(I245277), .Q(I245410) );
not I_14296 (I245248,I245410);
DFFARX1 I_14297  ( .D(I245393), .CLK(I2350), .RSTB(I245277), .Q(I245441) );
and I_14298 (I245242,I245328,I245441);
nand I_14299 (I245472,I136508,I136505);
and I_14300 (I245489,I245472,I136517);
DFFARX1 I_14301  ( .D(I245489), .CLK(I2350), .RSTB(I245277), .Q(I245506) );
nor I_14302 (I245523,I245506,I245345);
not I_14303 (I245540,I245506);
nand I_14304 (I245251,I245328,I245540);
DFFARX1 I_14305  ( .D(I136514), .CLK(I2350), .RSTB(I245277), .Q(I245571) );
and I_14306 (I245588,I245571,I136520);
nor I_14307 (I245605,I245588,I245506);
nor I_14308 (I245622,I245588,I245540);
nand I_14309 (I245257,I245376,I245622);
not I_14310 (I245260,I245588);
DFFARX1 I_14311  ( .D(I245588), .CLK(I2350), .RSTB(I245277), .Q(I245239) );
DFFARX1 I_14312  ( .D(I136496), .CLK(I2350), .RSTB(I245277), .Q(I245681) );
nand I_14313 (I245698,I245681,I245393);
and I_14314 (I245715,I245376,I245698);
DFFARX1 I_14315  ( .D(I245715), .CLK(I2350), .RSTB(I245277), .Q(I245269) );
nor I_14316 (I245266,I245681,I245588);
and I_14317 (I245760,I245681,I245523);
or I_14318 (I245777,I245376,I245760);
DFFARX1 I_14319  ( .D(I245777), .CLK(I2350), .RSTB(I245277), .Q(I245254) );
nand I_14320 (I245263,I245681,I245605);
not I_14321 (I245855,I2357);
nand I_14322 (I245872,I76331,I76313);
and I_14323 (I245889,I245872,I76325);
DFFARX1 I_14324  ( .D(I245889), .CLK(I2350), .RSTB(I245855), .Q(I245906) );
not I_14325 (I245923,I245906);
DFFARX1 I_14326  ( .D(I245906), .CLK(I2350), .RSTB(I245855), .Q(I245823) );
nor I_14327 (I245954,I76328,I76313);
DFFARX1 I_14328  ( .D(I76337), .CLK(I2350), .RSTB(I245855), .Q(I245971) );
DFFARX1 I_14329  ( .D(I245971), .CLK(I2350), .RSTB(I245855), .Q(I245988) );
not I_14330 (I245826,I245988);
DFFARX1 I_14331  ( .D(I245971), .CLK(I2350), .RSTB(I245855), .Q(I246019) );
and I_14332 (I245820,I245906,I246019);
nand I_14333 (I246050,I76316,I76340);
and I_14334 (I246067,I246050,I76319);
DFFARX1 I_14335  ( .D(I246067), .CLK(I2350), .RSTB(I245855), .Q(I246084) );
nor I_14336 (I246101,I246084,I245923);
not I_14337 (I246118,I246084);
nand I_14338 (I245829,I245906,I246118);
DFFARX1 I_14339  ( .D(I76322), .CLK(I2350), .RSTB(I245855), .Q(I246149) );
and I_14340 (I246166,I246149,I76334);
nor I_14341 (I246183,I246166,I246084);
nor I_14342 (I246200,I246166,I246118);
nand I_14343 (I245835,I245954,I246200);
not I_14344 (I245838,I246166);
DFFARX1 I_14345  ( .D(I246166), .CLK(I2350), .RSTB(I245855), .Q(I245817) );
DFFARX1 I_14346  ( .D(I76310), .CLK(I2350), .RSTB(I245855), .Q(I246259) );
nand I_14347 (I246276,I246259,I245971);
and I_14348 (I246293,I245954,I246276);
DFFARX1 I_14349  ( .D(I246293), .CLK(I2350), .RSTB(I245855), .Q(I245847) );
nor I_14350 (I245844,I246259,I246166);
and I_14351 (I246338,I246259,I246101);
or I_14352 (I246355,I245954,I246338);
DFFARX1 I_14353  ( .D(I246355), .CLK(I2350), .RSTB(I245855), .Q(I245832) );
nand I_14354 (I245841,I246259,I246183);
not I_14355 (I246433,I2357);
nand I_14356 (I246450,I148954,I148981);
and I_14357 (I246467,I246450,I148969);
DFFARX1 I_14358  ( .D(I246467), .CLK(I2350), .RSTB(I246433), .Q(I246484) );
not I_14359 (I246501,I246484);
DFFARX1 I_14360  ( .D(I246484), .CLK(I2350), .RSTB(I246433), .Q(I246401) );
nor I_14361 (I246532,I148957,I148981);
DFFARX1 I_14362  ( .D(I148972), .CLK(I2350), .RSTB(I246433), .Q(I246549) );
DFFARX1 I_14363  ( .D(I246549), .CLK(I2350), .RSTB(I246433), .Q(I246566) );
not I_14364 (I246404,I246566);
DFFARX1 I_14365  ( .D(I246549), .CLK(I2350), .RSTB(I246433), .Q(I246597) );
and I_14366 (I246398,I246484,I246597);
nand I_14367 (I246628,I148966,I148963);
and I_14368 (I246645,I246628,I148960);
DFFARX1 I_14369  ( .D(I246645), .CLK(I2350), .RSTB(I246433), .Q(I246662) );
nor I_14370 (I246679,I246662,I246501);
not I_14371 (I246696,I246662);
nand I_14372 (I246407,I246484,I246696);
DFFARX1 I_14373  ( .D(I148975), .CLK(I2350), .RSTB(I246433), .Q(I246727) );
and I_14374 (I246744,I246727,I148951);
nor I_14375 (I246761,I246744,I246662);
nor I_14376 (I246778,I246744,I246696);
nand I_14377 (I246413,I246532,I246778);
not I_14378 (I246416,I246744);
DFFARX1 I_14379  ( .D(I246744), .CLK(I2350), .RSTB(I246433), .Q(I246395) );
DFFARX1 I_14380  ( .D(I148978), .CLK(I2350), .RSTB(I246433), .Q(I246837) );
nand I_14381 (I246854,I246837,I246549);
and I_14382 (I246871,I246532,I246854);
DFFARX1 I_14383  ( .D(I246871), .CLK(I2350), .RSTB(I246433), .Q(I246425) );
nor I_14384 (I246422,I246837,I246744);
and I_14385 (I246916,I246837,I246679);
or I_14386 (I246933,I246532,I246916);
DFFARX1 I_14387  ( .D(I246933), .CLK(I2350), .RSTB(I246433), .Q(I246410) );
nand I_14388 (I246419,I246837,I246761);
not I_14389 (I247011,I2357);
nand I_14390 (I247028,I325471,I325468);
and I_14391 (I247045,I247028,I325462);
DFFARX1 I_14392  ( .D(I247045), .CLK(I2350), .RSTB(I247011), .Q(I247062) );
not I_14393 (I247079,I247062);
DFFARX1 I_14394  ( .D(I247062), .CLK(I2350), .RSTB(I247011), .Q(I246979) );
nor I_14395 (I247110,I325483,I325468);
DFFARX1 I_14396  ( .D(I325486), .CLK(I2350), .RSTB(I247011), .Q(I247127) );
DFFARX1 I_14397  ( .D(I247127), .CLK(I2350), .RSTB(I247011), .Q(I247144) );
not I_14398 (I246982,I247144);
DFFARX1 I_14399  ( .D(I247127), .CLK(I2350), .RSTB(I247011), .Q(I247175) );
and I_14400 (I246976,I247062,I247175);
nand I_14401 (I247206,I325489,I325480);
and I_14402 (I247223,I247206,I325492);
DFFARX1 I_14403  ( .D(I247223), .CLK(I2350), .RSTB(I247011), .Q(I247240) );
nor I_14404 (I247257,I247240,I247079);
not I_14405 (I247274,I247240);
nand I_14406 (I246985,I247062,I247274);
DFFARX1 I_14407  ( .D(I325465), .CLK(I2350), .RSTB(I247011), .Q(I247305) );
and I_14408 (I247322,I247305,I325474);
nor I_14409 (I247339,I247322,I247240);
nor I_14410 (I247356,I247322,I247274);
nand I_14411 (I246991,I247110,I247356);
not I_14412 (I246994,I247322);
DFFARX1 I_14413  ( .D(I247322), .CLK(I2350), .RSTB(I247011), .Q(I246973) );
DFFARX1 I_14414  ( .D(I325477), .CLK(I2350), .RSTB(I247011), .Q(I247415) );
nand I_14415 (I247432,I247415,I247127);
and I_14416 (I247449,I247110,I247432);
DFFARX1 I_14417  ( .D(I247449), .CLK(I2350), .RSTB(I247011), .Q(I247003) );
nor I_14418 (I247000,I247415,I247322);
and I_14419 (I247494,I247415,I247257);
or I_14420 (I247511,I247110,I247494);
DFFARX1 I_14421  ( .D(I247511), .CLK(I2350), .RSTB(I247011), .Q(I246988) );
nand I_14422 (I246997,I247415,I247339);
not I_14423 (I247589,I2357);
nand I_14424 (I247606,I148291,I148318);
and I_14425 (I247623,I247606,I148306);
DFFARX1 I_14426  ( .D(I247623), .CLK(I2350), .RSTB(I247589), .Q(I247640) );
not I_14427 (I247657,I247640);
DFFARX1 I_14428  ( .D(I247640), .CLK(I2350), .RSTB(I247589), .Q(I247557) );
nor I_14429 (I247688,I148294,I148318);
DFFARX1 I_14430  ( .D(I148309), .CLK(I2350), .RSTB(I247589), .Q(I247705) );
DFFARX1 I_14431  ( .D(I247705), .CLK(I2350), .RSTB(I247589), .Q(I247722) );
not I_14432 (I247560,I247722);
DFFARX1 I_14433  ( .D(I247705), .CLK(I2350), .RSTB(I247589), .Q(I247753) );
and I_14434 (I247554,I247640,I247753);
nand I_14435 (I247784,I148303,I148300);
and I_14436 (I247801,I247784,I148297);
DFFARX1 I_14437  ( .D(I247801), .CLK(I2350), .RSTB(I247589), .Q(I247818) );
nor I_14438 (I247835,I247818,I247657);
not I_14439 (I247852,I247818);
nand I_14440 (I247563,I247640,I247852);
DFFARX1 I_14441  ( .D(I148312), .CLK(I2350), .RSTB(I247589), .Q(I247883) );
and I_14442 (I247900,I247883,I148288);
nor I_14443 (I247917,I247900,I247818);
nor I_14444 (I247934,I247900,I247852);
nand I_14445 (I247569,I247688,I247934);
not I_14446 (I247572,I247900);
DFFARX1 I_14447  ( .D(I247900), .CLK(I2350), .RSTB(I247589), .Q(I247551) );
DFFARX1 I_14448  ( .D(I148315), .CLK(I2350), .RSTB(I247589), .Q(I247993) );
nand I_14449 (I248010,I247993,I247705);
and I_14450 (I248027,I247688,I248010);
DFFARX1 I_14451  ( .D(I248027), .CLK(I2350), .RSTB(I247589), .Q(I247581) );
nor I_14452 (I247578,I247993,I247900);
and I_14453 (I248072,I247993,I247835);
or I_14454 (I248089,I247688,I248072);
DFFARX1 I_14455  ( .D(I248089), .CLK(I2350), .RSTB(I247589), .Q(I247566) );
nand I_14456 (I247575,I247993,I247917);
not I_14457 (I248167,I2357);
nand I_14458 (I248184,I217918,I217915);
and I_14459 (I248201,I248184,I217927);
DFFARX1 I_14460  ( .D(I248201), .CLK(I2350), .RSTB(I248167), .Q(I248218) );
not I_14461 (I248235,I248218);
DFFARX1 I_14462  ( .D(I248218), .CLK(I2350), .RSTB(I248167), .Q(I248135) );
nor I_14463 (I248266,I217924,I217915);
DFFARX1 I_14464  ( .D(I217930), .CLK(I2350), .RSTB(I248167), .Q(I248283) );
DFFARX1 I_14465  ( .D(I248283), .CLK(I2350), .RSTB(I248167), .Q(I248300) );
not I_14466 (I248138,I248300);
DFFARX1 I_14467  ( .D(I248283), .CLK(I2350), .RSTB(I248167), .Q(I248331) );
and I_14468 (I248132,I248218,I248331);
nand I_14469 (I248362,I217906,I217909);
and I_14470 (I248379,I248362,I217933);
DFFARX1 I_14471  ( .D(I248379), .CLK(I2350), .RSTB(I248167), .Q(I248396) );
nor I_14472 (I248413,I248396,I248235);
not I_14473 (I248430,I248396);
nand I_14474 (I248141,I248218,I248430);
DFFARX1 I_14475  ( .D(I217912), .CLK(I2350), .RSTB(I248167), .Q(I248461) );
and I_14476 (I248478,I248461,I217903);
nor I_14477 (I248495,I248478,I248396);
nor I_14478 (I248512,I248478,I248430);
nand I_14479 (I248147,I248266,I248512);
not I_14480 (I248150,I248478);
DFFARX1 I_14481  ( .D(I248478), .CLK(I2350), .RSTB(I248167), .Q(I248129) );
DFFARX1 I_14482  ( .D(I217921), .CLK(I2350), .RSTB(I248167), .Q(I248571) );
nand I_14483 (I248588,I248571,I248283);
and I_14484 (I248605,I248266,I248588);
DFFARX1 I_14485  ( .D(I248605), .CLK(I2350), .RSTB(I248167), .Q(I248159) );
nor I_14486 (I248156,I248571,I248478);
and I_14487 (I248650,I248571,I248413);
or I_14488 (I248667,I248266,I248650);
DFFARX1 I_14489  ( .D(I248667), .CLK(I2350), .RSTB(I248167), .Q(I248144) );
nand I_14490 (I248153,I248571,I248495);
not I_14491 (I248745,I2357);
nand I_14492 (I248762,I394922,I394934);
and I_14493 (I248779,I248762,I394907);
DFFARX1 I_14494  ( .D(I248779), .CLK(I2350), .RSTB(I248745), .Q(I248796) );
not I_14495 (I248813,I248796);
DFFARX1 I_14496  ( .D(I248796), .CLK(I2350), .RSTB(I248745), .Q(I248713) );
nor I_14497 (I248844,I394925,I394934);
DFFARX1 I_14498  ( .D(I394916), .CLK(I2350), .RSTB(I248745), .Q(I248861) );
DFFARX1 I_14499  ( .D(I248861), .CLK(I2350), .RSTB(I248745), .Q(I248878) );
not I_14500 (I248716,I248878);
DFFARX1 I_14501  ( .D(I248861), .CLK(I2350), .RSTB(I248745), .Q(I248909) );
and I_14502 (I248710,I248796,I248909);
nand I_14503 (I248940,I394913,I394919);
and I_14504 (I248957,I248940,I394931);
DFFARX1 I_14505  ( .D(I248957), .CLK(I2350), .RSTB(I248745), .Q(I248974) );
nor I_14506 (I248991,I248974,I248813);
not I_14507 (I249008,I248974);
nand I_14508 (I248719,I248796,I249008);
DFFARX1 I_14509  ( .D(I394937), .CLK(I2350), .RSTB(I248745), .Q(I249039) );
and I_14510 (I249056,I249039,I394928);
nor I_14511 (I249073,I249056,I248974);
nor I_14512 (I249090,I249056,I249008);
nand I_14513 (I248725,I248844,I249090);
not I_14514 (I248728,I249056);
DFFARX1 I_14515  ( .D(I249056), .CLK(I2350), .RSTB(I248745), .Q(I248707) );
DFFARX1 I_14516  ( .D(I394910), .CLK(I2350), .RSTB(I248745), .Q(I249149) );
nand I_14517 (I249166,I249149,I248861);
and I_14518 (I249183,I248844,I249166);
DFFARX1 I_14519  ( .D(I249183), .CLK(I2350), .RSTB(I248745), .Q(I248737) );
nor I_14520 (I248734,I249149,I249056);
and I_14521 (I249228,I249149,I248991);
or I_14522 (I249245,I248844,I249228);
DFFARX1 I_14523  ( .D(I249245), .CLK(I2350), .RSTB(I248745), .Q(I248722) );
nand I_14524 (I248731,I249149,I249073);
not I_14525 (I249323,I2357);
nand I_14526 (I249340,I228254,I228251);
and I_14527 (I249357,I249340,I228263);
DFFARX1 I_14528  ( .D(I249357), .CLK(I2350), .RSTB(I249323), .Q(I249374) );
not I_14529 (I249391,I249374);
DFFARX1 I_14530  ( .D(I249374), .CLK(I2350), .RSTB(I249323), .Q(I249291) );
nor I_14531 (I249422,I228260,I228251);
DFFARX1 I_14532  ( .D(I228266), .CLK(I2350), .RSTB(I249323), .Q(I249439) );
DFFARX1 I_14533  ( .D(I249439), .CLK(I2350), .RSTB(I249323), .Q(I249456) );
not I_14534 (I249294,I249456);
DFFARX1 I_14535  ( .D(I249439), .CLK(I2350), .RSTB(I249323), .Q(I249487) );
and I_14536 (I249288,I249374,I249487);
nand I_14537 (I249518,I228242,I228245);
and I_14538 (I249535,I249518,I228269);
DFFARX1 I_14539  ( .D(I249535), .CLK(I2350), .RSTB(I249323), .Q(I249552) );
nor I_14540 (I249569,I249552,I249391);
not I_14541 (I249586,I249552);
nand I_14542 (I249297,I249374,I249586);
DFFARX1 I_14543  ( .D(I228248), .CLK(I2350), .RSTB(I249323), .Q(I249617) );
and I_14544 (I249634,I249617,I228239);
nor I_14545 (I249651,I249634,I249552);
nor I_14546 (I249668,I249634,I249586);
nand I_14547 (I249303,I249422,I249668);
not I_14548 (I249306,I249634);
DFFARX1 I_14549  ( .D(I249634), .CLK(I2350), .RSTB(I249323), .Q(I249285) );
DFFARX1 I_14550  ( .D(I228257), .CLK(I2350), .RSTB(I249323), .Q(I249727) );
nand I_14551 (I249744,I249727,I249439);
and I_14552 (I249761,I249422,I249744);
DFFARX1 I_14553  ( .D(I249761), .CLK(I2350), .RSTB(I249323), .Q(I249315) );
nor I_14554 (I249312,I249727,I249634);
and I_14555 (I249806,I249727,I249569);
or I_14556 (I249823,I249422,I249806);
DFFARX1 I_14557  ( .D(I249823), .CLK(I2350), .RSTB(I249323), .Q(I249300) );
nand I_14558 (I249309,I249727,I249651);
not I_14559 (I249901,I2357);
nand I_14560 (I249918,I138346,I138373);
and I_14561 (I249935,I249918,I138361);
DFFARX1 I_14562  ( .D(I249935), .CLK(I2350), .RSTB(I249901), .Q(I249952) );
not I_14563 (I249969,I249952);
DFFARX1 I_14564  ( .D(I249952), .CLK(I2350), .RSTB(I249901), .Q(I249869) );
nor I_14565 (I250000,I138349,I138373);
DFFARX1 I_14566  ( .D(I138364), .CLK(I2350), .RSTB(I249901), .Q(I250017) );
DFFARX1 I_14567  ( .D(I250017), .CLK(I2350), .RSTB(I249901), .Q(I250034) );
not I_14568 (I249872,I250034);
DFFARX1 I_14569  ( .D(I250017), .CLK(I2350), .RSTB(I249901), .Q(I250065) );
and I_14570 (I249866,I249952,I250065);
nand I_14571 (I250096,I138358,I138355);
and I_14572 (I250113,I250096,I138352);
DFFARX1 I_14573  ( .D(I250113), .CLK(I2350), .RSTB(I249901), .Q(I250130) );
nor I_14574 (I250147,I250130,I249969);
not I_14575 (I250164,I250130);
nand I_14576 (I249875,I249952,I250164);
DFFARX1 I_14577  ( .D(I138367), .CLK(I2350), .RSTB(I249901), .Q(I250195) );
and I_14578 (I250212,I250195,I138343);
nor I_14579 (I250229,I250212,I250130);
nor I_14580 (I250246,I250212,I250164);
nand I_14581 (I249881,I250000,I250246);
not I_14582 (I249884,I250212);
DFFARX1 I_14583  ( .D(I250212), .CLK(I2350), .RSTB(I249901), .Q(I249863) );
DFFARX1 I_14584  ( .D(I138370), .CLK(I2350), .RSTB(I249901), .Q(I250305) );
nand I_14585 (I250322,I250305,I250017);
and I_14586 (I250339,I250000,I250322);
DFFARX1 I_14587  ( .D(I250339), .CLK(I2350), .RSTB(I249901), .Q(I249893) );
nor I_14588 (I249890,I250305,I250212);
and I_14589 (I250384,I250305,I250147);
or I_14590 (I250401,I250000,I250384);
DFFARX1 I_14591  ( .D(I250401), .CLK(I2350), .RSTB(I249901), .Q(I249878) );
nand I_14592 (I249887,I250305,I250229);
not I_14593 (I250479,I2357);
nand I_14594 (I250496,I182767,I182794);
and I_14595 (I250513,I250496,I182782);
DFFARX1 I_14596  ( .D(I250513), .CLK(I2350), .RSTB(I250479), .Q(I250530) );
not I_14597 (I250547,I250530);
DFFARX1 I_14598  ( .D(I250530), .CLK(I2350), .RSTB(I250479), .Q(I250447) );
nor I_14599 (I250578,I182770,I182794);
DFFARX1 I_14600  ( .D(I182785), .CLK(I2350), .RSTB(I250479), .Q(I250595) );
DFFARX1 I_14601  ( .D(I250595), .CLK(I2350), .RSTB(I250479), .Q(I250612) );
not I_14602 (I250450,I250612);
DFFARX1 I_14603  ( .D(I250595), .CLK(I2350), .RSTB(I250479), .Q(I250643) );
and I_14604 (I250444,I250530,I250643);
nand I_14605 (I250674,I182779,I182776);
and I_14606 (I250691,I250674,I182773);
DFFARX1 I_14607  ( .D(I250691), .CLK(I2350), .RSTB(I250479), .Q(I250708) );
nor I_14608 (I250725,I250708,I250547);
not I_14609 (I250742,I250708);
nand I_14610 (I250453,I250530,I250742);
DFFARX1 I_14611  ( .D(I182788), .CLK(I2350), .RSTB(I250479), .Q(I250773) );
and I_14612 (I250790,I250773,I182764);
nor I_14613 (I250807,I250790,I250708);
nor I_14614 (I250824,I250790,I250742);
nand I_14615 (I250459,I250578,I250824);
not I_14616 (I250462,I250790);
DFFARX1 I_14617  ( .D(I250790), .CLK(I2350), .RSTB(I250479), .Q(I250441) );
DFFARX1 I_14618  ( .D(I182791), .CLK(I2350), .RSTB(I250479), .Q(I250883) );
nand I_14619 (I250900,I250883,I250595);
and I_14620 (I250917,I250578,I250900);
DFFARX1 I_14621  ( .D(I250917), .CLK(I2350), .RSTB(I250479), .Q(I250471) );
nor I_14622 (I250468,I250883,I250790);
and I_14623 (I250962,I250883,I250725);
or I_14624 (I250979,I250578,I250962);
DFFARX1 I_14625  ( .D(I250979), .CLK(I2350), .RSTB(I250479), .Q(I250456) );
nand I_14626 (I250465,I250883,I250807);
not I_14627 (I251057,I2357);
nand I_14628 (I251074,I340797,I340800);
and I_14629 (I251091,I251074,I340806);
DFFARX1 I_14630  ( .D(I251091), .CLK(I2350), .RSTB(I251057), .Q(I251108) );
not I_14631 (I251125,I251108);
DFFARX1 I_14632  ( .D(I251108), .CLK(I2350), .RSTB(I251057), .Q(I251025) );
nor I_14633 (I251156,I340803,I340800);
DFFARX1 I_14634  ( .D(I340782), .CLK(I2350), .RSTB(I251057), .Q(I251173) );
DFFARX1 I_14635  ( .D(I251173), .CLK(I2350), .RSTB(I251057), .Q(I251190) );
not I_14636 (I251028,I251190);
DFFARX1 I_14637  ( .D(I251173), .CLK(I2350), .RSTB(I251057), .Q(I251221) );
and I_14638 (I251022,I251108,I251221);
nand I_14639 (I251252,I340779,I340794);
and I_14640 (I251269,I251252,I340791);
DFFARX1 I_14641  ( .D(I251269), .CLK(I2350), .RSTB(I251057), .Q(I251286) );
nor I_14642 (I251303,I251286,I251125);
not I_14643 (I251320,I251286);
nand I_14644 (I251031,I251108,I251320);
DFFARX1 I_14645  ( .D(I340809), .CLK(I2350), .RSTB(I251057), .Q(I251351) );
and I_14646 (I251368,I251351,I340788);
nor I_14647 (I251385,I251368,I251286);
nor I_14648 (I251402,I251368,I251320);
nand I_14649 (I251037,I251156,I251402);
not I_14650 (I251040,I251368);
DFFARX1 I_14651  ( .D(I251368), .CLK(I2350), .RSTB(I251057), .Q(I251019) );
DFFARX1 I_14652  ( .D(I340785), .CLK(I2350), .RSTB(I251057), .Q(I251461) );
nand I_14653 (I251478,I251461,I251173);
and I_14654 (I251495,I251156,I251478);
DFFARX1 I_14655  ( .D(I251495), .CLK(I2350), .RSTB(I251057), .Q(I251049) );
nor I_14656 (I251046,I251461,I251368);
and I_14657 (I251540,I251461,I251303);
or I_14658 (I251557,I251156,I251540);
DFFARX1 I_14659  ( .D(I251557), .CLK(I2350), .RSTB(I251057), .Q(I251034) );
nand I_14660 (I251043,I251461,I251385);
not I_14661 (I251635,I2357);
nand I_14662 (I251652,I329636,I329633);
and I_14663 (I251669,I251652,I329627);
DFFARX1 I_14664  ( .D(I251669), .CLK(I2350), .RSTB(I251635), .Q(I251686) );
not I_14665 (I251703,I251686);
DFFARX1 I_14666  ( .D(I251686), .CLK(I2350), .RSTB(I251635), .Q(I251603) );
nor I_14667 (I251734,I329648,I329633);
DFFARX1 I_14668  ( .D(I329651), .CLK(I2350), .RSTB(I251635), .Q(I251751) );
DFFARX1 I_14669  ( .D(I251751), .CLK(I2350), .RSTB(I251635), .Q(I251768) );
not I_14670 (I251606,I251768);
DFFARX1 I_14671  ( .D(I251751), .CLK(I2350), .RSTB(I251635), .Q(I251799) );
and I_14672 (I251600,I251686,I251799);
nand I_14673 (I251830,I329654,I329645);
and I_14674 (I251847,I251830,I329657);
DFFARX1 I_14675  ( .D(I251847), .CLK(I2350), .RSTB(I251635), .Q(I251864) );
nor I_14676 (I251881,I251864,I251703);
not I_14677 (I251898,I251864);
nand I_14678 (I251609,I251686,I251898);
DFFARX1 I_14679  ( .D(I329630), .CLK(I2350), .RSTB(I251635), .Q(I251929) );
and I_14680 (I251946,I251929,I329639);
nor I_14681 (I251963,I251946,I251864);
nor I_14682 (I251980,I251946,I251898);
nand I_14683 (I251615,I251734,I251980);
not I_14684 (I251618,I251946);
DFFARX1 I_14685  ( .D(I251946), .CLK(I2350), .RSTB(I251635), .Q(I251597) );
DFFARX1 I_14686  ( .D(I329642), .CLK(I2350), .RSTB(I251635), .Q(I252039) );
nand I_14687 (I252056,I252039,I251751);
and I_14688 (I252073,I251734,I252056);
DFFARX1 I_14689  ( .D(I252073), .CLK(I2350), .RSTB(I251635), .Q(I251627) );
nor I_14690 (I251624,I252039,I251946);
and I_14691 (I252118,I252039,I251881);
or I_14692 (I252135,I251734,I252118);
DFFARX1 I_14693  ( .D(I252135), .CLK(I2350), .RSTB(I251635), .Q(I251612) );
nand I_14694 (I251621,I252039,I251963);
not I_14695 (I252213,I2357);
nand I_14696 (I252230,I115094,I115079);
and I_14697 (I252247,I252230,I115088);
DFFARX1 I_14698  ( .D(I252247), .CLK(I2350), .RSTB(I252213), .Q(I252264) );
not I_14699 (I252281,I252264);
DFFARX1 I_14700  ( .D(I252264), .CLK(I2350), .RSTB(I252213), .Q(I252181) );
nor I_14701 (I252312,I115097,I115079);
DFFARX1 I_14702  ( .D(I115076), .CLK(I2350), .RSTB(I252213), .Q(I252329) );
DFFARX1 I_14703  ( .D(I252329), .CLK(I2350), .RSTB(I252213), .Q(I252346) );
not I_14704 (I252184,I252346);
DFFARX1 I_14705  ( .D(I252329), .CLK(I2350), .RSTB(I252213), .Q(I252377) );
and I_14706 (I252178,I252264,I252377);
nand I_14707 (I252408,I115100,I115073);
and I_14708 (I252425,I252408,I115091);
DFFARX1 I_14709  ( .D(I252425), .CLK(I2350), .RSTB(I252213), .Q(I252442) );
nor I_14710 (I252459,I252442,I252281);
not I_14711 (I252476,I252442);
nand I_14712 (I252187,I252264,I252476);
DFFARX1 I_14713  ( .D(I115085), .CLK(I2350), .RSTB(I252213), .Q(I252507) );
and I_14714 (I252524,I252507,I115070);
nor I_14715 (I252541,I252524,I252442);
nor I_14716 (I252558,I252524,I252476);
nand I_14717 (I252193,I252312,I252558);
not I_14718 (I252196,I252524);
DFFARX1 I_14719  ( .D(I252524), .CLK(I2350), .RSTB(I252213), .Q(I252175) );
DFFARX1 I_14720  ( .D(I115082), .CLK(I2350), .RSTB(I252213), .Q(I252617) );
nand I_14721 (I252634,I252617,I252329);
and I_14722 (I252651,I252312,I252634);
DFFARX1 I_14723  ( .D(I252651), .CLK(I2350), .RSTB(I252213), .Q(I252205) );
nor I_14724 (I252202,I252617,I252524);
and I_14725 (I252696,I252617,I252459);
or I_14726 (I252713,I252312,I252696);
DFFARX1 I_14727  ( .D(I252713), .CLK(I2350), .RSTB(I252213), .Q(I252190) );
nand I_14728 (I252199,I252617,I252541);
not I_14729 (I252791,I2357);
nand I_14730 (I252808,I179452,I179479);
and I_14731 (I252825,I252808,I179467);
DFFARX1 I_14732  ( .D(I252825), .CLK(I2350), .RSTB(I252791), .Q(I252842) );
not I_14733 (I252859,I252842);
DFFARX1 I_14734  ( .D(I252842), .CLK(I2350), .RSTB(I252791), .Q(I252759) );
nor I_14735 (I252890,I179455,I179479);
DFFARX1 I_14736  ( .D(I179470), .CLK(I2350), .RSTB(I252791), .Q(I252907) );
DFFARX1 I_14737  ( .D(I252907), .CLK(I2350), .RSTB(I252791), .Q(I252924) );
not I_14738 (I252762,I252924);
DFFARX1 I_14739  ( .D(I252907), .CLK(I2350), .RSTB(I252791), .Q(I252955) );
and I_14740 (I252756,I252842,I252955);
nand I_14741 (I252986,I179464,I179461);
and I_14742 (I253003,I252986,I179458);
DFFARX1 I_14743  ( .D(I253003), .CLK(I2350), .RSTB(I252791), .Q(I253020) );
nor I_14744 (I253037,I253020,I252859);
not I_14745 (I253054,I253020);
nand I_14746 (I252765,I252842,I253054);
DFFARX1 I_14747  ( .D(I179473), .CLK(I2350), .RSTB(I252791), .Q(I253085) );
and I_14748 (I253102,I253085,I179449);
nor I_14749 (I253119,I253102,I253020);
nor I_14750 (I253136,I253102,I253054);
nand I_14751 (I252771,I252890,I253136);
not I_14752 (I252774,I253102);
DFFARX1 I_14753  ( .D(I253102), .CLK(I2350), .RSTB(I252791), .Q(I252753) );
DFFARX1 I_14754  ( .D(I179476), .CLK(I2350), .RSTB(I252791), .Q(I253195) );
nand I_14755 (I253212,I253195,I252907);
and I_14756 (I253229,I252890,I253212);
DFFARX1 I_14757  ( .D(I253229), .CLK(I2350), .RSTB(I252791), .Q(I252783) );
nor I_14758 (I252780,I253195,I253102);
and I_14759 (I253274,I253195,I253037);
or I_14760 (I253291,I252890,I253274);
DFFARX1 I_14761  ( .D(I253291), .CLK(I2350), .RSTB(I252791), .Q(I252768) );
nand I_14762 (I252777,I253195,I253119);
not I_14763 (I253369,I2357);
nand I_14764 (I253386,I6863,I6878);
and I_14765 (I253403,I253386,I6866);
DFFARX1 I_14766  ( .D(I253403), .CLK(I2350), .RSTB(I253369), .Q(I253420) );
not I_14767 (I253437,I253420);
DFFARX1 I_14768  ( .D(I253420), .CLK(I2350), .RSTB(I253369), .Q(I253337) );
nor I_14769 (I253468,I6875,I6878);
DFFARX1 I_14770  ( .D(I6860), .CLK(I2350), .RSTB(I253369), .Q(I253485) );
DFFARX1 I_14771  ( .D(I253485), .CLK(I2350), .RSTB(I253369), .Q(I253502) );
not I_14772 (I253340,I253502);
DFFARX1 I_14773  ( .D(I253485), .CLK(I2350), .RSTB(I253369), .Q(I253533) );
and I_14774 (I253334,I253420,I253533);
nand I_14775 (I253564,I6851,I6848);
and I_14776 (I253581,I253564,I6854);
DFFARX1 I_14777  ( .D(I253581), .CLK(I2350), .RSTB(I253369), .Q(I253598) );
nor I_14778 (I253615,I253598,I253437);
not I_14779 (I253632,I253598);
nand I_14780 (I253343,I253420,I253632);
DFFARX1 I_14781  ( .D(I6857), .CLK(I2350), .RSTB(I253369), .Q(I253663) );
and I_14782 (I253680,I253663,I6869);
nor I_14783 (I253697,I253680,I253598);
nor I_14784 (I253714,I253680,I253632);
nand I_14785 (I253349,I253468,I253714);
not I_14786 (I253352,I253680);
DFFARX1 I_14787  ( .D(I253680), .CLK(I2350), .RSTB(I253369), .Q(I253331) );
DFFARX1 I_14788  ( .D(I6872), .CLK(I2350), .RSTB(I253369), .Q(I253773) );
nand I_14789 (I253790,I253773,I253485);
and I_14790 (I253807,I253468,I253790);
DFFARX1 I_14791  ( .D(I253807), .CLK(I2350), .RSTB(I253369), .Q(I253361) );
nor I_14792 (I253358,I253773,I253680);
and I_14793 (I253852,I253773,I253615);
or I_14794 (I253869,I253468,I253852);
DFFARX1 I_14795  ( .D(I253869), .CLK(I2350), .RSTB(I253369), .Q(I253346) );
nand I_14796 (I253355,I253773,I253697);
not I_14797 (I253947,I2357);
nand I_14798 (I253964,I38217,I38199);
and I_14799 (I253981,I253964,I38211);
DFFARX1 I_14800  ( .D(I253981), .CLK(I2350), .RSTB(I253947), .Q(I253998) );
not I_14801 (I254015,I253998);
DFFARX1 I_14802  ( .D(I253998), .CLK(I2350), .RSTB(I253947), .Q(I253915) );
nor I_14803 (I254046,I38214,I38199);
DFFARX1 I_14804  ( .D(I38223), .CLK(I2350), .RSTB(I253947), .Q(I254063) );
DFFARX1 I_14805  ( .D(I254063), .CLK(I2350), .RSTB(I253947), .Q(I254080) );
not I_14806 (I253918,I254080);
DFFARX1 I_14807  ( .D(I254063), .CLK(I2350), .RSTB(I253947), .Q(I254111) );
and I_14808 (I253912,I253998,I254111);
nand I_14809 (I254142,I38202,I38226);
and I_14810 (I254159,I254142,I38205);
DFFARX1 I_14811  ( .D(I254159), .CLK(I2350), .RSTB(I253947), .Q(I254176) );
nor I_14812 (I254193,I254176,I254015);
not I_14813 (I254210,I254176);
nand I_14814 (I253921,I253998,I254210);
DFFARX1 I_14815  ( .D(I38208), .CLK(I2350), .RSTB(I253947), .Q(I254241) );
and I_14816 (I254258,I254241,I38220);
nor I_14817 (I254275,I254258,I254176);
nor I_14818 (I254292,I254258,I254210);
nand I_14819 (I253927,I254046,I254292);
not I_14820 (I253930,I254258);
DFFARX1 I_14821  ( .D(I254258), .CLK(I2350), .RSTB(I253947), .Q(I253909) );
DFFARX1 I_14822  ( .D(I38196), .CLK(I2350), .RSTB(I253947), .Q(I254351) );
nand I_14823 (I254368,I254351,I254063);
and I_14824 (I254385,I254046,I254368);
DFFARX1 I_14825  ( .D(I254385), .CLK(I2350), .RSTB(I253947), .Q(I253939) );
nor I_14826 (I253936,I254351,I254258);
and I_14827 (I254430,I254351,I254193);
or I_14828 (I254447,I254046,I254430);
DFFARX1 I_14829  ( .D(I254447), .CLK(I2350), .RSTB(I253947), .Q(I253924) );
nand I_14830 (I253933,I254351,I254275);
not I_14831 (I254525,I2357);
nand I_14832 (I254542,I5180,I5195);
and I_14833 (I254559,I254542,I5183);
DFFARX1 I_14834  ( .D(I254559), .CLK(I2350), .RSTB(I254525), .Q(I254576) );
not I_14835 (I254593,I254576);
DFFARX1 I_14836  ( .D(I254576), .CLK(I2350), .RSTB(I254525), .Q(I254493) );
nor I_14837 (I254624,I5192,I5195);
DFFARX1 I_14838  ( .D(I5177), .CLK(I2350), .RSTB(I254525), .Q(I254641) );
DFFARX1 I_14839  ( .D(I254641), .CLK(I2350), .RSTB(I254525), .Q(I254658) );
not I_14840 (I254496,I254658);
DFFARX1 I_14841  ( .D(I254641), .CLK(I2350), .RSTB(I254525), .Q(I254689) );
and I_14842 (I254490,I254576,I254689);
nand I_14843 (I254720,I5168,I5165);
and I_14844 (I254737,I254720,I5171);
DFFARX1 I_14845  ( .D(I254737), .CLK(I2350), .RSTB(I254525), .Q(I254754) );
nor I_14846 (I254771,I254754,I254593);
not I_14847 (I254788,I254754);
nand I_14848 (I254499,I254576,I254788);
DFFARX1 I_14849  ( .D(I5174), .CLK(I2350), .RSTB(I254525), .Q(I254819) );
and I_14850 (I254836,I254819,I5186);
nor I_14851 (I254853,I254836,I254754);
nor I_14852 (I254870,I254836,I254788);
nand I_14853 (I254505,I254624,I254870);
not I_14854 (I254508,I254836);
DFFARX1 I_14855  ( .D(I254836), .CLK(I2350), .RSTB(I254525), .Q(I254487) );
DFFARX1 I_14856  ( .D(I5189), .CLK(I2350), .RSTB(I254525), .Q(I254929) );
nand I_14857 (I254946,I254929,I254641);
and I_14858 (I254963,I254624,I254946);
DFFARX1 I_14859  ( .D(I254963), .CLK(I2350), .RSTB(I254525), .Q(I254517) );
nor I_14860 (I254514,I254929,I254836);
and I_14861 (I255008,I254929,I254771);
or I_14862 (I255025,I254624,I255008);
DFFARX1 I_14863  ( .D(I255025), .CLK(I2350), .RSTB(I254525), .Q(I254502) );
nand I_14864 (I254511,I254929,I254853);
not I_14865 (I255103,I2357);
nand I_14866 (I255120,I210166,I210163);
and I_14867 (I255137,I255120,I210175);
DFFARX1 I_14868  ( .D(I255137), .CLK(I2350), .RSTB(I255103), .Q(I255154) );
not I_14869 (I255171,I255154);
DFFARX1 I_14870  ( .D(I255154), .CLK(I2350), .RSTB(I255103), .Q(I255071) );
nor I_14871 (I255202,I210172,I210163);
DFFARX1 I_14872  ( .D(I210178), .CLK(I2350), .RSTB(I255103), .Q(I255219) );
DFFARX1 I_14873  ( .D(I255219), .CLK(I2350), .RSTB(I255103), .Q(I255236) );
not I_14874 (I255074,I255236);
DFFARX1 I_14875  ( .D(I255219), .CLK(I2350), .RSTB(I255103), .Q(I255267) );
and I_14876 (I255068,I255154,I255267);
nand I_14877 (I255298,I210154,I210157);
and I_14878 (I255315,I255298,I210181);
DFFARX1 I_14879  ( .D(I255315), .CLK(I2350), .RSTB(I255103), .Q(I255332) );
nor I_14880 (I255349,I255332,I255171);
not I_14881 (I255366,I255332);
nand I_14882 (I255077,I255154,I255366);
DFFARX1 I_14883  ( .D(I210160), .CLK(I2350), .RSTB(I255103), .Q(I255397) );
and I_14884 (I255414,I255397,I210151);
nor I_14885 (I255431,I255414,I255332);
nor I_14886 (I255448,I255414,I255366);
nand I_14887 (I255083,I255202,I255448);
not I_14888 (I255086,I255414);
DFFARX1 I_14889  ( .D(I255414), .CLK(I2350), .RSTB(I255103), .Q(I255065) );
DFFARX1 I_14890  ( .D(I210169), .CLK(I2350), .RSTB(I255103), .Q(I255507) );
nand I_14891 (I255524,I255507,I255219);
and I_14892 (I255541,I255202,I255524);
DFFARX1 I_14893  ( .D(I255541), .CLK(I2350), .RSTB(I255103), .Q(I255095) );
nor I_14894 (I255092,I255507,I255414);
and I_14895 (I255586,I255507,I255349);
or I_14896 (I255603,I255202,I255586);
DFFARX1 I_14897  ( .D(I255603), .CLK(I2350), .RSTB(I255103), .Q(I255080) );
nand I_14898 (I255089,I255507,I255431);
not I_14899 (I255681,I2357);
nand I_14900 (I255698,I137085,I137088);
and I_14901 (I255715,I255698,I137094);
DFFARX1 I_14902  ( .D(I255715), .CLK(I2350), .RSTB(I255681), .Q(I255732) );
not I_14903 (I255749,I255732);
DFFARX1 I_14904  ( .D(I255732), .CLK(I2350), .RSTB(I255681), .Q(I255649) );
nor I_14905 (I255780,I137106,I137088);
DFFARX1 I_14906  ( .D(I137097), .CLK(I2350), .RSTB(I255681), .Q(I255797) );
DFFARX1 I_14907  ( .D(I255797), .CLK(I2350), .RSTB(I255681), .Q(I255814) );
not I_14908 (I255652,I255814);
DFFARX1 I_14909  ( .D(I255797), .CLK(I2350), .RSTB(I255681), .Q(I255845) );
and I_14910 (I255646,I255732,I255845);
nand I_14911 (I255876,I137103,I137100);
and I_14912 (I255893,I255876,I137112);
DFFARX1 I_14913  ( .D(I255893), .CLK(I2350), .RSTB(I255681), .Q(I255910) );
nor I_14914 (I255927,I255910,I255749);
not I_14915 (I255944,I255910);
nand I_14916 (I255655,I255732,I255944);
DFFARX1 I_14917  ( .D(I137109), .CLK(I2350), .RSTB(I255681), .Q(I255975) );
and I_14918 (I255992,I255975,I137115);
nor I_14919 (I256009,I255992,I255910);
nor I_14920 (I256026,I255992,I255944);
nand I_14921 (I255661,I255780,I256026);
not I_14922 (I255664,I255992);
DFFARX1 I_14923  ( .D(I255992), .CLK(I2350), .RSTB(I255681), .Q(I255643) );
DFFARX1 I_14924  ( .D(I137091), .CLK(I2350), .RSTB(I255681), .Q(I256085) );
nand I_14925 (I256102,I256085,I255797);
and I_14926 (I256119,I255780,I256102);
DFFARX1 I_14927  ( .D(I256119), .CLK(I2350), .RSTB(I255681), .Q(I255673) );
nor I_14928 (I255670,I256085,I255992);
and I_14929 (I256164,I256085,I255927);
or I_14930 (I256181,I255780,I256164);
DFFARX1 I_14931  ( .D(I256181), .CLK(I2350), .RSTB(I255681), .Q(I255658) );
nand I_14932 (I255667,I256085,I256009);
not I_14933 (I256259,I2357);
nand I_14934 (I256276,I131730,I131733);
and I_14935 (I256293,I256276,I131739);
DFFARX1 I_14936  ( .D(I256293), .CLK(I2350), .RSTB(I256259), .Q(I256310) );
not I_14937 (I256327,I256310);
DFFARX1 I_14938  ( .D(I256310), .CLK(I2350), .RSTB(I256259), .Q(I256227) );
nor I_14939 (I256358,I131751,I131733);
DFFARX1 I_14940  ( .D(I131742), .CLK(I2350), .RSTB(I256259), .Q(I256375) );
DFFARX1 I_14941  ( .D(I256375), .CLK(I2350), .RSTB(I256259), .Q(I256392) );
not I_14942 (I256230,I256392);
DFFARX1 I_14943  ( .D(I256375), .CLK(I2350), .RSTB(I256259), .Q(I256423) );
and I_14944 (I256224,I256310,I256423);
nand I_14945 (I256454,I131748,I131745);
and I_14946 (I256471,I256454,I131757);
DFFARX1 I_14947  ( .D(I256471), .CLK(I2350), .RSTB(I256259), .Q(I256488) );
nor I_14948 (I256505,I256488,I256327);
not I_14949 (I256522,I256488);
nand I_14950 (I256233,I256310,I256522);
DFFARX1 I_14951  ( .D(I131754), .CLK(I2350), .RSTB(I256259), .Q(I256553) );
and I_14952 (I256570,I256553,I131760);
nor I_14953 (I256587,I256570,I256488);
nor I_14954 (I256604,I256570,I256522);
nand I_14955 (I256239,I256358,I256604);
not I_14956 (I256242,I256570);
DFFARX1 I_14957  ( .D(I256570), .CLK(I2350), .RSTB(I256259), .Q(I256221) );
DFFARX1 I_14958  ( .D(I131736), .CLK(I2350), .RSTB(I256259), .Q(I256663) );
nand I_14959 (I256680,I256663,I256375);
and I_14960 (I256697,I256358,I256680);
DFFARX1 I_14961  ( .D(I256697), .CLK(I2350), .RSTB(I256259), .Q(I256251) );
nor I_14962 (I256248,I256663,I256570);
and I_14963 (I256742,I256663,I256505);
or I_14964 (I256759,I256358,I256742);
DFFARX1 I_14965  ( .D(I256759), .CLK(I2350), .RSTB(I256259), .Q(I256236) );
nand I_14966 (I256245,I256663,I256587);
not I_14967 (I256837,I2357);
nand I_14968 (I256854,I311209,I311197);
and I_14969 (I256871,I256854,I311191);
DFFARX1 I_14970  ( .D(I256871), .CLK(I2350), .RSTB(I256837), .Q(I256888) );
not I_14971 (I256905,I256888);
DFFARX1 I_14972  ( .D(I256888), .CLK(I2350), .RSTB(I256837), .Q(I256805) );
nor I_14973 (I256936,I311188,I311197);
DFFARX1 I_14974  ( .D(I311182), .CLK(I2350), .RSTB(I256837), .Q(I256953) );
DFFARX1 I_14975  ( .D(I256953), .CLK(I2350), .RSTB(I256837), .Q(I256970) );
not I_14976 (I256808,I256970);
DFFARX1 I_14977  ( .D(I256953), .CLK(I2350), .RSTB(I256837), .Q(I257001) );
and I_14978 (I256802,I256888,I257001);
nand I_14979 (I257032,I311185,I311200);
and I_14980 (I257049,I257032,I311212);
DFFARX1 I_14981  ( .D(I257049), .CLK(I2350), .RSTB(I256837), .Q(I257066) );
nor I_14982 (I257083,I257066,I256905);
not I_14983 (I257100,I257066);
nand I_14984 (I256811,I256888,I257100);
DFFARX1 I_14985  ( .D(I311203), .CLK(I2350), .RSTB(I256837), .Q(I257131) );
and I_14986 (I257148,I257131,I311194);
nor I_14987 (I257165,I257148,I257066);
nor I_14988 (I257182,I257148,I257100);
nand I_14989 (I256817,I256936,I257182);
not I_14990 (I256820,I257148);
DFFARX1 I_14991  ( .D(I257148), .CLK(I2350), .RSTB(I256837), .Q(I256799) );
DFFARX1 I_14992  ( .D(I311206), .CLK(I2350), .RSTB(I256837), .Q(I257241) );
nand I_14993 (I257258,I257241,I256953);
and I_14994 (I257275,I256936,I257258);
DFFARX1 I_14995  ( .D(I257275), .CLK(I2350), .RSTB(I256837), .Q(I256829) );
nor I_14996 (I256826,I257241,I257148);
and I_14997 (I257320,I257241,I257083);
or I_14998 (I257337,I256936,I257320);
DFFARX1 I_14999  ( .D(I257337), .CLK(I2350), .RSTB(I256837), .Q(I256814) );
nand I_15000 (I256823,I257241,I257165);
not I_15001 (I257415,I2357);
nand I_15002 (I257432,I94017,I93996);
and I_15003 (I257449,I257432,I93993);
DFFARX1 I_15004  ( .D(I257449), .CLK(I2350), .RSTB(I257415), .Q(I257466) );
not I_15005 (I257483,I257466);
DFFARX1 I_15006  ( .D(I257466), .CLK(I2350), .RSTB(I257415), .Q(I257383) );
nor I_15007 (I257514,I94002,I93996);
DFFARX1 I_15008  ( .D(I93990), .CLK(I2350), .RSTB(I257415), .Q(I257531) );
DFFARX1 I_15009  ( .D(I257531), .CLK(I2350), .RSTB(I257415), .Q(I257548) );
not I_15010 (I257386,I257548);
DFFARX1 I_15011  ( .D(I257531), .CLK(I2350), .RSTB(I257415), .Q(I257579) );
and I_15012 (I257380,I257466,I257579);
nand I_15013 (I257610,I94020,I94011);
and I_15014 (I257627,I257610,I94008);
DFFARX1 I_15015  ( .D(I257627), .CLK(I2350), .RSTB(I257415), .Q(I257644) );
nor I_15016 (I257661,I257644,I257483);
not I_15017 (I257678,I257644);
nand I_15018 (I257389,I257466,I257678);
DFFARX1 I_15019  ( .D(I94005), .CLK(I2350), .RSTB(I257415), .Q(I257709) );
and I_15020 (I257726,I257709,I94014);
nor I_15021 (I257743,I257726,I257644);
nor I_15022 (I257760,I257726,I257678);
nand I_15023 (I257395,I257514,I257760);
not I_15024 (I257398,I257726);
DFFARX1 I_15025  ( .D(I257726), .CLK(I2350), .RSTB(I257415), .Q(I257377) );
DFFARX1 I_15026  ( .D(I93999), .CLK(I2350), .RSTB(I257415), .Q(I257819) );
nand I_15027 (I257836,I257819,I257531);
and I_15028 (I257853,I257514,I257836);
DFFARX1 I_15029  ( .D(I257853), .CLK(I2350), .RSTB(I257415), .Q(I257407) );
nor I_15030 (I257404,I257819,I257726);
and I_15031 (I257898,I257819,I257661);
or I_15032 (I257915,I257514,I257898);
DFFARX1 I_15033  ( .D(I257915), .CLK(I2350), .RSTB(I257415), .Q(I257392) );
nand I_15034 (I257401,I257819,I257743);
not I_15035 (I257993,I2357);
nand I_15036 (I258010,I74393,I74375);
and I_15037 (I258027,I258010,I74387);
DFFARX1 I_15038  ( .D(I258027), .CLK(I2350), .RSTB(I257993), .Q(I258044) );
not I_15039 (I258061,I258044);
DFFARX1 I_15040  ( .D(I258044), .CLK(I2350), .RSTB(I257993), .Q(I257961) );
nor I_15041 (I258092,I74390,I74375);
DFFARX1 I_15042  ( .D(I74399), .CLK(I2350), .RSTB(I257993), .Q(I258109) );
DFFARX1 I_15043  ( .D(I258109), .CLK(I2350), .RSTB(I257993), .Q(I258126) );
not I_15044 (I257964,I258126);
DFFARX1 I_15045  ( .D(I258109), .CLK(I2350), .RSTB(I257993), .Q(I258157) );
and I_15046 (I257958,I258044,I258157);
nand I_15047 (I258188,I74378,I74402);
and I_15048 (I258205,I258188,I74381);
DFFARX1 I_15049  ( .D(I258205), .CLK(I2350), .RSTB(I257993), .Q(I258222) );
nor I_15050 (I258239,I258222,I258061);
not I_15051 (I258256,I258222);
nand I_15052 (I257967,I258044,I258256);
DFFARX1 I_15053  ( .D(I74384), .CLK(I2350), .RSTB(I257993), .Q(I258287) );
and I_15054 (I258304,I258287,I74396);
nor I_15055 (I258321,I258304,I258222);
nor I_15056 (I258338,I258304,I258256);
nand I_15057 (I257973,I258092,I258338);
not I_15058 (I257976,I258304);
DFFARX1 I_15059  ( .D(I258304), .CLK(I2350), .RSTB(I257993), .Q(I257955) );
DFFARX1 I_15060  ( .D(I74372), .CLK(I2350), .RSTB(I257993), .Q(I258397) );
nand I_15061 (I258414,I258397,I258109);
and I_15062 (I258431,I258092,I258414);
DFFARX1 I_15063  ( .D(I258431), .CLK(I2350), .RSTB(I257993), .Q(I257985) );
nor I_15064 (I257982,I258397,I258304);
and I_15065 (I258476,I258397,I258239);
or I_15066 (I258493,I258092,I258476);
DFFARX1 I_15067  ( .D(I258493), .CLK(I2350), .RSTB(I257993), .Q(I257970) );
nand I_15068 (I257979,I258397,I258321);
not I_15069 (I258571,I2357);
nand I_15070 (I258588,I29173,I29155);
and I_15071 (I258605,I258588,I29167);
DFFARX1 I_15072  ( .D(I258605), .CLK(I2350), .RSTB(I258571), .Q(I258622) );
not I_15073 (I258639,I258622);
DFFARX1 I_15074  ( .D(I258622), .CLK(I2350), .RSTB(I258571), .Q(I258539) );
nor I_15075 (I258670,I29170,I29155);
DFFARX1 I_15076  ( .D(I29179), .CLK(I2350), .RSTB(I258571), .Q(I258687) );
DFFARX1 I_15077  ( .D(I258687), .CLK(I2350), .RSTB(I258571), .Q(I258704) );
not I_15078 (I258542,I258704);
DFFARX1 I_15079  ( .D(I258687), .CLK(I2350), .RSTB(I258571), .Q(I258735) );
and I_15080 (I258536,I258622,I258735);
nand I_15081 (I258766,I29158,I29182);
and I_15082 (I258783,I258766,I29161);
DFFARX1 I_15083  ( .D(I258783), .CLK(I2350), .RSTB(I258571), .Q(I258800) );
nor I_15084 (I258817,I258800,I258639);
not I_15085 (I258834,I258800);
nand I_15086 (I258545,I258622,I258834);
DFFARX1 I_15087  ( .D(I29164), .CLK(I2350), .RSTB(I258571), .Q(I258865) );
and I_15088 (I258882,I258865,I29176);
nor I_15089 (I258899,I258882,I258800);
nor I_15090 (I258916,I258882,I258834);
nand I_15091 (I258551,I258670,I258916);
not I_15092 (I258554,I258882);
DFFARX1 I_15093  ( .D(I258882), .CLK(I2350), .RSTB(I258571), .Q(I258533) );
DFFARX1 I_15094  ( .D(I29152), .CLK(I2350), .RSTB(I258571), .Q(I258975) );
nand I_15095 (I258992,I258975,I258687);
and I_15096 (I259009,I258670,I258992);
DFFARX1 I_15097  ( .D(I259009), .CLK(I2350), .RSTB(I258571), .Q(I258563) );
nor I_15098 (I258560,I258975,I258882);
and I_15099 (I259054,I258975,I258817);
or I_15100 (I259071,I258670,I259054);
DFFARX1 I_15101  ( .D(I259071), .CLK(I2350), .RSTB(I258571), .Q(I258548) );
nand I_15102 (I258557,I258975,I258899);
not I_15103 (I259149,I2357);
nand I_15104 (I259166,I283244,I283232);
and I_15105 (I259183,I259166,I283226);
DFFARX1 I_15106  ( .D(I259183), .CLK(I2350), .RSTB(I259149), .Q(I259200) );
not I_15107 (I259217,I259200);
DFFARX1 I_15108  ( .D(I259200), .CLK(I2350), .RSTB(I259149), .Q(I259117) );
nor I_15109 (I259248,I283223,I283232);
DFFARX1 I_15110  ( .D(I283217), .CLK(I2350), .RSTB(I259149), .Q(I259265) );
DFFARX1 I_15111  ( .D(I259265), .CLK(I2350), .RSTB(I259149), .Q(I259282) );
not I_15112 (I259120,I259282);
DFFARX1 I_15113  ( .D(I259265), .CLK(I2350), .RSTB(I259149), .Q(I259313) );
and I_15114 (I259114,I259200,I259313);
nand I_15115 (I259344,I283220,I283235);
and I_15116 (I259361,I259344,I283247);
DFFARX1 I_15117  ( .D(I259361), .CLK(I2350), .RSTB(I259149), .Q(I259378) );
nor I_15118 (I259395,I259378,I259217);
not I_15119 (I259412,I259378);
nand I_15120 (I259123,I259200,I259412);
DFFARX1 I_15121  ( .D(I283238), .CLK(I2350), .RSTB(I259149), .Q(I259443) );
and I_15122 (I259460,I259443,I283229);
nor I_15123 (I259477,I259460,I259378);
nor I_15124 (I259494,I259460,I259412);
nand I_15125 (I259129,I259248,I259494);
not I_15126 (I259132,I259460);
DFFARX1 I_15127  ( .D(I259460), .CLK(I2350), .RSTB(I259149), .Q(I259111) );
DFFARX1 I_15128  ( .D(I283241), .CLK(I2350), .RSTB(I259149), .Q(I259553) );
nand I_15129 (I259570,I259553,I259265);
and I_15130 (I259587,I259248,I259570);
DFFARX1 I_15131  ( .D(I259587), .CLK(I2350), .RSTB(I259149), .Q(I259141) );
nor I_15132 (I259138,I259553,I259460);
and I_15133 (I259632,I259553,I259395);
or I_15134 (I259649,I259248,I259632);
DFFARX1 I_15135  ( .D(I259649), .CLK(I2350), .RSTB(I259149), .Q(I259126) );
nand I_15136 (I259135,I259553,I259477);
not I_15137 (I259727,I2357);
nand I_15138 (I259744,I293359,I293347);
and I_15139 (I259761,I259744,I293341);
DFFARX1 I_15140  ( .D(I259761), .CLK(I2350), .RSTB(I259727), .Q(I259778) );
not I_15141 (I259795,I259778);
DFFARX1 I_15142  ( .D(I259778), .CLK(I2350), .RSTB(I259727), .Q(I259695) );
nor I_15143 (I259826,I293338,I293347);
DFFARX1 I_15144  ( .D(I293332), .CLK(I2350), .RSTB(I259727), .Q(I259843) );
DFFARX1 I_15145  ( .D(I259843), .CLK(I2350), .RSTB(I259727), .Q(I259860) );
not I_15146 (I259698,I259860);
DFFARX1 I_15147  ( .D(I259843), .CLK(I2350), .RSTB(I259727), .Q(I259891) );
and I_15148 (I259692,I259778,I259891);
nand I_15149 (I259922,I293335,I293350);
and I_15150 (I259939,I259922,I293362);
DFFARX1 I_15151  ( .D(I259939), .CLK(I2350), .RSTB(I259727), .Q(I259956) );
nor I_15152 (I259973,I259956,I259795);
not I_15153 (I259990,I259956);
nand I_15154 (I259701,I259778,I259990);
DFFARX1 I_15155  ( .D(I293353), .CLK(I2350), .RSTB(I259727), .Q(I260021) );
and I_15156 (I260038,I260021,I293344);
nor I_15157 (I260055,I260038,I259956);
nor I_15158 (I260072,I260038,I259990);
nand I_15159 (I259707,I259826,I260072);
not I_15160 (I259710,I260038);
DFFARX1 I_15161  ( .D(I260038), .CLK(I2350), .RSTB(I259727), .Q(I259689) );
DFFARX1 I_15162  ( .D(I293356), .CLK(I2350), .RSTB(I259727), .Q(I260131) );
nand I_15163 (I260148,I260131,I259843);
and I_15164 (I260165,I259826,I260148);
DFFARX1 I_15165  ( .D(I260165), .CLK(I2350), .RSTB(I259727), .Q(I259719) );
nor I_15166 (I259716,I260131,I260038);
and I_15167 (I260210,I260131,I259973);
or I_15168 (I260227,I259826,I260210);
DFFARX1 I_15169  ( .D(I260227), .CLK(I2350), .RSTB(I259727), .Q(I259704) );
nand I_15170 (I259713,I260131,I260055);
not I_15171 (I260305,I2357);
nand I_15172 (I260322,I118069,I118054);
and I_15173 (I260339,I260322,I118063);
DFFARX1 I_15174  ( .D(I260339), .CLK(I2350), .RSTB(I260305), .Q(I260356) );
not I_15175 (I260373,I260356);
DFFARX1 I_15176  ( .D(I260356), .CLK(I2350), .RSTB(I260305), .Q(I260273) );
nor I_15177 (I260404,I118072,I118054);
DFFARX1 I_15178  ( .D(I118051), .CLK(I2350), .RSTB(I260305), .Q(I260421) );
DFFARX1 I_15179  ( .D(I260421), .CLK(I2350), .RSTB(I260305), .Q(I260438) );
not I_15180 (I260276,I260438);
DFFARX1 I_15181  ( .D(I260421), .CLK(I2350), .RSTB(I260305), .Q(I260469) );
and I_15182 (I260270,I260356,I260469);
nand I_15183 (I260500,I118075,I118048);
and I_15184 (I260517,I260500,I118066);
DFFARX1 I_15185  ( .D(I260517), .CLK(I2350), .RSTB(I260305), .Q(I260534) );
nor I_15186 (I260551,I260534,I260373);
not I_15187 (I260568,I260534);
nand I_15188 (I260279,I260356,I260568);
DFFARX1 I_15189  ( .D(I118060), .CLK(I2350), .RSTB(I260305), .Q(I260599) );
and I_15190 (I260616,I260599,I118045);
nor I_15191 (I260633,I260616,I260534);
nor I_15192 (I260650,I260616,I260568);
nand I_15193 (I260285,I260404,I260650);
not I_15194 (I260288,I260616);
DFFARX1 I_15195  ( .D(I260616), .CLK(I2350), .RSTB(I260305), .Q(I260267) );
DFFARX1 I_15196  ( .D(I118057), .CLK(I2350), .RSTB(I260305), .Q(I260709) );
nand I_15197 (I260726,I260709,I260421);
and I_15198 (I260743,I260404,I260726);
DFFARX1 I_15199  ( .D(I260743), .CLK(I2350), .RSTB(I260305), .Q(I260297) );
nor I_15200 (I260294,I260709,I260616);
and I_15201 (I260788,I260709,I260551);
or I_15202 (I260805,I260404,I260788);
DFFARX1 I_15203  ( .D(I260805), .CLK(I2350), .RSTB(I260305), .Q(I260282) );
nand I_15204 (I260291,I260709,I260633);
not I_15205 (I260883,I2357);
nand I_15206 (I260900,I213396,I213393);
and I_15207 (I260917,I260900,I213405);
DFFARX1 I_15208  ( .D(I260917), .CLK(I2350), .RSTB(I260883), .Q(I260934) );
not I_15209 (I260951,I260934);
DFFARX1 I_15210  ( .D(I260934), .CLK(I2350), .RSTB(I260883), .Q(I260851) );
nor I_15211 (I260982,I213402,I213393);
DFFARX1 I_15212  ( .D(I213408), .CLK(I2350), .RSTB(I260883), .Q(I260999) );
DFFARX1 I_15213  ( .D(I260999), .CLK(I2350), .RSTB(I260883), .Q(I261016) );
not I_15214 (I260854,I261016);
DFFARX1 I_15215  ( .D(I260999), .CLK(I2350), .RSTB(I260883), .Q(I261047) );
and I_15216 (I260848,I260934,I261047);
nand I_15217 (I261078,I213384,I213387);
and I_15218 (I261095,I261078,I213411);
DFFARX1 I_15219  ( .D(I261095), .CLK(I2350), .RSTB(I260883), .Q(I261112) );
nor I_15220 (I261129,I261112,I260951);
not I_15221 (I261146,I261112);
nand I_15222 (I260857,I260934,I261146);
DFFARX1 I_15223  ( .D(I213390), .CLK(I2350), .RSTB(I260883), .Q(I261177) );
and I_15224 (I261194,I261177,I213381);
nor I_15225 (I261211,I261194,I261112);
nor I_15226 (I261228,I261194,I261146);
nand I_15227 (I260863,I260982,I261228);
not I_15228 (I260866,I261194);
DFFARX1 I_15229  ( .D(I261194), .CLK(I2350), .RSTB(I260883), .Q(I260845) );
DFFARX1 I_15230  ( .D(I213399), .CLK(I2350), .RSTB(I260883), .Q(I261287) );
nand I_15231 (I261304,I261287,I260999);
and I_15232 (I261321,I260982,I261304);
DFFARX1 I_15233  ( .D(I261321), .CLK(I2350), .RSTB(I260883), .Q(I260875) );
nor I_15234 (I260872,I261287,I261194);
and I_15235 (I261366,I261287,I261129);
or I_15236 (I261383,I260982,I261366);
DFFARX1 I_15237  ( .D(I261383), .CLK(I2350), .RSTB(I260883), .Q(I260860) );
nand I_15238 (I260869,I261287,I261211);
not I_15239 (I261461,I2357);
nand I_15240 (I261478,I176137,I176164);
and I_15241 (I261495,I261478,I176152);
DFFARX1 I_15242  ( .D(I261495), .CLK(I2350), .RSTB(I261461), .Q(I261512) );
not I_15243 (I261529,I261512);
DFFARX1 I_15244  ( .D(I261512), .CLK(I2350), .RSTB(I261461), .Q(I261429) );
nor I_15245 (I261560,I176140,I176164);
DFFARX1 I_15246  ( .D(I176155), .CLK(I2350), .RSTB(I261461), .Q(I261577) );
DFFARX1 I_15247  ( .D(I261577), .CLK(I2350), .RSTB(I261461), .Q(I261594) );
not I_15248 (I261432,I261594);
DFFARX1 I_15249  ( .D(I261577), .CLK(I2350), .RSTB(I261461), .Q(I261625) );
and I_15250 (I261426,I261512,I261625);
nand I_15251 (I261656,I176149,I176146);
and I_15252 (I261673,I261656,I176143);
DFFARX1 I_15253  ( .D(I261673), .CLK(I2350), .RSTB(I261461), .Q(I261690) );
nor I_15254 (I261707,I261690,I261529);
not I_15255 (I261724,I261690);
nand I_15256 (I261435,I261512,I261724);
DFFARX1 I_15257  ( .D(I176158), .CLK(I2350), .RSTB(I261461), .Q(I261755) );
and I_15258 (I261772,I261755,I176134);
nor I_15259 (I261789,I261772,I261690);
nor I_15260 (I261806,I261772,I261724);
nand I_15261 (I261441,I261560,I261806);
not I_15262 (I261444,I261772);
DFFARX1 I_15263  ( .D(I261772), .CLK(I2350), .RSTB(I261461), .Q(I261423) );
DFFARX1 I_15264  ( .D(I176161), .CLK(I2350), .RSTB(I261461), .Q(I261865) );
nand I_15265 (I261882,I261865,I261577);
and I_15266 (I261899,I261560,I261882);
DFFARX1 I_15267  ( .D(I261899), .CLK(I2350), .RSTB(I261461), .Q(I261453) );
nor I_15268 (I261450,I261865,I261772);
and I_15269 (I261944,I261865,I261707);
or I_15270 (I261961,I261560,I261944);
DFFARX1 I_15271  ( .D(I261961), .CLK(I2350), .RSTB(I261461), .Q(I261438) );
nand I_15272 (I261447,I261865,I261789);
not I_15273 (I262039,I2357);
nand I_15274 (I262056,I86061,I86040);
and I_15275 (I262073,I262056,I86037);
DFFARX1 I_15276  ( .D(I262073), .CLK(I2350), .RSTB(I262039), .Q(I262090) );
not I_15277 (I262107,I262090);
DFFARX1 I_15278  ( .D(I262090), .CLK(I2350), .RSTB(I262039), .Q(I262007) );
nor I_15279 (I262138,I86046,I86040);
DFFARX1 I_15280  ( .D(I86034), .CLK(I2350), .RSTB(I262039), .Q(I262155) );
DFFARX1 I_15281  ( .D(I262155), .CLK(I2350), .RSTB(I262039), .Q(I262172) );
not I_15282 (I262010,I262172);
DFFARX1 I_15283  ( .D(I262155), .CLK(I2350), .RSTB(I262039), .Q(I262203) );
and I_15284 (I262004,I262090,I262203);
nand I_15285 (I262234,I86064,I86055);
and I_15286 (I262251,I262234,I86052);
DFFARX1 I_15287  ( .D(I262251), .CLK(I2350), .RSTB(I262039), .Q(I262268) );
nor I_15288 (I262285,I262268,I262107);
not I_15289 (I262302,I262268);
nand I_15290 (I262013,I262090,I262302);
DFFARX1 I_15291  ( .D(I86049), .CLK(I2350), .RSTB(I262039), .Q(I262333) );
and I_15292 (I262350,I262333,I86058);
nor I_15293 (I262367,I262350,I262268);
nor I_15294 (I262384,I262350,I262302);
nand I_15295 (I262019,I262138,I262384);
not I_15296 (I262022,I262350);
DFFARX1 I_15297  ( .D(I262350), .CLK(I2350), .RSTB(I262039), .Q(I262001) );
DFFARX1 I_15298  ( .D(I86043), .CLK(I2350), .RSTB(I262039), .Q(I262443) );
nand I_15299 (I262460,I262443,I262155);
and I_15300 (I262477,I262138,I262460);
DFFARX1 I_15301  ( .D(I262477), .CLK(I2350), .RSTB(I262039), .Q(I262031) );
nor I_15302 (I262028,I262443,I262350);
and I_15303 (I262522,I262443,I262285);
or I_15304 (I262539,I262138,I262522);
DFFARX1 I_15305  ( .D(I262539), .CLK(I2350), .RSTB(I262039), .Q(I262016) );
nand I_15306 (I262025,I262443,I262367);
not I_15307 (I262617,I2357);
nand I_15308 (I262634,I212750,I212747);
and I_15309 (I262651,I262634,I212759);
DFFARX1 I_15310  ( .D(I262651), .CLK(I2350), .RSTB(I262617), .Q(I262668) );
not I_15311 (I262685,I262668);
DFFARX1 I_15312  ( .D(I262668), .CLK(I2350), .RSTB(I262617), .Q(I262585) );
nor I_15313 (I262716,I212756,I212747);
DFFARX1 I_15314  ( .D(I212762), .CLK(I2350), .RSTB(I262617), .Q(I262733) );
DFFARX1 I_15315  ( .D(I262733), .CLK(I2350), .RSTB(I262617), .Q(I262750) );
not I_15316 (I262588,I262750);
DFFARX1 I_15317  ( .D(I262733), .CLK(I2350), .RSTB(I262617), .Q(I262781) );
and I_15318 (I262582,I262668,I262781);
nand I_15319 (I262812,I212738,I212741);
and I_15320 (I262829,I262812,I212765);
DFFARX1 I_15321  ( .D(I262829), .CLK(I2350), .RSTB(I262617), .Q(I262846) );
nor I_15322 (I262863,I262846,I262685);
not I_15323 (I262880,I262846);
nand I_15324 (I262591,I262668,I262880);
DFFARX1 I_15325  ( .D(I212744), .CLK(I2350), .RSTB(I262617), .Q(I262911) );
and I_15326 (I262928,I262911,I212735);
nor I_15327 (I262945,I262928,I262846);
nor I_15328 (I262962,I262928,I262880);
nand I_15329 (I262597,I262716,I262962);
not I_15330 (I262600,I262928);
DFFARX1 I_15331  ( .D(I262928), .CLK(I2350), .RSTB(I262617), .Q(I262579) );
DFFARX1 I_15332  ( .D(I212753), .CLK(I2350), .RSTB(I262617), .Q(I263021) );
nand I_15333 (I263038,I263021,I262733);
and I_15334 (I263055,I262716,I263038);
DFFARX1 I_15335  ( .D(I263055), .CLK(I2350), .RSTB(I262617), .Q(I262609) );
nor I_15336 (I262606,I263021,I262928);
and I_15337 (I263100,I263021,I262863);
or I_15338 (I263117,I262716,I263100);
DFFARX1 I_15339  ( .D(I263117), .CLK(I2350), .RSTB(I262617), .Q(I262594) );
nand I_15340 (I262603,I263021,I262945);
not I_15341 (I263195,I2357);
nand I_15342 (I263212,I82791,I82773);
and I_15343 (I263229,I263212,I82785);
DFFARX1 I_15344  ( .D(I263229), .CLK(I2350), .RSTB(I263195), .Q(I263246) );
not I_15345 (I263263,I263246);
DFFARX1 I_15346  ( .D(I263246), .CLK(I2350), .RSTB(I263195), .Q(I263163) );
nor I_15347 (I263294,I82788,I82773);
DFFARX1 I_15348  ( .D(I82797), .CLK(I2350), .RSTB(I263195), .Q(I263311) );
DFFARX1 I_15349  ( .D(I263311), .CLK(I2350), .RSTB(I263195), .Q(I263328) );
not I_15350 (I263166,I263328);
DFFARX1 I_15351  ( .D(I263311), .CLK(I2350), .RSTB(I263195), .Q(I263359) );
and I_15352 (I263160,I263246,I263359);
nand I_15353 (I263390,I82776,I82800);
and I_15354 (I263407,I263390,I82779);
DFFARX1 I_15355  ( .D(I263407), .CLK(I2350), .RSTB(I263195), .Q(I263424) );
nor I_15356 (I263441,I263424,I263263);
not I_15357 (I263458,I263424);
nand I_15358 (I263169,I263246,I263458);
DFFARX1 I_15359  ( .D(I82782), .CLK(I2350), .RSTB(I263195), .Q(I263489) );
and I_15360 (I263506,I263489,I82794);
nor I_15361 (I263523,I263506,I263424);
nor I_15362 (I263540,I263506,I263458);
nand I_15363 (I263175,I263294,I263540);
not I_15364 (I263178,I263506);
DFFARX1 I_15365  ( .D(I263506), .CLK(I2350), .RSTB(I263195), .Q(I263157) );
DFFARX1 I_15366  ( .D(I82770), .CLK(I2350), .RSTB(I263195), .Q(I263599) );
nand I_15367 (I263616,I263599,I263311);
and I_15368 (I263633,I263294,I263616);
DFFARX1 I_15369  ( .D(I263633), .CLK(I2350), .RSTB(I263195), .Q(I263187) );
nor I_15370 (I263184,I263599,I263506);
and I_15371 (I263678,I263599,I263441);
or I_15372 (I263695,I263294,I263678);
DFFARX1 I_15373  ( .D(I263695), .CLK(I2350), .RSTB(I263195), .Q(I263172) );
nand I_15374 (I263181,I263599,I263523);
not I_15375 (I263773,I2357);
nand I_15376 (I263790,I75685,I75667);
and I_15377 (I263807,I263790,I75679);
DFFARX1 I_15378  ( .D(I263807), .CLK(I2350), .RSTB(I263773), .Q(I263824) );
not I_15379 (I263841,I263824);
DFFARX1 I_15380  ( .D(I263824), .CLK(I2350), .RSTB(I263773), .Q(I263741) );
nor I_15381 (I263872,I75682,I75667);
DFFARX1 I_15382  ( .D(I75691), .CLK(I2350), .RSTB(I263773), .Q(I263889) );
DFFARX1 I_15383  ( .D(I263889), .CLK(I2350), .RSTB(I263773), .Q(I263906) );
not I_15384 (I263744,I263906);
DFFARX1 I_15385  ( .D(I263889), .CLK(I2350), .RSTB(I263773), .Q(I263937) );
and I_15386 (I263738,I263824,I263937);
nand I_15387 (I263968,I75670,I75694);
and I_15388 (I263985,I263968,I75673);
DFFARX1 I_15389  ( .D(I263985), .CLK(I2350), .RSTB(I263773), .Q(I264002) );
nor I_15390 (I264019,I264002,I263841);
not I_15391 (I264036,I264002);
nand I_15392 (I263747,I263824,I264036);
DFFARX1 I_15393  ( .D(I75676), .CLK(I2350), .RSTB(I263773), .Q(I264067) );
and I_15394 (I264084,I264067,I75688);
nor I_15395 (I264101,I264084,I264002);
nor I_15396 (I264118,I264084,I264036);
nand I_15397 (I263753,I263872,I264118);
not I_15398 (I263756,I264084);
DFFARX1 I_15399  ( .D(I264084), .CLK(I2350), .RSTB(I263773), .Q(I263735) );
DFFARX1 I_15400  ( .D(I75664), .CLK(I2350), .RSTB(I263773), .Q(I264177) );
nand I_15401 (I264194,I264177,I263889);
and I_15402 (I264211,I263872,I264194);
DFFARX1 I_15403  ( .D(I264211), .CLK(I2350), .RSTB(I263773), .Q(I263765) );
nor I_15404 (I263762,I264177,I264084);
and I_15405 (I264256,I264177,I264019);
or I_15406 (I264273,I263872,I264256);
DFFARX1 I_15407  ( .D(I264273), .CLK(I2350), .RSTB(I263773), .Q(I263750) );
nand I_15408 (I263759,I264177,I264101);
not I_15409 (I264351,I2357);
nand I_15410 (I264368,I158236,I158263);
and I_15411 (I264385,I264368,I158251);
DFFARX1 I_15412  ( .D(I264385), .CLK(I2350), .RSTB(I264351), .Q(I264402) );
not I_15413 (I264419,I264402);
DFFARX1 I_15414  ( .D(I264402), .CLK(I2350), .RSTB(I264351), .Q(I264319) );
nor I_15415 (I264450,I158239,I158263);
DFFARX1 I_15416  ( .D(I158254), .CLK(I2350), .RSTB(I264351), .Q(I264467) );
DFFARX1 I_15417  ( .D(I264467), .CLK(I2350), .RSTB(I264351), .Q(I264484) );
not I_15418 (I264322,I264484);
DFFARX1 I_15419  ( .D(I264467), .CLK(I2350), .RSTB(I264351), .Q(I264515) );
and I_15420 (I264316,I264402,I264515);
nand I_15421 (I264546,I158248,I158245);
and I_15422 (I264563,I264546,I158242);
DFFARX1 I_15423  ( .D(I264563), .CLK(I2350), .RSTB(I264351), .Q(I264580) );
nor I_15424 (I264597,I264580,I264419);
not I_15425 (I264614,I264580);
nand I_15426 (I264325,I264402,I264614);
DFFARX1 I_15427  ( .D(I158257), .CLK(I2350), .RSTB(I264351), .Q(I264645) );
and I_15428 (I264662,I264645,I158233);
nor I_15429 (I264679,I264662,I264580);
nor I_15430 (I264696,I264662,I264614);
nand I_15431 (I264331,I264450,I264696);
not I_15432 (I264334,I264662);
DFFARX1 I_15433  ( .D(I264662), .CLK(I2350), .RSTB(I264351), .Q(I264313) );
DFFARX1 I_15434  ( .D(I158260), .CLK(I2350), .RSTB(I264351), .Q(I264755) );
nand I_15435 (I264772,I264755,I264467);
and I_15436 (I264789,I264450,I264772);
DFFARX1 I_15437  ( .D(I264789), .CLK(I2350), .RSTB(I264351), .Q(I264343) );
nor I_15438 (I264340,I264755,I264662);
and I_15439 (I264834,I264755,I264597);
or I_15440 (I264851,I264450,I264834);
DFFARX1 I_15441  ( .D(I264851), .CLK(I2350), .RSTB(I264351), .Q(I264328) );
nand I_15442 (I264337,I264755,I264679);
not I_15443 (I264929,I2357);
nand I_15444 (I264946,I114499,I114484);
and I_15445 (I264963,I264946,I114493);
DFFARX1 I_15446  ( .D(I264963), .CLK(I2350), .RSTB(I264929), .Q(I264980) );
not I_15447 (I264997,I264980);
DFFARX1 I_15448  ( .D(I264980), .CLK(I2350), .RSTB(I264929), .Q(I264897) );
nor I_15449 (I265028,I114502,I114484);
DFFARX1 I_15450  ( .D(I114481), .CLK(I2350), .RSTB(I264929), .Q(I265045) );
DFFARX1 I_15451  ( .D(I265045), .CLK(I2350), .RSTB(I264929), .Q(I265062) );
not I_15452 (I264900,I265062);
DFFARX1 I_15453  ( .D(I265045), .CLK(I2350), .RSTB(I264929), .Q(I265093) );
and I_15454 (I264894,I264980,I265093);
nand I_15455 (I265124,I114505,I114478);
and I_15456 (I265141,I265124,I114496);
DFFARX1 I_15457  ( .D(I265141), .CLK(I2350), .RSTB(I264929), .Q(I265158) );
nor I_15458 (I265175,I265158,I264997);
not I_15459 (I265192,I265158);
nand I_15460 (I264903,I264980,I265192);
DFFARX1 I_15461  ( .D(I114490), .CLK(I2350), .RSTB(I264929), .Q(I265223) );
and I_15462 (I265240,I265223,I114475);
nor I_15463 (I265257,I265240,I265158);
nor I_15464 (I265274,I265240,I265192);
nand I_15465 (I264909,I265028,I265274);
not I_15466 (I264912,I265240);
DFFARX1 I_15467  ( .D(I265240), .CLK(I2350), .RSTB(I264929), .Q(I264891) );
DFFARX1 I_15468  ( .D(I114487), .CLK(I2350), .RSTB(I264929), .Q(I265333) );
nand I_15469 (I265350,I265333,I265045);
and I_15470 (I265367,I265028,I265350);
DFFARX1 I_15471  ( .D(I265367), .CLK(I2350), .RSTB(I264929), .Q(I264921) );
nor I_15472 (I264918,I265333,I265240);
and I_15473 (I265412,I265333,I265175);
or I_15474 (I265429,I265028,I265412);
DFFARX1 I_15475  ( .D(I265429), .CLK(I2350), .RSTB(I264929), .Q(I264906) );
nand I_15476 (I264915,I265333,I265257);
not I_15477 (I265507,I2357);
nand I_15478 (I265524,I387408,I387420);
and I_15479 (I265541,I265524,I387393);
DFFARX1 I_15480  ( .D(I265541), .CLK(I2350), .RSTB(I265507), .Q(I265558) );
not I_15481 (I265575,I265558);
DFFARX1 I_15482  ( .D(I265558), .CLK(I2350), .RSTB(I265507), .Q(I265475) );
nor I_15483 (I265606,I387411,I387420);
DFFARX1 I_15484  ( .D(I387402), .CLK(I2350), .RSTB(I265507), .Q(I265623) );
DFFARX1 I_15485  ( .D(I265623), .CLK(I2350), .RSTB(I265507), .Q(I265640) );
not I_15486 (I265478,I265640);
DFFARX1 I_15487  ( .D(I265623), .CLK(I2350), .RSTB(I265507), .Q(I265671) );
and I_15488 (I265472,I265558,I265671);
nand I_15489 (I265702,I387399,I387405);
and I_15490 (I265719,I265702,I387417);
DFFARX1 I_15491  ( .D(I265719), .CLK(I2350), .RSTB(I265507), .Q(I265736) );
nor I_15492 (I265753,I265736,I265575);
not I_15493 (I265770,I265736);
nand I_15494 (I265481,I265558,I265770);
DFFARX1 I_15495  ( .D(I387423), .CLK(I2350), .RSTB(I265507), .Q(I265801) );
and I_15496 (I265818,I265801,I387414);
nor I_15497 (I265835,I265818,I265736);
nor I_15498 (I265852,I265818,I265770);
nand I_15499 (I265487,I265606,I265852);
not I_15500 (I265490,I265818);
DFFARX1 I_15501  ( .D(I265818), .CLK(I2350), .RSTB(I265507), .Q(I265469) );
DFFARX1 I_15502  ( .D(I387396), .CLK(I2350), .RSTB(I265507), .Q(I265911) );
nand I_15503 (I265928,I265911,I265623);
and I_15504 (I265945,I265606,I265928);
DFFARX1 I_15505  ( .D(I265945), .CLK(I2350), .RSTB(I265507), .Q(I265499) );
nor I_15506 (I265496,I265911,I265818);
and I_15507 (I265990,I265911,I265753);
or I_15508 (I266007,I265606,I265990);
DFFARX1 I_15509  ( .D(I266007), .CLK(I2350), .RSTB(I265507), .Q(I265484) );
nand I_15510 (I265493,I265911,I265835);
not I_15511 (I266085,I2357);
nand I_15512 (I266102,I188734,I188761);
and I_15513 (I266119,I266102,I188749);
DFFARX1 I_15514  ( .D(I266119), .CLK(I2350), .RSTB(I266085), .Q(I266136) );
not I_15515 (I266153,I266136);
DFFARX1 I_15516  ( .D(I266136), .CLK(I2350), .RSTB(I266085), .Q(I266053) );
nor I_15517 (I266184,I188737,I188761);
DFFARX1 I_15518  ( .D(I188752), .CLK(I2350), .RSTB(I266085), .Q(I266201) );
DFFARX1 I_15519  ( .D(I266201), .CLK(I2350), .RSTB(I266085), .Q(I266218) );
not I_15520 (I266056,I266218);
DFFARX1 I_15521  ( .D(I266201), .CLK(I2350), .RSTB(I266085), .Q(I266249) );
and I_15522 (I266050,I266136,I266249);
nand I_15523 (I266280,I188746,I188743);
and I_15524 (I266297,I266280,I188740);
DFFARX1 I_15525  ( .D(I266297), .CLK(I2350), .RSTB(I266085), .Q(I266314) );
nor I_15526 (I266331,I266314,I266153);
not I_15527 (I266348,I266314);
nand I_15528 (I266059,I266136,I266348);
DFFARX1 I_15529  ( .D(I188755), .CLK(I2350), .RSTB(I266085), .Q(I266379) );
and I_15530 (I266396,I266379,I188731);
nor I_15531 (I266413,I266396,I266314);
nor I_15532 (I266430,I266396,I266348);
nand I_15533 (I266065,I266184,I266430);
not I_15534 (I266068,I266396);
DFFARX1 I_15535  ( .D(I266396), .CLK(I2350), .RSTB(I266085), .Q(I266047) );
DFFARX1 I_15536  ( .D(I188758), .CLK(I2350), .RSTB(I266085), .Q(I266489) );
nand I_15537 (I266506,I266489,I266201);
and I_15538 (I266523,I266184,I266506);
DFFARX1 I_15539  ( .D(I266523), .CLK(I2350), .RSTB(I266085), .Q(I266077) );
nor I_15540 (I266074,I266489,I266396);
and I_15541 (I266568,I266489,I266331);
or I_15542 (I266585,I266184,I266568);
DFFARX1 I_15543  ( .D(I266585), .CLK(I2350), .RSTB(I266085), .Q(I266062) );
nand I_15544 (I266071,I266489,I266413);
not I_15545 (I266663,I2357);
or I_15546 (I266680,I214054,I214045);
or I_15547 (I266697,I214057,I214054);
nor I_15548 (I266714,I214030,I214051);
not I_15549 (I266731,I266714);
DFFARX1 I_15550  ( .D(I266714), .CLK(I2350), .RSTB(I266663), .Q(I266631) );
nand I_15551 (I266762,I266714,I266680);
not I_15552 (I266779,I214030);
and I_15553 (I266796,I266779,I214042);
nor I_15554 (I266813,I266796,I214045);
nor I_15555 (I266830,I214033,I214027);
DFFARX1 I_15556  ( .D(I266830), .CLK(I2350), .RSTB(I266663), .Q(I266847) );
nor I_15557 (I266864,I266847,I266731);
not I_15558 (I266881,I266847);
nand I_15559 (I266637,I266714,I266881);
DFFARX1 I_15560  ( .D(I266847), .CLK(I2350), .RSTB(I266663), .Q(I266628) );
nor I_15561 (I266926,I214033,I214057);
nand I_15562 (I266943,I266697,I266926);
nor I_15563 (I266652,I266680,I266926);
and I_15564 (I266974,I266926,I266864);
or I_15565 (I266991,I266813,I266974);
DFFARX1 I_15566  ( .D(I266991), .CLK(I2350), .RSTB(I266663), .Q(I266640) );
DFFARX1 I_15567  ( .D(I214036), .CLK(I2350), .RSTB(I266663), .Q(I267022) );
and I_15568 (I267039,I267022,I214048);
not I_15569 (I266646,I267039);
DFFARX1 I_15570  ( .D(I267039), .CLK(I2350), .RSTB(I266663), .Q(I267070) );
not I_15571 (I266634,I267070);
and I_15572 (I267101,I267039,I266762);
DFFARX1 I_15573  ( .D(I267101), .CLK(I2350), .RSTB(I266663), .Q(I266625) );
DFFARX1 I_15574  ( .D(I214039), .CLK(I2350), .RSTB(I266663), .Q(I267132) );
and I_15575 (I267149,I267132,I266943);
DFFARX1 I_15576  ( .D(I267149), .CLK(I2350), .RSTB(I266663), .Q(I266655) );
nor I_15577 (I267180,I267132,I267039);
nand I_15578 (I266649,I266813,I267180);
nor I_15579 (I267211,I267132,I266881);
nand I_15580 (I266643,I266697,I267211);
not I_15581 (I267275,I2357);
or I_15582 (I267292,I187408,I187405);
or I_15583 (I267309,I187420,I187408);
nor I_15584 (I267326,I187435,I187411);
not I_15585 (I267343,I267326);
DFFARX1 I_15586  ( .D(I267326), .CLK(I2350), .RSTB(I267275), .Q(I267243) );
nand I_15587 (I267374,I267326,I267292);
not I_15588 (I267391,I187435);
and I_15589 (I267408,I267391,I187429);
nor I_15590 (I267425,I267408,I187405);
nor I_15591 (I267442,I187423,I187432);
DFFARX1 I_15592  ( .D(I267442), .CLK(I2350), .RSTB(I267275), .Q(I267459) );
nor I_15593 (I267476,I267459,I267343);
not I_15594 (I267493,I267459);
nand I_15595 (I267249,I267326,I267493);
DFFARX1 I_15596  ( .D(I267459), .CLK(I2350), .RSTB(I267275), .Q(I267240) );
nor I_15597 (I267538,I187423,I187420);
nand I_15598 (I267555,I267309,I267538);
nor I_15599 (I267264,I267292,I267538);
and I_15600 (I267586,I267538,I267476);
or I_15601 (I267603,I267425,I267586);
DFFARX1 I_15602  ( .D(I267603), .CLK(I2350), .RSTB(I267275), .Q(I267252) );
DFFARX1 I_15603  ( .D(I187417), .CLK(I2350), .RSTB(I267275), .Q(I267634) );
and I_15604 (I267651,I267634,I187414);
not I_15605 (I267258,I267651);
DFFARX1 I_15606  ( .D(I267651), .CLK(I2350), .RSTB(I267275), .Q(I267682) );
not I_15607 (I267246,I267682);
and I_15608 (I267713,I267651,I267374);
DFFARX1 I_15609  ( .D(I267713), .CLK(I2350), .RSTB(I267275), .Q(I267237) );
DFFARX1 I_15610  ( .D(I187426), .CLK(I2350), .RSTB(I267275), .Q(I267744) );
and I_15611 (I267761,I267744,I267555);
DFFARX1 I_15612  ( .D(I267761), .CLK(I2350), .RSTB(I267275), .Q(I267267) );
nor I_15613 (I267792,I267744,I267651);
nand I_15614 (I267261,I267425,I267792);
nor I_15615 (I267823,I267744,I267493);
nand I_15616 (I267255,I267309,I267823);
not I_15617 (I267887,I2357);
or I_15618 (I267904,I337032,I337026);
or I_15619 (I267921,I337035,I337032);
nor I_15620 (I267938,I337029,I337011);
not I_15621 (I267955,I267938);
DFFARX1 I_15622  ( .D(I267938), .CLK(I2350), .RSTB(I267887), .Q(I267855) );
nand I_15623 (I267986,I267938,I267904);
not I_15624 (I268003,I337029);
and I_15625 (I268020,I268003,I337008);
nor I_15626 (I268037,I268020,I337026);
nor I_15627 (I268054,I337023,I337005);
DFFARX1 I_15628  ( .D(I268054), .CLK(I2350), .RSTB(I267887), .Q(I268071) );
nor I_15629 (I268088,I268071,I267955);
not I_15630 (I268105,I268071);
nand I_15631 (I267861,I267938,I268105);
DFFARX1 I_15632  ( .D(I268071), .CLK(I2350), .RSTB(I267887), .Q(I267852) );
nor I_15633 (I268150,I337023,I337035);
nand I_15634 (I268167,I267921,I268150);
nor I_15635 (I267876,I267904,I268150);
and I_15636 (I268198,I268150,I268088);
or I_15637 (I268215,I268037,I268198);
DFFARX1 I_15638  ( .D(I268215), .CLK(I2350), .RSTB(I267887), .Q(I267864) );
DFFARX1 I_15639  ( .D(I337017), .CLK(I2350), .RSTB(I267887), .Q(I268246) );
and I_15640 (I268263,I268246,I337020);
not I_15641 (I267870,I268263);
DFFARX1 I_15642  ( .D(I268263), .CLK(I2350), .RSTB(I267887), .Q(I268294) );
not I_15643 (I267858,I268294);
and I_15644 (I268325,I268263,I267986);
DFFARX1 I_15645  ( .D(I268325), .CLK(I2350), .RSTB(I267887), .Q(I267849) );
DFFARX1 I_15646  ( .D(I337014), .CLK(I2350), .RSTB(I267887), .Q(I268356) );
and I_15647 (I268373,I268356,I268167);
DFFARX1 I_15648  ( .D(I268373), .CLK(I2350), .RSTB(I267887), .Q(I267879) );
nor I_15649 (I268404,I268356,I268263);
nand I_15650 (I267873,I268037,I268404);
nor I_15651 (I268435,I268356,I268105);
nand I_15652 (I267867,I267921,I268435);
not I_15653 (I268499,I2357);
or I_15654 (I268516,I297521,I297527);
or I_15655 (I268533,I297524,I297521);
nor I_15656 (I268550,I297497,I297515);
not I_15657 (I268567,I268550);
DFFARX1 I_15658  ( .D(I268550), .CLK(I2350), .RSTB(I268499), .Q(I268467) );
nand I_15659 (I268598,I268550,I268516);
not I_15660 (I268615,I297497);
and I_15661 (I268632,I268615,I297509);
nor I_15662 (I268649,I268632,I297527);
nor I_15663 (I268666,I297512,I297500);
DFFARX1 I_15664  ( .D(I268666), .CLK(I2350), .RSTB(I268499), .Q(I268683) );
nor I_15665 (I268700,I268683,I268567);
not I_15666 (I268717,I268683);
nand I_15667 (I268473,I268550,I268717);
DFFARX1 I_15668  ( .D(I268683), .CLK(I2350), .RSTB(I268499), .Q(I268464) );
nor I_15669 (I268762,I297512,I297524);
nand I_15670 (I268779,I268533,I268762);
nor I_15671 (I268488,I268516,I268762);
and I_15672 (I268810,I268762,I268700);
or I_15673 (I268827,I268649,I268810);
DFFARX1 I_15674  ( .D(I268827), .CLK(I2350), .RSTB(I268499), .Q(I268476) );
DFFARX1 I_15675  ( .D(I297503), .CLK(I2350), .RSTB(I268499), .Q(I268858) );
and I_15676 (I268875,I268858,I297518);
not I_15677 (I268482,I268875);
DFFARX1 I_15678  ( .D(I268875), .CLK(I2350), .RSTB(I268499), .Q(I268906) );
not I_15679 (I268470,I268906);
and I_15680 (I268937,I268875,I268598);
DFFARX1 I_15681  ( .D(I268937), .CLK(I2350), .RSTB(I268499), .Q(I268461) );
DFFARX1 I_15682  ( .D(I297506), .CLK(I2350), .RSTB(I268499), .Q(I268968) );
and I_15683 (I268985,I268968,I268779);
DFFARX1 I_15684  ( .D(I268985), .CLK(I2350), .RSTB(I268499), .Q(I268491) );
nor I_15685 (I269016,I268968,I268875);
nand I_15686 (I268485,I268649,I269016);
nor I_15687 (I269047,I268968,I268717);
nand I_15688 (I268479,I268533,I269047);
not I_15689 (I269111,I2357);
or I_15690 (I269128,I388549,I388564);
or I_15691 (I269145,I388558,I388549);
nor I_15692 (I269162,I388555,I388552);
not I_15693 (I269179,I269162);
DFFARX1 I_15694  ( .D(I269162), .CLK(I2350), .RSTB(I269111), .Q(I269079) );
nand I_15695 (I269210,I269162,I269128);
not I_15696 (I269227,I388555);
and I_15697 (I269244,I269227,I388570);
nor I_15698 (I269261,I269244,I388564);
nor I_15699 (I269278,I388561,I388567);
DFFARX1 I_15700  ( .D(I269278), .CLK(I2350), .RSTB(I269111), .Q(I269295) );
nor I_15701 (I269312,I269295,I269179);
not I_15702 (I269329,I269295);
nand I_15703 (I269085,I269162,I269329);
DFFARX1 I_15704  ( .D(I269295), .CLK(I2350), .RSTB(I269111), .Q(I269076) );
nor I_15705 (I269374,I388561,I388558);
nand I_15706 (I269391,I269145,I269374);
nor I_15707 (I269100,I269128,I269374);
and I_15708 (I269422,I269374,I269312);
or I_15709 (I269439,I269261,I269422);
DFFARX1 I_15710  ( .D(I269439), .CLK(I2350), .RSTB(I269111), .Q(I269088) );
DFFARX1 I_15711  ( .D(I388579), .CLK(I2350), .RSTB(I269111), .Q(I269470) );
and I_15712 (I269487,I269470,I388576);
not I_15713 (I269094,I269487);
DFFARX1 I_15714  ( .D(I269487), .CLK(I2350), .RSTB(I269111), .Q(I269518) );
not I_15715 (I269082,I269518);
and I_15716 (I269549,I269487,I269210);
DFFARX1 I_15717  ( .D(I269549), .CLK(I2350), .RSTB(I269111), .Q(I269073) );
DFFARX1 I_15718  ( .D(I388573), .CLK(I2350), .RSTB(I269111), .Q(I269580) );
and I_15719 (I269597,I269580,I269391);
DFFARX1 I_15720  ( .D(I269597), .CLK(I2350), .RSTB(I269111), .Q(I269103) );
nor I_15721 (I269628,I269580,I269487);
nand I_15722 (I269097,I269261,I269628);
nor I_15723 (I269659,I269580,I269329);
nand I_15724 (I269091,I269145,I269659);
not I_15725 (I269723,I2357);
or I_15726 (I269740,I300496,I300502);
or I_15727 (I269757,I300499,I300496);
nor I_15728 (I269774,I300472,I300490);
not I_15729 (I269791,I269774);
DFFARX1 I_15730  ( .D(I269774), .CLK(I2350), .RSTB(I269723), .Q(I269691) );
nand I_15731 (I269822,I269774,I269740);
not I_15732 (I269839,I300472);
and I_15733 (I269856,I269839,I300484);
nor I_15734 (I269873,I269856,I300502);
nor I_15735 (I269890,I300487,I300475);
DFFARX1 I_15736  ( .D(I269890), .CLK(I2350), .RSTB(I269723), .Q(I269907) );
nor I_15737 (I269924,I269907,I269791);
not I_15738 (I269941,I269907);
nand I_15739 (I269697,I269774,I269941);
DFFARX1 I_15740  ( .D(I269907), .CLK(I2350), .RSTB(I269723), .Q(I269688) );
nor I_15741 (I269986,I300487,I300499);
nand I_15742 (I270003,I269757,I269986);
nor I_15743 (I269712,I269740,I269986);
and I_15744 (I270034,I269986,I269924);
or I_15745 (I270051,I269873,I270034);
DFFARX1 I_15746  ( .D(I270051), .CLK(I2350), .RSTB(I269723), .Q(I269700) );
DFFARX1 I_15747  ( .D(I300478), .CLK(I2350), .RSTB(I269723), .Q(I270082) );
and I_15748 (I270099,I270082,I300493);
not I_15749 (I269706,I270099);
DFFARX1 I_15750  ( .D(I270099), .CLK(I2350), .RSTB(I269723), .Q(I270130) );
not I_15751 (I269694,I270130);
and I_15752 (I270161,I270099,I269822);
DFFARX1 I_15753  ( .D(I270161), .CLK(I2350), .RSTB(I269723), .Q(I269685) );
DFFARX1 I_15754  ( .D(I300481), .CLK(I2350), .RSTB(I269723), .Q(I270192) );
and I_15755 (I270209,I270192,I270003);
DFFARX1 I_15756  ( .D(I270209), .CLK(I2350), .RSTB(I269723), .Q(I269715) );
nor I_15757 (I270240,I270192,I270099);
nand I_15758 (I269709,I269873,I270240);
nor I_15759 (I270271,I270192,I269941);
nand I_15760 (I269703,I269757,I270271);
not I_15761 (I270335,I2357);
or I_15762 (I270352,I32406,I32397);
or I_15763 (I270369,I32394,I32406);
nor I_15764 (I270386,I32391,I32409);
not I_15765 (I270403,I270386);
DFFARX1 I_15766  ( .D(I270386), .CLK(I2350), .RSTB(I270335), .Q(I270303) );
nand I_15767 (I270434,I270386,I270352);
not I_15768 (I270451,I32391);
and I_15769 (I270468,I270451,I32382);
nor I_15770 (I270485,I270468,I32397);
nor I_15771 (I270502,I32385,I32388);
DFFARX1 I_15772  ( .D(I270502), .CLK(I2350), .RSTB(I270335), .Q(I270519) );
nor I_15773 (I270536,I270519,I270403);
not I_15774 (I270553,I270519);
nand I_15775 (I270309,I270386,I270553);
DFFARX1 I_15776  ( .D(I270519), .CLK(I2350), .RSTB(I270335), .Q(I270300) );
nor I_15777 (I270598,I32385,I32394);
nand I_15778 (I270615,I270369,I270598);
nor I_15779 (I270324,I270352,I270598);
and I_15780 (I270646,I270598,I270536);
or I_15781 (I270663,I270485,I270646);
DFFARX1 I_15782  ( .D(I270663), .CLK(I2350), .RSTB(I270335), .Q(I270312) );
DFFARX1 I_15783  ( .D(I32400), .CLK(I2350), .RSTB(I270335), .Q(I270694) );
and I_15784 (I270711,I270694,I32412);
not I_15785 (I270318,I270711);
DFFARX1 I_15786  ( .D(I270711), .CLK(I2350), .RSTB(I270335), .Q(I270742) );
not I_15787 (I270306,I270742);
and I_15788 (I270773,I270711,I270434);
DFFARX1 I_15789  ( .D(I270773), .CLK(I2350), .RSTB(I270335), .Q(I270297) );
DFFARX1 I_15790  ( .D(I32403), .CLK(I2350), .RSTB(I270335), .Q(I270804) );
and I_15791 (I270821,I270804,I270615);
DFFARX1 I_15792  ( .D(I270821), .CLK(I2350), .RSTB(I270335), .Q(I270327) );
nor I_15793 (I270852,I270804,I270711);
nand I_15794 (I270321,I270485,I270852);
nor I_15795 (I270883,I270804,I270553);
nand I_15796 (I270315,I270369,I270883);
not I_15797 (I270947,I2357);
or I_15798 (I270964,I35636,I35627);
or I_15799 (I270981,I35624,I35636);
nor I_15800 (I270998,I35621,I35639);
not I_15801 (I271015,I270998);
DFFARX1 I_15802  ( .D(I270998), .CLK(I2350), .RSTB(I270947), .Q(I270915) );
nand I_15803 (I271046,I270998,I270964);
not I_15804 (I271063,I35621);
and I_15805 (I271080,I271063,I35612);
nor I_15806 (I271097,I271080,I35627);
nor I_15807 (I271114,I35615,I35618);
DFFARX1 I_15808  ( .D(I271114), .CLK(I2350), .RSTB(I270947), .Q(I271131) );
nor I_15809 (I271148,I271131,I271015);
not I_15810 (I271165,I271131);
nand I_15811 (I270921,I270998,I271165);
DFFARX1 I_15812  ( .D(I271131), .CLK(I2350), .RSTB(I270947), .Q(I270912) );
nor I_15813 (I271210,I35615,I35624);
nand I_15814 (I271227,I270981,I271210);
nor I_15815 (I270936,I270964,I271210);
and I_15816 (I271258,I271210,I271148);
or I_15817 (I271275,I271097,I271258);
DFFARX1 I_15818  ( .D(I271275), .CLK(I2350), .RSTB(I270947), .Q(I270924) );
DFFARX1 I_15819  ( .D(I35630), .CLK(I2350), .RSTB(I270947), .Q(I271306) );
and I_15820 (I271323,I271306,I35642);
not I_15821 (I270930,I271323);
DFFARX1 I_15822  ( .D(I271323), .CLK(I2350), .RSTB(I270947), .Q(I271354) );
not I_15823 (I270918,I271354);
and I_15824 (I271385,I271323,I271046);
DFFARX1 I_15825  ( .D(I271385), .CLK(I2350), .RSTB(I270947), .Q(I270909) );
DFFARX1 I_15826  ( .D(I35633), .CLK(I2350), .RSTB(I270947), .Q(I271416) );
and I_15827 (I271433,I271416,I271227);
DFFARX1 I_15828  ( .D(I271433), .CLK(I2350), .RSTB(I270947), .Q(I270939) );
nor I_15829 (I271464,I271416,I271323);
nand I_15830 (I270933,I271097,I271464);
nor I_15831 (I271495,I271416,I271165);
nand I_15832 (I270927,I270981,I271495);
not I_15833 (I271559,I2357);
or I_15834 (I271576,I287998,I287992);
or I_15835 (I271593,I287986,I287998);
nor I_15836 (I271610,I288007,I287995);
or I_15837 (I271548,I271610,I271576);
not I_15838 (I271641,I288007);
and I_15839 (I271658,I271641,I287980);
nor I_15840 (I271675,I271658,I287992);
not I_15841 (I271692,I271675);
nor I_15842 (I271709,I287983,I287977);
DFFARX1 I_15843  ( .D(I271709), .CLK(I2350), .RSTB(I271559), .Q(I271726) );
nor I_15844 (I271743,I271726,I271675);
nand I_15845 (I271533,I271576,I271743);
nor I_15846 (I271774,I271726,I271692);
not I_15847 (I271530,I271726);
nor I_15848 (I271805,I287983,I287986);
or I_15849 (I271542,I271576,I271805);
DFFARX1 I_15850  ( .D(I288004), .CLK(I2350), .RSTB(I271559), .Q(I271836) );
and I_15851 (I271853,I271836,I288001);
nor I_15852 (I271870,I271853,I271726);
DFFARX1 I_15853  ( .D(I271870), .CLK(I2350), .RSTB(I271559), .Q(I271536) );
nor I_15854 (I271551,I271853,I271805);
not I_15855 (I271915,I271853);
nor I_15856 (I271932,I271593,I271915);
nand I_15857 (I271521,I271853,I271692);
DFFARX1 I_15858  ( .D(I287989), .CLK(I2350), .RSTB(I271559), .Q(I271963) );
nor I_15859 (I271539,I271963,I271593);
not I_15860 (I271994,I271963);
and I_15861 (I272011,I271805,I271994);
nor I_15862 (I271545,I271610,I272011);
and I_15863 (I272042,I271963,I271932);
or I_15864 (I272059,I271610,I272042);
DFFARX1 I_15865  ( .D(I272059), .CLK(I2350), .RSTB(I271559), .Q(I271524) );
nand I_15866 (I271527,I271963,I271774);
not I_15867 (I272137,I2357);
or I_15868 (I272154,I79549,I79540);
or I_15869 (I272171,I79546,I79549);
nor I_15870 (I272188,I79555,I79564);
or I_15871 (I272126,I272188,I272154);
not I_15872 (I272219,I79555);
and I_15873 (I272236,I272219,I79567);
nor I_15874 (I272253,I272236,I79540);
not I_15875 (I272270,I272253);
nor I_15876 (I272287,I79558,I79561);
DFFARX1 I_15877  ( .D(I272287), .CLK(I2350), .RSTB(I272137), .Q(I272304) );
nor I_15878 (I272321,I272304,I272253);
nand I_15879 (I272111,I272154,I272321);
nor I_15880 (I272352,I272304,I272270);
not I_15881 (I272108,I272304);
nor I_15882 (I272383,I79558,I79546);
or I_15883 (I272120,I272154,I272383);
DFFARX1 I_15884  ( .D(I79543), .CLK(I2350), .RSTB(I272137), .Q(I272414) );
and I_15885 (I272431,I272414,I79552);
nor I_15886 (I272448,I272431,I272304);
DFFARX1 I_15887  ( .D(I272448), .CLK(I2350), .RSTB(I272137), .Q(I272114) );
nor I_15888 (I272129,I272431,I272383);
not I_15889 (I272493,I272431);
nor I_15890 (I272510,I272171,I272493);
nand I_15891 (I272099,I272431,I272270);
DFFARX1 I_15892  ( .D(I79570), .CLK(I2350), .RSTB(I272137), .Q(I272541) );
nor I_15893 (I272117,I272541,I272171);
not I_15894 (I272572,I272541);
and I_15895 (I272589,I272383,I272572);
nor I_15896 (I272123,I272188,I272589);
and I_15897 (I272620,I272541,I272510);
or I_15898 (I272637,I272188,I272620);
DFFARX1 I_15899  ( .D(I272637), .CLK(I2350), .RSTB(I272137), .Q(I272102) );
nand I_15900 (I272105,I272541,I272352);
not I_15901 (I272715,I2357);
or I_15902 (I272732,I194031,I194016);
or I_15903 (I272749,I194025,I194031);
nor I_15904 (I272766,I194019,I194007);
or I_15905 (I272704,I272766,I272732);
not I_15906 (I272797,I194019);
and I_15907 (I272814,I272797,I194028);
nor I_15908 (I272831,I272814,I194016);
not I_15909 (I272848,I272831);
nor I_15910 (I272865,I194013,I194004);
DFFARX1 I_15911  ( .D(I272865), .CLK(I2350), .RSTB(I272715), .Q(I272882) );
nor I_15912 (I272899,I272882,I272831);
nand I_15913 (I272689,I272732,I272899);
nor I_15914 (I272930,I272882,I272848);
not I_15915 (I272686,I272882);
nor I_15916 (I272961,I194013,I194025);
or I_15917 (I272698,I272732,I272961);
DFFARX1 I_15918  ( .D(I194022), .CLK(I2350), .RSTB(I272715), .Q(I272992) );
and I_15919 (I273009,I272992,I194001);
nor I_15920 (I273026,I273009,I272882);
DFFARX1 I_15921  ( .D(I273026), .CLK(I2350), .RSTB(I272715), .Q(I272692) );
nor I_15922 (I272707,I273009,I272961);
not I_15923 (I273071,I273009);
nor I_15924 (I273088,I272749,I273071);
nand I_15925 (I272677,I273009,I272848);
DFFARX1 I_15926  ( .D(I194010), .CLK(I2350), .RSTB(I272715), .Q(I273119) );
nor I_15927 (I272695,I273119,I272749);
not I_15928 (I273150,I273119);
and I_15929 (I273167,I272961,I273150);
nor I_15930 (I272701,I272766,I273167);
and I_15931 (I273198,I273119,I273088);
or I_15932 (I273215,I272766,I273198);
DFFARX1 I_15933  ( .D(I273215), .CLK(I2350), .RSTB(I272715), .Q(I272680) );
nand I_15934 (I272683,I273119,I272930);
not I_15935 (I273293,I2357);
or I_15936 (I273310,I337637,I337640);
or I_15937 (I273327,I337658,I337637);
nor I_15938 (I273344,I337652,I337661);
or I_15939 (I273282,I273344,I273310);
not I_15940 (I273375,I337652);
and I_15941 (I273392,I273375,I337664);
nor I_15942 (I273409,I273392,I337640);
not I_15943 (I273426,I273409);
nor I_15944 (I273443,I337649,I337634);
DFFARX1 I_15945  ( .D(I273443), .CLK(I2350), .RSTB(I273293), .Q(I273460) );
nor I_15946 (I273477,I273460,I273409);
nand I_15947 (I273267,I273310,I273477);
nor I_15948 (I273508,I273460,I273426);
not I_15949 (I273264,I273460);
nor I_15950 (I273539,I337649,I337658);
or I_15951 (I273276,I273310,I273539);
DFFARX1 I_15952  ( .D(I337646), .CLK(I2350), .RSTB(I273293), .Q(I273570) );
and I_15953 (I273587,I273570,I337655);
nor I_15954 (I273604,I273587,I273460);
DFFARX1 I_15955  ( .D(I273604), .CLK(I2350), .RSTB(I273293), .Q(I273270) );
nor I_15956 (I273285,I273587,I273539);
not I_15957 (I273649,I273587);
nor I_15958 (I273666,I273327,I273649);
nand I_15959 (I273255,I273587,I273426);
DFFARX1 I_15960  ( .D(I337643), .CLK(I2350), .RSTB(I273293), .Q(I273697) );
nor I_15961 (I273273,I273697,I273327);
not I_15962 (I273728,I273697);
and I_15963 (I273745,I273539,I273728);
nor I_15964 (I273279,I273344,I273745);
and I_15965 (I273776,I273697,I273666);
or I_15966 (I273793,I273344,I273776);
DFFARX1 I_15967  ( .D(I273793), .CLK(I2350), .RSTB(I273293), .Q(I273258) );
nand I_15968 (I273261,I273697,I273508);
not I_15969 (I273871,I2357);
or I_15970 (I273888,I122805,I122811);
or I_15971 (I273905,I122814,I122805);
nor I_15972 (I273922,I122829,I122817);
or I_15973 (I273860,I273922,I273888);
not I_15974 (I273953,I122829);
and I_15975 (I273970,I273953,I122808);
nor I_15976 (I273987,I273970,I122811);
not I_15977 (I274004,I273987);
nor I_15978 (I274021,I122823,I122832);
DFFARX1 I_15979  ( .D(I274021), .CLK(I2350), .RSTB(I273871), .Q(I274038) );
nor I_15980 (I274055,I274038,I273987);
nand I_15981 (I273845,I273888,I274055);
nor I_15982 (I274086,I274038,I274004);
not I_15983 (I273842,I274038);
nor I_15984 (I274117,I122823,I122814);
or I_15985 (I273854,I273888,I274117);
DFFARX1 I_15986  ( .D(I122820), .CLK(I2350), .RSTB(I273871), .Q(I274148) );
and I_15987 (I274165,I274148,I122835);
nor I_15988 (I274182,I274165,I274038);
DFFARX1 I_15989  ( .D(I274182), .CLK(I2350), .RSTB(I273871), .Q(I273848) );
nor I_15990 (I273863,I274165,I274117);
not I_15991 (I274227,I274165);
nor I_15992 (I274244,I273905,I274227);
nand I_15993 (I273833,I274165,I274004);
DFFARX1 I_15994  ( .D(I122826), .CLK(I2350), .RSTB(I273871), .Q(I274275) );
nor I_15995 (I273851,I274275,I273905);
not I_15996 (I274306,I274275);
and I_15997 (I274323,I274117,I274306);
nor I_15998 (I273857,I273922,I274323);
and I_15999 (I274354,I274275,I274244);
or I_16000 (I274371,I273922,I274354);
DFFARX1 I_16001  ( .D(I274371), .CLK(I2350), .RSTB(I273871), .Q(I273836) );
nand I_16002 (I273839,I274275,I274086);
not I_16003 (I274449,I2357);
or I_16004 (I274466,I120425,I120431);
or I_16005 (I274483,I120434,I120425);
nor I_16006 (I274500,I120449,I120437);
or I_16007 (I274438,I274500,I274466);
not I_16008 (I274531,I120449);
and I_16009 (I274548,I274531,I120428);
nor I_16010 (I274565,I274548,I120431);
not I_16011 (I274582,I274565);
nor I_16012 (I274599,I120443,I120452);
DFFARX1 I_16013  ( .D(I274599), .CLK(I2350), .RSTB(I274449), .Q(I274616) );
nor I_16014 (I274633,I274616,I274565);
nand I_16015 (I274423,I274466,I274633);
nor I_16016 (I274664,I274616,I274582);
not I_16017 (I274420,I274616);
nor I_16018 (I274695,I120443,I120434);
or I_16019 (I274432,I274466,I274695);
DFFARX1 I_16020  ( .D(I120440), .CLK(I2350), .RSTB(I274449), .Q(I274726) );
and I_16021 (I274743,I274726,I120455);
nor I_16022 (I274760,I274743,I274616);
DFFARX1 I_16023  ( .D(I274760), .CLK(I2350), .RSTB(I274449), .Q(I274426) );
nor I_16024 (I274441,I274743,I274695);
not I_16025 (I274805,I274743);
nor I_16026 (I274822,I274483,I274805);
nand I_16027 (I274411,I274743,I274582);
DFFARX1 I_16028  ( .D(I120446), .CLK(I2350), .RSTB(I274449), .Q(I274853) );
nor I_16029 (I274429,I274853,I274483);
not I_16030 (I274884,I274853);
and I_16031 (I274901,I274695,I274884);
nor I_16032 (I274435,I274500,I274901);
and I_16033 (I274932,I274853,I274822);
or I_16034 (I274949,I274500,I274932);
DFFARX1 I_16035  ( .D(I274949), .CLK(I2350), .RSTB(I274449), .Q(I274414) );
nand I_16036 (I274417,I274853,I274664);
not I_16037 (I275027,I2357);
or I_16038 (I275044,I357136,I357139);
or I_16039 (I275061,I357157,I357136);
nor I_16040 (I275078,I357151,I357160);
or I_16041 (I275016,I275078,I275044);
not I_16042 (I275109,I357151);
and I_16043 (I275126,I275109,I357163);
nor I_16044 (I275143,I275126,I357139);
not I_16045 (I275160,I275143);
nor I_16046 (I275177,I357148,I357133);
DFFARX1 I_16047  ( .D(I275177), .CLK(I2350), .RSTB(I275027), .Q(I275194) );
nor I_16048 (I275211,I275194,I275143);
nand I_16049 (I275001,I275044,I275211);
nor I_16050 (I275242,I275194,I275160);
not I_16051 (I274998,I275194);
nor I_16052 (I275273,I357148,I357157);
or I_16053 (I275010,I275044,I275273);
DFFARX1 I_16054  ( .D(I357145), .CLK(I2350), .RSTB(I275027), .Q(I275304) );
and I_16055 (I275321,I275304,I357154);
nor I_16056 (I275338,I275321,I275194);
DFFARX1 I_16057  ( .D(I275338), .CLK(I2350), .RSTB(I275027), .Q(I275004) );
nor I_16058 (I275019,I275321,I275273);
not I_16059 (I275383,I275321);
nor I_16060 (I275400,I275061,I275383);
nand I_16061 (I274989,I275321,I275160);
DFFARX1 I_16062  ( .D(I357142), .CLK(I2350), .RSTB(I275027), .Q(I275431) );
nor I_16063 (I275007,I275431,I275061);
not I_16064 (I275462,I275431);
and I_16065 (I275479,I275273,I275462);
nor I_16066 (I275013,I275078,I275479);
and I_16067 (I275510,I275431,I275400);
or I_16068 (I275527,I275078,I275510);
DFFARX1 I_16069  ( .D(I275527), .CLK(I2350), .RSTB(I275027), .Q(I274992) );
nand I_16070 (I274995,I275431,I275242);
not I_16071 (I275605,I2357);
or I_16072 (I275622,I215995,I215980);
or I_16073 (I275639,I215989,I215995);
nor I_16074 (I275656,I215983,I215971);
or I_16075 (I275594,I275656,I275622);
not I_16076 (I275687,I215983);
and I_16077 (I275704,I275687,I215992);
nor I_16078 (I275721,I275704,I215980);
not I_16079 (I275738,I275721);
nor I_16080 (I275755,I215977,I215968);
DFFARX1 I_16081  ( .D(I275755), .CLK(I2350), .RSTB(I275605), .Q(I275772) );
nor I_16082 (I275789,I275772,I275721);
nand I_16083 (I275579,I275622,I275789);
nor I_16084 (I275820,I275772,I275738);
not I_16085 (I275576,I275772);
nor I_16086 (I275851,I215977,I215989);
or I_16087 (I275588,I275622,I275851);
DFFARX1 I_16088  ( .D(I215986), .CLK(I2350), .RSTB(I275605), .Q(I275882) );
and I_16089 (I275899,I275882,I215965);
nor I_16090 (I275916,I275899,I275772);
DFFARX1 I_16091  ( .D(I275916), .CLK(I2350), .RSTB(I275605), .Q(I275582) );
nor I_16092 (I275597,I275899,I275851);
not I_16093 (I275961,I275899);
nor I_16094 (I275978,I275639,I275961);
nand I_16095 (I275567,I275899,I275738);
DFFARX1 I_16096  ( .D(I215974), .CLK(I2350), .RSTB(I275605), .Q(I276009) );
nor I_16097 (I275585,I276009,I275639);
not I_16098 (I276040,I276009);
and I_16099 (I276057,I275851,I276040);
nor I_16100 (I275591,I275656,I276057);
and I_16101 (I276088,I276009,I275978);
or I_16102 (I276105,I275656,I276088);
DFFARX1 I_16103  ( .D(I276105), .CLK(I2350), .RSTB(I275605), .Q(I275570) );
nand I_16104 (I275573,I276009,I275820);
not I_16105 (I276183,I2357);
or I_16106 (I276200,I386249,I386240);
or I_16107 (I276217,I386255,I386249);
nor I_16108 (I276234,I386246,I386243);
or I_16109 (I276172,I276234,I276200);
not I_16110 (I276265,I386246);
and I_16111 (I276282,I276265,I386237);
nor I_16112 (I276299,I276282,I386240);
not I_16113 (I276316,I276299);
nor I_16114 (I276333,I386258,I386264);
DFFARX1 I_16115  ( .D(I276333), .CLK(I2350), .RSTB(I276183), .Q(I276350) );
nor I_16116 (I276367,I276350,I276299);
nand I_16117 (I276157,I276200,I276367);
nor I_16118 (I276398,I276350,I276316);
not I_16119 (I276154,I276350);
nor I_16120 (I276429,I386258,I386255);
or I_16121 (I276166,I276200,I276429);
DFFARX1 I_16122  ( .D(I386252), .CLK(I2350), .RSTB(I276183), .Q(I276460) );
and I_16123 (I276477,I276460,I386261);
nor I_16124 (I276494,I276477,I276350);
DFFARX1 I_16125  ( .D(I276494), .CLK(I2350), .RSTB(I276183), .Q(I276160) );
nor I_16126 (I276175,I276477,I276429);
not I_16127 (I276539,I276477);
nor I_16128 (I276556,I276217,I276539);
nand I_16129 (I276145,I276477,I276316);
DFFARX1 I_16130  ( .D(I386267), .CLK(I2350), .RSTB(I276183), .Q(I276587) );
nor I_16131 (I276163,I276587,I276217);
not I_16132 (I276618,I276587);
and I_16133 (I276635,I276429,I276618);
nor I_16134 (I276169,I276234,I276635);
and I_16135 (I276666,I276587,I276556);
or I_16136 (I276683,I276234,I276666);
DFFARX1 I_16137  ( .D(I276683), .CLK(I2350), .RSTB(I276183), .Q(I276148) );
nand I_16138 (I276151,I276587,I276398);
not I_16139 (I276761,I2357);
or I_16140 (I276778,I350217,I350220);
or I_16141 (I276795,I350238,I350217);
nor I_16142 (I276812,I350232,I350241);
or I_16143 (I276750,I276812,I276778);
not I_16144 (I276843,I350232);
and I_16145 (I276860,I276843,I350244);
nor I_16146 (I276877,I276860,I350220);
not I_16147 (I276894,I276877);
nor I_16148 (I276911,I350229,I350214);
DFFARX1 I_16149  ( .D(I276911), .CLK(I2350), .RSTB(I276761), .Q(I276928) );
nor I_16150 (I276945,I276928,I276877);
nand I_16151 (I276735,I276778,I276945);
nor I_16152 (I276976,I276928,I276894);
not I_16153 (I276732,I276928);
nor I_16154 (I277007,I350229,I350238);
or I_16155 (I276744,I276778,I277007);
DFFARX1 I_16156  ( .D(I350226), .CLK(I2350), .RSTB(I276761), .Q(I277038) );
and I_16157 (I277055,I277038,I350235);
nor I_16158 (I277072,I277055,I276928);
DFFARX1 I_16159  ( .D(I277072), .CLK(I2350), .RSTB(I276761), .Q(I276738) );
nor I_16160 (I276753,I277055,I277007);
not I_16161 (I277117,I277055);
nor I_16162 (I277134,I276795,I277117);
nand I_16163 (I276723,I277055,I276894);
DFFARX1 I_16164  ( .D(I350223), .CLK(I2350), .RSTB(I276761), .Q(I277165) );
nor I_16165 (I276741,I277165,I276795);
not I_16166 (I277196,I277165);
and I_16167 (I277213,I277007,I277196);
nor I_16168 (I276747,I276812,I277213);
and I_16169 (I277244,I277165,I277134);
or I_16170 (I277261,I276812,I277244);
DFFARX1 I_16171  ( .D(I277261), .CLK(I2350), .RSTB(I276761), .Q(I276726) );
nand I_16172 (I276729,I277165,I276976);
not I_16173 (I277339,I2357);
or I_16174 (I277356,I347072,I347075);
or I_16175 (I277373,I347093,I347072);
nor I_16176 (I277390,I347087,I347096);
or I_16177 (I277328,I277390,I277356);
not I_16178 (I277421,I347087);
and I_16179 (I277438,I277421,I347099);
nor I_16180 (I277455,I277438,I347075);
not I_16181 (I277472,I277455);
nor I_16182 (I277489,I347084,I347069);
DFFARX1 I_16183  ( .D(I277489), .CLK(I2350), .RSTB(I277339), .Q(I277506) );
nor I_16184 (I277523,I277506,I277455);
nand I_16185 (I277313,I277356,I277523);
nor I_16186 (I277554,I277506,I277472);
not I_16187 (I277310,I277506);
nor I_16188 (I277585,I347084,I347093);
or I_16189 (I277322,I277356,I277585);
DFFARX1 I_16190  ( .D(I347081), .CLK(I2350), .RSTB(I277339), .Q(I277616) );
and I_16191 (I277633,I277616,I347090);
nor I_16192 (I277650,I277633,I277506);
DFFARX1 I_16193  ( .D(I277650), .CLK(I2350), .RSTB(I277339), .Q(I277316) );
nor I_16194 (I277331,I277633,I277585);
not I_16195 (I277695,I277633);
nor I_16196 (I277712,I277373,I277695);
nand I_16197 (I277301,I277633,I277472);
DFFARX1 I_16198  ( .D(I347078), .CLK(I2350), .RSTB(I277339), .Q(I277743) );
nor I_16199 (I277319,I277743,I277373);
not I_16200 (I277774,I277743);
and I_16201 (I277791,I277585,I277774);
nor I_16202 (I277325,I277390,I277791);
and I_16203 (I277822,I277743,I277712);
or I_16204 (I277839,I277390,I277822);
DFFARX1 I_16205  ( .D(I277839), .CLK(I2350), .RSTB(I277339), .Q(I277304) );
nand I_16206 (I277307,I277743,I277554);
not I_16207 (I277917,I2357);
or I_16208 (I277934,I191392,I191386);
or I_16209 (I277951,I191404,I191392);
nor I_16210 (I277968,I191383,I191410);
or I_16211 (I277906,I277968,I277934);
not I_16212 (I277999,I191383);
and I_16213 (I278016,I277999,I191407);
nor I_16214 (I278033,I278016,I191386);
not I_16215 (I278050,I278033);
nor I_16216 (I278067,I191398,I191413);
DFFARX1 I_16217  ( .D(I278067), .CLK(I2350), .RSTB(I277917), .Q(I278084) );
nor I_16218 (I278101,I278084,I278033);
nand I_16219 (I277891,I277934,I278101);
nor I_16220 (I278132,I278084,I278050);
not I_16221 (I277888,I278084);
nor I_16222 (I278163,I191398,I191404);
or I_16223 (I277900,I277934,I278163);
DFFARX1 I_16224  ( .D(I191395), .CLK(I2350), .RSTB(I277917), .Q(I278194) );
and I_16225 (I278211,I278194,I191401);
nor I_16226 (I278228,I278211,I278084);
DFFARX1 I_16227  ( .D(I278228), .CLK(I2350), .RSTB(I277917), .Q(I277894) );
nor I_16228 (I277909,I278211,I278163);
not I_16229 (I278273,I278211);
nor I_16230 (I278290,I277951,I278273);
nand I_16231 (I277879,I278211,I278050);
DFFARX1 I_16232  ( .D(I191389), .CLK(I2350), .RSTB(I277917), .Q(I278321) );
nor I_16233 (I277897,I278321,I277951);
not I_16234 (I278352,I278321);
and I_16235 (I278369,I278163,I278352);
nor I_16236 (I277903,I277968,I278369);
and I_16237 (I278400,I278321,I278290);
or I_16238 (I278417,I277968,I278400);
DFFARX1 I_16239  ( .D(I278417), .CLK(I2350), .RSTB(I277917), .Q(I277882) );
nand I_16240 (I277885,I278321,I278132);
not I_16241 (I278495,I2357);
nand I_16242 (I278512,I137698,I137704);
and I_16243 (I278529,I278512,I137686);
DFFARX1 I_16244  ( .D(I278529), .CLK(I2350), .RSTB(I278495), .Q(I278546) );
nor I_16245 (I278563,I137680,I137704);
nor I_16246 (I278580,I278563,I278546);
not I_16247 (I278478,I278563);
DFFARX1 I_16248  ( .D(I137710), .CLK(I2350), .RSTB(I278495), .Q(I278611) );
not I_16249 (I278628,I278611);
nor I_16250 (I278645,I278563,I278628);
nand I_16251 (I278481,I278611,I278580);
DFFARX1 I_16252  ( .D(I278611), .CLK(I2350), .RSTB(I278495), .Q(I278463) );
nand I_16253 (I278690,I137701,I137692);
and I_16254 (I278707,I278690,I137695);
DFFARX1 I_16255  ( .D(I278707), .CLK(I2350), .RSTB(I278495), .Q(I278724) );
nor I_16256 (I278484,I278724,I278546);
nand I_16257 (I278475,I278724,I278645);
DFFARX1 I_16258  ( .D(I137707), .CLK(I2350), .RSTB(I278495), .Q(I278769) );
and I_16259 (I278786,I278769,I137683);
DFFARX1 I_16260  ( .D(I278786), .CLK(I2350), .RSTB(I278495), .Q(I278803) );
not I_16261 (I278466,I278803);
nand I_16262 (I278834,I278786,I278724);
and I_16263 (I278851,I278546,I278834);
DFFARX1 I_16264  ( .D(I278851), .CLK(I2350), .RSTB(I278495), .Q(I278457) );
DFFARX1 I_16265  ( .D(I137689), .CLK(I2350), .RSTB(I278495), .Q(I278882) );
nand I_16266 (I278899,I278882,I278546);
and I_16267 (I278916,I278724,I278899);
DFFARX1 I_16268  ( .D(I278916), .CLK(I2350), .RSTB(I278495), .Q(I278487) );
not I_16269 (I278947,I278882);
nor I_16270 (I278964,I278563,I278947);
and I_16271 (I278981,I278882,I278964);
or I_16272 (I278998,I278786,I278981);
DFFARX1 I_16273  ( .D(I278998), .CLK(I2350), .RSTB(I278495), .Q(I278472) );
nand I_16274 (I278469,I278882,I278628);
DFFARX1 I_16275  ( .D(I278882), .CLK(I2350), .RSTB(I278495), .Q(I278460) );
not I_16276 (I279090,I2357);
nand I_16277 (I279107,I375392,I375383);
and I_16278 (I279124,I279107,I375401);
DFFARX1 I_16279  ( .D(I279124), .CLK(I2350), .RSTB(I279090), .Q(I279141) );
nor I_16280 (I279158,I375398,I375383);
nor I_16281 (I279175,I279158,I279141);
not I_16282 (I279073,I279158);
DFFARX1 I_16283  ( .D(I375380), .CLK(I2350), .RSTB(I279090), .Q(I279206) );
not I_16284 (I279223,I279206);
nor I_16285 (I279240,I279158,I279223);
nand I_16286 (I279076,I279206,I279175);
DFFARX1 I_16287  ( .D(I279206), .CLK(I2350), .RSTB(I279090), .Q(I279058) );
nand I_16288 (I279285,I375389,I375404);
and I_16289 (I279302,I279285,I375395);
DFFARX1 I_16290  ( .D(I279302), .CLK(I2350), .RSTB(I279090), .Q(I279319) );
nor I_16291 (I279079,I279319,I279141);
nand I_16292 (I279070,I279319,I279240);
DFFARX1 I_16293  ( .D(I375377), .CLK(I2350), .RSTB(I279090), .Q(I279364) );
and I_16294 (I279381,I279364,I375386);
DFFARX1 I_16295  ( .D(I279381), .CLK(I2350), .RSTB(I279090), .Q(I279398) );
not I_16296 (I279061,I279398);
nand I_16297 (I279429,I279381,I279319);
and I_16298 (I279446,I279141,I279429);
DFFARX1 I_16299  ( .D(I279446), .CLK(I2350), .RSTB(I279090), .Q(I279052) );
DFFARX1 I_16300  ( .D(I375374), .CLK(I2350), .RSTB(I279090), .Q(I279477) );
nand I_16301 (I279494,I279477,I279141);
and I_16302 (I279511,I279319,I279494);
DFFARX1 I_16303  ( .D(I279511), .CLK(I2350), .RSTB(I279090), .Q(I279082) );
not I_16304 (I279542,I279477);
nor I_16305 (I279559,I279158,I279542);
and I_16306 (I279576,I279477,I279559);
or I_16307 (I279593,I279381,I279576);
DFFARX1 I_16308  ( .D(I279593), .CLK(I2350), .RSTB(I279090), .Q(I279067) );
nand I_16309 (I279064,I279477,I279223);
DFFARX1 I_16310  ( .D(I279477), .CLK(I2350), .RSTB(I279090), .Q(I279055) );
not I_16311 (I279685,I2357);
nand I_16312 (I279702,I176815,I176821);
and I_16313 (I279719,I279702,I176803);
DFFARX1 I_16314  ( .D(I279719), .CLK(I2350), .RSTB(I279685), .Q(I279736) );
nor I_16315 (I279753,I176797,I176821);
nor I_16316 (I279770,I279753,I279736);
not I_16317 (I279668,I279753);
DFFARX1 I_16318  ( .D(I176827), .CLK(I2350), .RSTB(I279685), .Q(I279801) );
not I_16319 (I279818,I279801);
nor I_16320 (I279835,I279753,I279818);
nand I_16321 (I279671,I279801,I279770);
DFFARX1 I_16322  ( .D(I279801), .CLK(I2350), .RSTB(I279685), .Q(I279653) );
nand I_16323 (I279880,I176818,I176809);
and I_16324 (I279897,I279880,I176812);
DFFARX1 I_16325  ( .D(I279897), .CLK(I2350), .RSTB(I279685), .Q(I279914) );
nor I_16326 (I279674,I279914,I279736);
nand I_16327 (I279665,I279914,I279835);
DFFARX1 I_16328  ( .D(I176824), .CLK(I2350), .RSTB(I279685), .Q(I279959) );
and I_16329 (I279976,I279959,I176800);
DFFARX1 I_16330  ( .D(I279976), .CLK(I2350), .RSTB(I279685), .Q(I279993) );
not I_16331 (I279656,I279993);
nand I_16332 (I280024,I279976,I279914);
and I_16333 (I280041,I279736,I280024);
DFFARX1 I_16334  ( .D(I280041), .CLK(I2350), .RSTB(I279685), .Q(I279647) );
DFFARX1 I_16335  ( .D(I176806), .CLK(I2350), .RSTB(I279685), .Q(I280072) );
nand I_16336 (I280089,I280072,I279736);
and I_16337 (I280106,I279914,I280089);
DFFARX1 I_16338  ( .D(I280106), .CLK(I2350), .RSTB(I279685), .Q(I279677) );
not I_16339 (I280137,I280072);
nor I_16340 (I280154,I279753,I280137);
and I_16341 (I280171,I280072,I280154);
or I_16342 (I280188,I279976,I280171);
DFFARX1 I_16343  ( .D(I280188), .CLK(I2350), .RSTB(I279685), .Q(I279662) );
nand I_16344 (I279659,I280072,I279818);
DFFARX1 I_16345  ( .D(I280072), .CLK(I2350), .RSTB(I279685), .Q(I279650) );
not I_16346 (I280280,I2357);
nand I_16347 (I280297,I101964,I101976);
and I_16348 (I280314,I280297,I101955);
DFFARX1 I_16349  ( .D(I280314), .CLK(I2350), .RSTB(I280280), .Q(I280331) );
nor I_16350 (I280348,I101946,I101976);
nor I_16351 (I280365,I280348,I280331);
not I_16352 (I280263,I280348);
DFFARX1 I_16353  ( .D(I101958), .CLK(I2350), .RSTB(I280280), .Q(I280396) );
not I_16354 (I280413,I280396);
nor I_16355 (I280430,I280348,I280413);
nand I_16356 (I280266,I280396,I280365);
DFFARX1 I_16357  ( .D(I280396), .CLK(I2350), .RSTB(I280280), .Q(I280248) );
nand I_16358 (I280475,I101973,I101961);
and I_16359 (I280492,I280475,I101949);
DFFARX1 I_16360  ( .D(I280492), .CLK(I2350), .RSTB(I280280), .Q(I280509) );
nor I_16361 (I280269,I280509,I280331);
nand I_16362 (I280260,I280509,I280430);
DFFARX1 I_16363  ( .D(I101967), .CLK(I2350), .RSTB(I280280), .Q(I280554) );
and I_16364 (I280571,I280554,I101952);
DFFARX1 I_16365  ( .D(I280571), .CLK(I2350), .RSTB(I280280), .Q(I280588) );
not I_16366 (I280251,I280588);
nand I_16367 (I280619,I280571,I280509);
and I_16368 (I280636,I280331,I280619);
DFFARX1 I_16369  ( .D(I280636), .CLK(I2350), .RSTB(I280280), .Q(I280242) );
DFFARX1 I_16370  ( .D(I101970), .CLK(I2350), .RSTB(I280280), .Q(I280667) );
nand I_16371 (I280684,I280667,I280331);
and I_16372 (I280701,I280509,I280684);
DFFARX1 I_16373  ( .D(I280701), .CLK(I2350), .RSTB(I280280), .Q(I280272) );
not I_16374 (I280732,I280667);
nor I_16375 (I280749,I280348,I280732);
and I_16376 (I280766,I280667,I280749);
or I_16377 (I280783,I280571,I280766);
DFFARX1 I_16378  ( .D(I280783), .CLK(I2350), .RSTB(I280280), .Q(I280257) );
nand I_16379 (I280254,I280667,I280413);
DFFARX1 I_16380  ( .D(I280667), .CLK(I2350), .RSTB(I280280), .Q(I280245) );
not I_16381 (I280875,I2357);
nand I_16382 (I280892,I225673,I225685);
and I_16383 (I280909,I280892,I225667);
DFFARX1 I_16384  ( .D(I280909), .CLK(I2350), .RSTB(I280875), .Q(I280926) );
nor I_16385 (I280943,I225679,I225685);
nor I_16386 (I280960,I280943,I280926);
not I_16387 (I280858,I280943);
DFFARX1 I_16388  ( .D(I225664), .CLK(I2350), .RSTB(I280875), .Q(I280991) );
not I_16389 (I281008,I280991);
nor I_16390 (I281025,I280943,I281008);
nand I_16391 (I280861,I280991,I280960);
DFFARX1 I_16392  ( .D(I280991), .CLK(I2350), .RSTB(I280875), .Q(I280843) );
nand I_16393 (I281070,I225655,I225670);
and I_16394 (I281087,I281070,I225661);
DFFARX1 I_16395  ( .D(I281087), .CLK(I2350), .RSTB(I280875), .Q(I281104) );
nor I_16396 (I280864,I281104,I280926);
nand I_16397 (I280855,I281104,I281025);
DFFARX1 I_16398  ( .D(I225682), .CLK(I2350), .RSTB(I280875), .Q(I281149) );
and I_16399 (I281166,I281149,I225676);
DFFARX1 I_16400  ( .D(I281166), .CLK(I2350), .RSTB(I280875), .Q(I281183) );
not I_16401 (I280846,I281183);
nand I_16402 (I281214,I281166,I281104);
and I_16403 (I281231,I280926,I281214);
DFFARX1 I_16404  ( .D(I281231), .CLK(I2350), .RSTB(I280875), .Q(I280837) );
DFFARX1 I_16405  ( .D(I225658), .CLK(I2350), .RSTB(I280875), .Q(I281262) );
nand I_16406 (I281279,I281262,I280926);
and I_16407 (I281296,I281104,I281279);
DFFARX1 I_16408  ( .D(I281296), .CLK(I2350), .RSTB(I280875), .Q(I280867) );
not I_16409 (I281327,I281262);
nor I_16410 (I281344,I280943,I281327);
and I_16411 (I281361,I281262,I281344);
or I_16412 (I281378,I281166,I281361);
DFFARX1 I_16413  ( .D(I281378), .CLK(I2350), .RSTB(I280875), .Q(I280852) );
nand I_16414 (I280849,I281262,I281008);
DFFARX1 I_16415  ( .D(I281262), .CLK(I2350), .RSTB(I280875), .Q(I280840) );
not I_16416 (I281470,I2357);
nand I_16417 (I281487,I110583,I110595);
and I_16418 (I281504,I281487,I110574);
DFFARX1 I_16419  ( .D(I281504), .CLK(I2350), .RSTB(I281470), .Q(I281521) );
nor I_16420 (I281538,I110565,I110595);
nor I_16421 (I281555,I281538,I281521);
not I_16422 (I281453,I281538);
DFFARX1 I_16423  ( .D(I110577), .CLK(I2350), .RSTB(I281470), .Q(I281586) );
not I_16424 (I281603,I281586);
nor I_16425 (I281620,I281538,I281603);
nand I_16426 (I281456,I281586,I281555);
DFFARX1 I_16427  ( .D(I281586), .CLK(I2350), .RSTB(I281470), .Q(I281438) );
nand I_16428 (I281665,I110592,I110580);
and I_16429 (I281682,I281665,I110568);
DFFARX1 I_16430  ( .D(I281682), .CLK(I2350), .RSTB(I281470), .Q(I281699) );
nor I_16431 (I281459,I281699,I281521);
nand I_16432 (I281450,I281699,I281620);
DFFARX1 I_16433  ( .D(I110586), .CLK(I2350), .RSTB(I281470), .Q(I281744) );
and I_16434 (I281761,I281744,I110571);
DFFARX1 I_16435  ( .D(I281761), .CLK(I2350), .RSTB(I281470), .Q(I281778) );
not I_16436 (I281441,I281778);
nand I_16437 (I281809,I281761,I281699);
and I_16438 (I281826,I281521,I281809);
DFFARX1 I_16439  ( .D(I281826), .CLK(I2350), .RSTB(I281470), .Q(I281432) );
DFFARX1 I_16440  ( .D(I110589), .CLK(I2350), .RSTB(I281470), .Q(I281857) );
nand I_16441 (I281874,I281857,I281521);
and I_16442 (I281891,I281699,I281874);
DFFARX1 I_16443  ( .D(I281891), .CLK(I2350), .RSTB(I281470), .Q(I281462) );
not I_16444 (I281922,I281857);
nor I_16445 (I281939,I281538,I281922);
and I_16446 (I281956,I281857,I281939);
or I_16447 (I281973,I281761,I281956);
DFFARX1 I_16448  ( .D(I281973), .CLK(I2350), .RSTB(I281470), .Q(I281447) );
nand I_16449 (I281444,I281857,I281603);
DFFARX1 I_16450  ( .D(I281857), .CLK(I2350), .RSTB(I281470), .Q(I281435) );
not I_16451 (I282065,I2357);
nand I_16452 (I282082,I219859,I219871);
and I_16453 (I282099,I282082,I219853);
DFFARX1 I_16454  ( .D(I282099), .CLK(I2350), .RSTB(I282065), .Q(I282116) );
nor I_16455 (I282133,I219865,I219871);
nor I_16456 (I282150,I282133,I282116);
not I_16457 (I282048,I282133);
DFFARX1 I_16458  ( .D(I219850), .CLK(I2350), .RSTB(I282065), .Q(I282181) );
not I_16459 (I282198,I282181);
nor I_16460 (I282215,I282133,I282198);
nand I_16461 (I282051,I282181,I282150);
DFFARX1 I_16462  ( .D(I282181), .CLK(I2350), .RSTB(I282065), .Q(I282033) );
nand I_16463 (I282260,I219841,I219856);
and I_16464 (I282277,I282260,I219847);
DFFARX1 I_16465  ( .D(I282277), .CLK(I2350), .RSTB(I282065), .Q(I282294) );
nor I_16466 (I282054,I282294,I282116);
nand I_16467 (I282045,I282294,I282215);
DFFARX1 I_16468  ( .D(I219868), .CLK(I2350), .RSTB(I282065), .Q(I282339) );
and I_16469 (I282356,I282339,I219862);
DFFARX1 I_16470  ( .D(I282356), .CLK(I2350), .RSTB(I282065), .Q(I282373) );
not I_16471 (I282036,I282373);
nand I_16472 (I282404,I282356,I282294);
and I_16473 (I282421,I282116,I282404);
DFFARX1 I_16474  ( .D(I282421), .CLK(I2350), .RSTB(I282065), .Q(I282027) );
DFFARX1 I_16475  ( .D(I219844), .CLK(I2350), .RSTB(I282065), .Q(I282452) );
nand I_16476 (I282469,I282452,I282116);
and I_16477 (I282486,I282294,I282469);
DFFARX1 I_16478  ( .D(I282486), .CLK(I2350), .RSTB(I282065), .Q(I282057) );
not I_16479 (I282517,I282452);
nor I_16480 (I282534,I282133,I282517);
and I_16481 (I282551,I282452,I282534);
or I_16482 (I282568,I282356,I282551);
DFFARX1 I_16483  ( .D(I282568), .CLK(I2350), .RSTB(I282065), .Q(I282042) );
nand I_16484 (I282039,I282452,I282198);
DFFARX1 I_16485  ( .D(I282452), .CLK(I2350), .RSTB(I282065), .Q(I282030) );
not I_16486 (I282660,I2357);
nand I_16487 (I282677,I24803,I24809);
and I_16488 (I282694,I282677,I24806);
DFFARX1 I_16489  ( .D(I282694), .CLK(I2350), .RSTB(I282660), .Q(I282711) );
nor I_16490 (I282728,I24830,I24809);
nor I_16491 (I282745,I282728,I282711);
not I_16492 (I282643,I282728);
DFFARX1 I_16493  ( .D(I24821), .CLK(I2350), .RSTB(I282660), .Q(I282776) );
not I_16494 (I282793,I282776);
nor I_16495 (I282810,I282728,I282793);
nand I_16496 (I282646,I282776,I282745);
DFFARX1 I_16497  ( .D(I282776), .CLK(I2350), .RSTB(I282660), .Q(I282628) );
nand I_16498 (I282855,I24824,I24827);
and I_16499 (I282872,I282855,I24800);
DFFARX1 I_16500  ( .D(I282872), .CLK(I2350), .RSTB(I282660), .Q(I282889) );
nor I_16501 (I282649,I282889,I282711);
nand I_16502 (I282640,I282889,I282810);
DFFARX1 I_16503  ( .D(I24818), .CLK(I2350), .RSTB(I282660), .Q(I282934) );
and I_16504 (I282951,I282934,I24812);
DFFARX1 I_16505  ( .D(I282951), .CLK(I2350), .RSTB(I282660), .Q(I282968) );
not I_16506 (I282631,I282968);
nand I_16507 (I282999,I282951,I282889);
and I_16508 (I283016,I282711,I282999);
DFFARX1 I_16509  ( .D(I283016), .CLK(I2350), .RSTB(I282660), .Q(I282622) );
DFFARX1 I_16510  ( .D(I24815), .CLK(I2350), .RSTB(I282660), .Q(I283047) );
nand I_16511 (I283064,I283047,I282711);
and I_16512 (I283081,I282889,I283064);
DFFARX1 I_16513  ( .D(I283081), .CLK(I2350), .RSTB(I282660), .Q(I282652) );
not I_16514 (I283112,I283047);
nor I_16515 (I283129,I282728,I283112);
and I_16516 (I283146,I283047,I283129);
or I_16517 (I283163,I282951,I283146);
DFFARX1 I_16518  ( .D(I283163), .CLK(I2350), .RSTB(I282660), .Q(I282637) );
nand I_16519 (I282634,I283047,I282793);
DFFARX1 I_16520  ( .D(I283047), .CLK(I2350), .RSTB(I282660), .Q(I282625) );
not I_16521 (I283255,I2357);
nand I_16522 (I283272,I269100,I269073);
and I_16523 (I283289,I283272,I269076);
DFFARX1 I_16524  ( .D(I283289), .CLK(I2350), .RSTB(I283255), .Q(I283306) );
nor I_16525 (I283323,I269085,I269073);
nor I_16526 (I283340,I283323,I283306);
not I_16527 (I283238,I283323);
DFFARX1 I_16528  ( .D(I269082), .CLK(I2350), .RSTB(I283255), .Q(I283371) );
not I_16529 (I283388,I283371);
nor I_16530 (I283405,I283323,I283388);
nand I_16531 (I283241,I283371,I283340);
DFFARX1 I_16532  ( .D(I283371), .CLK(I2350), .RSTB(I283255), .Q(I283223) );
nand I_16533 (I283450,I269079,I269088);
and I_16534 (I283467,I283450,I269097);
DFFARX1 I_16535  ( .D(I283467), .CLK(I2350), .RSTB(I283255), .Q(I283484) );
nor I_16536 (I283244,I283484,I283306);
nand I_16537 (I283235,I283484,I283405);
DFFARX1 I_16538  ( .D(I269103), .CLK(I2350), .RSTB(I283255), .Q(I283529) );
and I_16539 (I283546,I283529,I269094);
DFFARX1 I_16540  ( .D(I283546), .CLK(I2350), .RSTB(I283255), .Q(I283563) );
not I_16541 (I283226,I283563);
nand I_16542 (I283594,I283546,I283484);
and I_16543 (I283611,I283306,I283594);
DFFARX1 I_16544  ( .D(I283611), .CLK(I2350), .RSTB(I283255), .Q(I283217) );
DFFARX1 I_16545  ( .D(I269091), .CLK(I2350), .RSTB(I283255), .Q(I283642) );
nand I_16546 (I283659,I283642,I283306);
and I_16547 (I283676,I283484,I283659);
DFFARX1 I_16548  ( .D(I283676), .CLK(I2350), .RSTB(I283255), .Q(I283247) );
not I_16549 (I283707,I283642);
nor I_16550 (I283724,I283323,I283707);
and I_16551 (I283741,I283642,I283724);
or I_16552 (I283758,I283546,I283741);
DFFARX1 I_16553  ( .D(I283758), .CLK(I2350), .RSTB(I283255), .Q(I283232) );
nand I_16554 (I283229,I283642,I283388);
DFFARX1 I_16555  ( .D(I283642), .CLK(I2350), .RSTB(I283255), .Q(I283220) );
not I_16556 (I283850,I2357);
nand I_16557 (I283867,I394341,I394347);
and I_16558 (I283884,I283867,I394338);
DFFARX1 I_16559  ( .D(I283884), .CLK(I2350), .RSTB(I283850), .Q(I283901) );
nor I_16560 (I283918,I394350,I394347);
nor I_16561 (I283935,I283918,I283901);
not I_16562 (I283833,I283918);
DFFARX1 I_16563  ( .D(I394329), .CLK(I2350), .RSTB(I283850), .Q(I283966) );
not I_16564 (I283983,I283966);
nor I_16565 (I284000,I283918,I283983);
nand I_16566 (I283836,I283966,I283935);
DFFARX1 I_16567  ( .D(I283966), .CLK(I2350), .RSTB(I283850), .Q(I283818) );
nand I_16568 (I284045,I394353,I394335);
and I_16569 (I284062,I284045,I394344);
DFFARX1 I_16570  ( .D(I284062), .CLK(I2350), .RSTB(I283850), .Q(I284079) );
nor I_16571 (I283839,I284079,I283901);
nand I_16572 (I283830,I284079,I284000);
DFFARX1 I_16573  ( .D(I394359), .CLK(I2350), .RSTB(I283850), .Q(I284124) );
and I_16574 (I284141,I284124,I394332);
DFFARX1 I_16575  ( .D(I284141), .CLK(I2350), .RSTB(I283850), .Q(I284158) );
not I_16576 (I283821,I284158);
nand I_16577 (I284189,I284141,I284079);
and I_16578 (I284206,I283901,I284189);
DFFARX1 I_16579  ( .D(I284206), .CLK(I2350), .RSTB(I283850), .Q(I283812) );
DFFARX1 I_16580  ( .D(I394356), .CLK(I2350), .RSTB(I283850), .Q(I284237) );
nand I_16581 (I284254,I284237,I283901);
and I_16582 (I284271,I284079,I284254);
DFFARX1 I_16583  ( .D(I284271), .CLK(I2350), .RSTB(I283850), .Q(I283842) );
not I_16584 (I284302,I284237);
nor I_16585 (I284319,I283918,I284302);
and I_16586 (I284336,I284237,I284319);
or I_16587 (I284353,I284141,I284336);
DFFARX1 I_16588  ( .D(I284353), .CLK(I2350), .RSTB(I283850), .Q(I283827) );
nand I_16589 (I283824,I284237,I283983);
DFFARX1 I_16590  ( .D(I284237), .CLK(I2350), .RSTB(I283850), .Q(I283815) );
not I_16591 (I284445,I2357);
nand I_16592 (I284462,I44019,I44031);
and I_16593 (I284479,I284462,I44040);
DFFARX1 I_16594  ( .D(I284479), .CLK(I2350), .RSTB(I284445), .Q(I284496) );
nor I_16595 (I284513,I44034,I44031);
nor I_16596 (I284530,I284513,I284496);
not I_16597 (I284428,I284513);
DFFARX1 I_16598  ( .D(I44028), .CLK(I2350), .RSTB(I284445), .Q(I284561) );
not I_16599 (I284578,I284561);
nor I_16600 (I284595,I284513,I284578);
nand I_16601 (I284431,I284561,I284530);
DFFARX1 I_16602  ( .D(I284561), .CLK(I2350), .RSTB(I284445), .Q(I284413) );
nand I_16603 (I284640,I44025,I44022);
and I_16604 (I284657,I284640,I44013);
DFFARX1 I_16605  ( .D(I284657), .CLK(I2350), .RSTB(I284445), .Q(I284674) );
nor I_16606 (I284434,I284674,I284496);
nand I_16607 (I284425,I284674,I284595);
DFFARX1 I_16608  ( .D(I44037), .CLK(I2350), .RSTB(I284445), .Q(I284719) );
and I_16609 (I284736,I284719,I44016);
DFFARX1 I_16610  ( .D(I284736), .CLK(I2350), .RSTB(I284445), .Q(I284753) );
not I_16611 (I284416,I284753);
nand I_16612 (I284784,I284736,I284674);
and I_16613 (I284801,I284496,I284784);
DFFARX1 I_16614  ( .D(I284801), .CLK(I2350), .RSTB(I284445), .Q(I284407) );
DFFARX1 I_16615  ( .D(I44010), .CLK(I2350), .RSTB(I284445), .Q(I284832) );
nand I_16616 (I284849,I284832,I284496);
and I_16617 (I284866,I284674,I284849);
DFFARX1 I_16618  ( .D(I284866), .CLK(I2350), .RSTB(I284445), .Q(I284437) );
not I_16619 (I284897,I284832);
nor I_16620 (I284914,I284513,I284897);
and I_16621 (I284931,I284832,I284914);
or I_16622 (I284948,I284736,I284931);
DFFARX1 I_16623  ( .D(I284948), .CLK(I2350), .RSTB(I284445), .Q(I284422) );
nand I_16624 (I284419,I284832,I284578);
DFFARX1 I_16625  ( .D(I284832), .CLK(I2350), .RSTB(I284445), .Q(I284410) );
not I_16626 (I285040,I2357);
nand I_16627 (I285057,I276175,I276163);
and I_16628 (I285074,I285057,I276160);
DFFARX1 I_16629  ( .D(I285074), .CLK(I2350), .RSTB(I285040), .Q(I285091) );
nor I_16630 (I285108,I276154,I276163);
nor I_16631 (I285125,I285108,I285091);
not I_16632 (I285023,I285108);
DFFARX1 I_16633  ( .D(I276169), .CLK(I2350), .RSTB(I285040), .Q(I285156) );
not I_16634 (I285173,I285156);
nor I_16635 (I285190,I285108,I285173);
nand I_16636 (I285026,I285156,I285125);
DFFARX1 I_16637  ( .D(I285156), .CLK(I2350), .RSTB(I285040), .Q(I285008) );
nand I_16638 (I285235,I276166,I276172);
and I_16639 (I285252,I285235,I276157);
DFFARX1 I_16640  ( .D(I285252), .CLK(I2350), .RSTB(I285040), .Q(I285269) );
nor I_16641 (I285029,I285269,I285091);
nand I_16642 (I285020,I285269,I285190);
DFFARX1 I_16643  ( .D(I276145), .CLK(I2350), .RSTB(I285040), .Q(I285314) );
and I_16644 (I285331,I285314,I276148);
DFFARX1 I_16645  ( .D(I285331), .CLK(I2350), .RSTB(I285040), .Q(I285348) );
not I_16646 (I285011,I285348);
nand I_16647 (I285379,I285331,I285269);
and I_16648 (I285396,I285091,I285379);
DFFARX1 I_16649  ( .D(I285396), .CLK(I2350), .RSTB(I285040), .Q(I285002) );
DFFARX1 I_16650  ( .D(I276151), .CLK(I2350), .RSTB(I285040), .Q(I285427) );
nand I_16651 (I285444,I285427,I285091);
and I_16652 (I285461,I285269,I285444);
DFFARX1 I_16653  ( .D(I285461), .CLK(I2350), .RSTB(I285040), .Q(I285032) );
not I_16654 (I285492,I285427);
nor I_16655 (I285509,I285108,I285492);
and I_16656 (I285526,I285427,I285509);
or I_16657 (I285543,I285331,I285526);
DFFARX1 I_16658  ( .D(I285543), .CLK(I2350), .RSTB(I285040), .Q(I285017) );
nand I_16659 (I285014,I285427,I285173);
DFFARX1 I_16660  ( .D(I285427), .CLK(I2350), .RSTB(I285040), .Q(I285005) );
not I_16661 (I285635,I2357);
nand I_16662 (I285652,I55001,I55013);
and I_16663 (I285669,I285652,I55022);
DFFARX1 I_16664  ( .D(I285669), .CLK(I2350), .RSTB(I285635), .Q(I285686) );
nor I_16665 (I285703,I55016,I55013);
nor I_16666 (I285720,I285703,I285686);
not I_16667 (I285618,I285703);
DFFARX1 I_16668  ( .D(I55010), .CLK(I2350), .RSTB(I285635), .Q(I285751) );
not I_16669 (I285768,I285751);
nor I_16670 (I285785,I285703,I285768);
nand I_16671 (I285621,I285751,I285720);
DFFARX1 I_16672  ( .D(I285751), .CLK(I2350), .RSTB(I285635), .Q(I285603) );
nand I_16673 (I285830,I55007,I55004);
and I_16674 (I285847,I285830,I54995);
DFFARX1 I_16675  ( .D(I285847), .CLK(I2350), .RSTB(I285635), .Q(I285864) );
nor I_16676 (I285624,I285864,I285686);
nand I_16677 (I285615,I285864,I285785);
DFFARX1 I_16678  ( .D(I55019), .CLK(I2350), .RSTB(I285635), .Q(I285909) );
and I_16679 (I285926,I285909,I54998);
DFFARX1 I_16680  ( .D(I285926), .CLK(I2350), .RSTB(I285635), .Q(I285943) );
not I_16681 (I285606,I285943);
nand I_16682 (I285974,I285926,I285864);
and I_16683 (I285991,I285686,I285974);
DFFARX1 I_16684  ( .D(I285991), .CLK(I2350), .RSTB(I285635), .Q(I285597) );
DFFARX1 I_16685  ( .D(I54992), .CLK(I2350), .RSTB(I285635), .Q(I286022) );
nand I_16686 (I286039,I286022,I285686);
and I_16687 (I286056,I285864,I286039);
DFFARX1 I_16688  ( .D(I286056), .CLK(I2350), .RSTB(I285635), .Q(I285627) );
not I_16689 (I286087,I286022);
nor I_16690 (I286104,I285703,I286087);
and I_16691 (I286121,I286022,I286104);
or I_16692 (I286138,I285926,I286121);
DFFARX1 I_16693  ( .D(I286138), .CLK(I2350), .RSTB(I285635), .Q(I285612) );
nand I_16694 (I285609,I286022,I285768);
DFFARX1 I_16695  ( .D(I286022), .CLK(I2350), .RSTB(I285635), .Q(I285600) );
not I_16696 (I286230,I2357);
nand I_16697 (I286247,I63399,I63411);
and I_16698 (I286264,I286247,I63420);
DFFARX1 I_16699  ( .D(I286264), .CLK(I2350), .RSTB(I286230), .Q(I286281) );
nor I_16700 (I286298,I63414,I63411);
nor I_16701 (I286315,I286298,I286281);
not I_16702 (I286213,I286298);
DFFARX1 I_16703  ( .D(I63408), .CLK(I2350), .RSTB(I286230), .Q(I286346) );
not I_16704 (I286363,I286346);
nor I_16705 (I286380,I286298,I286363);
nand I_16706 (I286216,I286346,I286315);
DFFARX1 I_16707  ( .D(I286346), .CLK(I2350), .RSTB(I286230), .Q(I286198) );
nand I_16708 (I286425,I63405,I63402);
and I_16709 (I286442,I286425,I63393);
DFFARX1 I_16710  ( .D(I286442), .CLK(I2350), .RSTB(I286230), .Q(I286459) );
nor I_16711 (I286219,I286459,I286281);
nand I_16712 (I286210,I286459,I286380);
DFFARX1 I_16713  ( .D(I63417), .CLK(I2350), .RSTB(I286230), .Q(I286504) );
and I_16714 (I286521,I286504,I63396);
DFFARX1 I_16715  ( .D(I286521), .CLK(I2350), .RSTB(I286230), .Q(I286538) );
not I_16716 (I286201,I286538);
nand I_16717 (I286569,I286521,I286459);
and I_16718 (I286586,I286281,I286569);
DFFARX1 I_16719  ( .D(I286586), .CLK(I2350), .RSTB(I286230), .Q(I286192) );
DFFARX1 I_16720  ( .D(I63390), .CLK(I2350), .RSTB(I286230), .Q(I286617) );
nand I_16721 (I286634,I286617,I286281);
and I_16722 (I286651,I286459,I286634);
DFFARX1 I_16723  ( .D(I286651), .CLK(I2350), .RSTB(I286230), .Q(I286222) );
not I_16724 (I286682,I286617);
nor I_16725 (I286699,I286298,I286682);
and I_16726 (I286716,I286617,I286699);
or I_16727 (I286733,I286521,I286716);
DFFARX1 I_16728  ( .D(I286733), .CLK(I2350), .RSTB(I286230), .Q(I286207) );
nand I_16729 (I286204,I286617,I286363);
DFFARX1 I_16730  ( .D(I286617), .CLK(I2350), .RSTB(I286230), .Q(I286195) );
not I_16731 (I286825,I2357);
nand I_16732 (I286842,I160903,I160909);
and I_16733 (I286859,I286842,I160891);
DFFARX1 I_16734  ( .D(I286859), .CLK(I2350), .RSTB(I286825), .Q(I286876) );
nor I_16735 (I286893,I160885,I160909);
nor I_16736 (I286910,I286893,I286876);
not I_16737 (I286808,I286893);
DFFARX1 I_16738  ( .D(I160915), .CLK(I2350), .RSTB(I286825), .Q(I286941) );
not I_16739 (I286958,I286941);
nor I_16740 (I286975,I286893,I286958);
nand I_16741 (I286811,I286941,I286910);
DFFARX1 I_16742  ( .D(I286941), .CLK(I2350), .RSTB(I286825), .Q(I286793) );
nand I_16743 (I287020,I160906,I160897);
and I_16744 (I287037,I287020,I160900);
DFFARX1 I_16745  ( .D(I287037), .CLK(I2350), .RSTB(I286825), .Q(I287054) );
nor I_16746 (I286814,I287054,I286876);
nand I_16747 (I286805,I287054,I286975);
DFFARX1 I_16748  ( .D(I160912), .CLK(I2350), .RSTB(I286825), .Q(I287099) );
and I_16749 (I287116,I287099,I160888);
DFFARX1 I_16750  ( .D(I287116), .CLK(I2350), .RSTB(I286825), .Q(I287133) );
not I_16751 (I286796,I287133);
nand I_16752 (I287164,I287116,I287054);
and I_16753 (I287181,I286876,I287164);
DFFARX1 I_16754  ( .D(I287181), .CLK(I2350), .RSTB(I286825), .Q(I286787) );
DFFARX1 I_16755  ( .D(I160894), .CLK(I2350), .RSTB(I286825), .Q(I287212) );
nand I_16756 (I287229,I287212,I286876);
and I_16757 (I287246,I287054,I287229);
DFFARX1 I_16758  ( .D(I287246), .CLK(I2350), .RSTB(I286825), .Q(I286817) );
not I_16759 (I287277,I287212);
nor I_16760 (I287294,I286893,I287277);
and I_16761 (I287311,I287212,I287294);
or I_16762 (I287328,I287116,I287311);
DFFARX1 I_16763  ( .D(I287328), .CLK(I2350), .RSTB(I286825), .Q(I286802) );
nand I_16764 (I286799,I287212,I286958);
DFFARX1 I_16765  ( .D(I287212), .CLK(I2350), .RSTB(I286825), .Q(I286790) );
not I_16766 (I287420,I2357);
nand I_16767 (I287437,I341426,I341417);
and I_16768 (I287454,I287437,I341435);
DFFARX1 I_16769  ( .D(I287454), .CLK(I2350), .RSTB(I287420), .Q(I287471) );
nor I_16770 (I287488,I341432,I341417);
nor I_16771 (I287505,I287488,I287471);
not I_16772 (I287403,I287488);
DFFARX1 I_16773  ( .D(I341414), .CLK(I2350), .RSTB(I287420), .Q(I287536) );
not I_16774 (I287553,I287536);
nor I_16775 (I287570,I287488,I287553);
nand I_16776 (I287406,I287536,I287505);
DFFARX1 I_16777  ( .D(I287536), .CLK(I2350), .RSTB(I287420), .Q(I287388) );
nand I_16778 (I287615,I341423,I341438);
and I_16779 (I287632,I287615,I341429);
DFFARX1 I_16780  ( .D(I287632), .CLK(I2350), .RSTB(I287420), .Q(I287649) );
nor I_16781 (I287409,I287649,I287471);
nand I_16782 (I287400,I287649,I287570);
DFFARX1 I_16783  ( .D(I341411), .CLK(I2350), .RSTB(I287420), .Q(I287694) );
and I_16784 (I287711,I287694,I341420);
DFFARX1 I_16785  ( .D(I287711), .CLK(I2350), .RSTB(I287420), .Q(I287728) );
not I_16786 (I287391,I287728);
nand I_16787 (I287759,I287711,I287649);
and I_16788 (I287776,I287471,I287759);
DFFARX1 I_16789  ( .D(I287776), .CLK(I2350), .RSTB(I287420), .Q(I287382) );
DFFARX1 I_16790  ( .D(I341408), .CLK(I2350), .RSTB(I287420), .Q(I287807) );
nand I_16791 (I287824,I287807,I287471);
and I_16792 (I287841,I287649,I287824);
DFFARX1 I_16793  ( .D(I287841), .CLK(I2350), .RSTB(I287420), .Q(I287412) );
not I_16794 (I287872,I287807);
nor I_16795 (I287889,I287488,I287872);
and I_16796 (I287906,I287807,I287889);
or I_16797 (I287923,I287711,I287906);
DFFARX1 I_16798  ( .D(I287923), .CLK(I2350), .RSTB(I287420), .Q(I287397) );
nand I_16799 (I287394,I287807,I287553);
DFFARX1 I_16800  ( .D(I287807), .CLK(I2350), .RSTB(I287420), .Q(I287385) );
not I_16801 (I288015,I2357);
nand I_16802 (I288032,I259716,I259719);
and I_16803 (I288049,I288032,I259713);
DFFARX1 I_16804  ( .D(I288049), .CLK(I2350), .RSTB(I288015), .Q(I288066) );
nor I_16805 (I288083,I259710,I259719);
nor I_16806 (I288100,I288083,I288066);
not I_16807 (I287998,I288083);
DFFARX1 I_16808  ( .D(I259692), .CLK(I2350), .RSTB(I288015), .Q(I288131) );
not I_16809 (I288148,I288131);
nor I_16810 (I288165,I288083,I288148);
nand I_16811 (I288001,I288131,I288100);
DFFARX1 I_16812  ( .D(I288131), .CLK(I2350), .RSTB(I288015), .Q(I287983) );
nand I_16813 (I288210,I259701,I259698);
and I_16814 (I288227,I288210,I259707);
DFFARX1 I_16815  ( .D(I288227), .CLK(I2350), .RSTB(I288015), .Q(I288244) );
nor I_16816 (I288004,I288244,I288066);
nand I_16817 (I287995,I288244,I288165);
DFFARX1 I_16818  ( .D(I259689), .CLK(I2350), .RSTB(I288015), .Q(I288289) );
and I_16819 (I288306,I288289,I259704);
DFFARX1 I_16820  ( .D(I288306), .CLK(I2350), .RSTB(I288015), .Q(I288323) );
not I_16821 (I287986,I288323);
nand I_16822 (I288354,I288306,I288244);
and I_16823 (I288371,I288066,I288354);
DFFARX1 I_16824  ( .D(I288371), .CLK(I2350), .RSTB(I288015), .Q(I287977) );
DFFARX1 I_16825  ( .D(I259695), .CLK(I2350), .RSTB(I288015), .Q(I288402) );
nand I_16826 (I288419,I288402,I288066);
and I_16827 (I288436,I288244,I288419);
DFFARX1 I_16828  ( .D(I288436), .CLK(I2350), .RSTB(I288015), .Q(I288007) );
not I_16829 (I288467,I288402);
nor I_16830 (I288484,I288083,I288467);
and I_16831 (I288501,I288402,I288484);
or I_16832 (I288518,I288306,I288501);
DFFARX1 I_16833  ( .D(I288518), .CLK(I2350), .RSTB(I288015), .Q(I287992) );
nand I_16834 (I287989,I288402,I288148);
DFFARX1 I_16835  ( .D(I288402), .CLK(I2350), .RSTB(I288015), .Q(I287980) );
not I_16836 (I288610,I2357);
nand I_16837 (I288627,I272129,I272117);
and I_16838 (I288644,I288627,I272114);
DFFARX1 I_16839  ( .D(I288644), .CLK(I2350), .RSTB(I288610), .Q(I288661) );
nor I_16840 (I288678,I272108,I272117);
nor I_16841 (I288695,I288678,I288661);
not I_16842 (I288593,I288678);
DFFARX1 I_16843  ( .D(I272123), .CLK(I2350), .RSTB(I288610), .Q(I288726) );
not I_16844 (I288743,I288726);
nor I_16845 (I288760,I288678,I288743);
nand I_16846 (I288596,I288726,I288695);
DFFARX1 I_16847  ( .D(I288726), .CLK(I2350), .RSTB(I288610), .Q(I288578) );
nand I_16848 (I288805,I272120,I272126);
and I_16849 (I288822,I288805,I272111);
DFFARX1 I_16850  ( .D(I288822), .CLK(I2350), .RSTB(I288610), .Q(I288839) );
nor I_16851 (I288599,I288839,I288661);
nand I_16852 (I288590,I288839,I288760);
DFFARX1 I_16853  ( .D(I272099), .CLK(I2350), .RSTB(I288610), .Q(I288884) );
and I_16854 (I288901,I288884,I272102);
DFFARX1 I_16855  ( .D(I288901), .CLK(I2350), .RSTB(I288610), .Q(I288918) );
not I_16856 (I288581,I288918);
nand I_16857 (I288949,I288901,I288839);
and I_16858 (I288966,I288661,I288949);
DFFARX1 I_16859  ( .D(I288966), .CLK(I2350), .RSTB(I288610), .Q(I288572) );
DFFARX1 I_16860  ( .D(I272105), .CLK(I2350), .RSTB(I288610), .Q(I288997) );
nand I_16861 (I289014,I288997,I288661);
and I_16862 (I289031,I288839,I289014);
DFFARX1 I_16863  ( .D(I289031), .CLK(I2350), .RSTB(I288610), .Q(I288602) );
not I_16864 (I289062,I288997);
nor I_16865 (I289079,I288678,I289062);
and I_16866 (I289096,I288997,I289079);
or I_16867 (I289113,I288901,I289096);
DFFARX1 I_16868  ( .D(I289113), .CLK(I2350), .RSTB(I288610), .Q(I288587) );
nand I_16869 (I288584,I288997,I288743);
DFFARX1 I_16870  ( .D(I288997), .CLK(I2350), .RSTB(I288610), .Q(I288575) );
not I_16871 (I289205,I2357);
nand I_16872 (I289222,I318932,I318923);
and I_16873 (I289239,I289222,I318941);
DFFARX1 I_16874  ( .D(I289239), .CLK(I2350), .RSTB(I289205), .Q(I289256) );
nor I_16875 (I289273,I318920,I318923);
nor I_16876 (I289290,I289273,I289256);
not I_16877 (I289188,I289273);
DFFARX1 I_16878  ( .D(I318929), .CLK(I2350), .RSTB(I289205), .Q(I289321) );
not I_16879 (I289338,I289321);
nor I_16880 (I289355,I289273,I289338);
nand I_16881 (I289191,I289321,I289290);
DFFARX1 I_16882  ( .D(I289321), .CLK(I2350), .RSTB(I289205), .Q(I289173) );
nand I_16883 (I289400,I318944,I318926);
and I_16884 (I289417,I289400,I318947);
DFFARX1 I_16885  ( .D(I289417), .CLK(I2350), .RSTB(I289205), .Q(I289434) );
nor I_16886 (I289194,I289434,I289256);
nand I_16887 (I289185,I289434,I289355);
DFFARX1 I_16888  ( .D(I318935), .CLK(I2350), .RSTB(I289205), .Q(I289479) );
and I_16889 (I289496,I289479,I318917);
DFFARX1 I_16890  ( .D(I289496), .CLK(I2350), .RSTB(I289205), .Q(I289513) );
not I_16891 (I289176,I289513);
nand I_16892 (I289544,I289496,I289434);
and I_16893 (I289561,I289256,I289544);
DFFARX1 I_16894  ( .D(I289561), .CLK(I2350), .RSTB(I289205), .Q(I289167) );
DFFARX1 I_16895  ( .D(I318938), .CLK(I2350), .RSTB(I289205), .Q(I289592) );
nand I_16896 (I289609,I289592,I289256);
and I_16897 (I289626,I289434,I289609);
DFFARX1 I_16898  ( .D(I289626), .CLK(I2350), .RSTB(I289205), .Q(I289197) );
not I_16899 (I289657,I289592);
nor I_16900 (I289674,I289273,I289657);
and I_16901 (I289691,I289592,I289674);
or I_16902 (I289708,I289496,I289691);
DFFARX1 I_16903  ( .D(I289708), .CLK(I2350), .RSTB(I289205), .Q(I289182) );
nand I_16904 (I289179,I289592,I289338);
DFFARX1 I_16905  ( .D(I289592), .CLK(I2350), .RSTB(I289205), .Q(I289170) );
not I_16906 (I289800,I2357);
nand I_16907 (I289817,I322502,I322493);
and I_16908 (I289834,I289817,I322511);
DFFARX1 I_16909  ( .D(I289834), .CLK(I2350), .RSTB(I289800), .Q(I289851) );
nor I_16910 (I289868,I322490,I322493);
nor I_16911 (I289885,I289868,I289851);
not I_16912 (I289783,I289868);
DFFARX1 I_16913  ( .D(I322499), .CLK(I2350), .RSTB(I289800), .Q(I289916) );
not I_16914 (I289933,I289916);
nor I_16915 (I289950,I289868,I289933);
nand I_16916 (I289786,I289916,I289885);
DFFARX1 I_16917  ( .D(I289916), .CLK(I2350), .RSTB(I289800), .Q(I289768) );
nand I_16918 (I289995,I322514,I322496);
and I_16919 (I290012,I289995,I322517);
DFFARX1 I_16920  ( .D(I290012), .CLK(I2350), .RSTB(I289800), .Q(I290029) );
nor I_16921 (I289789,I290029,I289851);
nand I_16922 (I289780,I290029,I289950);
DFFARX1 I_16923  ( .D(I322505), .CLK(I2350), .RSTB(I289800), .Q(I290074) );
and I_16924 (I290091,I290074,I322487);
DFFARX1 I_16925  ( .D(I290091), .CLK(I2350), .RSTB(I289800), .Q(I290108) );
not I_16926 (I289771,I290108);
nand I_16927 (I290139,I290091,I290029);
and I_16928 (I290156,I289851,I290139);
DFFARX1 I_16929  ( .D(I290156), .CLK(I2350), .RSTB(I289800), .Q(I289762) );
DFFARX1 I_16930  ( .D(I322508), .CLK(I2350), .RSTB(I289800), .Q(I290187) );
nand I_16931 (I290204,I290187,I289851);
and I_16932 (I290221,I290029,I290204);
DFFARX1 I_16933  ( .D(I290221), .CLK(I2350), .RSTB(I289800), .Q(I289792) );
not I_16934 (I290252,I290187);
nor I_16935 (I290269,I289868,I290252);
and I_16936 (I290286,I290187,I290269);
or I_16937 (I290303,I290091,I290286);
DFFARX1 I_16938  ( .D(I290303), .CLK(I2350), .RSTB(I289800), .Q(I289777) );
nand I_16939 (I289774,I290187,I289933);
DFFARX1 I_16940  ( .D(I290187), .CLK(I2350), .RSTB(I289800), .Q(I289765) );
not I_16941 (I290395,I2357);
nand I_16942 (I290412,I126390,I126387);
and I_16943 (I290429,I290412,I126384);
DFFARX1 I_16944  ( .D(I290429), .CLK(I2350), .RSTB(I290395), .Q(I290446) );
nor I_16945 (I290463,I126375,I126387);
nor I_16946 (I290480,I290463,I290446);
not I_16947 (I290378,I290463);
DFFARX1 I_16948  ( .D(I126393), .CLK(I2350), .RSTB(I290395), .Q(I290511) );
not I_16949 (I290528,I290511);
nor I_16950 (I290545,I290463,I290528);
nand I_16951 (I290381,I290511,I290480);
DFFARX1 I_16952  ( .D(I290511), .CLK(I2350), .RSTB(I290395), .Q(I290363) );
nand I_16953 (I290590,I126378,I126402);
and I_16954 (I290607,I290590,I126381);
DFFARX1 I_16955  ( .D(I290607), .CLK(I2350), .RSTB(I290395), .Q(I290624) );
nor I_16956 (I290384,I290624,I290446);
nand I_16957 (I290375,I290624,I290545);
DFFARX1 I_16958  ( .D(I126399), .CLK(I2350), .RSTB(I290395), .Q(I290669) );
and I_16959 (I290686,I290669,I126396);
DFFARX1 I_16960  ( .D(I290686), .CLK(I2350), .RSTB(I290395), .Q(I290703) );
not I_16961 (I290366,I290703);
nand I_16962 (I290734,I290686,I290624);
and I_16963 (I290751,I290446,I290734);
DFFARX1 I_16964  ( .D(I290751), .CLK(I2350), .RSTB(I290395), .Q(I290357) );
DFFARX1 I_16965  ( .D(I126405), .CLK(I2350), .RSTB(I290395), .Q(I290782) );
nand I_16966 (I290799,I290782,I290446);
and I_16967 (I290816,I290624,I290799);
DFFARX1 I_16968  ( .D(I290816), .CLK(I2350), .RSTB(I290395), .Q(I290387) );
not I_16969 (I290847,I290782);
nor I_16970 (I290864,I290463,I290847);
and I_16971 (I290881,I290782,I290864);
or I_16972 (I290898,I290686,I290881);
DFFARX1 I_16973  ( .D(I290898), .CLK(I2350), .RSTB(I290395), .Q(I290372) );
nand I_16974 (I290369,I290782,I290528);
DFFARX1 I_16975  ( .D(I290782), .CLK(I2350), .RSTB(I290395), .Q(I290360) );
not I_16976 (I290990,I2357);
nand I_16977 (I291007,I263762,I263765);
and I_16978 (I291024,I291007,I263759);
DFFARX1 I_16979  ( .D(I291024), .CLK(I2350), .RSTB(I290990), .Q(I291041) );
nor I_16980 (I291058,I263756,I263765);
nor I_16981 (I291075,I291058,I291041);
not I_16982 (I290973,I291058);
DFFARX1 I_16983  ( .D(I263738), .CLK(I2350), .RSTB(I290990), .Q(I291106) );
not I_16984 (I291123,I291106);
nor I_16985 (I291140,I291058,I291123);
nand I_16986 (I290976,I291106,I291075);
DFFARX1 I_16987  ( .D(I291106), .CLK(I2350), .RSTB(I290990), .Q(I290958) );
nand I_16988 (I291185,I263747,I263744);
and I_16989 (I291202,I291185,I263753);
DFFARX1 I_16990  ( .D(I291202), .CLK(I2350), .RSTB(I290990), .Q(I291219) );
nor I_16991 (I290979,I291219,I291041);
nand I_16992 (I290970,I291219,I291140);
DFFARX1 I_16993  ( .D(I263735), .CLK(I2350), .RSTB(I290990), .Q(I291264) );
and I_16994 (I291281,I291264,I263750);
DFFARX1 I_16995  ( .D(I291281), .CLK(I2350), .RSTB(I290990), .Q(I291298) );
not I_16996 (I290961,I291298);
nand I_16997 (I291329,I291281,I291219);
and I_16998 (I291346,I291041,I291329);
DFFARX1 I_16999  ( .D(I291346), .CLK(I2350), .RSTB(I290990), .Q(I290952) );
DFFARX1 I_17000  ( .D(I263741), .CLK(I2350), .RSTB(I290990), .Q(I291377) );
nand I_17001 (I291394,I291377,I291041);
and I_17002 (I291411,I291219,I291394);
DFFARX1 I_17003  ( .D(I291411), .CLK(I2350), .RSTB(I290990), .Q(I290982) );
not I_17004 (I291442,I291377);
nor I_17005 (I291459,I291058,I291442);
and I_17006 (I291476,I291377,I291459);
or I_17007 (I291493,I291281,I291476);
DFFARX1 I_17008  ( .D(I291493), .CLK(I2350), .RSTB(I290990), .Q(I290967) );
nand I_17009 (I290964,I291377,I291123);
DFFARX1 I_17010  ( .D(I291377), .CLK(I2350), .RSTB(I290990), .Q(I290955) );
not I_17011 (I291585,I2357);
nand I_17012 (I291602,I372876,I372867);
and I_17013 (I291619,I291602,I372885);
DFFARX1 I_17014  ( .D(I291619), .CLK(I2350), .RSTB(I291585), .Q(I291636) );
nor I_17015 (I291653,I372882,I372867);
nor I_17016 (I291670,I291653,I291636);
not I_17017 (I291568,I291653);
DFFARX1 I_17018  ( .D(I372864), .CLK(I2350), .RSTB(I291585), .Q(I291701) );
not I_17019 (I291718,I291701);
nor I_17020 (I291735,I291653,I291718);
nand I_17021 (I291571,I291701,I291670);
DFFARX1 I_17022  ( .D(I291701), .CLK(I2350), .RSTB(I291585), .Q(I291553) );
nand I_17023 (I291780,I372873,I372888);
and I_17024 (I291797,I291780,I372879);
DFFARX1 I_17025  ( .D(I291797), .CLK(I2350), .RSTB(I291585), .Q(I291814) );
nor I_17026 (I291574,I291814,I291636);
nand I_17027 (I291565,I291814,I291735);
DFFARX1 I_17028  ( .D(I372861), .CLK(I2350), .RSTB(I291585), .Q(I291859) );
and I_17029 (I291876,I291859,I372870);
DFFARX1 I_17030  ( .D(I291876), .CLK(I2350), .RSTB(I291585), .Q(I291893) );
not I_17031 (I291556,I291893);
nand I_17032 (I291924,I291876,I291814);
and I_17033 (I291941,I291636,I291924);
DFFARX1 I_17034  ( .D(I291941), .CLK(I2350), .RSTB(I291585), .Q(I291547) );
DFFARX1 I_17035  ( .D(I372858), .CLK(I2350), .RSTB(I291585), .Q(I291972) );
nand I_17036 (I291989,I291972,I291636);
and I_17037 (I292006,I291814,I291989);
DFFARX1 I_17038  ( .D(I292006), .CLK(I2350), .RSTB(I291585), .Q(I291577) );
not I_17039 (I292037,I291972);
nor I_17040 (I292054,I291653,I292037);
and I_17041 (I292071,I291972,I292054);
or I_17042 (I292088,I291876,I292071);
DFFARX1 I_17043  ( .D(I292088), .CLK(I2350), .RSTB(I291585), .Q(I291562) );
nand I_17044 (I291559,I291972,I291718);
DFFARX1 I_17045  ( .D(I291972), .CLK(I2350), .RSTB(I291585), .Q(I291550) );
not I_17046 (I292180,I2357);
nand I_17047 (I292197,I92682,I92694);
and I_17048 (I292214,I292197,I92673);
DFFARX1 I_17049  ( .D(I292214), .CLK(I2350), .RSTB(I292180), .Q(I292231) );
nor I_17050 (I292248,I92664,I92694);
nor I_17051 (I292265,I292248,I292231);
not I_17052 (I292163,I292248);
DFFARX1 I_17053  ( .D(I92676), .CLK(I2350), .RSTB(I292180), .Q(I292296) );
not I_17054 (I292313,I292296);
nor I_17055 (I292330,I292248,I292313);
nand I_17056 (I292166,I292296,I292265);
DFFARX1 I_17057  ( .D(I292296), .CLK(I2350), .RSTB(I292180), .Q(I292148) );
nand I_17058 (I292375,I92691,I92679);
and I_17059 (I292392,I292375,I92667);
DFFARX1 I_17060  ( .D(I292392), .CLK(I2350), .RSTB(I292180), .Q(I292409) );
nor I_17061 (I292169,I292409,I292231);
nand I_17062 (I292160,I292409,I292330);
DFFARX1 I_17063  ( .D(I92685), .CLK(I2350), .RSTB(I292180), .Q(I292454) );
and I_17064 (I292471,I292454,I92670);
DFFARX1 I_17065  ( .D(I292471), .CLK(I2350), .RSTB(I292180), .Q(I292488) );
not I_17066 (I292151,I292488);
nand I_17067 (I292519,I292471,I292409);
and I_17068 (I292536,I292231,I292519);
DFFARX1 I_17069  ( .D(I292536), .CLK(I2350), .RSTB(I292180), .Q(I292142) );
DFFARX1 I_17070  ( .D(I92688), .CLK(I2350), .RSTB(I292180), .Q(I292567) );
nand I_17071 (I292584,I292567,I292231);
and I_17072 (I292601,I292409,I292584);
DFFARX1 I_17073  ( .D(I292601), .CLK(I2350), .RSTB(I292180), .Q(I292172) );
not I_17074 (I292632,I292567);
nor I_17075 (I292649,I292248,I292632);
and I_17076 (I292666,I292567,I292649);
or I_17077 (I292683,I292471,I292666);
DFFARX1 I_17078  ( .D(I292683), .CLK(I2350), .RSTB(I292180), .Q(I292157) );
nand I_17079 (I292154,I292567,I292313);
DFFARX1 I_17080  ( .D(I292567), .CLK(I2350), .RSTB(I292180), .Q(I292145) );
not I_17081 (I292775,I2357);
nand I_17082 (I292792,I267876,I267849);
and I_17083 (I292809,I292792,I267852);
DFFARX1 I_17084  ( .D(I292809), .CLK(I2350), .RSTB(I292775), .Q(I292826) );
nor I_17085 (I292843,I267861,I267849);
nor I_17086 (I292860,I292843,I292826);
not I_17087 (I292758,I292843);
DFFARX1 I_17088  ( .D(I267858), .CLK(I2350), .RSTB(I292775), .Q(I292891) );
not I_17089 (I292908,I292891);
nor I_17090 (I292925,I292843,I292908);
nand I_17091 (I292761,I292891,I292860);
DFFARX1 I_17092  ( .D(I292891), .CLK(I2350), .RSTB(I292775), .Q(I292743) );
nand I_17093 (I292970,I267855,I267864);
and I_17094 (I292987,I292970,I267873);
DFFARX1 I_17095  ( .D(I292987), .CLK(I2350), .RSTB(I292775), .Q(I293004) );
nor I_17096 (I292764,I293004,I292826);
nand I_17097 (I292755,I293004,I292925);
DFFARX1 I_17098  ( .D(I267879), .CLK(I2350), .RSTB(I292775), .Q(I293049) );
and I_17099 (I293066,I293049,I267870);
DFFARX1 I_17100  ( .D(I293066), .CLK(I2350), .RSTB(I292775), .Q(I293083) );
not I_17101 (I292746,I293083);
nand I_17102 (I293114,I293066,I293004);
and I_17103 (I293131,I292826,I293114);
DFFARX1 I_17104  ( .D(I293131), .CLK(I2350), .RSTB(I292775), .Q(I292737) );
DFFARX1 I_17105  ( .D(I267867), .CLK(I2350), .RSTB(I292775), .Q(I293162) );
nand I_17106 (I293179,I293162,I292826);
and I_17107 (I293196,I293004,I293179);
DFFARX1 I_17108  ( .D(I293196), .CLK(I2350), .RSTB(I292775), .Q(I292767) );
not I_17109 (I293227,I293162);
nor I_17110 (I293244,I292843,I293227);
and I_17111 (I293261,I293162,I293244);
or I_17112 (I293278,I293066,I293261);
DFFARX1 I_17113  ( .D(I293278), .CLK(I2350), .RSTB(I292775), .Q(I292752) );
nand I_17114 (I292749,I293162,I292908);
DFFARX1 I_17115  ( .D(I293162), .CLK(I2350), .RSTB(I292775), .Q(I292740) );
not I_17116 (I293370,I2357);
nand I_17117 (I293387,I374763,I374754);
and I_17118 (I293404,I293387,I374772);
DFFARX1 I_17119  ( .D(I293404), .CLK(I2350), .RSTB(I293370), .Q(I293421) );
nor I_17120 (I293438,I374769,I374754);
nor I_17121 (I293455,I293438,I293421);
not I_17122 (I293353,I293438);
DFFARX1 I_17123  ( .D(I374751), .CLK(I2350), .RSTB(I293370), .Q(I293486) );
not I_17124 (I293503,I293486);
nor I_17125 (I293520,I293438,I293503);
nand I_17126 (I293356,I293486,I293455);
DFFARX1 I_17127  ( .D(I293486), .CLK(I2350), .RSTB(I293370), .Q(I293338) );
nand I_17128 (I293565,I374760,I374775);
and I_17129 (I293582,I293565,I374766);
DFFARX1 I_17130  ( .D(I293582), .CLK(I2350), .RSTB(I293370), .Q(I293599) );
nor I_17131 (I293359,I293599,I293421);
nand I_17132 (I293350,I293599,I293520);
DFFARX1 I_17133  ( .D(I374748), .CLK(I2350), .RSTB(I293370), .Q(I293644) );
and I_17134 (I293661,I293644,I374757);
DFFARX1 I_17135  ( .D(I293661), .CLK(I2350), .RSTB(I293370), .Q(I293678) );
not I_17136 (I293341,I293678);
nand I_17137 (I293709,I293661,I293599);
and I_17138 (I293726,I293421,I293709);
DFFARX1 I_17139  ( .D(I293726), .CLK(I2350), .RSTB(I293370), .Q(I293332) );
DFFARX1 I_17140  ( .D(I374745), .CLK(I2350), .RSTB(I293370), .Q(I293757) );
nand I_17141 (I293774,I293757,I293421);
and I_17142 (I293791,I293599,I293774);
DFFARX1 I_17143  ( .D(I293791), .CLK(I2350), .RSTB(I293370), .Q(I293362) );
not I_17144 (I293822,I293757);
nor I_17145 (I293839,I293438,I293822);
and I_17146 (I293856,I293757,I293839);
or I_17147 (I293873,I293661,I293856);
DFFARX1 I_17148  ( .D(I293873), .CLK(I2350), .RSTB(I293370), .Q(I293347) );
nand I_17149 (I293344,I293757,I293503);
DFFARX1 I_17150  ( .D(I293757), .CLK(I2350), .RSTB(I293370), .Q(I293335) );
not I_17151 (I293965,I2357);
nand I_17152 (I293982,I391451,I391457);
and I_17153 (I293999,I293982,I391448);
DFFARX1 I_17154  ( .D(I293999), .CLK(I2350), .RSTB(I293965), .Q(I294016) );
nor I_17155 (I294033,I391460,I391457);
nor I_17156 (I294050,I294033,I294016);
not I_17157 (I293948,I294033);
DFFARX1 I_17158  ( .D(I391439), .CLK(I2350), .RSTB(I293965), .Q(I294081) );
not I_17159 (I294098,I294081);
nor I_17160 (I294115,I294033,I294098);
nand I_17161 (I293951,I294081,I294050);
DFFARX1 I_17162  ( .D(I294081), .CLK(I2350), .RSTB(I293965), .Q(I293933) );
nand I_17163 (I294160,I391463,I391445);
and I_17164 (I294177,I294160,I391454);
DFFARX1 I_17165  ( .D(I294177), .CLK(I2350), .RSTB(I293965), .Q(I294194) );
nor I_17166 (I293954,I294194,I294016);
nand I_17167 (I293945,I294194,I294115);
DFFARX1 I_17168  ( .D(I391469), .CLK(I2350), .RSTB(I293965), .Q(I294239) );
and I_17169 (I294256,I294239,I391442);
DFFARX1 I_17170  ( .D(I294256), .CLK(I2350), .RSTB(I293965), .Q(I294273) );
not I_17171 (I293936,I294273);
nand I_17172 (I294304,I294256,I294194);
and I_17173 (I294321,I294016,I294304);
DFFARX1 I_17174  ( .D(I294321), .CLK(I2350), .RSTB(I293965), .Q(I293927) );
DFFARX1 I_17175  ( .D(I391466), .CLK(I2350), .RSTB(I293965), .Q(I294352) );
nand I_17176 (I294369,I294352,I294016);
and I_17177 (I294386,I294194,I294369);
DFFARX1 I_17178  ( .D(I294386), .CLK(I2350), .RSTB(I293965), .Q(I293957) );
not I_17179 (I294417,I294352);
nor I_17180 (I294434,I294033,I294417);
and I_17181 (I294451,I294352,I294434);
or I_17182 (I294468,I294256,I294451);
DFFARX1 I_17183  ( .D(I294468), .CLK(I2350), .RSTB(I293965), .Q(I293942) );
nand I_17184 (I293939,I294352,I294098);
DFFARX1 I_17185  ( .D(I294352), .CLK(I2350), .RSTB(I293965), .Q(I293930) );
not I_17186 (I294560,I2357);
nand I_17187 (I294577,I335765,I335756);
and I_17188 (I294594,I294577,I335774);
DFFARX1 I_17189  ( .D(I294594), .CLK(I2350), .RSTB(I294560), .Q(I294611) );
nor I_17190 (I294628,I335771,I335756);
nor I_17191 (I294645,I294628,I294611);
not I_17192 (I294543,I294628);
DFFARX1 I_17193  ( .D(I335753), .CLK(I2350), .RSTB(I294560), .Q(I294676) );
not I_17194 (I294693,I294676);
nor I_17195 (I294710,I294628,I294693);
nand I_17196 (I294546,I294676,I294645);
DFFARX1 I_17197  ( .D(I294676), .CLK(I2350), .RSTB(I294560), .Q(I294528) );
nand I_17198 (I294755,I335762,I335777);
and I_17199 (I294772,I294755,I335768);
DFFARX1 I_17200  ( .D(I294772), .CLK(I2350), .RSTB(I294560), .Q(I294789) );
nor I_17201 (I294549,I294789,I294611);
nand I_17202 (I294540,I294789,I294710);
DFFARX1 I_17203  ( .D(I335750), .CLK(I2350), .RSTB(I294560), .Q(I294834) );
and I_17204 (I294851,I294834,I335759);
DFFARX1 I_17205  ( .D(I294851), .CLK(I2350), .RSTB(I294560), .Q(I294868) );
not I_17206 (I294531,I294868);
nand I_17207 (I294899,I294851,I294789);
and I_17208 (I294916,I294611,I294899);
DFFARX1 I_17209  ( .D(I294916), .CLK(I2350), .RSTB(I294560), .Q(I294522) );
DFFARX1 I_17210  ( .D(I335747), .CLK(I2350), .RSTB(I294560), .Q(I294947) );
nand I_17211 (I294964,I294947,I294611);
and I_17212 (I294981,I294789,I294964);
DFFARX1 I_17213  ( .D(I294981), .CLK(I2350), .RSTB(I294560), .Q(I294552) );
not I_17214 (I295012,I294947);
nor I_17215 (I295029,I294628,I295012);
and I_17216 (I295046,I294947,I295029);
or I_17217 (I295063,I294851,I295046);
DFFARX1 I_17218  ( .D(I295063), .CLK(I2350), .RSTB(I294560), .Q(I294537) );
nand I_17219 (I294534,I294947,I294693);
DFFARX1 I_17220  ( .D(I294947), .CLK(I2350), .RSTB(I294560), .Q(I294525) );
not I_17221 (I295155,I2357);
nand I_17222 (I295172,I331427,I331418);
and I_17223 (I295189,I295172,I331436);
DFFARX1 I_17224  ( .D(I295189), .CLK(I2350), .RSTB(I295155), .Q(I295206) );
nor I_17225 (I295223,I331415,I331418);
nor I_17226 (I295240,I295223,I295206);
not I_17227 (I295138,I295223);
DFFARX1 I_17228  ( .D(I331424), .CLK(I2350), .RSTB(I295155), .Q(I295271) );
not I_17229 (I295288,I295271);
nor I_17230 (I295305,I295223,I295288);
nand I_17231 (I295141,I295271,I295240);
DFFARX1 I_17232  ( .D(I295271), .CLK(I2350), .RSTB(I295155), .Q(I295123) );
nand I_17233 (I295350,I331439,I331421);
and I_17234 (I295367,I295350,I331442);
DFFARX1 I_17235  ( .D(I295367), .CLK(I2350), .RSTB(I295155), .Q(I295384) );
nor I_17236 (I295144,I295384,I295206);
nand I_17237 (I295135,I295384,I295305);
DFFARX1 I_17238  ( .D(I331430), .CLK(I2350), .RSTB(I295155), .Q(I295429) );
and I_17239 (I295446,I295429,I331412);
DFFARX1 I_17240  ( .D(I295446), .CLK(I2350), .RSTB(I295155), .Q(I295463) );
not I_17241 (I295126,I295463);
nand I_17242 (I295494,I295446,I295384);
and I_17243 (I295511,I295206,I295494);
DFFARX1 I_17244  ( .D(I295511), .CLK(I2350), .RSTB(I295155), .Q(I295117) );
DFFARX1 I_17245  ( .D(I331433), .CLK(I2350), .RSTB(I295155), .Q(I295542) );
nand I_17246 (I295559,I295542,I295206);
and I_17247 (I295576,I295384,I295559);
DFFARX1 I_17248  ( .D(I295576), .CLK(I2350), .RSTB(I295155), .Q(I295147) );
not I_17249 (I295607,I295542);
nor I_17250 (I295624,I295223,I295607);
and I_17251 (I295641,I295542,I295624);
or I_17252 (I295658,I295446,I295641);
DFFARX1 I_17253  ( .D(I295658), .CLK(I2350), .RSTB(I295155), .Q(I295132) );
nand I_17254 (I295129,I295542,I295288);
DFFARX1 I_17255  ( .D(I295542), .CLK(I2350), .RSTB(I295155), .Q(I295120) );
not I_17256 (I295750,I2357);
nand I_17257 (I295767,I182119,I182125);
and I_17258 (I295784,I295767,I182107);
DFFARX1 I_17259  ( .D(I295784), .CLK(I2350), .RSTB(I295750), .Q(I295801) );
nor I_17260 (I295818,I182101,I182125);
nor I_17261 (I295835,I295818,I295801);
not I_17262 (I295733,I295818);
DFFARX1 I_17263  ( .D(I182131), .CLK(I2350), .RSTB(I295750), .Q(I295866) );
not I_17264 (I295883,I295866);
nor I_17265 (I295900,I295818,I295883);
nand I_17266 (I295736,I295866,I295835);
DFFARX1 I_17267  ( .D(I295866), .CLK(I2350), .RSTB(I295750), .Q(I295718) );
nand I_17268 (I295945,I182122,I182113);
and I_17269 (I295962,I295945,I182116);
DFFARX1 I_17270  ( .D(I295962), .CLK(I2350), .RSTB(I295750), .Q(I295979) );
nor I_17271 (I295739,I295979,I295801);
nand I_17272 (I295730,I295979,I295900);
DFFARX1 I_17273  ( .D(I182128), .CLK(I2350), .RSTB(I295750), .Q(I296024) );
and I_17274 (I296041,I296024,I182104);
DFFARX1 I_17275  ( .D(I296041), .CLK(I2350), .RSTB(I295750), .Q(I296058) );
not I_17276 (I295721,I296058);
nand I_17277 (I296089,I296041,I295979);
and I_17278 (I296106,I295801,I296089);
DFFARX1 I_17279  ( .D(I296106), .CLK(I2350), .RSTB(I295750), .Q(I295712) );
DFFARX1 I_17280  ( .D(I182110), .CLK(I2350), .RSTB(I295750), .Q(I296137) );
nand I_17281 (I296154,I296137,I295801);
and I_17282 (I296171,I295979,I296154);
DFFARX1 I_17283  ( .D(I296171), .CLK(I2350), .RSTB(I295750), .Q(I295742) );
not I_17284 (I296202,I296137);
nor I_17285 (I296219,I295818,I296202);
and I_17286 (I296236,I296137,I296219);
or I_17287 (I296253,I296041,I296236);
DFFARX1 I_17288  ( .D(I296253), .CLK(I2350), .RSTB(I295750), .Q(I295727) );
nand I_17289 (I295724,I296137,I295883);
DFFARX1 I_17290  ( .D(I296137), .CLK(I2350), .RSTB(I295750), .Q(I295715) );
not I_17291 (I296345,I2357);
nand I_17292 (I296362,I260294,I260297);
and I_17293 (I296379,I296362,I260291);
DFFARX1 I_17294  ( .D(I296379), .CLK(I2350), .RSTB(I296345), .Q(I296396) );
nor I_17295 (I296413,I260288,I260297);
nor I_17296 (I296430,I296413,I296396);
not I_17297 (I296328,I296413);
DFFARX1 I_17298  ( .D(I260270), .CLK(I2350), .RSTB(I296345), .Q(I296461) );
not I_17299 (I296478,I296461);
nor I_17300 (I296495,I296413,I296478);
nand I_17301 (I296331,I296461,I296430);
DFFARX1 I_17302  ( .D(I296461), .CLK(I2350), .RSTB(I296345), .Q(I296313) );
nand I_17303 (I296540,I260279,I260276);
and I_17304 (I296557,I296540,I260285);
DFFARX1 I_17305  ( .D(I296557), .CLK(I2350), .RSTB(I296345), .Q(I296574) );
nor I_17306 (I296334,I296574,I296396);
nand I_17307 (I296325,I296574,I296495);
DFFARX1 I_17308  ( .D(I260267), .CLK(I2350), .RSTB(I296345), .Q(I296619) );
and I_17309 (I296636,I296619,I260282);
DFFARX1 I_17310  ( .D(I296636), .CLK(I2350), .RSTB(I296345), .Q(I296653) );
not I_17311 (I296316,I296653);
nand I_17312 (I296684,I296636,I296574);
and I_17313 (I296701,I296396,I296684);
DFFARX1 I_17314  ( .D(I296701), .CLK(I2350), .RSTB(I296345), .Q(I296307) );
DFFARX1 I_17315  ( .D(I260273), .CLK(I2350), .RSTB(I296345), .Q(I296732) );
nand I_17316 (I296749,I296732,I296396);
and I_17317 (I296766,I296574,I296749);
DFFARX1 I_17318  ( .D(I296766), .CLK(I2350), .RSTB(I296345), .Q(I296337) );
not I_17319 (I296797,I296732);
nor I_17320 (I296814,I296413,I296797);
and I_17321 (I296831,I296732,I296814);
or I_17322 (I296848,I296636,I296831);
DFFARX1 I_17323  ( .D(I296848), .CLK(I2350), .RSTB(I296345), .Q(I296322) );
nand I_17324 (I296319,I296732,I296478);
DFFARX1 I_17325  ( .D(I296732), .CLK(I2350), .RSTB(I296345), .Q(I296310) );
not I_17326 (I296940,I2357);
nand I_17327 (I296957,I107268,I107280);
and I_17328 (I296974,I296957,I107259);
DFFARX1 I_17329  ( .D(I296974), .CLK(I2350), .RSTB(I296940), .Q(I296991) );
nor I_17330 (I297008,I107250,I107280);
nor I_17331 (I297025,I297008,I296991);
not I_17332 (I296923,I297008);
DFFARX1 I_17333  ( .D(I107262), .CLK(I2350), .RSTB(I296940), .Q(I297056) );
not I_17334 (I297073,I297056);
nor I_17335 (I297090,I297008,I297073);
nand I_17336 (I296926,I297056,I297025);
DFFARX1 I_17337  ( .D(I297056), .CLK(I2350), .RSTB(I296940), .Q(I296908) );
nand I_17338 (I297135,I107277,I107265);
and I_17339 (I297152,I297135,I107253);
DFFARX1 I_17340  ( .D(I297152), .CLK(I2350), .RSTB(I296940), .Q(I297169) );
nor I_17341 (I296929,I297169,I296991);
nand I_17342 (I296920,I297169,I297090);
DFFARX1 I_17343  ( .D(I107271), .CLK(I2350), .RSTB(I296940), .Q(I297214) );
and I_17344 (I297231,I297214,I107256);
DFFARX1 I_17345  ( .D(I297231), .CLK(I2350), .RSTB(I296940), .Q(I297248) );
not I_17346 (I296911,I297248);
nand I_17347 (I297279,I297231,I297169);
and I_17348 (I297296,I296991,I297279);
DFFARX1 I_17349  ( .D(I297296), .CLK(I2350), .RSTB(I296940), .Q(I296902) );
DFFARX1 I_17350  ( .D(I107274), .CLK(I2350), .RSTB(I296940), .Q(I297327) );
nand I_17351 (I297344,I297327,I296991);
and I_17352 (I297361,I297169,I297344);
DFFARX1 I_17353  ( .D(I297361), .CLK(I2350), .RSTB(I296940), .Q(I296932) );
not I_17354 (I297392,I297327);
nor I_17355 (I297409,I297008,I297392);
and I_17356 (I297426,I297327,I297409);
or I_17357 (I297443,I297231,I297426);
DFFARX1 I_17358  ( .D(I297443), .CLK(I2350), .RSTB(I296940), .Q(I296917) );
nand I_17359 (I296914,I297327,I297073);
DFFARX1 I_17360  ( .D(I297327), .CLK(I2350), .RSTB(I296940), .Q(I296905) );
not I_17361 (I297535,I2357);
nand I_17362 (I297552,I55647,I55659);
and I_17363 (I297569,I297552,I55668);
DFFARX1 I_17364  ( .D(I297569), .CLK(I2350), .RSTB(I297535), .Q(I297586) );
nor I_17365 (I297603,I55662,I55659);
nor I_17366 (I297620,I297603,I297586);
not I_17367 (I297518,I297603);
DFFARX1 I_17368  ( .D(I55656), .CLK(I2350), .RSTB(I297535), .Q(I297651) );
not I_17369 (I297668,I297651);
nor I_17370 (I297685,I297603,I297668);
nand I_17371 (I297521,I297651,I297620);
DFFARX1 I_17372  ( .D(I297651), .CLK(I2350), .RSTB(I297535), .Q(I297503) );
nand I_17373 (I297730,I55653,I55650);
and I_17374 (I297747,I297730,I55641);
DFFARX1 I_17375  ( .D(I297747), .CLK(I2350), .RSTB(I297535), .Q(I297764) );
nor I_17376 (I297524,I297764,I297586);
nand I_17377 (I297515,I297764,I297685);
DFFARX1 I_17378  ( .D(I55665), .CLK(I2350), .RSTB(I297535), .Q(I297809) );
and I_17379 (I297826,I297809,I55644);
DFFARX1 I_17380  ( .D(I297826), .CLK(I2350), .RSTB(I297535), .Q(I297843) );
not I_17381 (I297506,I297843);
nand I_17382 (I297874,I297826,I297764);
and I_17383 (I297891,I297586,I297874);
DFFARX1 I_17384  ( .D(I297891), .CLK(I2350), .RSTB(I297535), .Q(I297497) );
DFFARX1 I_17385  ( .D(I55638), .CLK(I2350), .RSTB(I297535), .Q(I297922) );
nand I_17386 (I297939,I297922,I297586);
and I_17387 (I297956,I297764,I297939);
DFFARX1 I_17388  ( .D(I297956), .CLK(I2350), .RSTB(I297535), .Q(I297527) );
not I_17389 (I297987,I297922);
nor I_17390 (I298004,I297603,I297987);
and I_17391 (I298021,I297922,I298004);
or I_17392 (I298038,I297826,I298021);
DFFARX1 I_17393  ( .D(I298038), .CLK(I2350), .RSTB(I297535), .Q(I297512) );
nand I_17394 (I297509,I297922,I297668);
DFFARX1 I_17395  ( .D(I297922), .CLK(I2350), .RSTB(I297535), .Q(I297500) );
not I_17396 (I298130,I2357);
nand I_17397 (I298147,I98649,I98661);
and I_17398 (I298164,I298147,I98640);
DFFARX1 I_17399  ( .D(I298164), .CLK(I2350), .RSTB(I298130), .Q(I298181) );
nor I_17400 (I298198,I98631,I98661);
nor I_17401 (I298215,I298198,I298181);
not I_17402 (I298113,I298198);
DFFARX1 I_17403  ( .D(I98643), .CLK(I2350), .RSTB(I298130), .Q(I298246) );
not I_17404 (I298263,I298246);
nor I_17405 (I298280,I298198,I298263);
nand I_17406 (I298116,I298246,I298215);
DFFARX1 I_17407  ( .D(I298246), .CLK(I2350), .RSTB(I298130), .Q(I298098) );
nand I_17408 (I298325,I98658,I98646);
and I_17409 (I298342,I298325,I98634);
DFFARX1 I_17410  ( .D(I298342), .CLK(I2350), .RSTB(I298130), .Q(I298359) );
nor I_17411 (I298119,I298359,I298181);
nand I_17412 (I298110,I298359,I298280);
DFFARX1 I_17413  ( .D(I98652), .CLK(I2350), .RSTB(I298130), .Q(I298404) );
and I_17414 (I298421,I298404,I98637);
DFFARX1 I_17415  ( .D(I298421), .CLK(I2350), .RSTB(I298130), .Q(I298438) );
not I_17416 (I298101,I298438);
nand I_17417 (I298469,I298421,I298359);
and I_17418 (I298486,I298181,I298469);
DFFARX1 I_17419  ( .D(I298486), .CLK(I2350), .RSTB(I298130), .Q(I298092) );
DFFARX1 I_17420  ( .D(I98655), .CLK(I2350), .RSTB(I298130), .Q(I298517) );
nand I_17421 (I298534,I298517,I298181);
and I_17422 (I298551,I298359,I298534);
DFFARX1 I_17423  ( .D(I298551), .CLK(I2350), .RSTB(I298130), .Q(I298122) );
not I_17424 (I298582,I298517);
nor I_17425 (I298599,I298198,I298582);
and I_17426 (I298616,I298517,I298599);
or I_17427 (I298633,I298421,I298616);
DFFARX1 I_17428  ( .D(I298633), .CLK(I2350), .RSTB(I298130), .Q(I298107) );
nand I_17429 (I298104,I298517,I298263);
DFFARX1 I_17430  ( .D(I298517), .CLK(I2350), .RSTB(I298130), .Q(I298095) );
not I_17431 (I298725,I2357);
nand I_17432 (I298742,I180130,I180136);
and I_17433 (I298759,I298742,I180118);
DFFARX1 I_17434  ( .D(I298759), .CLK(I2350), .RSTB(I298725), .Q(I298776) );
nor I_17435 (I298793,I180112,I180136);
nor I_17436 (I298810,I298793,I298776);
not I_17437 (I298708,I298793);
DFFARX1 I_17438  ( .D(I180142), .CLK(I2350), .RSTB(I298725), .Q(I298841) );
not I_17439 (I298858,I298841);
nor I_17440 (I298875,I298793,I298858);
nand I_17441 (I298711,I298841,I298810);
DFFARX1 I_17442  ( .D(I298841), .CLK(I2350), .RSTB(I298725), .Q(I298693) );
nand I_17443 (I298920,I180133,I180124);
and I_17444 (I298937,I298920,I180127);
DFFARX1 I_17445  ( .D(I298937), .CLK(I2350), .RSTB(I298725), .Q(I298954) );
nor I_17446 (I298714,I298954,I298776);
nand I_17447 (I298705,I298954,I298875);
DFFARX1 I_17448  ( .D(I180139), .CLK(I2350), .RSTB(I298725), .Q(I298999) );
and I_17449 (I299016,I298999,I180115);
DFFARX1 I_17450  ( .D(I299016), .CLK(I2350), .RSTB(I298725), .Q(I299033) );
not I_17451 (I298696,I299033);
nand I_17452 (I299064,I299016,I298954);
and I_17453 (I299081,I298776,I299064);
DFFARX1 I_17454  ( .D(I299081), .CLK(I2350), .RSTB(I298725), .Q(I298687) );
DFFARX1 I_17455  ( .D(I180121), .CLK(I2350), .RSTB(I298725), .Q(I299112) );
nand I_17456 (I299129,I299112,I298776);
and I_17457 (I299146,I298954,I299129);
DFFARX1 I_17458  ( .D(I299146), .CLK(I2350), .RSTB(I298725), .Q(I298717) );
not I_17459 (I299177,I299112);
nor I_17460 (I299194,I298793,I299177);
and I_17461 (I299211,I299112,I299194);
or I_17462 (I299228,I299016,I299211);
DFFARX1 I_17463  ( .D(I299228), .CLK(I2350), .RSTB(I298725), .Q(I298702) );
nand I_17464 (I298699,I299112,I298858);
DFFARX1 I_17465  ( .D(I299112), .CLK(I2350), .RSTB(I298725), .Q(I298690) );
not I_17466 (I299320,I2357);
nand I_17467 (I299337,I143002,I143008);
and I_17468 (I299354,I299337,I142990);
DFFARX1 I_17469  ( .D(I299354), .CLK(I2350), .RSTB(I299320), .Q(I299371) );
nor I_17470 (I299388,I142984,I143008);
nor I_17471 (I299405,I299388,I299371);
not I_17472 (I299303,I299388);
DFFARX1 I_17473  ( .D(I143014), .CLK(I2350), .RSTB(I299320), .Q(I299436) );
not I_17474 (I299453,I299436);
nor I_17475 (I299470,I299388,I299453);
nand I_17476 (I299306,I299436,I299405);
DFFARX1 I_17477  ( .D(I299436), .CLK(I2350), .RSTB(I299320), .Q(I299288) );
nand I_17478 (I299515,I143005,I142996);
and I_17479 (I299532,I299515,I142999);
DFFARX1 I_17480  ( .D(I299532), .CLK(I2350), .RSTB(I299320), .Q(I299549) );
nor I_17481 (I299309,I299549,I299371);
nand I_17482 (I299300,I299549,I299470);
DFFARX1 I_17483  ( .D(I143011), .CLK(I2350), .RSTB(I299320), .Q(I299594) );
and I_17484 (I299611,I299594,I142987);
DFFARX1 I_17485  ( .D(I299611), .CLK(I2350), .RSTB(I299320), .Q(I299628) );
not I_17486 (I299291,I299628);
nand I_17487 (I299659,I299611,I299549);
and I_17488 (I299676,I299371,I299659);
DFFARX1 I_17489  ( .D(I299676), .CLK(I2350), .RSTB(I299320), .Q(I299282) );
DFFARX1 I_17490  ( .D(I142993), .CLK(I2350), .RSTB(I299320), .Q(I299707) );
nand I_17491 (I299724,I299707,I299371);
and I_17492 (I299741,I299549,I299724);
DFFARX1 I_17493  ( .D(I299741), .CLK(I2350), .RSTB(I299320), .Q(I299312) );
not I_17494 (I299772,I299707);
nor I_17495 (I299789,I299388,I299772);
and I_17496 (I299806,I299707,I299789);
or I_17497 (I299823,I299611,I299806);
DFFARX1 I_17498  ( .D(I299823), .CLK(I2350), .RSTB(I299320), .Q(I299297) );
nand I_17499 (I299294,I299707,I299453);
DFFARX1 I_17500  ( .D(I299707), .CLK(I2350), .RSTB(I299320), .Q(I299285) );
not I_17501 (I299915,I2357);
nand I_17502 (I299932,I265496,I265499);
and I_17503 (I299949,I299932,I265493);
DFFARX1 I_17504  ( .D(I299949), .CLK(I2350), .RSTB(I299915), .Q(I299966) );
nor I_17505 (I299983,I265490,I265499);
nor I_17506 (I300000,I299983,I299966);
not I_17507 (I299898,I299983);
DFFARX1 I_17508  ( .D(I265472), .CLK(I2350), .RSTB(I299915), .Q(I300031) );
not I_17509 (I300048,I300031);
nor I_17510 (I300065,I299983,I300048);
nand I_17511 (I299901,I300031,I300000);
DFFARX1 I_17512  ( .D(I300031), .CLK(I2350), .RSTB(I299915), .Q(I299883) );
nand I_17513 (I300110,I265481,I265478);
and I_17514 (I300127,I300110,I265487);
DFFARX1 I_17515  ( .D(I300127), .CLK(I2350), .RSTB(I299915), .Q(I300144) );
nor I_17516 (I299904,I300144,I299966);
nand I_17517 (I299895,I300144,I300065);
DFFARX1 I_17518  ( .D(I265469), .CLK(I2350), .RSTB(I299915), .Q(I300189) );
and I_17519 (I300206,I300189,I265484);
DFFARX1 I_17520  ( .D(I300206), .CLK(I2350), .RSTB(I299915), .Q(I300223) );
not I_17521 (I299886,I300223);
nand I_17522 (I300254,I300206,I300144);
and I_17523 (I300271,I299966,I300254);
DFFARX1 I_17524  ( .D(I300271), .CLK(I2350), .RSTB(I299915), .Q(I299877) );
DFFARX1 I_17525  ( .D(I265475), .CLK(I2350), .RSTB(I299915), .Q(I300302) );
nand I_17526 (I300319,I300302,I299966);
and I_17527 (I300336,I300144,I300319);
DFFARX1 I_17528  ( .D(I300336), .CLK(I2350), .RSTB(I299915), .Q(I299907) );
not I_17529 (I300367,I300302);
nor I_17530 (I300384,I299983,I300367);
and I_17531 (I300401,I300302,I300384);
or I_17532 (I300418,I300206,I300401);
DFFARX1 I_17533  ( .D(I300418), .CLK(I2350), .RSTB(I299915), .Q(I299892) );
nand I_17534 (I299889,I300302,I300048);
DFFARX1 I_17535  ( .D(I300302), .CLK(I2350), .RSTB(I299915), .Q(I299880) );
not I_17536 (I300510,I2357);
nand I_17537 (I300527,I370360,I370351);
and I_17538 (I300544,I300527,I370369);
DFFARX1 I_17539  ( .D(I300544), .CLK(I2350), .RSTB(I300510), .Q(I300561) );
nor I_17540 (I300578,I370366,I370351);
nor I_17541 (I300595,I300578,I300561);
not I_17542 (I300493,I300578);
DFFARX1 I_17543  ( .D(I370348), .CLK(I2350), .RSTB(I300510), .Q(I300626) );
not I_17544 (I300643,I300626);
nor I_17545 (I300660,I300578,I300643);
nand I_17546 (I300496,I300626,I300595);
DFFARX1 I_17547  ( .D(I300626), .CLK(I2350), .RSTB(I300510), .Q(I300478) );
nand I_17548 (I300705,I370357,I370372);
and I_17549 (I300722,I300705,I370363);
DFFARX1 I_17550  ( .D(I300722), .CLK(I2350), .RSTB(I300510), .Q(I300739) );
nor I_17551 (I300499,I300739,I300561);
nand I_17552 (I300490,I300739,I300660);
DFFARX1 I_17553  ( .D(I370345), .CLK(I2350), .RSTB(I300510), .Q(I300784) );
and I_17554 (I300801,I300784,I370354);
DFFARX1 I_17555  ( .D(I300801), .CLK(I2350), .RSTB(I300510), .Q(I300818) );
not I_17556 (I300481,I300818);
nand I_17557 (I300849,I300801,I300739);
and I_17558 (I300866,I300561,I300849);
DFFARX1 I_17559  ( .D(I300866), .CLK(I2350), .RSTB(I300510), .Q(I300472) );
DFFARX1 I_17560  ( .D(I370342), .CLK(I2350), .RSTB(I300510), .Q(I300897) );
nand I_17561 (I300914,I300897,I300561);
and I_17562 (I300931,I300739,I300914);
DFFARX1 I_17563  ( .D(I300931), .CLK(I2350), .RSTB(I300510), .Q(I300502) );
not I_17564 (I300962,I300897);
nor I_17565 (I300979,I300578,I300962);
and I_17566 (I300996,I300897,I300979);
or I_17567 (I301013,I300801,I300996);
DFFARX1 I_17568  ( .D(I301013), .CLK(I2350), .RSTB(I300510), .Q(I300487) );
nand I_17569 (I300484,I300897,I300643);
DFFARX1 I_17570  ( .D(I300897), .CLK(I2350), .RSTB(I300510), .Q(I300475) );
not I_17571 (I301105,I2357);
nand I_17572 (I301122,I378537,I378528);
and I_17573 (I301139,I301122,I378546);
DFFARX1 I_17574  ( .D(I301139), .CLK(I2350), .RSTB(I301105), .Q(I301156) );
nor I_17575 (I301173,I378543,I378528);
nor I_17576 (I301190,I301173,I301156);
not I_17577 (I301088,I301173);
DFFARX1 I_17578  ( .D(I378525), .CLK(I2350), .RSTB(I301105), .Q(I301221) );
not I_17579 (I301238,I301221);
nor I_17580 (I301255,I301173,I301238);
nand I_17581 (I301091,I301221,I301190);
DFFARX1 I_17582  ( .D(I301221), .CLK(I2350), .RSTB(I301105), .Q(I301073) );
nand I_17583 (I301300,I378534,I378549);
and I_17584 (I301317,I301300,I378540);
DFFARX1 I_17585  ( .D(I301317), .CLK(I2350), .RSTB(I301105), .Q(I301334) );
nor I_17586 (I301094,I301334,I301156);
nand I_17587 (I301085,I301334,I301255);
DFFARX1 I_17588  ( .D(I378522), .CLK(I2350), .RSTB(I301105), .Q(I301379) );
and I_17589 (I301396,I301379,I378531);
DFFARX1 I_17590  ( .D(I301396), .CLK(I2350), .RSTB(I301105), .Q(I301413) );
not I_17591 (I301076,I301413);
nand I_17592 (I301444,I301396,I301334);
and I_17593 (I301461,I301156,I301444);
DFFARX1 I_17594  ( .D(I301461), .CLK(I2350), .RSTB(I301105), .Q(I301067) );
DFFARX1 I_17595  ( .D(I378519), .CLK(I2350), .RSTB(I301105), .Q(I301492) );
nand I_17596 (I301509,I301492,I301156);
and I_17597 (I301526,I301334,I301509);
DFFARX1 I_17598  ( .D(I301526), .CLK(I2350), .RSTB(I301105), .Q(I301097) );
not I_17599 (I301557,I301492);
nor I_17600 (I301574,I301173,I301557);
and I_17601 (I301591,I301492,I301574);
or I_17602 (I301608,I301396,I301591);
DFFARX1 I_17603  ( .D(I301608), .CLK(I2350), .RSTB(I301105), .Q(I301082) );
nand I_17604 (I301079,I301492,I301238);
DFFARX1 I_17605  ( .D(I301492), .CLK(I2350), .RSTB(I301105), .Q(I301070) );
not I_17606 (I301700,I2357);
nand I_17607 (I301717,I124605,I124602);
and I_17608 (I301734,I301717,I124599);
DFFARX1 I_17609  ( .D(I301734), .CLK(I2350), .RSTB(I301700), .Q(I301751) );
nor I_17610 (I301768,I124590,I124602);
nor I_17611 (I301785,I301768,I301751);
not I_17612 (I301683,I301768);
DFFARX1 I_17613  ( .D(I124608), .CLK(I2350), .RSTB(I301700), .Q(I301816) );
not I_17614 (I301833,I301816);
nor I_17615 (I301850,I301768,I301833);
nand I_17616 (I301686,I301816,I301785);
DFFARX1 I_17617  ( .D(I301816), .CLK(I2350), .RSTB(I301700), .Q(I301668) );
nand I_17618 (I301895,I124593,I124617);
and I_17619 (I301912,I301895,I124596);
DFFARX1 I_17620  ( .D(I301912), .CLK(I2350), .RSTB(I301700), .Q(I301929) );
nor I_17621 (I301689,I301929,I301751);
nand I_17622 (I301680,I301929,I301850);
DFFARX1 I_17623  ( .D(I124614), .CLK(I2350), .RSTB(I301700), .Q(I301974) );
and I_17624 (I301991,I301974,I124611);
DFFARX1 I_17625  ( .D(I301991), .CLK(I2350), .RSTB(I301700), .Q(I302008) );
not I_17626 (I301671,I302008);
nand I_17627 (I302039,I301991,I301929);
and I_17628 (I302056,I301751,I302039);
DFFARX1 I_17629  ( .D(I302056), .CLK(I2350), .RSTB(I301700), .Q(I301662) );
DFFARX1 I_17630  ( .D(I124620), .CLK(I2350), .RSTB(I301700), .Q(I302087) );
nand I_17631 (I302104,I302087,I301751);
and I_17632 (I302121,I301929,I302104);
DFFARX1 I_17633  ( .D(I302121), .CLK(I2350), .RSTB(I301700), .Q(I301692) );
not I_17634 (I302152,I302087);
nor I_17635 (I302169,I301768,I302152);
and I_17636 (I302186,I302087,I302169);
or I_17637 (I302203,I301991,I302186);
DFFARX1 I_17638  ( .D(I302203), .CLK(I2350), .RSTB(I301700), .Q(I301677) );
nand I_17639 (I301674,I302087,I301833);
DFFARX1 I_17640  ( .D(I302087), .CLK(I2350), .RSTB(I301700), .Q(I301665) );
not I_17641 (I302295,I2357);
nand I_17642 (I302312,I11900,I11906);
and I_17643 (I302329,I302312,I11903);
DFFARX1 I_17644  ( .D(I302329), .CLK(I2350), .RSTB(I302295), .Q(I302346) );
nor I_17645 (I302363,I11927,I11906);
nor I_17646 (I302380,I302363,I302346);
not I_17647 (I302278,I302363);
DFFARX1 I_17648  ( .D(I11918), .CLK(I2350), .RSTB(I302295), .Q(I302411) );
not I_17649 (I302428,I302411);
nor I_17650 (I302445,I302363,I302428);
nand I_17651 (I302281,I302411,I302380);
DFFARX1 I_17652  ( .D(I302411), .CLK(I2350), .RSTB(I302295), .Q(I302263) );
nand I_17653 (I302490,I11921,I11924);
and I_17654 (I302507,I302490,I11897);
DFFARX1 I_17655  ( .D(I302507), .CLK(I2350), .RSTB(I302295), .Q(I302524) );
nor I_17656 (I302284,I302524,I302346);
nand I_17657 (I302275,I302524,I302445);
DFFARX1 I_17658  ( .D(I11915), .CLK(I2350), .RSTB(I302295), .Q(I302569) );
and I_17659 (I302586,I302569,I11909);
DFFARX1 I_17660  ( .D(I302586), .CLK(I2350), .RSTB(I302295), .Q(I302603) );
not I_17661 (I302266,I302603);
nand I_17662 (I302634,I302586,I302524);
and I_17663 (I302651,I302346,I302634);
DFFARX1 I_17664  ( .D(I302651), .CLK(I2350), .RSTB(I302295), .Q(I302257) );
DFFARX1 I_17665  ( .D(I11912), .CLK(I2350), .RSTB(I302295), .Q(I302682) );
nand I_17666 (I302699,I302682,I302346);
and I_17667 (I302716,I302524,I302699);
DFFARX1 I_17668  ( .D(I302716), .CLK(I2350), .RSTB(I302295), .Q(I302287) );
not I_17669 (I302747,I302682);
nor I_17670 (I302764,I302363,I302747);
and I_17671 (I302781,I302682,I302764);
or I_17672 (I302798,I302586,I302781);
DFFARX1 I_17673  ( .D(I302798), .CLK(I2350), .RSTB(I302295), .Q(I302272) );
nand I_17674 (I302269,I302682,I302428);
DFFARX1 I_17675  ( .D(I302682), .CLK(I2350), .RSTB(I302295), .Q(I302260) );
not I_17676 (I302890,I2357);
nand I_17677 (I302907,I220505,I220517);
and I_17678 (I302924,I302907,I220499);
DFFARX1 I_17679  ( .D(I302924), .CLK(I2350), .RSTB(I302890), .Q(I302941) );
nor I_17680 (I302958,I220511,I220517);
nor I_17681 (I302975,I302958,I302941);
not I_17682 (I302873,I302958);
DFFARX1 I_17683  ( .D(I220496), .CLK(I2350), .RSTB(I302890), .Q(I303006) );
not I_17684 (I303023,I303006);
nor I_17685 (I303040,I302958,I303023);
nand I_17686 (I302876,I303006,I302975);
DFFARX1 I_17687  ( .D(I303006), .CLK(I2350), .RSTB(I302890), .Q(I302858) );
nand I_17688 (I303085,I220487,I220502);
and I_17689 (I303102,I303085,I220493);
DFFARX1 I_17690  ( .D(I303102), .CLK(I2350), .RSTB(I302890), .Q(I303119) );
nor I_17691 (I302879,I303119,I302941);
nand I_17692 (I302870,I303119,I303040);
DFFARX1 I_17693  ( .D(I220514), .CLK(I2350), .RSTB(I302890), .Q(I303164) );
and I_17694 (I303181,I303164,I220508);
DFFARX1 I_17695  ( .D(I303181), .CLK(I2350), .RSTB(I302890), .Q(I303198) );
not I_17696 (I302861,I303198);
nand I_17697 (I303229,I303181,I303119);
and I_17698 (I303246,I302941,I303229);
DFFARX1 I_17699  ( .D(I303246), .CLK(I2350), .RSTB(I302890), .Q(I302852) );
DFFARX1 I_17700  ( .D(I220490), .CLK(I2350), .RSTB(I302890), .Q(I303277) );
nand I_17701 (I303294,I303277,I302941);
and I_17702 (I303311,I303119,I303294);
DFFARX1 I_17703  ( .D(I303311), .CLK(I2350), .RSTB(I302890), .Q(I302882) );
not I_17704 (I303342,I303277);
nor I_17705 (I303359,I302958,I303342);
and I_17706 (I303376,I303277,I303359);
or I_17707 (I303393,I303181,I303376);
DFFARX1 I_17708  ( .D(I303393), .CLK(I2350), .RSTB(I302890), .Q(I302867) );
nand I_17709 (I302864,I303277,I303023);
DFFARX1 I_17710  ( .D(I303277), .CLK(I2350), .RSTB(I302890), .Q(I302855) );
not I_17711 (I303485,I2357);
nand I_17712 (I303502,I72443,I72455);
and I_17713 (I303519,I303502,I72464);
DFFARX1 I_17714  ( .D(I303519), .CLK(I2350), .RSTB(I303485), .Q(I303536) );
nor I_17715 (I303553,I72458,I72455);
nor I_17716 (I303570,I303553,I303536);
not I_17717 (I303468,I303553);
DFFARX1 I_17718  ( .D(I72452), .CLK(I2350), .RSTB(I303485), .Q(I303601) );
not I_17719 (I303618,I303601);
nor I_17720 (I303635,I303553,I303618);
nand I_17721 (I303471,I303601,I303570);
DFFARX1 I_17722  ( .D(I303601), .CLK(I2350), .RSTB(I303485), .Q(I303453) );
nand I_17723 (I303680,I72449,I72446);
and I_17724 (I303697,I303680,I72437);
DFFARX1 I_17725  ( .D(I303697), .CLK(I2350), .RSTB(I303485), .Q(I303714) );
nor I_17726 (I303474,I303714,I303536);
nand I_17727 (I303465,I303714,I303635);
DFFARX1 I_17728  ( .D(I72461), .CLK(I2350), .RSTB(I303485), .Q(I303759) );
and I_17729 (I303776,I303759,I72440);
DFFARX1 I_17730  ( .D(I303776), .CLK(I2350), .RSTB(I303485), .Q(I303793) );
not I_17731 (I303456,I303793);
nand I_17732 (I303824,I303776,I303714);
and I_17733 (I303841,I303536,I303824);
DFFARX1 I_17734  ( .D(I303841), .CLK(I2350), .RSTB(I303485), .Q(I303447) );
DFFARX1 I_17735  ( .D(I72434), .CLK(I2350), .RSTB(I303485), .Q(I303872) );
nand I_17736 (I303889,I303872,I303536);
and I_17737 (I303906,I303714,I303889);
DFFARX1 I_17738  ( .D(I303906), .CLK(I2350), .RSTB(I303485), .Q(I303477) );
not I_17739 (I303937,I303872);
nor I_17740 (I303954,I303553,I303937);
and I_17741 (I303971,I303872,I303954);
or I_17742 (I303988,I303776,I303971);
DFFARX1 I_17743  ( .D(I303988), .CLK(I2350), .RSTB(I303485), .Q(I303462) );
nand I_17744 (I303459,I303872,I303618);
DFFARX1 I_17745  ( .D(I303872), .CLK(I2350), .RSTB(I303485), .Q(I303450) );
not I_17746 (I304080,I2357);
nand I_17747 (I304097,I185434,I185440);
and I_17748 (I304114,I304097,I185422);
DFFARX1 I_17749  ( .D(I304114), .CLK(I2350), .RSTB(I304080), .Q(I304131) );
nor I_17750 (I304148,I185416,I185440);
nor I_17751 (I304165,I304148,I304131);
not I_17752 (I304063,I304148);
DFFARX1 I_17753  ( .D(I185446), .CLK(I2350), .RSTB(I304080), .Q(I304196) );
not I_17754 (I304213,I304196);
nor I_17755 (I304230,I304148,I304213);
nand I_17756 (I304066,I304196,I304165);
DFFARX1 I_17757  ( .D(I304196), .CLK(I2350), .RSTB(I304080), .Q(I304048) );
nand I_17758 (I304275,I185437,I185428);
and I_17759 (I304292,I304275,I185431);
DFFARX1 I_17760  ( .D(I304292), .CLK(I2350), .RSTB(I304080), .Q(I304309) );
nor I_17761 (I304069,I304309,I304131);
nand I_17762 (I304060,I304309,I304230);
DFFARX1 I_17763  ( .D(I185443), .CLK(I2350), .RSTB(I304080), .Q(I304354) );
and I_17764 (I304371,I304354,I185419);
DFFARX1 I_17765  ( .D(I304371), .CLK(I2350), .RSTB(I304080), .Q(I304388) );
not I_17766 (I304051,I304388);
nand I_17767 (I304419,I304371,I304309);
and I_17768 (I304436,I304131,I304419);
DFFARX1 I_17769  ( .D(I304436), .CLK(I2350), .RSTB(I304080), .Q(I304042) );
DFFARX1 I_17770  ( .D(I185425), .CLK(I2350), .RSTB(I304080), .Q(I304467) );
nand I_17771 (I304484,I304467,I304131);
and I_17772 (I304501,I304309,I304484);
DFFARX1 I_17773  ( .D(I304501), .CLK(I2350), .RSTB(I304080), .Q(I304072) );
not I_17774 (I304532,I304467);
nor I_17775 (I304549,I304148,I304532);
and I_17776 (I304566,I304467,I304549);
or I_17777 (I304583,I304371,I304566);
DFFARX1 I_17778  ( .D(I304583), .CLK(I2350), .RSTB(I304080), .Q(I304057) );
nand I_17779 (I304054,I304467,I304213);
DFFARX1 I_17780  ( .D(I304467), .CLK(I2350), .RSTB(I304080), .Q(I304045) );
not I_17781 (I304675,I2357);
nand I_17782 (I304692,I369731,I369722);
and I_17783 (I304709,I304692,I369740);
DFFARX1 I_17784  ( .D(I304709), .CLK(I2350), .RSTB(I304675), .Q(I304726) );
nor I_17785 (I304743,I369737,I369722);
nor I_17786 (I304760,I304743,I304726);
not I_17787 (I304658,I304743);
DFFARX1 I_17788  ( .D(I369719), .CLK(I2350), .RSTB(I304675), .Q(I304791) );
not I_17789 (I304808,I304791);
nor I_17790 (I304825,I304743,I304808);
nand I_17791 (I304661,I304791,I304760);
DFFARX1 I_17792  ( .D(I304791), .CLK(I2350), .RSTB(I304675), .Q(I304643) );
nand I_17793 (I304870,I369728,I369743);
and I_17794 (I304887,I304870,I369734);
DFFARX1 I_17795  ( .D(I304887), .CLK(I2350), .RSTB(I304675), .Q(I304904) );
nor I_17796 (I304664,I304904,I304726);
nand I_17797 (I304655,I304904,I304825);
DFFARX1 I_17798  ( .D(I369716), .CLK(I2350), .RSTB(I304675), .Q(I304949) );
and I_17799 (I304966,I304949,I369725);
DFFARX1 I_17800  ( .D(I304966), .CLK(I2350), .RSTB(I304675), .Q(I304983) );
not I_17801 (I304646,I304983);
nand I_17802 (I305014,I304966,I304904);
and I_17803 (I305031,I304726,I305014);
DFFARX1 I_17804  ( .D(I305031), .CLK(I2350), .RSTB(I304675), .Q(I304637) );
DFFARX1 I_17805  ( .D(I369713), .CLK(I2350), .RSTB(I304675), .Q(I305062) );
nand I_17806 (I305079,I305062,I304726);
and I_17807 (I305096,I304904,I305079);
DFFARX1 I_17808  ( .D(I305096), .CLK(I2350), .RSTB(I304675), .Q(I304667) );
not I_17809 (I305127,I305062);
nor I_17810 (I305144,I304743,I305127);
and I_17811 (I305161,I305062,I305144);
or I_17812 (I305178,I304966,I305161);
DFFARX1 I_17813  ( .D(I305178), .CLK(I2350), .RSTB(I304675), .Q(I304652) );
nand I_17814 (I304649,I305062,I304808);
DFFARX1 I_17815  ( .D(I305062), .CLK(I2350), .RSTB(I304675), .Q(I304640) );
not I_17816 (I305270,I2357);
nand I_17817 (I305287,I46603,I46615);
and I_17818 (I305304,I305287,I46624);
DFFARX1 I_17819  ( .D(I305304), .CLK(I2350), .RSTB(I305270), .Q(I305321) );
nor I_17820 (I305338,I46618,I46615);
nor I_17821 (I305355,I305338,I305321);
not I_17822 (I305253,I305338);
DFFARX1 I_17823  ( .D(I46612), .CLK(I2350), .RSTB(I305270), .Q(I305386) );
not I_17824 (I305403,I305386);
nor I_17825 (I305420,I305338,I305403);
nand I_17826 (I305256,I305386,I305355);
DFFARX1 I_17827  ( .D(I305386), .CLK(I2350), .RSTB(I305270), .Q(I305238) );
nand I_17828 (I305465,I46609,I46606);
and I_17829 (I305482,I305465,I46597);
DFFARX1 I_17830  ( .D(I305482), .CLK(I2350), .RSTB(I305270), .Q(I305499) );
nor I_17831 (I305259,I305499,I305321);
nand I_17832 (I305250,I305499,I305420);
DFFARX1 I_17833  ( .D(I46621), .CLK(I2350), .RSTB(I305270), .Q(I305544) );
and I_17834 (I305561,I305544,I46600);
DFFARX1 I_17835  ( .D(I305561), .CLK(I2350), .RSTB(I305270), .Q(I305578) );
not I_17836 (I305241,I305578);
nand I_17837 (I305609,I305561,I305499);
and I_17838 (I305626,I305321,I305609);
DFFARX1 I_17839  ( .D(I305626), .CLK(I2350), .RSTB(I305270), .Q(I305232) );
DFFARX1 I_17840  ( .D(I46594), .CLK(I2350), .RSTB(I305270), .Q(I305657) );
nand I_17841 (I305674,I305657,I305321);
and I_17842 (I305691,I305499,I305674);
DFFARX1 I_17843  ( .D(I305691), .CLK(I2350), .RSTB(I305270), .Q(I305262) );
not I_17844 (I305722,I305657);
nor I_17845 (I305739,I305338,I305722);
and I_17846 (I305756,I305657,I305739);
or I_17847 (I305773,I305561,I305756);
DFFARX1 I_17848  ( .D(I305773), .CLK(I2350), .RSTB(I305270), .Q(I305247) );
nand I_17849 (I305244,I305657,I305403);
DFFARX1 I_17850  ( .D(I305657), .CLK(I2350), .RSTB(I305270), .Q(I305235) );
not I_17851 (I305865,I2357);
nand I_17852 (I305882,I60169,I60181);
and I_17853 (I305899,I305882,I60190);
DFFARX1 I_17854  ( .D(I305899), .CLK(I2350), .RSTB(I305865), .Q(I305916) );
nor I_17855 (I305933,I60184,I60181);
nor I_17856 (I305950,I305933,I305916);
not I_17857 (I305848,I305933);
DFFARX1 I_17858  ( .D(I60178), .CLK(I2350), .RSTB(I305865), .Q(I305981) );
not I_17859 (I305998,I305981);
nor I_17860 (I306015,I305933,I305998);
nand I_17861 (I305851,I305981,I305950);
DFFARX1 I_17862  ( .D(I305981), .CLK(I2350), .RSTB(I305865), .Q(I305833) );
nand I_17863 (I306060,I60175,I60172);
and I_17864 (I306077,I306060,I60163);
DFFARX1 I_17865  ( .D(I306077), .CLK(I2350), .RSTB(I305865), .Q(I306094) );
nor I_17866 (I305854,I306094,I305916);
nand I_17867 (I305845,I306094,I306015);
DFFARX1 I_17868  ( .D(I60187), .CLK(I2350), .RSTB(I305865), .Q(I306139) );
and I_17869 (I306156,I306139,I60166);
DFFARX1 I_17870  ( .D(I306156), .CLK(I2350), .RSTB(I305865), .Q(I306173) );
not I_17871 (I305836,I306173);
nand I_17872 (I306204,I306156,I306094);
and I_17873 (I306221,I305916,I306204);
DFFARX1 I_17874  ( .D(I306221), .CLK(I2350), .RSTB(I305865), .Q(I305827) );
DFFARX1 I_17875  ( .D(I60160), .CLK(I2350), .RSTB(I305865), .Q(I306252) );
nand I_17876 (I306269,I306252,I305916);
and I_17877 (I306286,I306094,I306269);
DFFARX1 I_17878  ( .D(I306286), .CLK(I2350), .RSTB(I305865), .Q(I305857) );
not I_17879 (I306317,I306252);
nor I_17880 (I306334,I305933,I306317);
and I_17881 (I306351,I306252,I306334);
or I_17882 (I306368,I306156,I306351);
DFFARX1 I_17883  ( .D(I306368), .CLK(I2350), .RSTB(I305865), .Q(I305842) );
nand I_17884 (I305839,I306252,I305998);
DFFARX1 I_17885  ( .D(I306252), .CLK(I2350), .RSTB(I305865), .Q(I305830) );
not I_17886 (I306460,I2357);
nand I_17887 (I306477,I40143,I40155);
and I_17888 (I306494,I306477,I40164);
DFFARX1 I_17889  ( .D(I306494), .CLK(I2350), .RSTB(I306460), .Q(I306511) );
nor I_17890 (I306528,I40158,I40155);
nor I_17891 (I306545,I306528,I306511);
not I_17892 (I306443,I306528);
DFFARX1 I_17893  ( .D(I40152), .CLK(I2350), .RSTB(I306460), .Q(I306576) );
not I_17894 (I306593,I306576);
nor I_17895 (I306610,I306528,I306593);
nand I_17896 (I306446,I306576,I306545);
DFFARX1 I_17897  ( .D(I306576), .CLK(I2350), .RSTB(I306460), .Q(I306428) );
nand I_17898 (I306655,I40149,I40146);
and I_17899 (I306672,I306655,I40137);
DFFARX1 I_17900  ( .D(I306672), .CLK(I2350), .RSTB(I306460), .Q(I306689) );
nor I_17901 (I306449,I306689,I306511);
nand I_17902 (I306440,I306689,I306610);
DFFARX1 I_17903  ( .D(I40161), .CLK(I2350), .RSTB(I306460), .Q(I306734) );
and I_17904 (I306751,I306734,I40140);
DFFARX1 I_17905  ( .D(I306751), .CLK(I2350), .RSTB(I306460), .Q(I306768) );
not I_17906 (I306431,I306768);
nand I_17907 (I306799,I306751,I306689);
and I_17908 (I306816,I306511,I306799);
DFFARX1 I_17909  ( .D(I306816), .CLK(I2350), .RSTB(I306460), .Q(I306422) );
DFFARX1 I_17910  ( .D(I40134), .CLK(I2350), .RSTB(I306460), .Q(I306847) );
nand I_17911 (I306864,I306847,I306511);
and I_17912 (I306881,I306689,I306864);
DFFARX1 I_17913  ( .D(I306881), .CLK(I2350), .RSTB(I306460), .Q(I306452) );
not I_17914 (I306912,I306847);
nor I_17915 (I306929,I306528,I306912);
and I_17916 (I306946,I306847,I306929);
or I_17917 (I306963,I306751,I306946);
DFFARX1 I_17918  ( .D(I306963), .CLK(I2350), .RSTB(I306460), .Q(I306437) );
nand I_17919 (I306434,I306847,I306593);
DFFARX1 I_17920  ( .D(I306847), .CLK(I2350), .RSTB(I306460), .Q(I306425) );
not I_17921 (I307055,I2357);
nand I_17922 (I307072,I339539,I339530);
and I_17923 (I307089,I307072,I339548);
DFFARX1 I_17924  ( .D(I307089), .CLK(I2350), .RSTB(I307055), .Q(I307106) );
nor I_17925 (I307123,I339545,I339530);
nor I_17926 (I307140,I307123,I307106);
not I_17927 (I307038,I307123);
DFFARX1 I_17928  ( .D(I339527), .CLK(I2350), .RSTB(I307055), .Q(I307171) );
not I_17929 (I307188,I307171);
nor I_17930 (I307205,I307123,I307188);
nand I_17931 (I307041,I307171,I307140);
DFFARX1 I_17932  ( .D(I307171), .CLK(I2350), .RSTB(I307055), .Q(I307023) );
nand I_17933 (I307250,I339536,I339551);
and I_17934 (I307267,I307250,I339542);
DFFARX1 I_17935  ( .D(I307267), .CLK(I2350), .RSTB(I307055), .Q(I307284) );
nor I_17936 (I307044,I307284,I307106);
nand I_17937 (I307035,I307284,I307205);
DFFARX1 I_17938  ( .D(I339524), .CLK(I2350), .RSTB(I307055), .Q(I307329) );
and I_17939 (I307346,I307329,I339533);
DFFARX1 I_17940  ( .D(I307346), .CLK(I2350), .RSTB(I307055), .Q(I307363) );
not I_17941 (I307026,I307363);
nand I_17942 (I307394,I307346,I307284);
and I_17943 (I307411,I307106,I307394);
DFFARX1 I_17944  ( .D(I307411), .CLK(I2350), .RSTB(I307055), .Q(I307017) );
DFFARX1 I_17945  ( .D(I339521), .CLK(I2350), .RSTB(I307055), .Q(I307442) );
nand I_17946 (I307459,I307442,I307106);
and I_17947 (I307476,I307284,I307459);
DFFARX1 I_17948  ( .D(I307476), .CLK(I2350), .RSTB(I307055), .Q(I307047) );
not I_17949 (I307507,I307442);
nor I_17950 (I307524,I307123,I307507);
and I_17951 (I307541,I307442,I307524);
or I_17952 (I307558,I307346,I307541);
DFFARX1 I_17953  ( .D(I307558), .CLK(I2350), .RSTB(I307055), .Q(I307032) );
nand I_17954 (I307029,I307442,I307188);
DFFARX1 I_17955  ( .D(I307442), .CLK(I2350), .RSTB(I307055), .Q(I307020) );
not I_17956 (I307650,I2357);
nand I_17957 (I307667,I184771,I184777);
and I_17958 (I307684,I307667,I184759);
DFFARX1 I_17959  ( .D(I307684), .CLK(I2350), .RSTB(I307650), .Q(I307701) );
nor I_17960 (I307718,I184753,I184777);
nor I_17961 (I307735,I307718,I307701);
not I_17962 (I307633,I307718);
DFFARX1 I_17963  ( .D(I184783), .CLK(I2350), .RSTB(I307650), .Q(I307766) );
not I_17964 (I307783,I307766);
nor I_17965 (I307800,I307718,I307783);
nand I_17966 (I307636,I307766,I307735);
DFFARX1 I_17967  ( .D(I307766), .CLK(I2350), .RSTB(I307650), .Q(I307618) );
nand I_17968 (I307845,I184774,I184765);
and I_17969 (I307862,I307845,I184768);
DFFARX1 I_17970  ( .D(I307862), .CLK(I2350), .RSTB(I307650), .Q(I307879) );
nor I_17971 (I307639,I307879,I307701);
nand I_17972 (I307630,I307879,I307800);
DFFARX1 I_17973  ( .D(I184780), .CLK(I2350), .RSTB(I307650), .Q(I307924) );
and I_17974 (I307941,I307924,I184756);
DFFARX1 I_17975  ( .D(I307941), .CLK(I2350), .RSTB(I307650), .Q(I307958) );
not I_17976 (I307621,I307958);
nand I_17977 (I307989,I307941,I307879);
and I_17978 (I308006,I307701,I307989);
DFFARX1 I_17979  ( .D(I308006), .CLK(I2350), .RSTB(I307650), .Q(I307612) );
DFFARX1 I_17980  ( .D(I184762), .CLK(I2350), .RSTB(I307650), .Q(I308037) );
nand I_17981 (I308054,I308037,I307701);
and I_17982 (I308071,I307879,I308054);
DFFARX1 I_17983  ( .D(I308071), .CLK(I2350), .RSTB(I307650), .Q(I307642) );
not I_17984 (I308102,I308037);
nor I_17985 (I308119,I307718,I308102);
and I_17986 (I308136,I308037,I308119);
or I_17987 (I308153,I307941,I308136);
DFFARX1 I_17988  ( .D(I308153), .CLK(I2350), .RSTB(I307650), .Q(I307627) );
nand I_17989 (I307624,I308037,I307783);
DFFARX1 I_17990  ( .D(I308037), .CLK(I2350), .RSTB(I307650), .Q(I307615) );
not I_17991 (I308245,I2357);
nand I_17992 (I308262,I97323,I97335);
and I_17993 (I308279,I308262,I97314);
DFFARX1 I_17994  ( .D(I308279), .CLK(I2350), .RSTB(I308245), .Q(I308296) );
nor I_17995 (I308313,I97305,I97335);
nor I_17996 (I308330,I308313,I308296);
not I_17997 (I308228,I308313);
DFFARX1 I_17998  ( .D(I97317), .CLK(I2350), .RSTB(I308245), .Q(I308361) );
not I_17999 (I308378,I308361);
nor I_18000 (I308395,I308313,I308378);
nand I_18001 (I308231,I308361,I308330);
DFFARX1 I_18002  ( .D(I308361), .CLK(I2350), .RSTB(I308245), .Q(I308213) );
nand I_18003 (I308440,I97332,I97320);
and I_18004 (I308457,I308440,I97308);
DFFARX1 I_18005  ( .D(I308457), .CLK(I2350), .RSTB(I308245), .Q(I308474) );
nor I_18006 (I308234,I308474,I308296);
nand I_18007 (I308225,I308474,I308395);
DFFARX1 I_18008  ( .D(I97326), .CLK(I2350), .RSTB(I308245), .Q(I308519) );
and I_18009 (I308536,I308519,I97311);
DFFARX1 I_18010  ( .D(I308536), .CLK(I2350), .RSTB(I308245), .Q(I308553) );
not I_18011 (I308216,I308553);
nand I_18012 (I308584,I308536,I308474);
and I_18013 (I308601,I308296,I308584);
DFFARX1 I_18014  ( .D(I308601), .CLK(I2350), .RSTB(I308245), .Q(I308207) );
DFFARX1 I_18015  ( .D(I97329), .CLK(I2350), .RSTB(I308245), .Q(I308632) );
nand I_18016 (I308649,I308632,I308296);
and I_18017 (I308666,I308474,I308649);
DFFARX1 I_18018  ( .D(I308666), .CLK(I2350), .RSTB(I308245), .Q(I308237) );
not I_18019 (I308697,I308632);
nor I_18020 (I308714,I308313,I308697);
and I_18021 (I308731,I308632,I308714);
or I_18022 (I308748,I308536,I308731);
DFFARX1 I_18023  ( .D(I308748), .CLK(I2350), .RSTB(I308245), .Q(I308222) );
nand I_18024 (I308219,I308632,I308378);
DFFARX1 I_18025  ( .D(I308632), .CLK(I2350), .RSTB(I308245), .Q(I308210) );
not I_18026 (I308840,I2357);
nand I_18027 (I308857,I262028,I262031);
and I_18028 (I308874,I308857,I262025);
DFFARX1 I_18029  ( .D(I308874), .CLK(I2350), .RSTB(I308840), .Q(I308891) );
nor I_18030 (I308908,I262022,I262031);
nor I_18031 (I308925,I308908,I308891);
not I_18032 (I308823,I308908);
DFFARX1 I_18033  ( .D(I262004), .CLK(I2350), .RSTB(I308840), .Q(I308956) );
not I_18034 (I308973,I308956);
nor I_18035 (I308990,I308908,I308973);
nand I_18036 (I308826,I308956,I308925);
DFFARX1 I_18037  ( .D(I308956), .CLK(I2350), .RSTB(I308840), .Q(I308808) );
nand I_18038 (I309035,I262013,I262010);
and I_18039 (I309052,I309035,I262019);
DFFARX1 I_18040  ( .D(I309052), .CLK(I2350), .RSTB(I308840), .Q(I309069) );
nor I_18041 (I308829,I309069,I308891);
nand I_18042 (I308820,I309069,I308990);
DFFARX1 I_18043  ( .D(I262001), .CLK(I2350), .RSTB(I308840), .Q(I309114) );
and I_18044 (I309131,I309114,I262016);
DFFARX1 I_18045  ( .D(I309131), .CLK(I2350), .RSTB(I308840), .Q(I309148) );
not I_18046 (I308811,I309148);
nand I_18047 (I309179,I309131,I309069);
and I_18048 (I309196,I308891,I309179);
DFFARX1 I_18049  ( .D(I309196), .CLK(I2350), .RSTB(I308840), .Q(I308802) );
DFFARX1 I_18050  ( .D(I262007), .CLK(I2350), .RSTB(I308840), .Q(I309227) );
nand I_18051 (I309244,I309227,I308891);
and I_18052 (I309261,I309069,I309244);
DFFARX1 I_18053  ( .D(I309261), .CLK(I2350), .RSTB(I308840), .Q(I308832) );
not I_18054 (I309292,I309227);
nor I_18055 (I309309,I308908,I309292);
and I_18056 (I309326,I309227,I309309);
or I_18057 (I309343,I309131,I309326);
DFFARX1 I_18058  ( .D(I309343), .CLK(I2350), .RSTB(I308840), .Q(I308817) );
nand I_18059 (I308814,I309227,I308973);
DFFARX1 I_18060  ( .D(I309227), .CLK(I2350), .RSTB(I308840), .Q(I308805) );
not I_18061 (I309435,I2357);
nand I_18062 (I309452,I1879,I1327);
and I_18063 (I309469,I309452,I1375);
DFFARX1 I_18064  ( .D(I309469), .CLK(I2350), .RSTB(I309435), .Q(I309486) );
nor I_18065 (I309503,I1551,I1327);
nor I_18066 (I309520,I309503,I309486);
not I_18067 (I309418,I309503);
DFFARX1 I_18068  ( .D(I1431), .CLK(I2350), .RSTB(I309435), .Q(I309551) );
not I_18069 (I309568,I309551);
nor I_18070 (I309585,I309503,I309568);
nand I_18071 (I309421,I309551,I309520);
DFFARX1 I_18072  ( .D(I309551), .CLK(I2350), .RSTB(I309435), .Q(I309403) );
nand I_18073 (I309630,I1871,I1607);
and I_18074 (I309647,I309630,I2055);
DFFARX1 I_18075  ( .D(I309647), .CLK(I2350), .RSTB(I309435), .Q(I309664) );
nor I_18076 (I309424,I309664,I309486);
nand I_18077 (I309415,I309664,I309585);
DFFARX1 I_18078  ( .D(I1239), .CLK(I2350), .RSTB(I309435), .Q(I309709) );
and I_18079 (I309726,I309709,I1767);
DFFARX1 I_18080  ( .D(I309726), .CLK(I2350), .RSTB(I309435), .Q(I309743) );
not I_18081 (I309406,I309743);
nand I_18082 (I309774,I309726,I309664);
and I_18083 (I309791,I309486,I309774);
DFFARX1 I_18084  ( .D(I309791), .CLK(I2350), .RSTB(I309435), .Q(I309397) );
DFFARX1 I_18085  ( .D(I1287), .CLK(I2350), .RSTB(I309435), .Q(I309822) );
nand I_18086 (I309839,I309822,I309486);
and I_18087 (I309856,I309664,I309839);
DFFARX1 I_18088  ( .D(I309856), .CLK(I2350), .RSTB(I309435), .Q(I309427) );
not I_18089 (I309887,I309822);
nor I_18090 (I309904,I309503,I309887);
and I_18091 (I309921,I309822,I309904);
or I_18092 (I309938,I309726,I309921);
DFFARX1 I_18093  ( .D(I309938), .CLK(I2350), .RSTB(I309435), .Q(I309412) );
nand I_18094 (I309409,I309822,I309568);
DFFARX1 I_18095  ( .D(I309822), .CLK(I2350), .RSTB(I309435), .Q(I309400) );
not I_18096 (I310030,I2357);
nand I_18097 (I310047,I43373,I43385);
and I_18098 (I310064,I310047,I43394);
DFFARX1 I_18099  ( .D(I310064), .CLK(I2350), .RSTB(I310030), .Q(I310081) );
nor I_18100 (I310098,I43388,I43385);
nor I_18101 (I310115,I310098,I310081);
not I_18102 (I310013,I310098);
DFFARX1 I_18103  ( .D(I43382), .CLK(I2350), .RSTB(I310030), .Q(I310146) );
not I_18104 (I310163,I310146);
nor I_18105 (I310180,I310098,I310163);
nand I_18106 (I310016,I310146,I310115);
DFFARX1 I_18107  ( .D(I310146), .CLK(I2350), .RSTB(I310030), .Q(I309998) );
nand I_18108 (I310225,I43379,I43376);
and I_18109 (I310242,I310225,I43367);
DFFARX1 I_18110  ( .D(I310242), .CLK(I2350), .RSTB(I310030), .Q(I310259) );
nor I_18111 (I310019,I310259,I310081);
nand I_18112 (I310010,I310259,I310180);
DFFARX1 I_18113  ( .D(I43391), .CLK(I2350), .RSTB(I310030), .Q(I310304) );
and I_18114 (I310321,I310304,I43370);
DFFARX1 I_18115  ( .D(I310321), .CLK(I2350), .RSTB(I310030), .Q(I310338) );
not I_18116 (I310001,I310338);
nand I_18117 (I310369,I310321,I310259);
and I_18118 (I310386,I310081,I310369);
DFFARX1 I_18119  ( .D(I310386), .CLK(I2350), .RSTB(I310030), .Q(I309992) );
DFFARX1 I_18120  ( .D(I43364), .CLK(I2350), .RSTB(I310030), .Q(I310417) );
nand I_18121 (I310434,I310417,I310081);
and I_18122 (I310451,I310259,I310434);
DFFARX1 I_18123  ( .D(I310451), .CLK(I2350), .RSTB(I310030), .Q(I310022) );
not I_18124 (I310482,I310417);
nor I_18125 (I310499,I310098,I310482);
and I_18126 (I310516,I310417,I310499);
or I_18127 (I310533,I310321,I310516);
DFFARX1 I_18128  ( .D(I310533), .CLK(I2350), .RSTB(I310030), .Q(I310007) );
nand I_18129 (I310004,I310417,I310163);
DFFARX1 I_18130  ( .D(I310417), .CLK(I2350), .RSTB(I310030), .Q(I309995) );
not I_18131 (I310625,I2357);
nand I_18132 (I310642,I235851,I235839);
and I_18133 (I310659,I310642,I235845);
DFFARX1 I_18134  ( .D(I310659), .CLK(I2350), .RSTB(I310625), .Q(I310676) );
nor I_18135 (I310693,I235836,I235839);
nor I_18136 (I310710,I310693,I310676);
not I_18137 (I310608,I310693);
DFFARX1 I_18138  ( .D(I235821), .CLK(I2350), .RSTB(I310625), .Q(I310741) );
not I_18139 (I310758,I310741);
nor I_18140 (I310775,I310693,I310758);
nand I_18141 (I310611,I310741,I310710);
DFFARX1 I_18142  ( .D(I310741), .CLK(I2350), .RSTB(I310625), .Q(I310593) );
nand I_18143 (I310820,I235830,I235848);
and I_18144 (I310837,I310820,I235842);
DFFARX1 I_18145  ( .D(I310837), .CLK(I2350), .RSTB(I310625), .Q(I310854) );
nor I_18146 (I310614,I310854,I310676);
nand I_18147 (I310605,I310854,I310775);
DFFARX1 I_18148  ( .D(I235833), .CLK(I2350), .RSTB(I310625), .Q(I310899) );
and I_18149 (I310916,I310899,I235827);
DFFARX1 I_18150  ( .D(I310916), .CLK(I2350), .RSTB(I310625), .Q(I310933) );
not I_18151 (I310596,I310933);
nand I_18152 (I310964,I310916,I310854);
and I_18153 (I310981,I310676,I310964);
DFFARX1 I_18154  ( .D(I310981), .CLK(I2350), .RSTB(I310625), .Q(I310587) );
DFFARX1 I_18155  ( .D(I235824), .CLK(I2350), .RSTB(I310625), .Q(I311012) );
nand I_18156 (I311029,I311012,I310676);
and I_18157 (I311046,I310854,I311029);
DFFARX1 I_18158  ( .D(I311046), .CLK(I2350), .RSTB(I310625), .Q(I310617) );
not I_18159 (I311077,I311012);
nor I_18160 (I311094,I310693,I311077);
and I_18161 (I311111,I311012,I311094);
or I_18162 (I311128,I310916,I311111);
DFFARX1 I_18163  ( .D(I311128), .CLK(I2350), .RSTB(I310625), .Q(I310602) );
nand I_18164 (I310599,I311012,I310758);
DFFARX1 I_18165  ( .D(I311012), .CLK(I2350), .RSTB(I310625), .Q(I310590) );
not I_18166 (I311220,I2357);
nand I_18167 (I311237,I109257,I109269);
and I_18168 (I311254,I311237,I109248);
DFFARX1 I_18169  ( .D(I311254), .CLK(I2350), .RSTB(I311220), .Q(I311271) );
nor I_18170 (I311288,I109239,I109269);
nor I_18171 (I311305,I311288,I311271);
not I_18172 (I311203,I311288);
DFFARX1 I_18173  ( .D(I109251), .CLK(I2350), .RSTB(I311220), .Q(I311336) );
not I_18174 (I311353,I311336);
nor I_18175 (I311370,I311288,I311353);
nand I_18176 (I311206,I311336,I311305);
DFFARX1 I_18177  ( .D(I311336), .CLK(I2350), .RSTB(I311220), .Q(I311188) );
nand I_18178 (I311415,I109266,I109254);
and I_18179 (I311432,I311415,I109242);
DFFARX1 I_18180  ( .D(I311432), .CLK(I2350), .RSTB(I311220), .Q(I311449) );
nor I_18181 (I311209,I311449,I311271);
nand I_18182 (I311200,I311449,I311370);
DFFARX1 I_18183  ( .D(I109260), .CLK(I2350), .RSTB(I311220), .Q(I311494) );
and I_18184 (I311511,I311494,I109245);
DFFARX1 I_18185  ( .D(I311511), .CLK(I2350), .RSTB(I311220), .Q(I311528) );
not I_18186 (I311191,I311528);
nand I_18187 (I311559,I311511,I311449);
and I_18188 (I311576,I311271,I311559);
DFFARX1 I_18189  ( .D(I311576), .CLK(I2350), .RSTB(I311220), .Q(I311182) );
DFFARX1 I_18190  ( .D(I109263), .CLK(I2350), .RSTB(I311220), .Q(I311607) );
nand I_18191 (I311624,I311607,I311271);
and I_18192 (I311641,I311449,I311624);
DFFARX1 I_18193  ( .D(I311641), .CLK(I2350), .RSTB(I311220), .Q(I311212) );
not I_18194 (I311672,I311607);
nor I_18195 (I311689,I311288,I311672);
and I_18196 (I311706,I311607,I311689);
or I_18197 (I311723,I311511,I311706);
DFFARX1 I_18198  ( .D(I311723), .CLK(I2350), .RSTB(I311220), .Q(I311197) );
nand I_18199 (I311194,I311607,I311353);
DFFARX1 I_18200  ( .D(I311607), .CLK(I2350), .RSTB(I311220), .Q(I311185) );
not I_18201 (I311815,I2357);
nand I_18202 (I311832,I330832,I330823);
and I_18203 (I311849,I311832,I330841);
DFFARX1 I_18204  ( .D(I311849), .CLK(I2350), .RSTB(I311815), .Q(I311866) );
nor I_18205 (I311883,I330820,I330823);
nor I_18206 (I311900,I311883,I311866);
not I_18207 (I311798,I311883);
DFFARX1 I_18208  ( .D(I330829), .CLK(I2350), .RSTB(I311815), .Q(I311931) );
not I_18209 (I311948,I311931);
nor I_18210 (I311965,I311883,I311948);
nand I_18211 (I311801,I311931,I311900);
DFFARX1 I_18212  ( .D(I311931), .CLK(I2350), .RSTB(I311815), .Q(I311783) );
nand I_18213 (I312010,I330844,I330826);
and I_18214 (I312027,I312010,I330847);
DFFARX1 I_18215  ( .D(I312027), .CLK(I2350), .RSTB(I311815), .Q(I312044) );
nor I_18216 (I311804,I312044,I311866);
nand I_18217 (I311795,I312044,I311965);
DFFARX1 I_18218  ( .D(I330835), .CLK(I2350), .RSTB(I311815), .Q(I312089) );
and I_18219 (I312106,I312089,I330817);
DFFARX1 I_18220  ( .D(I312106), .CLK(I2350), .RSTB(I311815), .Q(I312123) );
not I_18221 (I311786,I312123);
nand I_18222 (I312154,I312106,I312044);
and I_18223 (I312171,I311866,I312154);
DFFARX1 I_18224  ( .D(I312171), .CLK(I2350), .RSTB(I311815), .Q(I311777) );
DFFARX1 I_18225  ( .D(I330838), .CLK(I2350), .RSTB(I311815), .Q(I312202) );
nand I_18226 (I312219,I312202,I311866);
and I_18227 (I312236,I312044,I312219);
DFFARX1 I_18228  ( .D(I312236), .CLK(I2350), .RSTB(I311815), .Q(I311807) );
not I_18229 (I312267,I312202);
nor I_18230 (I312284,I311883,I312267);
and I_18231 (I312301,I312202,I312284);
or I_18232 (I312318,I312106,I312301);
DFFARX1 I_18233  ( .D(I312318), .CLK(I2350), .RSTB(I311815), .Q(I311792) );
nand I_18234 (I311789,I312202,I311948);
DFFARX1 I_18235  ( .D(I312202), .CLK(I2350), .RSTB(I311815), .Q(I311780) );
not I_18236 (I312410,I2357);
nand I_18237 (I312427,I100638,I100650);
and I_18238 (I312444,I312427,I100629);
DFFARX1 I_18239  ( .D(I312444), .CLK(I2350), .RSTB(I312410), .Q(I312461) );
nor I_18240 (I312478,I100620,I100650);
nor I_18241 (I312495,I312478,I312461);
not I_18242 (I312393,I312478);
DFFARX1 I_18243  ( .D(I100632), .CLK(I2350), .RSTB(I312410), .Q(I312526) );
not I_18244 (I312543,I312526);
nor I_18245 (I312560,I312478,I312543);
nand I_18246 (I312396,I312526,I312495);
DFFARX1 I_18247  ( .D(I312526), .CLK(I2350), .RSTB(I312410), .Q(I312378) );
nand I_18248 (I312605,I100647,I100635);
and I_18249 (I312622,I312605,I100623);
DFFARX1 I_18250  ( .D(I312622), .CLK(I2350), .RSTB(I312410), .Q(I312639) );
nor I_18251 (I312399,I312639,I312461);
nand I_18252 (I312390,I312639,I312560);
DFFARX1 I_18253  ( .D(I100641), .CLK(I2350), .RSTB(I312410), .Q(I312684) );
and I_18254 (I312701,I312684,I100626);
DFFARX1 I_18255  ( .D(I312701), .CLK(I2350), .RSTB(I312410), .Q(I312718) );
not I_18256 (I312381,I312718);
nand I_18257 (I312749,I312701,I312639);
and I_18258 (I312766,I312461,I312749);
DFFARX1 I_18259  ( .D(I312766), .CLK(I2350), .RSTB(I312410), .Q(I312372) );
DFFARX1 I_18260  ( .D(I100644), .CLK(I2350), .RSTB(I312410), .Q(I312797) );
nand I_18261 (I312814,I312797,I312461);
and I_18262 (I312831,I312639,I312814);
DFFARX1 I_18263  ( .D(I312831), .CLK(I2350), .RSTB(I312410), .Q(I312402) );
not I_18264 (I312862,I312797);
nor I_18265 (I312879,I312478,I312862);
and I_18266 (I312896,I312797,I312879);
or I_18267 (I312913,I312701,I312896);
DFFARX1 I_18268  ( .D(I312913), .CLK(I2350), .RSTB(I312410), .Q(I312387) );
nand I_18269 (I312384,I312797,I312543);
DFFARX1 I_18270  ( .D(I312797), .CLK(I2350), .RSTB(I312410), .Q(I312375) );
not I_18271 (I313005,I2357);
nand I_18272 (I313022,I275597,I275585);
and I_18273 (I313039,I313022,I275582);
DFFARX1 I_18274  ( .D(I313039), .CLK(I2350), .RSTB(I313005), .Q(I313056) );
nor I_18275 (I313073,I275576,I275585);
nor I_18276 (I313090,I313073,I313056);
not I_18277 (I312988,I313073);
DFFARX1 I_18278  ( .D(I275591), .CLK(I2350), .RSTB(I313005), .Q(I313121) );
not I_18279 (I313138,I313121);
nor I_18280 (I313155,I313073,I313138);
nand I_18281 (I312991,I313121,I313090);
DFFARX1 I_18282  ( .D(I313121), .CLK(I2350), .RSTB(I313005), .Q(I312973) );
nand I_18283 (I313200,I275588,I275594);
and I_18284 (I313217,I313200,I275579);
DFFARX1 I_18285  ( .D(I313217), .CLK(I2350), .RSTB(I313005), .Q(I313234) );
nor I_18286 (I312994,I313234,I313056);
nand I_18287 (I312985,I313234,I313155);
DFFARX1 I_18288  ( .D(I275567), .CLK(I2350), .RSTB(I313005), .Q(I313279) );
and I_18289 (I313296,I313279,I275570);
DFFARX1 I_18290  ( .D(I313296), .CLK(I2350), .RSTB(I313005), .Q(I313313) );
not I_18291 (I312976,I313313);
nand I_18292 (I313344,I313296,I313234);
and I_18293 (I313361,I313056,I313344);
DFFARX1 I_18294  ( .D(I313361), .CLK(I2350), .RSTB(I313005), .Q(I312967) );
DFFARX1 I_18295  ( .D(I275573), .CLK(I2350), .RSTB(I313005), .Q(I313392) );
nand I_18296 (I313409,I313392,I313056);
and I_18297 (I313426,I313234,I313409);
DFFARX1 I_18298  ( .D(I313426), .CLK(I2350), .RSTB(I313005), .Q(I312997) );
not I_18299 (I313457,I313392);
nor I_18300 (I313474,I313073,I313457);
and I_18301 (I313491,I313392,I313474);
or I_18302 (I313508,I313296,I313491);
DFFARX1 I_18303  ( .D(I313508), .CLK(I2350), .RSTB(I313005), .Q(I312982) );
nand I_18304 (I312979,I313392,I313138);
DFFARX1 I_18305  ( .D(I313392), .CLK(I2350), .RSTB(I313005), .Q(I312970) );
not I_18306 (I313600,I2357);
nand I_18307 (I313617,I113910,I113895);
and I_18308 (I313634,I313617,I113907);
DFFARX1 I_18309  ( .D(I313634), .CLK(I2350), .RSTB(I313600), .Q(I313651) );
nor I_18310 (I313668,I113898,I113895);
DFFARX1 I_18311  ( .D(I113889), .CLK(I2350), .RSTB(I313600), .Q(I313685) );
nand I_18312 (I313702,I313685,I313668);
DFFARX1 I_18313  ( .D(I313685), .CLK(I2350), .RSTB(I313600), .Q(I313571) );
nand I_18314 (I313733,I113880,I113904);
and I_18315 (I313750,I313733,I113883);
DFFARX1 I_18316  ( .D(I313750), .CLK(I2350), .RSTB(I313600), .Q(I313767) );
not I_18317 (I313784,I313767);
nor I_18318 (I313801,I313651,I313784);
and I_18319 (I313818,I313668,I313801);
and I_18320 (I313835,I313767,I313702);
DFFARX1 I_18321  ( .D(I313835), .CLK(I2350), .RSTB(I313600), .Q(I313568) );
DFFARX1 I_18322  ( .D(I313767), .CLK(I2350), .RSTB(I313600), .Q(I313562) );
DFFARX1 I_18323  ( .D(I113901), .CLK(I2350), .RSTB(I313600), .Q(I313880) );
and I_18324 (I313897,I313880,I113886);
nand I_18325 (I313914,I313897,I313767);
nor I_18326 (I313589,I313897,I313668);
not I_18327 (I313945,I313897);
nor I_18328 (I313962,I313651,I313945);
nand I_18329 (I313580,I313685,I313962);
nand I_18330 (I313574,I313767,I313945);
or I_18331 (I314007,I313897,I313818);
DFFARX1 I_18332  ( .D(I314007), .CLK(I2350), .RSTB(I313600), .Q(I313577) );
DFFARX1 I_18333  ( .D(I113892), .CLK(I2350), .RSTB(I313600), .Q(I314038) );
and I_18334 (I314055,I314038,I313914);
DFFARX1 I_18335  ( .D(I314055), .CLK(I2350), .RSTB(I313600), .Q(I313592) );
nor I_18336 (I314086,I314038,I313651);
nand I_18337 (I313586,I313897,I314086);
not I_18338 (I313583,I314038);
DFFARX1 I_18339  ( .D(I314038), .CLK(I2350), .RSTB(I313600), .Q(I314131) );
and I_18340 (I313565,I314038,I314131);
not I_18341 (I314195,I2357);
nand I_18342 (I314212,I118670,I118655);
and I_18343 (I314229,I314212,I118667);
DFFARX1 I_18344  ( .D(I314229), .CLK(I2350), .RSTB(I314195), .Q(I314246) );
nor I_18345 (I314263,I118658,I118655);
DFFARX1 I_18346  ( .D(I118649), .CLK(I2350), .RSTB(I314195), .Q(I314280) );
nand I_18347 (I314297,I314280,I314263);
DFFARX1 I_18348  ( .D(I314280), .CLK(I2350), .RSTB(I314195), .Q(I314166) );
nand I_18349 (I314328,I118640,I118664);
and I_18350 (I314345,I314328,I118643);
DFFARX1 I_18351  ( .D(I314345), .CLK(I2350), .RSTB(I314195), .Q(I314362) );
not I_18352 (I314379,I314362);
nor I_18353 (I314396,I314246,I314379);
and I_18354 (I314413,I314263,I314396);
and I_18355 (I314430,I314362,I314297);
DFFARX1 I_18356  ( .D(I314430), .CLK(I2350), .RSTB(I314195), .Q(I314163) );
DFFARX1 I_18357  ( .D(I314362), .CLK(I2350), .RSTB(I314195), .Q(I314157) );
DFFARX1 I_18358  ( .D(I118661), .CLK(I2350), .RSTB(I314195), .Q(I314475) );
and I_18359 (I314492,I314475,I118646);
nand I_18360 (I314509,I314492,I314362);
nor I_18361 (I314184,I314492,I314263);
not I_18362 (I314540,I314492);
nor I_18363 (I314557,I314246,I314540);
nand I_18364 (I314175,I314280,I314557);
nand I_18365 (I314169,I314362,I314540);
or I_18366 (I314602,I314492,I314413);
DFFARX1 I_18367  ( .D(I314602), .CLK(I2350), .RSTB(I314195), .Q(I314172) );
DFFARX1 I_18368  ( .D(I118652), .CLK(I2350), .RSTB(I314195), .Q(I314633) );
and I_18369 (I314650,I314633,I314509);
DFFARX1 I_18370  ( .D(I314650), .CLK(I2350), .RSTB(I314195), .Q(I314187) );
nor I_18371 (I314681,I314633,I314246);
nand I_18372 (I314181,I314492,I314681);
not I_18373 (I314178,I314633);
DFFARX1 I_18374  ( .D(I314633), .CLK(I2350), .RSTB(I314195), .Q(I314726) );
and I_18375 (I314160,I314633,I314726);
not I_18376 (I314790,I2357);
nand I_18377 (I314807,I219213,I219225);
and I_18378 (I314824,I314807,I219216);
DFFARX1 I_18379  ( .D(I314824), .CLK(I2350), .RSTB(I314790), .Q(I314841) );
nor I_18380 (I314858,I219210,I219225);
DFFARX1 I_18381  ( .D(I219201), .CLK(I2350), .RSTB(I314790), .Q(I314875) );
nand I_18382 (I314892,I314875,I314858);
DFFARX1 I_18383  ( .D(I314875), .CLK(I2350), .RSTB(I314790), .Q(I314761) );
nand I_18384 (I314923,I219207,I219198);
and I_18385 (I314940,I314923,I219204);
DFFARX1 I_18386  ( .D(I314940), .CLK(I2350), .RSTB(I314790), .Q(I314957) );
not I_18387 (I314974,I314957);
nor I_18388 (I314991,I314841,I314974);
and I_18389 (I315008,I314858,I314991);
and I_18390 (I315025,I314957,I314892);
DFFARX1 I_18391  ( .D(I315025), .CLK(I2350), .RSTB(I314790), .Q(I314758) );
DFFARX1 I_18392  ( .D(I314957), .CLK(I2350), .RSTB(I314790), .Q(I314752) );
DFFARX1 I_18393  ( .D(I219219), .CLK(I2350), .RSTB(I314790), .Q(I315070) );
and I_18394 (I315087,I315070,I219195);
nand I_18395 (I315104,I315087,I314957);
nor I_18396 (I314779,I315087,I314858);
not I_18397 (I315135,I315087);
nor I_18398 (I315152,I314841,I315135);
nand I_18399 (I314770,I314875,I315152);
nand I_18400 (I314764,I314957,I315135);
or I_18401 (I315197,I315087,I315008);
DFFARX1 I_18402  ( .D(I315197), .CLK(I2350), .RSTB(I314790), .Q(I314767) );
DFFARX1 I_18403  ( .D(I219222), .CLK(I2350), .RSTB(I314790), .Q(I315228) );
and I_18404 (I315245,I315228,I315104);
DFFARX1 I_18405  ( .D(I315245), .CLK(I2350), .RSTB(I314790), .Q(I314782) );
nor I_18406 (I315276,I315228,I314841);
nand I_18407 (I314776,I315087,I315276);
not I_18408 (I314773,I315228);
DFFARX1 I_18409  ( .D(I315228), .CLK(I2350), .RSTB(I314790), .Q(I315321) );
and I_18410 (I314755,I315228,I315321);
not I_18411 (I315385,I2357);
nand I_18412 (I315402,I66001,I65977);
and I_18413 (I315419,I315402,I65986);
DFFARX1 I_18414  ( .D(I315419), .CLK(I2350), .RSTB(I315385), .Q(I315436) );
nor I_18415 (I315453,I65980,I65977);
DFFARX1 I_18416  ( .D(I65995), .CLK(I2350), .RSTB(I315385), .Q(I315470) );
nand I_18417 (I315487,I315470,I315453);
DFFARX1 I_18418  ( .D(I315470), .CLK(I2350), .RSTB(I315385), .Q(I315356) );
nand I_18419 (I315518,I65989,I66004);
and I_18420 (I315535,I315518,I65983);
DFFARX1 I_18421  ( .D(I315535), .CLK(I2350), .RSTB(I315385), .Q(I315552) );
not I_18422 (I315569,I315552);
nor I_18423 (I315586,I315436,I315569);
and I_18424 (I315603,I315453,I315586);
and I_18425 (I315620,I315552,I315487);
DFFARX1 I_18426  ( .D(I315620), .CLK(I2350), .RSTB(I315385), .Q(I315353) );
DFFARX1 I_18427  ( .D(I315552), .CLK(I2350), .RSTB(I315385), .Q(I315347) );
DFFARX1 I_18428  ( .D(I65974), .CLK(I2350), .RSTB(I315385), .Q(I315665) );
and I_18429 (I315682,I315665,I65992);
nand I_18430 (I315699,I315682,I315552);
nor I_18431 (I315374,I315682,I315453);
not I_18432 (I315730,I315682);
nor I_18433 (I315747,I315436,I315730);
nand I_18434 (I315365,I315470,I315747);
nand I_18435 (I315359,I315552,I315730);
or I_18436 (I315792,I315682,I315603);
DFFARX1 I_18437  ( .D(I315792), .CLK(I2350), .RSTB(I315385), .Q(I315362) );
DFFARX1 I_18438  ( .D(I65998), .CLK(I2350), .RSTB(I315385), .Q(I315823) );
and I_18439 (I315840,I315823,I315699);
DFFARX1 I_18440  ( .D(I315840), .CLK(I2350), .RSTB(I315385), .Q(I315377) );
nor I_18441 (I315871,I315823,I315436);
nand I_18442 (I315371,I315682,I315871);
not I_18443 (I315368,I315823);
DFFARX1 I_18444  ( .D(I315823), .CLK(I2350), .RSTB(I315385), .Q(I315916) );
and I_18445 (I315350,I315823,I315916);
not I_18446 (I315980,I2357);
nand I_18447 (I315997,I367856,I367844);
and I_18448 (I316014,I315997,I367829);
DFFARX1 I_18449  ( .D(I316014), .CLK(I2350), .RSTB(I315980), .Q(I316031) );
nor I_18450 (I316048,I367841,I367844);
DFFARX1 I_18451  ( .D(I367853), .CLK(I2350), .RSTB(I315980), .Q(I316065) );
nand I_18452 (I316082,I316065,I316048);
DFFARX1 I_18453  ( .D(I316065), .CLK(I2350), .RSTB(I315980), .Q(I315951) );
nand I_18454 (I316113,I367826,I367850);
and I_18455 (I316130,I316113,I367835);
DFFARX1 I_18456  ( .D(I316130), .CLK(I2350), .RSTB(I315980), .Q(I316147) );
not I_18457 (I316164,I316147);
nor I_18458 (I316181,I316031,I316164);
and I_18459 (I316198,I316048,I316181);
and I_18460 (I316215,I316147,I316082);
DFFARX1 I_18461  ( .D(I316215), .CLK(I2350), .RSTB(I315980), .Q(I315948) );
DFFARX1 I_18462  ( .D(I316147), .CLK(I2350), .RSTB(I315980), .Q(I315942) );
DFFARX1 I_18463  ( .D(I367838), .CLK(I2350), .RSTB(I315980), .Q(I316260) );
and I_18464 (I316277,I316260,I367847);
nand I_18465 (I316294,I316277,I316147);
nor I_18466 (I315969,I316277,I316048);
not I_18467 (I316325,I316277);
nor I_18468 (I316342,I316031,I316325);
nand I_18469 (I315960,I316065,I316342);
nand I_18470 (I315954,I316147,I316325);
or I_18471 (I316387,I316277,I316198);
DFFARX1 I_18472  ( .D(I316387), .CLK(I2350), .RSTB(I315980), .Q(I315957) );
DFFARX1 I_18473  ( .D(I367832), .CLK(I2350), .RSTB(I315980), .Q(I316418) );
and I_18474 (I316435,I316418,I316294);
DFFARX1 I_18475  ( .D(I316435), .CLK(I2350), .RSTB(I315980), .Q(I315972) );
nor I_18476 (I316466,I316418,I316031);
nand I_18477 (I315966,I316277,I316466);
not I_18478 (I315963,I316418);
DFFARX1 I_18479  ( .D(I316418), .CLK(I2350), .RSTB(I315980), .Q(I316511) );
and I_18480 (I315945,I316418,I316511);
not I_18481 (I316575,I2357);
nand I_18482 (I316592,I289182,I289167);
and I_18483 (I316609,I316592,I289173);
DFFARX1 I_18484  ( .D(I316609), .CLK(I2350), .RSTB(I316575), .Q(I316626) );
nor I_18485 (I316643,I289176,I289167);
DFFARX1 I_18486  ( .D(I289188), .CLK(I2350), .RSTB(I316575), .Q(I316660) );
nand I_18487 (I316677,I316660,I316643);
DFFARX1 I_18488  ( .D(I316660), .CLK(I2350), .RSTB(I316575), .Q(I316546) );
nand I_18489 (I316708,I289179,I289170);
and I_18490 (I316725,I316708,I289197);
DFFARX1 I_18491  ( .D(I316725), .CLK(I2350), .RSTB(I316575), .Q(I316742) );
not I_18492 (I316759,I316742);
nor I_18493 (I316776,I316626,I316759);
and I_18494 (I316793,I316643,I316776);
and I_18495 (I316810,I316742,I316677);
DFFARX1 I_18496  ( .D(I316810), .CLK(I2350), .RSTB(I316575), .Q(I316543) );
DFFARX1 I_18497  ( .D(I316742), .CLK(I2350), .RSTB(I316575), .Q(I316537) );
DFFARX1 I_18498  ( .D(I289185), .CLK(I2350), .RSTB(I316575), .Q(I316855) );
and I_18499 (I316872,I316855,I289191);
nand I_18500 (I316889,I316872,I316742);
nor I_18501 (I316564,I316872,I316643);
not I_18502 (I316920,I316872);
nor I_18503 (I316937,I316626,I316920);
nand I_18504 (I316555,I316660,I316937);
nand I_18505 (I316549,I316742,I316920);
or I_18506 (I316982,I316872,I316793);
DFFARX1 I_18507  ( .D(I316982), .CLK(I2350), .RSTB(I316575), .Q(I316552) );
DFFARX1 I_18508  ( .D(I289194), .CLK(I2350), .RSTB(I316575), .Q(I317013) );
and I_18509 (I317030,I317013,I316889);
DFFARX1 I_18510  ( .D(I317030), .CLK(I2350), .RSTB(I316575), .Q(I316567) );
nor I_18511 (I317061,I317013,I316626);
nand I_18512 (I316561,I316872,I317061);
not I_18513 (I316558,I317013);
DFFARX1 I_18514  ( .D(I317013), .CLK(I2350), .RSTB(I316575), .Q(I317106) );
and I_18515 (I316540,I317013,I317106);
not I_18516 (I317170,I2357);
nand I_18517 (I317187,I181468,I181438);
and I_18518 (I317204,I317187,I181456);
DFFARX1 I_18519  ( .D(I317204), .CLK(I2350), .RSTB(I317170), .Q(I317221) );
nor I_18520 (I317238,I181450,I181438);
DFFARX1 I_18521  ( .D(I181447), .CLK(I2350), .RSTB(I317170), .Q(I317255) );
nand I_18522 (I317272,I317255,I317238);
DFFARX1 I_18523  ( .D(I317255), .CLK(I2350), .RSTB(I317170), .Q(I317141) );
nand I_18524 (I317303,I181441,I181444);
and I_18525 (I317320,I317303,I181462);
DFFARX1 I_18526  ( .D(I317320), .CLK(I2350), .RSTB(I317170), .Q(I317337) );
not I_18527 (I317354,I317337);
nor I_18528 (I317371,I317221,I317354);
and I_18529 (I317388,I317238,I317371);
and I_18530 (I317405,I317337,I317272);
DFFARX1 I_18531  ( .D(I317405), .CLK(I2350), .RSTB(I317170), .Q(I317138) );
DFFARX1 I_18532  ( .D(I317337), .CLK(I2350), .RSTB(I317170), .Q(I317132) );
DFFARX1 I_18533  ( .D(I181465), .CLK(I2350), .RSTB(I317170), .Q(I317450) );
and I_18534 (I317467,I317450,I181459);
nand I_18535 (I317484,I317467,I317337);
nor I_18536 (I317159,I317467,I317238);
not I_18537 (I317515,I317467);
nor I_18538 (I317532,I317221,I317515);
nand I_18539 (I317150,I317255,I317532);
nand I_18540 (I317144,I317337,I317515);
or I_18541 (I317577,I317467,I317388);
DFFARX1 I_18542  ( .D(I317577), .CLK(I2350), .RSTB(I317170), .Q(I317147) );
DFFARX1 I_18543  ( .D(I181453), .CLK(I2350), .RSTB(I317170), .Q(I317608) );
and I_18544 (I317625,I317608,I317484);
DFFARX1 I_18545  ( .D(I317625), .CLK(I2350), .RSTB(I317170), .Q(I317162) );
nor I_18546 (I317656,I317608,I317221);
nand I_18547 (I317156,I317467,I317656);
not I_18548 (I317153,I317608);
DFFARX1 I_18549  ( .D(I317608), .CLK(I2350), .RSTB(I317170), .Q(I317701) );
and I_18550 (I317135,I317608,I317701);
not I_18551 (I317765,I2357);
nand I_18552 (I317782,I9656,I9671);
and I_18553 (I317799,I317782,I9677);
DFFARX1 I_18554  ( .D(I317799), .CLK(I2350), .RSTB(I317765), .Q(I317816) );
nor I_18555 (I317833,I9665,I9671);
DFFARX1 I_18556  ( .D(I9653), .CLK(I2350), .RSTB(I317765), .Q(I317850) );
nand I_18557 (I317867,I317850,I317833);
DFFARX1 I_18558  ( .D(I317850), .CLK(I2350), .RSTB(I317765), .Q(I317736) );
nand I_18559 (I317898,I9659,I9662);
and I_18560 (I317915,I317898,I9668);
DFFARX1 I_18561  ( .D(I317915), .CLK(I2350), .RSTB(I317765), .Q(I317932) );
not I_18562 (I317949,I317932);
nor I_18563 (I317966,I317816,I317949);
and I_18564 (I317983,I317833,I317966);
and I_18565 (I318000,I317932,I317867);
DFFARX1 I_18566  ( .D(I318000), .CLK(I2350), .RSTB(I317765), .Q(I317733) );
DFFARX1 I_18567  ( .D(I317932), .CLK(I2350), .RSTB(I317765), .Q(I317727) );
DFFARX1 I_18568  ( .D(I9674), .CLK(I2350), .RSTB(I317765), .Q(I318045) );
and I_18569 (I318062,I318045,I9683);
nand I_18570 (I318079,I318062,I317932);
nor I_18571 (I317754,I318062,I317833);
not I_18572 (I318110,I318062);
nor I_18573 (I318127,I317816,I318110);
nand I_18574 (I317745,I317850,I318127);
nand I_18575 (I317739,I317932,I318110);
or I_18576 (I318172,I318062,I317983);
DFFARX1 I_18577  ( .D(I318172), .CLK(I2350), .RSTB(I317765), .Q(I317742) );
DFFARX1 I_18578  ( .D(I9680), .CLK(I2350), .RSTB(I317765), .Q(I318203) );
and I_18579 (I318220,I318203,I318079);
DFFARX1 I_18580  ( .D(I318220), .CLK(I2350), .RSTB(I317765), .Q(I317757) );
nor I_18581 (I318251,I318203,I317816);
nand I_18582 (I317751,I318062,I318251);
not I_18583 (I317748,I318203);
DFFARX1 I_18584  ( .D(I318203), .CLK(I2350), .RSTB(I317765), .Q(I318296) );
and I_18585 (I317730,I318203,I318296);
not I_18586 (I318360,I2357);
nand I_18587 (I318377,I223735,I223747);
and I_18588 (I318394,I318377,I223738);
DFFARX1 I_18589  ( .D(I318394), .CLK(I2350), .RSTB(I318360), .Q(I318411) );
nor I_18590 (I318428,I223732,I223747);
DFFARX1 I_18591  ( .D(I223723), .CLK(I2350), .RSTB(I318360), .Q(I318445) );
nand I_18592 (I318462,I318445,I318428);
DFFARX1 I_18593  ( .D(I318445), .CLK(I2350), .RSTB(I318360), .Q(I318331) );
nand I_18594 (I318493,I223729,I223720);
and I_18595 (I318510,I318493,I223726);
DFFARX1 I_18596  ( .D(I318510), .CLK(I2350), .RSTB(I318360), .Q(I318527) );
not I_18597 (I318544,I318527);
nor I_18598 (I318561,I318411,I318544);
and I_18599 (I318578,I318428,I318561);
and I_18600 (I318595,I318527,I318462);
DFFARX1 I_18601  ( .D(I318595), .CLK(I2350), .RSTB(I318360), .Q(I318328) );
DFFARX1 I_18602  ( .D(I318527), .CLK(I2350), .RSTB(I318360), .Q(I318322) );
DFFARX1 I_18603  ( .D(I223741), .CLK(I2350), .RSTB(I318360), .Q(I318640) );
and I_18604 (I318657,I318640,I223717);
nand I_18605 (I318674,I318657,I318527);
nor I_18606 (I318349,I318657,I318428);
not I_18607 (I318705,I318657);
nor I_18608 (I318722,I318411,I318705);
nand I_18609 (I318340,I318445,I318722);
nand I_18610 (I318334,I318527,I318705);
or I_18611 (I318767,I318657,I318578);
DFFARX1 I_18612  ( .D(I318767), .CLK(I2350), .RSTB(I318360), .Q(I318337) );
DFFARX1 I_18613  ( .D(I223744), .CLK(I2350), .RSTB(I318360), .Q(I318798) );
and I_18614 (I318815,I318798,I318674);
DFFARX1 I_18615  ( .D(I318815), .CLK(I2350), .RSTB(I318360), .Q(I318352) );
nor I_18616 (I318846,I318798,I318411);
nand I_18617 (I318346,I318657,I318846);
not I_18618 (I318343,I318798);
DFFARX1 I_18619  ( .D(I318798), .CLK(I2350), .RSTB(I318360), .Q(I318891) );
and I_18620 (I318325,I318798,I318891);
not I_18621 (I318955,I2357);
nand I_18622 (I318972,I397219,I397222);
and I_18623 (I318989,I318972,I397231);
DFFARX1 I_18624  ( .D(I318989), .CLK(I2350), .RSTB(I318955), .Q(I319006) );
nor I_18625 (I319023,I397225,I397222);
DFFARX1 I_18626  ( .D(I397246), .CLK(I2350), .RSTB(I318955), .Q(I319040) );
nand I_18627 (I319057,I319040,I319023);
DFFARX1 I_18628  ( .D(I319040), .CLK(I2350), .RSTB(I318955), .Q(I318926) );
nand I_18629 (I319088,I397243,I397249);
and I_18630 (I319105,I319088,I397234);
DFFARX1 I_18631  ( .D(I319105), .CLK(I2350), .RSTB(I318955), .Q(I319122) );
not I_18632 (I319139,I319122);
nor I_18633 (I319156,I319006,I319139);
and I_18634 (I319173,I319023,I319156);
and I_18635 (I319190,I319122,I319057);
DFFARX1 I_18636  ( .D(I319190), .CLK(I2350), .RSTB(I318955), .Q(I318923) );
DFFARX1 I_18637  ( .D(I319122), .CLK(I2350), .RSTB(I318955), .Q(I318917) );
DFFARX1 I_18638  ( .D(I397237), .CLK(I2350), .RSTB(I318955), .Q(I319235) );
and I_18639 (I319252,I319235,I397240);
nand I_18640 (I319269,I319252,I319122);
nor I_18641 (I318944,I319252,I319023);
not I_18642 (I319300,I319252);
nor I_18643 (I319317,I319006,I319300);
nand I_18644 (I318935,I319040,I319317);
nand I_18645 (I318929,I319122,I319300);
or I_18646 (I319362,I319252,I319173);
DFFARX1 I_18647  ( .D(I319362), .CLK(I2350), .RSTB(I318955), .Q(I318932) );
DFFARX1 I_18648  ( .D(I397228), .CLK(I2350), .RSTB(I318955), .Q(I319393) );
and I_18649 (I319410,I319393,I319269);
DFFARX1 I_18650  ( .D(I319410), .CLK(I2350), .RSTB(I318955), .Q(I318947) );
nor I_18651 (I319441,I319393,I319006);
nand I_18652 (I318941,I319252,I319441);
not I_18653 (I318938,I319393);
DFFARX1 I_18654  ( .D(I319393), .CLK(I2350), .RSTB(I318955), .Q(I319486) );
and I_18655 (I318920,I319393,I319486);
not I_18656 (I319550,I2357);
nand I_18657 (I319567,I129948,I129945);
and I_18658 (I319584,I319567,I129972);
DFFARX1 I_18659  ( .D(I319584), .CLK(I2350), .RSTB(I319550), .Q(I319601) );
nor I_18660 (I319618,I129975,I129945);
DFFARX1 I_18661  ( .D(I129963), .CLK(I2350), .RSTB(I319550), .Q(I319635) );
nand I_18662 (I319652,I319635,I319618);
DFFARX1 I_18663  ( .D(I319635), .CLK(I2350), .RSTB(I319550), .Q(I319521) );
nand I_18664 (I319683,I129969,I129954);
and I_18665 (I319700,I319683,I129960);
DFFARX1 I_18666  ( .D(I319700), .CLK(I2350), .RSTB(I319550), .Q(I319717) );
not I_18667 (I319734,I319717);
nor I_18668 (I319751,I319601,I319734);
and I_18669 (I319768,I319618,I319751);
and I_18670 (I319785,I319717,I319652);
DFFARX1 I_18671  ( .D(I319785), .CLK(I2350), .RSTB(I319550), .Q(I319518) );
DFFARX1 I_18672  ( .D(I319717), .CLK(I2350), .RSTB(I319550), .Q(I319512) );
DFFARX1 I_18673  ( .D(I129951), .CLK(I2350), .RSTB(I319550), .Q(I319830) );
and I_18674 (I319847,I319830,I129957);
nand I_18675 (I319864,I319847,I319717);
nor I_18676 (I319539,I319847,I319618);
not I_18677 (I319895,I319847);
nor I_18678 (I319912,I319601,I319895);
nand I_18679 (I319530,I319635,I319912);
nand I_18680 (I319524,I319717,I319895);
or I_18681 (I319957,I319847,I319768);
DFFARX1 I_18682  ( .D(I319957), .CLK(I2350), .RSTB(I319550), .Q(I319527) );
DFFARX1 I_18683  ( .D(I129966), .CLK(I2350), .RSTB(I319550), .Q(I319988) );
and I_18684 (I320005,I319988,I319864);
DFFARX1 I_18685  ( .D(I320005), .CLK(I2350), .RSTB(I319550), .Q(I319542) );
nor I_18686 (I320036,I319988,I319601);
nand I_18687 (I319536,I319847,I320036);
not I_18688 (I319533,I319988);
DFFARX1 I_18689  ( .D(I319988), .CLK(I2350), .RSTB(I319550), .Q(I320081) );
and I_18690 (I319515,I319988,I320081);
not I_18691 (I320145,I2357);
nand I_18692 (I320162,I250453,I250468);
and I_18693 (I320179,I320162,I250465);
DFFARX1 I_18694  ( .D(I320179), .CLK(I2350), .RSTB(I320145), .Q(I320196) );
nor I_18695 (I320213,I250441,I250468);
DFFARX1 I_18696  ( .D(I250459), .CLK(I2350), .RSTB(I320145), .Q(I320230) );
nand I_18697 (I320247,I320230,I320213);
DFFARX1 I_18698  ( .D(I320230), .CLK(I2350), .RSTB(I320145), .Q(I320116) );
nand I_18699 (I320278,I250462,I250450);
and I_18700 (I320295,I320278,I250456);
DFFARX1 I_18701  ( .D(I320295), .CLK(I2350), .RSTB(I320145), .Q(I320312) );
not I_18702 (I320329,I320312);
nor I_18703 (I320346,I320196,I320329);
and I_18704 (I320363,I320213,I320346);
and I_18705 (I320380,I320312,I320247);
DFFARX1 I_18706  ( .D(I320380), .CLK(I2350), .RSTB(I320145), .Q(I320113) );
DFFARX1 I_18707  ( .D(I320312), .CLK(I2350), .RSTB(I320145), .Q(I320107) );
DFFARX1 I_18708  ( .D(I250447), .CLK(I2350), .RSTB(I320145), .Q(I320425) );
and I_18709 (I320442,I320425,I250471);
nand I_18710 (I320459,I320442,I320312);
nor I_18711 (I320134,I320442,I320213);
not I_18712 (I320490,I320442);
nor I_18713 (I320507,I320196,I320490);
nand I_18714 (I320125,I320230,I320507);
nand I_18715 (I320119,I320312,I320490);
or I_18716 (I320552,I320442,I320363);
DFFARX1 I_18717  ( .D(I320552), .CLK(I2350), .RSTB(I320145), .Q(I320122) );
DFFARX1 I_18718  ( .D(I250444), .CLK(I2350), .RSTB(I320145), .Q(I320583) );
and I_18719 (I320600,I320583,I320459);
DFFARX1 I_18720  ( .D(I320600), .CLK(I2350), .RSTB(I320145), .Q(I320137) );
nor I_18721 (I320631,I320583,I320196);
nand I_18722 (I320131,I320442,I320631);
not I_18723 (I320128,I320583);
DFFARX1 I_18724  ( .D(I320583), .CLK(I2350), .RSTB(I320145), .Q(I320676) );
and I_18725 (I320110,I320583,I320676);
not I_18726 (I320740,I2357);
nand I_18727 (I320757,I130543,I130540);
and I_18728 (I320774,I320757,I130567);
DFFARX1 I_18729  ( .D(I320774), .CLK(I2350), .RSTB(I320740), .Q(I320791) );
nor I_18730 (I320808,I130570,I130540);
DFFARX1 I_18731  ( .D(I130558), .CLK(I2350), .RSTB(I320740), .Q(I320825) );
nand I_18732 (I320842,I320825,I320808);
DFFARX1 I_18733  ( .D(I320825), .CLK(I2350), .RSTB(I320740), .Q(I320711) );
nand I_18734 (I320873,I130564,I130549);
and I_18735 (I320890,I320873,I130555);
DFFARX1 I_18736  ( .D(I320890), .CLK(I2350), .RSTB(I320740), .Q(I320907) );
not I_18737 (I320924,I320907);
nor I_18738 (I320941,I320791,I320924);
and I_18739 (I320958,I320808,I320941);
and I_18740 (I320975,I320907,I320842);
DFFARX1 I_18741  ( .D(I320975), .CLK(I2350), .RSTB(I320740), .Q(I320708) );
DFFARX1 I_18742  ( .D(I320907), .CLK(I2350), .RSTB(I320740), .Q(I320702) );
DFFARX1 I_18743  ( .D(I130546), .CLK(I2350), .RSTB(I320740), .Q(I321020) );
and I_18744 (I321037,I321020,I130552);
nand I_18745 (I321054,I321037,I320907);
nor I_18746 (I320729,I321037,I320808);
not I_18747 (I321085,I321037);
nor I_18748 (I321102,I320791,I321085);
nand I_18749 (I320720,I320825,I321102);
nand I_18750 (I320714,I320907,I321085);
or I_18751 (I321147,I321037,I320958);
DFFARX1 I_18752  ( .D(I321147), .CLK(I2350), .RSTB(I320740), .Q(I320717) );
DFFARX1 I_18753  ( .D(I130561), .CLK(I2350), .RSTB(I320740), .Q(I321178) );
and I_18754 (I321195,I321178,I321054);
DFFARX1 I_18755  ( .D(I321195), .CLK(I2350), .RSTB(I320740), .Q(I320732) );
nor I_18756 (I321226,I321178,I320791);
nand I_18757 (I320726,I321037,I321226);
not I_18758 (I320723,I321178);
DFFARX1 I_18759  ( .D(I321178), .CLK(I2350), .RSTB(I320740), .Q(I321271) );
and I_18760 (I320705,I321178,I321271);
not I_18761 (I321335,I2357);
nand I_18762 (I321352,I150307,I150277);
and I_18763 (I321369,I321352,I150295);
DFFARX1 I_18764  ( .D(I321369), .CLK(I2350), .RSTB(I321335), .Q(I321386) );
nor I_18765 (I321403,I150289,I150277);
DFFARX1 I_18766  ( .D(I150286), .CLK(I2350), .RSTB(I321335), .Q(I321420) );
nand I_18767 (I321437,I321420,I321403);
DFFARX1 I_18768  ( .D(I321420), .CLK(I2350), .RSTB(I321335), .Q(I321306) );
nand I_18769 (I321468,I150280,I150283);
and I_18770 (I321485,I321468,I150301);
DFFARX1 I_18771  ( .D(I321485), .CLK(I2350), .RSTB(I321335), .Q(I321502) );
not I_18772 (I321519,I321502);
nor I_18773 (I321536,I321386,I321519);
and I_18774 (I321553,I321403,I321536);
and I_18775 (I321570,I321502,I321437);
DFFARX1 I_18776  ( .D(I321570), .CLK(I2350), .RSTB(I321335), .Q(I321303) );
DFFARX1 I_18777  ( .D(I321502), .CLK(I2350), .RSTB(I321335), .Q(I321297) );
DFFARX1 I_18778  ( .D(I150304), .CLK(I2350), .RSTB(I321335), .Q(I321615) );
and I_18779 (I321632,I321615,I150298);
nand I_18780 (I321649,I321632,I321502);
nor I_18781 (I321324,I321632,I321403);
not I_18782 (I321680,I321632);
nor I_18783 (I321697,I321386,I321680);
nand I_18784 (I321315,I321420,I321697);
nand I_18785 (I321309,I321502,I321680);
or I_18786 (I321742,I321632,I321553);
DFFARX1 I_18787  ( .D(I321742), .CLK(I2350), .RSTB(I321335), .Q(I321312) );
DFFARX1 I_18788  ( .D(I150292), .CLK(I2350), .RSTB(I321335), .Q(I321773) );
and I_18789 (I321790,I321773,I321649);
DFFARX1 I_18790  ( .D(I321790), .CLK(I2350), .RSTB(I321335), .Q(I321327) );
nor I_18791 (I321821,I321773,I321386);
nand I_18792 (I321321,I321632,I321821);
not I_18793 (I321318,I321773);
DFFARX1 I_18794  ( .D(I321773), .CLK(I2350), .RSTB(I321335), .Q(I321866) );
and I_18795 (I321300,I321773,I321866);
not I_18796 (I321930,I2357);
nand I_18797 (I321947,I284422,I284407);
and I_18798 (I321964,I321947,I284413);
DFFARX1 I_18799  ( .D(I321964), .CLK(I2350), .RSTB(I321930), .Q(I321981) );
nor I_18800 (I321998,I284416,I284407);
DFFARX1 I_18801  ( .D(I284428), .CLK(I2350), .RSTB(I321930), .Q(I322015) );
nand I_18802 (I322032,I322015,I321998);
DFFARX1 I_18803  ( .D(I322015), .CLK(I2350), .RSTB(I321930), .Q(I321901) );
nand I_18804 (I322063,I284419,I284410);
and I_18805 (I322080,I322063,I284437);
DFFARX1 I_18806  ( .D(I322080), .CLK(I2350), .RSTB(I321930), .Q(I322097) );
not I_18807 (I322114,I322097);
nor I_18808 (I322131,I321981,I322114);
and I_18809 (I322148,I321998,I322131);
and I_18810 (I322165,I322097,I322032);
DFFARX1 I_18811  ( .D(I322165), .CLK(I2350), .RSTB(I321930), .Q(I321898) );
DFFARX1 I_18812  ( .D(I322097), .CLK(I2350), .RSTB(I321930), .Q(I321892) );
DFFARX1 I_18813  ( .D(I284425), .CLK(I2350), .RSTB(I321930), .Q(I322210) );
and I_18814 (I322227,I322210,I284431);
nand I_18815 (I322244,I322227,I322097);
nor I_18816 (I321919,I322227,I321998);
not I_18817 (I322275,I322227);
nor I_18818 (I322292,I321981,I322275);
nand I_18819 (I321910,I322015,I322292);
nand I_18820 (I321904,I322097,I322275);
or I_18821 (I322337,I322227,I322148);
DFFARX1 I_18822  ( .D(I322337), .CLK(I2350), .RSTB(I321930), .Q(I321907) );
DFFARX1 I_18823  ( .D(I284434), .CLK(I2350), .RSTB(I321930), .Q(I322368) );
and I_18824 (I322385,I322368,I322244);
DFFARX1 I_18825  ( .D(I322385), .CLK(I2350), .RSTB(I321930), .Q(I321922) );
nor I_18826 (I322416,I322368,I321981);
nand I_18827 (I321916,I322227,I322416);
not I_18828 (I321913,I322368);
DFFARX1 I_18829  ( .D(I322368), .CLK(I2350), .RSTB(I321930), .Q(I322461) );
and I_18830 (I321895,I322368,I322461);
not I_18831 (I322525,I2357);
nand I_18832 (I322542,I386815,I386818);
and I_18833 (I322559,I322542,I386827);
DFFARX1 I_18834  ( .D(I322559), .CLK(I2350), .RSTB(I322525), .Q(I322576) );
nor I_18835 (I322593,I386821,I386818);
DFFARX1 I_18836  ( .D(I386842), .CLK(I2350), .RSTB(I322525), .Q(I322610) );
nand I_18837 (I322627,I322610,I322593);
DFFARX1 I_18838  ( .D(I322610), .CLK(I2350), .RSTB(I322525), .Q(I322496) );
nand I_18839 (I322658,I386839,I386845);
and I_18840 (I322675,I322658,I386830);
DFFARX1 I_18841  ( .D(I322675), .CLK(I2350), .RSTB(I322525), .Q(I322692) );
not I_18842 (I322709,I322692);
nor I_18843 (I322726,I322576,I322709);
and I_18844 (I322743,I322593,I322726);
and I_18845 (I322760,I322692,I322627);
DFFARX1 I_18846  ( .D(I322760), .CLK(I2350), .RSTB(I322525), .Q(I322493) );
DFFARX1 I_18847  ( .D(I322692), .CLK(I2350), .RSTB(I322525), .Q(I322487) );
DFFARX1 I_18848  ( .D(I386833), .CLK(I2350), .RSTB(I322525), .Q(I322805) );
and I_18849 (I322822,I322805,I386836);
nand I_18850 (I322839,I322822,I322692);
nor I_18851 (I322514,I322822,I322593);
not I_18852 (I322870,I322822);
nor I_18853 (I322887,I322576,I322870);
nand I_18854 (I322505,I322610,I322887);
nand I_18855 (I322499,I322692,I322870);
or I_18856 (I322932,I322822,I322743);
DFFARX1 I_18857  ( .D(I322932), .CLK(I2350), .RSTB(I322525), .Q(I322502) );
DFFARX1 I_18858  ( .D(I386824), .CLK(I2350), .RSTB(I322525), .Q(I322963) );
and I_18859 (I322980,I322963,I322839);
DFFARX1 I_18860  ( .D(I322980), .CLK(I2350), .RSTB(I322525), .Q(I322517) );
nor I_18861 (I323011,I322963,I322576);
nand I_18862 (I322511,I322822,I323011);
not I_18863 (I322508,I322963);
DFFARX1 I_18864  ( .D(I322963), .CLK(I2350), .RSTB(I322525), .Q(I323056) );
and I_18865 (I322490,I322963,I323056);
not I_18866 (I323120,I2357);
nand I_18867 (I323137,I62771,I62747);
and I_18868 (I323154,I323137,I62756);
DFFARX1 I_18869  ( .D(I323154), .CLK(I2350), .RSTB(I323120), .Q(I323171) );
nor I_18870 (I323188,I62750,I62747);
DFFARX1 I_18871  ( .D(I62765), .CLK(I2350), .RSTB(I323120), .Q(I323205) );
nand I_18872 (I323222,I323205,I323188);
DFFARX1 I_18873  ( .D(I323205), .CLK(I2350), .RSTB(I323120), .Q(I323091) );
nand I_18874 (I323253,I62759,I62774);
and I_18875 (I323270,I323253,I62753);
DFFARX1 I_18876  ( .D(I323270), .CLK(I2350), .RSTB(I323120), .Q(I323287) );
not I_18877 (I323304,I323287);
nor I_18878 (I323321,I323171,I323304);
and I_18879 (I323338,I323188,I323321);
and I_18880 (I323355,I323287,I323222);
DFFARX1 I_18881  ( .D(I323355), .CLK(I2350), .RSTB(I323120), .Q(I323088) );
DFFARX1 I_18882  ( .D(I323287), .CLK(I2350), .RSTB(I323120), .Q(I323082) );
DFFARX1 I_18883  ( .D(I62744), .CLK(I2350), .RSTB(I323120), .Q(I323400) );
and I_18884 (I323417,I323400,I62762);
nand I_18885 (I323434,I323417,I323287);
nor I_18886 (I323109,I323417,I323188);
not I_18887 (I323465,I323417);
nor I_18888 (I323482,I323171,I323465);
nand I_18889 (I323100,I323205,I323482);
nand I_18890 (I323094,I323287,I323465);
or I_18891 (I323527,I323417,I323338);
DFFARX1 I_18892  ( .D(I323527), .CLK(I2350), .RSTB(I323120), .Q(I323097) );
DFFARX1 I_18893  ( .D(I62768), .CLK(I2350), .RSTB(I323120), .Q(I323558) );
and I_18894 (I323575,I323558,I323434);
DFFARX1 I_18895  ( .D(I323575), .CLK(I2350), .RSTB(I323120), .Q(I323112) );
nor I_18896 (I323606,I323558,I323171);
nand I_18897 (I323106,I323417,I323606);
not I_18898 (I323103,I323558);
DFFARX1 I_18899  ( .D(I323558), .CLK(I2350), .RSTB(I323120), .Q(I323651) );
and I_18900 (I323085,I323558,I323651);
not I_18901 (I323715,I2357);
nand I_18902 (I323732,I334519,I334507);
and I_18903 (I323749,I323732,I334492);
DFFARX1 I_18904  ( .D(I323749), .CLK(I2350), .RSTB(I323715), .Q(I323766) );
nor I_18905 (I323783,I334504,I334507);
DFFARX1 I_18906  ( .D(I334516), .CLK(I2350), .RSTB(I323715), .Q(I323800) );
nand I_18907 (I323817,I323800,I323783);
DFFARX1 I_18908  ( .D(I323800), .CLK(I2350), .RSTB(I323715), .Q(I323686) );
nand I_18909 (I323848,I334489,I334513);
and I_18910 (I323865,I323848,I334498);
DFFARX1 I_18911  ( .D(I323865), .CLK(I2350), .RSTB(I323715), .Q(I323882) );
not I_18912 (I323899,I323882);
nor I_18913 (I323916,I323766,I323899);
and I_18914 (I323933,I323783,I323916);
and I_18915 (I323950,I323882,I323817);
DFFARX1 I_18916  ( .D(I323950), .CLK(I2350), .RSTB(I323715), .Q(I323683) );
DFFARX1 I_18917  ( .D(I323882), .CLK(I2350), .RSTB(I323715), .Q(I323677) );
DFFARX1 I_18918  ( .D(I334501), .CLK(I2350), .RSTB(I323715), .Q(I323995) );
and I_18919 (I324012,I323995,I334510);
nand I_18920 (I324029,I324012,I323882);
nor I_18921 (I323704,I324012,I323783);
not I_18922 (I324060,I324012);
nor I_18923 (I324077,I323766,I324060);
nand I_18924 (I323695,I323800,I324077);
nand I_18925 (I323689,I323882,I324060);
or I_18926 (I324122,I324012,I323933);
DFFARX1 I_18927  ( .D(I324122), .CLK(I2350), .RSTB(I323715), .Q(I323692) );
DFFARX1 I_18928  ( .D(I334495), .CLK(I2350), .RSTB(I323715), .Q(I324153) );
and I_18929 (I324170,I324153,I324029);
DFFARX1 I_18930  ( .D(I324170), .CLK(I2350), .RSTB(I323715), .Q(I323707) );
nor I_18931 (I324201,I324153,I323766);
nand I_18932 (I323701,I324012,I324201);
not I_18933 (I323698,I324153);
DFFARX1 I_18934  ( .D(I324153), .CLK(I2350), .RSTB(I323715), .Q(I324246) );
and I_18935 (I323680,I324153,I324246);
not I_18936 (I324310,I2357);
nand I_18937 (I324327,I128190,I128175);
and I_18938 (I324344,I324327,I128187);
DFFARX1 I_18939  ( .D(I324344), .CLK(I2350), .RSTB(I324310), .Q(I324361) );
nor I_18940 (I324378,I128178,I128175);
DFFARX1 I_18941  ( .D(I128169), .CLK(I2350), .RSTB(I324310), .Q(I324395) );
nand I_18942 (I324412,I324395,I324378);
DFFARX1 I_18943  ( .D(I324395), .CLK(I2350), .RSTB(I324310), .Q(I324281) );
nand I_18944 (I324443,I128160,I128184);
and I_18945 (I324460,I324443,I128163);
DFFARX1 I_18946  ( .D(I324460), .CLK(I2350), .RSTB(I324310), .Q(I324477) );
not I_18947 (I324494,I324477);
nor I_18948 (I324511,I324361,I324494);
and I_18949 (I324528,I324378,I324511);
and I_18950 (I324545,I324477,I324412);
DFFARX1 I_18951  ( .D(I324545), .CLK(I2350), .RSTB(I324310), .Q(I324278) );
DFFARX1 I_18952  ( .D(I324477), .CLK(I2350), .RSTB(I324310), .Q(I324272) );
DFFARX1 I_18953  ( .D(I128181), .CLK(I2350), .RSTB(I324310), .Q(I324590) );
and I_18954 (I324607,I324590,I128166);
nand I_18955 (I324624,I324607,I324477);
nor I_18956 (I324299,I324607,I324378);
not I_18957 (I324655,I324607);
nor I_18958 (I324672,I324361,I324655);
nand I_18959 (I324290,I324395,I324672);
nand I_18960 (I324284,I324477,I324655);
or I_18961 (I324717,I324607,I324528);
DFFARX1 I_18962  ( .D(I324717), .CLK(I2350), .RSTB(I324310), .Q(I324287) );
DFFARX1 I_18963  ( .D(I128172), .CLK(I2350), .RSTB(I324310), .Q(I324748) );
and I_18964 (I324765,I324748,I324624);
DFFARX1 I_18965  ( .D(I324765), .CLK(I2350), .RSTB(I324310), .Q(I324302) );
nor I_18966 (I324796,I324748,I324361);
nand I_18967 (I324296,I324607,I324796);
not I_18968 (I324293,I324748);
DFFARX1 I_18969  ( .D(I324748), .CLK(I2350), .RSTB(I324310), .Q(I324841) );
and I_18970 (I324275,I324748,I324841);
not I_18971 (I324905,I2357);
nand I_18972 (I324922,I41453,I41429);
and I_18973 (I324939,I324922,I41438);
DFFARX1 I_18974  ( .D(I324939), .CLK(I2350), .RSTB(I324905), .Q(I324956) );
nor I_18975 (I324973,I41432,I41429);
DFFARX1 I_18976  ( .D(I41447), .CLK(I2350), .RSTB(I324905), .Q(I324990) );
nand I_18977 (I325007,I324990,I324973);
DFFARX1 I_18978  ( .D(I324990), .CLK(I2350), .RSTB(I324905), .Q(I324876) );
nand I_18979 (I325038,I41441,I41456);
and I_18980 (I325055,I325038,I41435);
DFFARX1 I_18981  ( .D(I325055), .CLK(I2350), .RSTB(I324905), .Q(I325072) );
not I_18982 (I325089,I325072);
nor I_18983 (I325106,I324956,I325089);
and I_18984 (I325123,I324973,I325106);
and I_18985 (I325140,I325072,I325007);
DFFARX1 I_18986  ( .D(I325140), .CLK(I2350), .RSTB(I324905), .Q(I324873) );
DFFARX1 I_18987  ( .D(I325072), .CLK(I2350), .RSTB(I324905), .Q(I324867) );
DFFARX1 I_18988  ( .D(I41426), .CLK(I2350), .RSTB(I324905), .Q(I325185) );
and I_18989 (I325202,I325185,I41444);
nand I_18990 (I325219,I325202,I325072);
nor I_18991 (I324894,I325202,I324973);
not I_18992 (I325250,I325202);
nor I_18993 (I325267,I324956,I325250);
nand I_18994 (I324885,I324990,I325267);
nand I_18995 (I324879,I325072,I325250);
or I_18996 (I325312,I325202,I325123);
DFFARX1 I_18997  ( .D(I325312), .CLK(I2350), .RSTB(I324905), .Q(I324882) );
DFFARX1 I_18998  ( .D(I41450), .CLK(I2350), .RSTB(I324905), .Q(I325343) );
and I_18999 (I325360,I325343,I325219);
DFFARX1 I_19000  ( .D(I325360), .CLK(I2350), .RSTB(I324905), .Q(I324897) );
nor I_19001 (I325391,I325343,I324956);
nand I_19002 (I324891,I325202,I325391);
not I_19003 (I324888,I325343);
DFFARX1 I_19004  ( .D(I325343), .CLK(I2350), .RSTB(I324905), .Q(I325436) );
and I_19005 (I324870,I325343,I325436);
not I_19006 (I325500,I2357);
nand I_19007 (I325517,I257967,I257982);
and I_19008 (I325534,I325517,I257979);
DFFARX1 I_19009  ( .D(I325534), .CLK(I2350), .RSTB(I325500), .Q(I325551) );
nor I_19010 (I325568,I257955,I257982);
DFFARX1 I_19011  ( .D(I257973), .CLK(I2350), .RSTB(I325500), .Q(I325585) );
nand I_19012 (I325602,I325585,I325568);
DFFARX1 I_19013  ( .D(I325585), .CLK(I2350), .RSTB(I325500), .Q(I325471) );
nand I_19014 (I325633,I257976,I257964);
and I_19015 (I325650,I325633,I257970);
DFFARX1 I_19016  ( .D(I325650), .CLK(I2350), .RSTB(I325500), .Q(I325667) );
not I_19017 (I325684,I325667);
nor I_19018 (I325701,I325551,I325684);
and I_19019 (I325718,I325568,I325701);
and I_19020 (I325735,I325667,I325602);
DFFARX1 I_19021  ( .D(I325735), .CLK(I2350), .RSTB(I325500), .Q(I325468) );
DFFARX1 I_19022  ( .D(I325667), .CLK(I2350), .RSTB(I325500), .Q(I325462) );
DFFARX1 I_19023  ( .D(I257961), .CLK(I2350), .RSTB(I325500), .Q(I325780) );
and I_19024 (I325797,I325780,I257985);
nand I_19025 (I325814,I325797,I325667);
nor I_19026 (I325489,I325797,I325568);
not I_19027 (I325845,I325797);
nor I_19028 (I325862,I325551,I325845);
nand I_19029 (I325480,I325585,I325862);
nand I_19030 (I325474,I325667,I325845);
or I_19031 (I325907,I325797,I325718);
DFFARX1 I_19032  ( .D(I325907), .CLK(I2350), .RSTB(I325500), .Q(I325477) );
DFFARX1 I_19033  ( .D(I257958), .CLK(I2350), .RSTB(I325500), .Q(I325938) );
and I_19034 (I325955,I325938,I325814);
DFFARX1 I_19035  ( .D(I325955), .CLK(I2350), .RSTB(I325500), .Q(I325492) );
nor I_19036 (I325986,I325938,I325551);
nand I_19037 (I325486,I325797,I325986);
not I_19038 (I325483,I325938);
DFFARX1 I_19039  ( .D(I325938), .CLK(I2350), .RSTB(I325500), .Q(I326031) );
and I_19040 (I325465,I325938,I326031);
not I_19041 (I326095,I2357);
nand I_19042 (I326112,I349615,I349603);
and I_19043 (I326129,I326112,I349588);
DFFARX1 I_19044  ( .D(I326129), .CLK(I2350), .RSTB(I326095), .Q(I326146) );
nor I_19045 (I326163,I349600,I349603);
DFFARX1 I_19046  ( .D(I349612), .CLK(I2350), .RSTB(I326095), .Q(I326180) );
nand I_19047 (I326197,I326180,I326163);
DFFARX1 I_19048  ( .D(I326180), .CLK(I2350), .RSTB(I326095), .Q(I326066) );
nand I_19049 (I326228,I349585,I349609);
and I_19050 (I326245,I326228,I349594);
DFFARX1 I_19051  ( .D(I326245), .CLK(I2350), .RSTB(I326095), .Q(I326262) );
not I_19052 (I326279,I326262);
nor I_19053 (I326296,I326146,I326279);
and I_19054 (I326313,I326163,I326296);
and I_19055 (I326330,I326262,I326197);
DFFARX1 I_19056  ( .D(I326330), .CLK(I2350), .RSTB(I326095), .Q(I326063) );
DFFARX1 I_19057  ( .D(I326262), .CLK(I2350), .RSTB(I326095), .Q(I326057) );
DFFARX1 I_19058  ( .D(I349597), .CLK(I2350), .RSTB(I326095), .Q(I326375) );
and I_19059 (I326392,I326375,I349606);
nand I_19060 (I326409,I326392,I326262);
nor I_19061 (I326084,I326392,I326163);
not I_19062 (I326440,I326392);
nor I_19063 (I326457,I326146,I326440);
nand I_19064 (I326075,I326180,I326457);
nand I_19065 (I326069,I326262,I326440);
or I_19066 (I326502,I326392,I326313);
DFFARX1 I_19067  ( .D(I326502), .CLK(I2350), .RSTB(I326095), .Q(I326072) );
DFFARX1 I_19068  ( .D(I349591), .CLK(I2350), .RSTB(I326095), .Q(I326533) );
and I_19069 (I326550,I326533,I326409);
DFFARX1 I_19070  ( .D(I326550), .CLK(I2350), .RSTB(I326095), .Q(I326087) );
nor I_19071 (I326581,I326533,I326146);
nand I_19072 (I326081,I326392,I326581);
not I_19073 (I326078,I326533);
DFFARX1 I_19074  ( .D(I326533), .CLK(I2350), .RSTB(I326095), .Q(I326626) );
and I_19075 (I326060,I326533,I326626);
not I_19076 (I326690,I2357);
nand I_19077 (I326707,I240049,I240064);
and I_19078 (I326724,I326707,I240061);
DFFARX1 I_19079  ( .D(I326724), .CLK(I2350), .RSTB(I326690), .Q(I326741) );
nor I_19080 (I326758,I240037,I240064);
DFFARX1 I_19081  ( .D(I240055), .CLK(I2350), .RSTB(I326690), .Q(I326775) );
nand I_19082 (I326792,I326775,I326758);
DFFARX1 I_19083  ( .D(I326775), .CLK(I2350), .RSTB(I326690), .Q(I326661) );
nand I_19084 (I326823,I240058,I240046);
and I_19085 (I326840,I326823,I240052);
DFFARX1 I_19086  ( .D(I326840), .CLK(I2350), .RSTB(I326690), .Q(I326857) );
not I_19087 (I326874,I326857);
nor I_19088 (I326891,I326741,I326874);
and I_19089 (I326908,I326758,I326891);
and I_19090 (I326925,I326857,I326792);
DFFARX1 I_19091  ( .D(I326925), .CLK(I2350), .RSTB(I326690), .Q(I326658) );
DFFARX1 I_19092  ( .D(I326857), .CLK(I2350), .RSTB(I326690), .Q(I326652) );
DFFARX1 I_19093  ( .D(I240043), .CLK(I2350), .RSTB(I326690), .Q(I326970) );
and I_19094 (I326987,I326970,I240067);
nand I_19095 (I327004,I326987,I326857);
nor I_19096 (I326679,I326987,I326758);
not I_19097 (I327035,I326987);
nor I_19098 (I327052,I326741,I327035);
nand I_19099 (I326670,I326775,I327052);
nand I_19100 (I326664,I326857,I327035);
or I_19101 (I327097,I326987,I326908);
DFFARX1 I_19102  ( .D(I327097), .CLK(I2350), .RSTB(I326690), .Q(I326667) );
DFFARX1 I_19103  ( .D(I240040), .CLK(I2350), .RSTB(I326690), .Q(I327128) );
and I_19104 (I327145,I327128,I327004);
DFFARX1 I_19105  ( .D(I327145), .CLK(I2350), .RSTB(I326690), .Q(I326682) );
nor I_19106 (I327176,I327128,I326741);
nand I_19107 (I326676,I326987,I327176);
not I_19108 (I326673,I327128);
DFFARX1 I_19109  ( .D(I327128), .CLK(I2350), .RSTB(I326690), .Q(I327221) );
and I_19110 (I326655,I327128,I327221);
not I_19111 (I327285,I2357);
nand I_19112 (I327302,I133518,I133515);
and I_19113 (I327319,I327302,I133542);
DFFARX1 I_19114  ( .D(I327319), .CLK(I2350), .RSTB(I327285), .Q(I327336) );
nor I_19115 (I327353,I133545,I133515);
DFFARX1 I_19116  ( .D(I133533), .CLK(I2350), .RSTB(I327285), .Q(I327370) );
nand I_19117 (I327387,I327370,I327353);
DFFARX1 I_19118  ( .D(I327370), .CLK(I2350), .RSTB(I327285), .Q(I327256) );
nand I_19119 (I327418,I133539,I133524);
and I_19120 (I327435,I327418,I133530);
DFFARX1 I_19121  ( .D(I327435), .CLK(I2350), .RSTB(I327285), .Q(I327452) );
not I_19122 (I327469,I327452);
nor I_19123 (I327486,I327336,I327469);
and I_19124 (I327503,I327353,I327486);
and I_19125 (I327520,I327452,I327387);
DFFARX1 I_19126  ( .D(I327520), .CLK(I2350), .RSTB(I327285), .Q(I327253) );
DFFARX1 I_19127  ( .D(I327452), .CLK(I2350), .RSTB(I327285), .Q(I327247) );
DFFARX1 I_19128  ( .D(I133521), .CLK(I2350), .RSTB(I327285), .Q(I327565) );
and I_19129 (I327582,I327565,I133527);
nand I_19130 (I327599,I327582,I327452);
nor I_19131 (I327274,I327582,I327353);
not I_19132 (I327630,I327582);
nor I_19133 (I327647,I327336,I327630);
nand I_19134 (I327265,I327370,I327647);
nand I_19135 (I327259,I327452,I327630);
or I_19136 (I327692,I327582,I327503);
DFFARX1 I_19137  ( .D(I327692), .CLK(I2350), .RSTB(I327285), .Q(I327262) );
DFFARX1 I_19138  ( .D(I133536), .CLK(I2350), .RSTB(I327285), .Q(I327723) );
and I_19139 (I327740,I327723,I327599);
DFFARX1 I_19140  ( .D(I327740), .CLK(I2350), .RSTB(I327285), .Q(I327277) );
nor I_19141 (I327771,I327723,I327336);
nand I_19142 (I327271,I327582,I327771);
not I_19143 (I327268,I327723);
DFFARX1 I_19144  ( .D(I327723), .CLK(I2350), .RSTB(I327285), .Q(I327816) );
and I_19145 (I327250,I327723,I327816);
not I_19146 (I327880,I2357);
nand I_19147 (I327897,I40807,I40783);
and I_19148 (I327914,I327897,I40792);
DFFARX1 I_19149  ( .D(I327914), .CLK(I2350), .RSTB(I327880), .Q(I327931) );
nor I_19150 (I327948,I40786,I40783);
DFFARX1 I_19151  ( .D(I40801), .CLK(I2350), .RSTB(I327880), .Q(I327965) );
nand I_19152 (I327982,I327965,I327948);
DFFARX1 I_19153  ( .D(I327965), .CLK(I2350), .RSTB(I327880), .Q(I327851) );
nand I_19154 (I328013,I40795,I40810);
and I_19155 (I328030,I328013,I40789);
DFFARX1 I_19156  ( .D(I328030), .CLK(I2350), .RSTB(I327880), .Q(I328047) );
not I_19157 (I328064,I328047);
nor I_19158 (I328081,I327931,I328064);
and I_19159 (I328098,I327948,I328081);
and I_19160 (I328115,I328047,I327982);
DFFARX1 I_19161  ( .D(I328115), .CLK(I2350), .RSTB(I327880), .Q(I327848) );
DFFARX1 I_19162  ( .D(I328047), .CLK(I2350), .RSTB(I327880), .Q(I327842) );
DFFARX1 I_19163  ( .D(I40780), .CLK(I2350), .RSTB(I327880), .Q(I328160) );
and I_19164 (I328177,I328160,I40798);
nand I_19165 (I328194,I328177,I328047);
nor I_19166 (I327869,I328177,I327948);
not I_19167 (I328225,I328177);
nor I_19168 (I328242,I327931,I328225);
nand I_19169 (I327860,I327965,I328242);
nand I_19170 (I327854,I328047,I328225);
or I_19171 (I328287,I328177,I328098);
DFFARX1 I_19172  ( .D(I328287), .CLK(I2350), .RSTB(I327880), .Q(I327857) );
DFFARX1 I_19173  ( .D(I40804), .CLK(I2350), .RSTB(I327880), .Q(I328318) );
and I_19174 (I328335,I328318,I328194);
DFFARX1 I_19175  ( .D(I328335), .CLK(I2350), .RSTB(I327880), .Q(I327872) );
nor I_19176 (I328366,I328318,I327931);
nand I_19177 (I327866,I328177,I328366);
not I_19178 (I327863,I328318);
DFFARX1 I_19179  ( .D(I328318), .CLK(I2350), .RSTB(I327880), .Q(I328411) );
and I_19180 (I327845,I328318,I328411);
not I_19181 (I328475,I2357);
nand I_19182 (I328492,I296322,I296307);
and I_19183 (I328509,I328492,I296313);
DFFARX1 I_19184  ( .D(I328509), .CLK(I2350), .RSTB(I328475), .Q(I328526) );
nor I_19185 (I328543,I296316,I296307);
DFFARX1 I_19186  ( .D(I296328), .CLK(I2350), .RSTB(I328475), .Q(I328560) );
nand I_19187 (I328577,I328560,I328543);
DFFARX1 I_19188  ( .D(I328560), .CLK(I2350), .RSTB(I328475), .Q(I328446) );
nand I_19189 (I328608,I296319,I296310);
and I_19190 (I328625,I328608,I296337);
DFFARX1 I_19191  ( .D(I328625), .CLK(I2350), .RSTB(I328475), .Q(I328642) );
not I_19192 (I328659,I328642);
nor I_19193 (I328676,I328526,I328659);
and I_19194 (I328693,I328543,I328676);
and I_19195 (I328710,I328642,I328577);
DFFARX1 I_19196  ( .D(I328710), .CLK(I2350), .RSTB(I328475), .Q(I328443) );
DFFARX1 I_19197  ( .D(I328642), .CLK(I2350), .RSTB(I328475), .Q(I328437) );
DFFARX1 I_19198  ( .D(I296325), .CLK(I2350), .RSTB(I328475), .Q(I328755) );
and I_19199 (I328772,I328755,I296331);
nand I_19200 (I328789,I328772,I328642);
nor I_19201 (I328464,I328772,I328543);
not I_19202 (I328820,I328772);
nor I_19203 (I328837,I328526,I328820);
nand I_19204 (I328455,I328560,I328837);
nand I_19205 (I328449,I328642,I328820);
or I_19206 (I328882,I328772,I328693);
DFFARX1 I_19207  ( .D(I328882), .CLK(I2350), .RSTB(I328475), .Q(I328452) );
DFFARX1 I_19208  ( .D(I296334), .CLK(I2350), .RSTB(I328475), .Q(I328913) );
and I_19209 (I328930,I328913,I328789);
DFFARX1 I_19210  ( .D(I328930), .CLK(I2350), .RSTB(I328475), .Q(I328467) );
nor I_19211 (I328961,I328913,I328526);
nand I_19212 (I328461,I328772,I328961);
not I_19213 (I328458,I328913);
DFFARX1 I_19214  ( .D(I328913), .CLK(I2350), .RSTB(I328475), .Q(I329006) );
and I_19215 (I328440,I328913,I329006);
not I_19216 (I329070,I2357);
nand I_19217 (I329087,I212107,I212119);
and I_19218 (I329104,I329087,I212110);
DFFARX1 I_19219  ( .D(I329104), .CLK(I2350), .RSTB(I329070), .Q(I329121) );
nor I_19220 (I329138,I212104,I212119);
DFFARX1 I_19221  ( .D(I212095), .CLK(I2350), .RSTB(I329070), .Q(I329155) );
nand I_19222 (I329172,I329155,I329138);
DFFARX1 I_19223  ( .D(I329155), .CLK(I2350), .RSTB(I329070), .Q(I329041) );
nand I_19224 (I329203,I212101,I212092);
and I_19225 (I329220,I329203,I212098);
DFFARX1 I_19226  ( .D(I329220), .CLK(I2350), .RSTB(I329070), .Q(I329237) );
not I_19227 (I329254,I329237);
nor I_19228 (I329271,I329121,I329254);
and I_19229 (I329288,I329138,I329271);
and I_19230 (I329305,I329237,I329172);
DFFARX1 I_19231  ( .D(I329305), .CLK(I2350), .RSTB(I329070), .Q(I329038) );
DFFARX1 I_19232  ( .D(I329237), .CLK(I2350), .RSTB(I329070), .Q(I329032) );
DFFARX1 I_19233  ( .D(I212113), .CLK(I2350), .RSTB(I329070), .Q(I329350) );
and I_19234 (I329367,I329350,I212089);
nand I_19235 (I329384,I329367,I329237);
nor I_19236 (I329059,I329367,I329138);
not I_19237 (I329415,I329367);
nor I_19238 (I329432,I329121,I329415);
nand I_19239 (I329050,I329155,I329432);
nand I_19240 (I329044,I329237,I329415);
or I_19241 (I329477,I329367,I329288);
DFFARX1 I_19242  ( .D(I329477), .CLK(I2350), .RSTB(I329070), .Q(I329047) );
DFFARX1 I_19243  ( .D(I212116), .CLK(I2350), .RSTB(I329070), .Q(I329508) );
and I_19244 (I329525,I329508,I329384);
DFFARX1 I_19245  ( .D(I329525), .CLK(I2350), .RSTB(I329070), .Q(I329062) );
nor I_19246 (I329556,I329508,I329121);
nand I_19247 (I329056,I329367,I329556);
not I_19248 (I329053,I329508);
DFFARX1 I_19249  ( .D(I329508), .CLK(I2350), .RSTB(I329070), .Q(I329601) );
and I_19250 (I329035,I329508,I329601);
not I_19251 (I329665,I2357);
nand I_19252 (I329682,I350873,I350861);
and I_19253 (I329699,I329682,I350846);
DFFARX1 I_19254  ( .D(I329699), .CLK(I2350), .RSTB(I329665), .Q(I329716) );
nor I_19255 (I329733,I350858,I350861);
DFFARX1 I_19256  ( .D(I350870), .CLK(I2350), .RSTB(I329665), .Q(I329750) );
nand I_19257 (I329767,I329750,I329733);
DFFARX1 I_19258  ( .D(I329750), .CLK(I2350), .RSTB(I329665), .Q(I329636) );
nand I_19259 (I329798,I350843,I350867);
and I_19260 (I329815,I329798,I350852);
DFFARX1 I_19261  ( .D(I329815), .CLK(I2350), .RSTB(I329665), .Q(I329832) );
not I_19262 (I329849,I329832);
nor I_19263 (I329866,I329716,I329849);
and I_19264 (I329883,I329733,I329866);
and I_19265 (I329900,I329832,I329767);
DFFARX1 I_19266  ( .D(I329900), .CLK(I2350), .RSTB(I329665), .Q(I329633) );
DFFARX1 I_19267  ( .D(I329832), .CLK(I2350), .RSTB(I329665), .Q(I329627) );
DFFARX1 I_19268  ( .D(I350855), .CLK(I2350), .RSTB(I329665), .Q(I329945) );
and I_19269 (I329962,I329945,I350864);
nand I_19270 (I329979,I329962,I329832);
nor I_19271 (I329654,I329962,I329733);
not I_19272 (I330010,I329962);
nor I_19273 (I330027,I329716,I330010);
nand I_19274 (I329645,I329750,I330027);
nand I_19275 (I329639,I329832,I330010);
or I_19276 (I330072,I329962,I329883);
DFFARX1 I_19277  ( .D(I330072), .CLK(I2350), .RSTB(I329665), .Q(I329642) );
DFFARX1 I_19278  ( .D(I350849), .CLK(I2350), .RSTB(I329665), .Q(I330103) );
and I_19279 (I330120,I330103,I329979);
DFFARX1 I_19280  ( .D(I330120), .CLK(I2350), .RSTB(I329665), .Q(I329657) );
nor I_19281 (I330151,I330103,I329716);
nand I_19282 (I329651,I329962,I330151);
not I_19283 (I329648,I330103);
DFFARX1 I_19284  ( .D(I330103), .CLK(I2350), .RSTB(I329665), .Q(I330196) );
and I_19285 (I329630,I330103,I330196);
not I_19286 (I330260,I2357);
nand I_19287 (I330277,I389705,I389708);
and I_19288 (I330294,I330277,I389717);
DFFARX1 I_19289  ( .D(I330294), .CLK(I2350), .RSTB(I330260), .Q(I330311) );
nor I_19290 (I330328,I389711,I389708);
DFFARX1 I_19291  ( .D(I389732), .CLK(I2350), .RSTB(I330260), .Q(I330345) );
nand I_19292 (I330362,I330345,I330328);
DFFARX1 I_19293  ( .D(I330345), .CLK(I2350), .RSTB(I330260), .Q(I330231) );
nand I_19294 (I330393,I389729,I389735);
and I_19295 (I330410,I330393,I389720);
DFFARX1 I_19296  ( .D(I330410), .CLK(I2350), .RSTB(I330260), .Q(I330427) );
not I_19297 (I330444,I330427);
nor I_19298 (I330461,I330311,I330444);
and I_19299 (I330478,I330328,I330461);
and I_19300 (I330495,I330427,I330362);
DFFARX1 I_19301  ( .D(I330495), .CLK(I2350), .RSTB(I330260), .Q(I330228) );
DFFARX1 I_19302  ( .D(I330427), .CLK(I2350), .RSTB(I330260), .Q(I330222) );
DFFARX1 I_19303  ( .D(I389723), .CLK(I2350), .RSTB(I330260), .Q(I330540) );
and I_19304 (I330557,I330540,I389726);
nand I_19305 (I330574,I330557,I330427);
nor I_19306 (I330249,I330557,I330328);
not I_19307 (I330605,I330557);
nor I_19308 (I330622,I330311,I330605);
nand I_19309 (I330240,I330345,I330622);
nand I_19310 (I330234,I330427,I330605);
or I_19311 (I330667,I330557,I330478);
DFFARX1 I_19312  ( .D(I330667), .CLK(I2350), .RSTB(I330260), .Q(I330237) );
DFFARX1 I_19313  ( .D(I389714), .CLK(I2350), .RSTB(I330260), .Q(I330698) );
and I_19314 (I330715,I330698,I330574);
DFFARX1 I_19315  ( .D(I330715), .CLK(I2350), .RSTB(I330260), .Q(I330252) );
nor I_19316 (I330746,I330698,I330311);
nand I_19317 (I330246,I330557,I330746);
not I_19318 (I330243,I330698);
DFFARX1 I_19319  ( .D(I330698), .CLK(I2350), .RSTB(I330260), .Q(I330791) );
and I_19320 (I330225,I330698,I330791);
not I_19321 (I330855,I2357);
nand I_19322 (I330872,I228903,I228915);
and I_19323 (I330889,I330872,I228906);
DFFARX1 I_19324  ( .D(I330889), .CLK(I2350), .RSTB(I330855), .Q(I330906) );
nor I_19325 (I330923,I228900,I228915);
DFFARX1 I_19326  ( .D(I228891), .CLK(I2350), .RSTB(I330855), .Q(I330940) );
nand I_19327 (I330957,I330940,I330923);
DFFARX1 I_19328  ( .D(I330940), .CLK(I2350), .RSTB(I330855), .Q(I330826) );
nand I_19329 (I330988,I228897,I228888);
and I_19330 (I331005,I330988,I228894);
DFFARX1 I_19331  ( .D(I331005), .CLK(I2350), .RSTB(I330855), .Q(I331022) );
not I_19332 (I331039,I331022);
nor I_19333 (I331056,I330906,I331039);
and I_19334 (I331073,I330923,I331056);
and I_19335 (I331090,I331022,I330957);
DFFARX1 I_19336  ( .D(I331090), .CLK(I2350), .RSTB(I330855), .Q(I330823) );
DFFARX1 I_19337  ( .D(I331022), .CLK(I2350), .RSTB(I330855), .Q(I330817) );
DFFARX1 I_19338  ( .D(I228909), .CLK(I2350), .RSTB(I330855), .Q(I331135) );
and I_19339 (I331152,I331135,I228885);
nand I_19340 (I331169,I331152,I331022);
nor I_19341 (I330844,I331152,I330923);
not I_19342 (I331200,I331152);
nor I_19343 (I331217,I330906,I331200);
nand I_19344 (I330835,I330940,I331217);
nand I_19345 (I330829,I331022,I331200);
or I_19346 (I331262,I331152,I331073);
DFFARX1 I_19347  ( .D(I331262), .CLK(I2350), .RSTB(I330855), .Q(I330832) );
DFFARX1 I_19348  ( .D(I228912), .CLK(I2350), .RSTB(I330855), .Q(I331293) );
and I_19349 (I331310,I331293,I331169);
DFFARX1 I_19350  ( .D(I331310), .CLK(I2350), .RSTB(I330855), .Q(I330847) );
nor I_19351 (I331341,I331293,I330906);
nand I_19352 (I330841,I331152,I331341);
not I_19353 (I330838,I331293);
DFFARX1 I_19354  ( .D(I331293), .CLK(I2350), .RSTB(I330855), .Q(I331386) );
and I_19355 (I330820,I331293,I331386);
not I_19356 (I331450,I2357);
nand I_19357 (I331467,I82151,I82127);
and I_19358 (I331484,I331467,I82136);
DFFARX1 I_19359  ( .D(I331484), .CLK(I2350), .RSTB(I331450), .Q(I331501) );
nor I_19360 (I331518,I82130,I82127);
DFFARX1 I_19361  ( .D(I82145), .CLK(I2350), .RSTB(I331450), .Q(I331535) );
nand I_19362 (I331552,I331535,I331518);
DFFARX1 I_19363  ( .D(I331535), .CLK(I2350), .RSTB(I331450), .Q(I331421) );
nand I_19364 (I331583,I82139,I82154);
and I_19365 (I331600,I331583,I82133);
DFFARX1 I_19366  ( .D(I331600), .CLK(I2350), .RSTB(I331450), .Q(I331617) );
not I_19367 (I331634,I331617);
nor I_19368 (I331651,I331501,I331634);
and I_19369 (I331668,I331518,I331651);
and I_19370 (I331685,I331617,I331552);
DFFARX1 I_19371  ( .D(I331685), .CLK(I2350), .RSTB(I331450), .Q(I331418) );
DFFARX1 I_19372  ( .D(I331617), .CLK(I2350), .RSTB(I331450), .Q(I331412) );
DFFARX1 I_19373  ( .D(I82124), .CLK(I2350), .RSTB(I331450), .Q(I331730) );
and I_19374 (I331747,I331730,I82142);
nand I_19375 (I331764,I331747,I331617);
nor I_19376 (I331439,I331747,I331518);
not I_19377 (I331795,I331747);
nor I_19378 (I331812,I331501,I331795);
nand I_19379 (I331430,I331535,I331812);
nand I_19380 (I331424,I331617,I331795);
or I_19381 (I331857,I331747,I331668);
DFFARX1 I_19382  ( .D(I331857), .CLK(I2350), .RSTB(I331450), .Q(I331427) );
DFFARX1 I_19383  ( .D(I82148), .CLK(I2350), .RSTB(I331450), .Q(I331888) );
and I_19384 (I331905,I331888,I331764);
DFFARX1 I_19385  ( .D(I331905), .CLK(I2350), .RSTB(I331450), .Q(I331442) );
nor I_19386 (I331936,I331888,I331501);
nand I_19387 (I331436,I331747,I331936);
not I_19388 (I331433,I331888);
DFFARX1 I_19389  ( .D(I331888), .CLK(I2350), .RSTB(I331450), .Q(I331981) );
and I_19390 (I331415,I331888,I331981);
not I_19391 (I332045,I2357);
nand I_19392 (I332062,I207585,I207597);
and I_19393 (I332079,I332062,I207588);
DFFARX1 I_19394  ( .D(I332079), .CLK(I2350), .RSTB(I332045), .Q(I332096) );
nor I_19395 (I332113,I207582,I207597);
DFFARX1 I_19396  ( .D(I207573), .CLK(I2350), .RSTB(I332045), .Q(I332130) );
nand I_19397 (I332147,I332130,I332113);
DFFARX1 I_19398  ( .D(I332130), .CLK(I2350), .RSTB(I332045), .Q(I332016) );
nand I_19399 (I332178,I207579,I207570);
and I_19400 (I332195,I332178,I207576);
DFFARX1 I_19401  ( .D(I332195), .CLK(I2350), .RSTB(I332045), .Q(I332212) );
not I_19402 (I332229,I332212);
nor I_19403 (I332246,I332096,I332229);
and I_19404 (I332263,I332113,I332246);
and I_19405 (I332280,I332212,I332147);
DFFARX1 I_19406  ( .D(I332280), .CLK(I2350), .RSTB(I332045), .Q(I332013) );
DFFARX1 I_19407  ( .D(I332212), .CLK(I2350), .RSTB(I332045), .Q(I332007) );
DFFARX1 I_19408  ( .D(I207591), .CLK(I2350), .RSTB(I332045), .Q(I332325) );
and I_19409 (I332342,I332325,I207567);
nand I_19410 (I332359,I332342,I332212);
nor I_19411 (I332034,I332342,I332113);
not I_19412 (I332390,I332342);
nor I_19413 (I332407,I332096,I332390);
nand I_19414 (I332025,I332130,I332407);
nand I_19415 (I332019,I332212,I332390);
or I_19416 (I332452,I332342,I332263);
DFFARX1 I_19417  ( .D(I332452), .CLK(I2350), .RSTB(I332045), .Q(I332022) );
DFFARX1 I_19418  ( .D(I207594), .CLK(I2350), .RSTB(I332045), .Q(I332483) );
and I_19419 (I332500,I332483,I332359);
DFFARX1 I_19420  ( .D(I332500), .CLK(I2350), .RSTB(I332045), .Q(I332037) );
nor I_19421 (I332531,I332483,I332096);
nand I_19422 (I332031,I332342,I332531);
not I_19423 (I332028,I332483);
DFFARX1 I_19424  ( .D(I332483), .CLK(I2350), .RSTB(I332045), .Q(I332576) );
and I_19425 (I332010,I332483,I332576);
not I_19426 (I332640,I2357);
not I_19427 (I332657,I2924);
nor I_19428 (I332674,I2927,I2936);
nand I_19429 (I332691,I332674,I2951);
nor I_19430 (I332708,I332657,I2927);
nand I_19431 (I332725,I332708,I2930);
not I_19432 (I332742,I2927);
not I_19433 (I332759,I332742);
not I_19434 (I332776,I2921);
nor I_19435 (I332793,I332776,I2945);
and I_19436 (I332810,I332793,I2933);
or I_19437 (I332827,I332810,I2939);
DFFARX1 I_19438  ( .D(I332827), .CLK(I2350), .RSTB(I332640), .Q(I332844) );
nand I_19439 (I332861,I332657,I2921);
or I_19440 (I332629,I332861,I332844);
not I_19441 (I332892,I332861);
nor I_19442 (I332909,I332844,I332892);
and I_19443 (I332926,I332742,I332909);
nand I_19444 (I332602,I332861,I332759);
DFFARX1 I_19445  ( .D(I2942), .CLK(I2350), .RSTB(I332640), .Q(I332957) );
or I_19446 (I332623,I332957,I332844);
nor I_19447 (I332988,I332957,I332725);
nor I_19448 (I333005,I332957,I332759);
nand I_19449 (I332608,I332691,I333005);
or I_19450 (I333036,I332957,I332926);
DFFARX1 I_19451  ( .D(I333036), .CLK(I2350), .RSTB(I332640), .Q(I332605) );
not I_19452 (I332611,I332957);
DFFARX1 I_19453  ( .D(I2948), .CLK(I2350), .RSTB(I332640), .Q(I333081) );
not I_19454 (I333098,I333081);
nor I_19455 (I333115,I333098,I332691);
DFFARX1 I_19456  ( .D(I333115), .CLK(I2350), .RSTB(I332640), .Q(I332617) );
nor I_19457 (I332632,I332957,I333098);
nor I_19458 (I332620,I333098,I332861);
not I_19459 (I333174,I333098);
and I_19460 (I333191,I332725,I333174);
nor I_19461 (I332626,I332861,I333191);
nand I_19462 (I332614,I333098,I332988);
not I_19463 (I333269,I2357);
not I_19464 (I333286,I162229);
nor I_19465 (I333303,I162235,I162214);
nand I_19466 (I333320,I333303,I162220);
nor I_19467 (I333337,I333286,I162235);
nand I_19468 (I333354,I333337,I162226);
not I_19469 (I333371,I162235);
not I_19470 (I333388,I333371);
not I_19471 (I333405,I162223);
nor I_19472 (I333422,I333405,I162241);
and I_19473 (I333439,I333422,I162232);
or I_19474 (I333456,I333439,I162211);
DFFARX1 I_19475  ( .D(I333456), .CLK(I2350), .RSTB(I333269), .Q(I333473) );
nand I_19476 (I333490,I333286,I162223);
or I_19477 (I333258,I333490,I333473);
not I_19478 (I333521,I333490);
nor I_19479 (I333538,I333473,I333521);
and I_19480 (I333555,I333371,I333538);
nand I_19481 (I333231,I333490,I333388);
DFFARX1 I_19482  ( .D(I162238), .CLK(I2350), .RSTB(I333269), .Q(I333586) );
or I_19483 (I333252,I333586,I333473);
nor I_19484 (I333617,I333586,I333354);
nor I_19485 (I333634,I333586,I333388);
nand I_19486 (I333237,I333320,I333634);
or I_19487 (I333665,I333586,I333555);
DFFARX1 I_19488  ( .D(I333665), .CLK(I2350), .RSTB(I333269), .Q(I333234) );
not I_19489 (I333240,I333586);
DFFARX1 I_19490  ( .D(I162217), .CLK(I2350), .RSTB(I333269), .Q(I333710) );
not I_19491 (I333727,I333710);
nor I_19492 (I333744,I333727,I333320);
DFFARX1 I_19493  ( .D(I333744), .CLK(I2350), .RSTB(I333269), .Q(I333246) );
nor I_19494 (I333261,I333586,I333727);
nor I_19495 (I333249,I333727,I333490);
not I_19496 (I333803,I333727);
and I_19497 (I333820,I333354,I333803);
nor I_19498 (I333255,I333490,I333820);
nand I_19499 (I333243,I333727,I333617);
not I_19500 (I333898,I2357);
not I_19501 (I333915,I205001);
nor I_19502 (I333932,I205010,I205013);
nand I_19503 (I333949,I333932,I204998);
nor I_19504 (I333966,I333915,I205010);
nand I_19505 (I333983,I333966,I204995);
not I_19506 (I334000,I205010);
not I_19507 (I334017,I334000);
not I_19508 (I334034,I204983);
nor I_19509 (I334051,I334034,I204989);
and I_19510 (I334068,I334051,I204986);
or I_19511 (I334085,I334068,I205007);
DFFARX1 I_19512  ( .D(I334085), .CLK(I2350), .RSTB(I333898), .Q(I334102) );
nand I_19513 (I334119,I333915,I204983);
or I_19514 (I333887,I334119,I334102);
not I_19515 (I334150,I334119);
nor I_19516 (I334167,I334102,I334150);
and I_19517 (I334184,I334000,I334167);
nand I_19518 (I333860,I334119,I334017);
DFFARX1 I_19519  ( .D(I204992), .CLK(I2350), .RSTB(I333898), .Q(I334215) );
or I_19520 (I333881,I334215,I334102);
nor I_19521 (I334246,I334215,I333983);
nor I_19522 (I334263,I334215,I334017);
nand I_19523 (I333866,I333949,I334263);
or I_19524 (I334294,I334215,I334184);
DFFARX1 I_19525  ( .D(I334294), .CLK(I2350), .RSTB(I333898), .Q(I333863) );
not I_19526 (I333869,I334215);
DFFARX1 I_19527  ( .D(I205004), .CLK(I2350), .RSTB(I333898), .Q(I334339) );
not I_19528 (I334356,I334339);
nor I_19529 (I334373,I334356,I333949);
DFFARX1 I_19530  ( .D(I334373), .CLK(I2350), .RSTB(I333898), .Q(I333875) );
nor I_19531 (I333890,I334215,I334356);
nor I_19532 (I333878,I334356,I334119);
not I_19533 (I334432,I334356);
and I_19534 (I334449,I333983,I334432);
nor I_19535 (I333884,I334119,I334449);
nand I_19536 (I333872,I334356,I334246);
not I_19537 (I334527,I2357);
not I_19538 (I334544,I293933);
nor I_19539 (I334561,I293951,I293930);
nand I_19540 (I334578,I334561,I293954);
nor I_19541 (I334595,I334544,I293951);
nand I_19542 (I334612,I334595,I293948);
not I_19543 (I334629,I293951);
not I_19544 (I334646,I334629);
not I_19545 (I334663,I293939);
nor I_19546 (I334680,I334663,I293927);
and I_19547 (I334697,I334680,I293945);
or I_19548 (I334714,I334697,I293957);
DFFARX1 I_19549  ( .D(I334714), .CLK(I2350), .RSTB(I334527), .Q(I334731) );
nand I_19550 (I334748,I334544,I293939);
or I_19551 (I334516,I334748,I334731);
not I_19552 (I334779,I334748);
nor I_19553 (I334796,I334731,I334779);
and I_19554 (I334813,I334629,I334796);
nand I_19555 (I334489,I334748,I334646);
DFFARX1 I_19556  ( .D(I293936), .CLK(I2350), .RSTB(I334527), .Q(I334844) );
or I_19557 (I334510,I334844,I334731);
nor I_19558 (I334875,I334844,I334612);
nor I_19559 (I334892,I334844,I334646);
nand I_19560 (I334495,I334578,I334892);
or I_19561 (I334923,I334844,I334813);
DFFARX1 I_19562  ( .D(I334923), .CLK(I2350), .RSTB(I334527), .Q(I334492) );
not I_19563 (I334498,I334844);
DFFARX1 I_19564  ( .D(I293942), .CLK(I2350), .RSTB(I334527), .Q(I334968) );
not I_19565 (I334985,I334968);
nor I_19566 (I335002,I334985,I334578);
DFFARX1 I_19567  ( .D(I335002), .CLK(I2350), .RSTB(I334527), .Q(I334504) );
nor I_19568 (I334519,I334844,I334985);
nor I_19569 (I334507,I334985,I334748);
not I_19570 (I335061,I334985);
and I_19571 (I335078,I334612,I335061);
nor I_19572 (I334513,I334748,I335078);
nand I_19573 (I334501,I334985,I334875);
not I_19574 (I335156,I2357);
not I_19575 (I335173,I139687);
nor I_19576 (I335190,I139693,I139672);
nand I_19577 (I335207,I335190,I139678);
nor I_19578 (I335224,I335173,I139693);
nand I_19579 (I335241,I335224,I139684);
not I_19580 (I335258,I139693);
not I_19581 (I335275,I335258);
not I_19582 (I335292,I139681);
nor I_19583 (I335309,I335292,I139699);
and I_19584 (I335326,I335309,I139690);
or I_19585 (I335343,I335326,I139669);
DFFARX1 I_19586  ( .D(I335343), .CLK(I2350), .RSTB(I335156), .Q(I335360) );
nand I_19587 (I335377,I335173,I139681);
or I_19588 (I335145,I335377,I335360);
not I_19589 (I335408,I335377);
nor I_19590 (I335425,I335360,I335408);
and I_19591 (I335442,I335258,I335425);
nand I_19592 (I335118,I335377,I335275);
DFFARX1 I_19593  ( .D(I139696), .CLK(I2350), .RSTB(I335156), .Q(I335473) );
or I_19594 (I335139,I335473,I335360);
nor I_19595 (I335504,I335473,I335241);
nor I_19596 (I335521,I335473,I335275);
nand I_19597 (I335124,I335207,I335521);
or I_19598 (I335552,I335473,I335442);
DFFARX1 I_19599  ( .D(I335552), .CLK(I2350), .RSTB(I335156), .Q(I335121) );
not I_19600 (I335127,I335473);
DFFARX1 I_19601  ( .D(I139675), .CLK(I2350), .RSTB(I335156), .Q(I335597) );
not I_19602 (I335614,I335597);
nor I_19603 (I335631,I335614,I335207);
DFFARX1 I_19604  ( .D(I335631), .CLK(I2350), .RSTB(I335156), .Q(I335133) );
nor I_19605 (I335148,I335473,I335614);
nor I_19606 (I335136,I335614,I335377);
not I_19607 (I335690,I335614);
and I_19608 (I335707,I335241,I335690);
nor I_19609 (I335142,I335377,I335707);
nand I_19610 (I335130,I335614,I335504);
not I_19611 (I335785,I2357);
not I_19612 (I335802,I303453);
nor I_19613 (I335819,I303471,I303450);
nand I_19614 (I335836,I335819,I303474);
nor I_19615 (I335853,I335802,I303471);
nand I_19616 (I335870,I335853,I303468);
not I_19617 (I335887,I303471);
not I_19618 (I335904,I335887);
not I_19619 (I335921,I303459);
nor I_19620 (I335938,I335921,I303447);
and I_19621 (I335955,I335938,I303465);
or I_19622 (I335972,I335955,I303477);
DFFARX1 I_19623  ( .D(I335972), .CLK(I2350), .RSTB(I335785), .Q(I335989) );
nand I_19624 (I336006,I335802,I303459);
or I_19625 (I335774,I336006,I335989);
not I_19626 (I336037,I336006);
nor I_19627 (I336054,I335989,I336037);
and I_19628 (I336071,I335887,I336054);
nand I_19629 (I335747,I336006,I335904);
DFFARX1 I_19630  ( .D(I303456), .CLK(I2350), .RSTB(I335785), .Q(I336102) );
or I_19631 (I335768,I336102,I335989);
nor I_19632 (I336133,I336102,I335870);
nor I_19633 (I336150,I336102,I335904);
nand I_19634 (I335753,I335836,I336150);
or I_19635 (I336181,I336102,I336071);
DFFARX1 I_19636  ( .D(I336181), .CLK(I2350), .RSTB(I335785), .Q(I335750) );
not I_19637 (I335756,I336102);
DFFARX1 I_19638  ( .D(I303462), .CLK(I2350), .RSTB(I335785), .Q(I336226) );
not I_19639 (I336243,I336226);
nor I_19640 (I336260,I336243,I335836);
DFFARX1 I_19641  ( .D(I336260), .CLK(I2350), .RSTB(I335785), .Q(I335762) );
nor I_19642 (I335777,I336102,I336243);
nor I_19643 (I335765,I336243,I336006);
not I_19644 (I336319,I336243);
and I_19645 (I336336,I335870,I336319);
nor I_19646 (I335771,I336006,I336336);
nand I_19647 (I335759,I336243,I336133);
not I_19648 (I336414,I2357);
not I_19649 (I336431,I115695);
nor I_19650 (I336448,I115671,I115686);
nand I_19651 (I336465,I336448,I115668);
nor I_19652 (I336482,I336431,I115671);
nand I_19653 (I336499,I336482,I115683);
not I_19654 (I336516,I115671);
not I_19655 (I336533,I336516);
not I_19656 (I336550,I115674);
nor I_19657 (I336567,I336550,I115689);
and I_19658 (I336584,I336567,I115680);
or I_19659 (I336601,I336584,I115665);
DFFARX1 I_19660  ( .D(I336601), .CLK(I2350), .RSTB(I336414), .Q(I336618) );
nand I_19661 (I336635,I336431,I115674);
or I_19662 (I336403,I336635,I336618);
not I_19663 (I336666,I336635);
nor I_19664 (I336683,I336618,I336666);
and I_19665 (I336700,I336516,I336683);
nand I_19666 (I336376,I336635,I336533);
DFFARX1 I_19667  ( .D(I115677), .CLK(I2350), .RSTB(I336414), .Q(I336731) );
or I_19668 (I336397,I336731,I336618);
nor I_19669 (I336762,I336731,I336499);
nor I_19670 (I336779,I336731,I336533);
nand I_19671 (I336382,I336465,I336779);
or I_19672 (I336810,I336731,I336700);
DFFARX1 I_19673  ( .D(I336810), .CLK(I2350), .RSTB(I336414), .Q(I336379) );
not I_19674 (I336385,I336731);
DFFARX1 I_19675  ( .D(I115692), .CLK(I2350), .RSTB(I336414), .Q(I336855) );
not I_19676 (I336872,I336855);
nor I_19677 (I336889,I336872,I336465);
DFFARX1 I_19678  ( .D(I336889), .CLK(I2350), .RSTB(I336414), .Q(I336391) );
nor I_19679 (I336406,I336731,I336872);
nor I_19680 (I336394,I336872,I336635);
not I_19681 (I336948,I336872);
and I_19682 (I336965,I336499,I336948);
nor I_19683 (I336400,I336635,I336965);
nand I_19684 (I336388,I336872,I336762);
not I_19685 (I337043,I2357);
not I_19686 (I337060,I192727);
nor I_19687 (I337077,I192736,I192739);
nand I_19688 (I337094,I337077,I192724);
nor I_19689 (I337111,I337060,I192736);
nand I_19690 (I337128,I337111,I192721);
not I_19691 (I337145,I192736);
not I_19692 (I337162,I337145);
not I_19693 (I337179,I192709);
nor I_19694 (I337196,I337179,I192715);
and I_19695 (I337213,I337196,I192712);
or I_19696 (I337230,I337213,I192733);
DFFARX1 I_19697  ( .D(I337230), .CLK(I2350), .RSTB(I337043), .Q(I337247) );
nand I_19698 (I337264,I337060,I192709);
or I_19699 (I337032,I337264,I337247);
not I_19700 (I337295,I337264);
nor I_19701 (I337312,I337247,I337295);
and I_19702 (I337329,I337145,I337312);
nand I_19703 (I337005,I337264,I337162);
DFFARX1 I_19704  ( .D(I192718), .CLK(I2350), .RSTB(I337043), .Q(I337360) );
or I_19705 (I337026,I337360,I337247);
nor I_19706 (I337391,I337360,I337128);
nor I_19707 (I337408,I337360,I337162);
nand I_19708 (I337011,I337094,I337408);
or I_19709 (I337439,I337360,I337329);
DFFARX1 I_19710  ( .D(I337439), .CLK(I2350), .RSTB(I337043), .Q(I337008) );
not I_19711 (I337014,I337360);
DFFARX1 I_19712  ( .D(I192730), .CLK(I2350), .RSTB(I337043), .Q(I337484) );
not I_19713 (I337501,I337484);
nor I_19714 (I337518,I337501,I337094);
DFFARX1 I_19715  ( .D(I337518), .CLK(I2350), .RSTB(I337043), .Q(I337020) );
nor I_19716 (I337035,I337360,I337501);
nor I_19717 (I337023,I337501,I337264);
not I_19718 (I337577,I337501);
and I_19719 (I337594,I337128,I337577);
nor I_19720 (I337029,I337264,I337594);
nand I_19721 (I337017,I337501,I337391);
not I_19722 (I337672,I2357);
not I_19723 (I337689,I384509);
nor I_19724 (I337706,I384533,I384518);
nand I_19725 (I337723,I337706,I384503);
nor I_19726 (I337740,I337689,I384533);
nand I_19727 (I337757,I337740,I384530);
not I_19728 (I337774,I384533);
not I_19729 (I337791,I337774);
not I_19730 (I337808,I384512);
nor I_19731 (I337825,I337808,I384506);
and I_19732 (I337842,I337825,I384527);
or I_19733 (I337859,I337842,I384515);
DFFARX1 I_19734  ( .D(I337859), .CLK(I2350), .RSTB(I337672), .Q(I337876) );
nand I_19735 (I337893,I337689,I384512);
or I_19736 (I337661,I337893,I337876);
not I_19737 (I337924,I337893);
nor I_19738 (I337941,I337876,I337924);
and I_19739 (I337958,I337774,I337941);
nand I_19740 (I337634,I337893,I337791);
DFFARX1 I_19741  ( .D(I384524), .CLK(I2350), .RSTB(I337672), .Q(I337989) );
or I_19742 (I337655,I337989,I337876);
nor I_19743 (I338020,I337989,I337757);
nor I_19744 (I338037,I337989,I337791);
nand I_19745 (I337640,I337723,I338037);
or I_19746 (I338068,I337989,I337958);
DFFARX1 I_19747  ( .D(I338068), .CLK(I2350), .RSTB(I337672), .Q(I337637) );
not I_19748 (I337643,I337989);
DFFARX1 I_19749  ( .D(I384521), .CLK(I2350), .RSTB(I337672), .Q(I338113) );
not I_19750 (I338130,I338113);
nor I_19751 (I338147,I338130,I337723);
DFFARX1 I_19752  ( .D(I338147), .CLK(I2350), .RSTB(I337672), .Q(I337649) );
nor I_19753 (I337664,I337989,I338130);
nor I_19754 (I337652,I338130,I337893);
not I_19755 (I338206,I338130);
and I_19756 (I338223,I337757,I338206);
nor I_19757 (I337658,I337893,I338223);
nand I_19758 (I337646,I338130,I338020);
not I_19759 (I338301,I2357);
not I_19760 (I338318,I14144);
nor I_19761 (I338335,I14147,I14156);
nand I_19762 (I338352,I338335,I14171);
nor I_19763 (I338369,I338318,I14147);
nand I_19764 (I338386,I338369,I14150);
not I_19765 (I338403,I14147);
not I_19766 (I338420,I338403);
not I_19767 (I338437,I14141);
nor I_19768 (I338454,I338437,I14165);
and I_19769 (I338471,I338454,I14153);
or I_19770 (I338488,I338471,I14159);
DFFARX1 I_19771  ( .D(I338488), .CLK(I2350), .RSTB(I338301), .Q(I338505) );
nand I_19772 (I338522,I338318,I14141);
or I_19773 (I338290,I338522,I338505);
not I_19774 (I338553,I338522);
nor I_19775 (I338570,I338505,I338553);
and I_19776 (I338587,I338403,I338570);
nand I_19777 (I338263,I338522,I338420);
DFFARX1 I_19778  ( .D(I14162), .CLK(I2350), .RSTB(I338301), .Q(I338618) );
or I_19779 (I338284,I338618,I338505);
nor I_19780 (I338649,I338618,I338386);
nor I_19781 (I338666,I338618,I338420);
nand I_19782 (I338269,I338352,I338666);
or I_19783 (I338697,I338618,I338587);
DFFARX1 I_19784  ( .D(I338697), .CLK(I2350), .RSTB(I338301), .Q(I338266) );
not I_19785 (I338272,I338618);
DFFARX1 I_19786  ( .D(I14168), .CLK(I2350), .RSTB(I338301), .Q(I338742) );
not I_19787 (I338759,I338742);
nor I_19788 (I338776,I338759,I338352);
DFFARX1 I_19789  ( .D(I338776), .CLK(I2350), .RSTB(I338301), .Q(I338278) );
nor I_19790 (I338293,I338618,I338759);
nor I_19791 (I338281,I338759,I338522);
not I_19792 (I338835,I338759);
and I_19793 (I338852,I338386,I338835);
nor I_19794 (I338287,I338522,I338852);
nand I_19795 (I338275,I338759,I338649);
not I_19796 (I338930,I2357);
not I_19797 (I338947,I396647);
nor I_19798 (I338964,I396671,I396656);
nand I_19799 (I338981,I338964,I396641);
nor I_19800 (I338998,I338947,I396671);
nand I_19801 (I339015,I338998,I396668);
not I_19802 (I339032,I396671);
not I_19803 (I339049,I339032);
not I_19804 (I339066,I396650);
nor I_19805 (I339083,I339066,I396644);
and I_19806 (I339100,I339083,I396665);
or I_19807 (I339117,I339100,I396653);
DFFARX1 I_19808  ( .D(I339117), .CLK(I2350), .RSTB(I338930), .Q(I339134) );
nand I_19809 (I339151,I338947,I396650);
or I_19810 (I338919,I339151,I339134);
not I_19811 (I339182,I339151);
nor I_19812 (I339199,I339134,I339182);
and I_19813 (I339216,I339032,I339199);
nand I_19814 (I338892,I339151,I339049);
DFFARX1 I_19815  ( .D(I396662), .CLK(I2350), .RSTB(I338930), .Q(I339247) );
or I_19816 (I338913,I339247,I339134);
nor I_19817 (I339278,I339247,I339015);
nor I_19818 (I339295,I339247,I339049);
nand I_19819 (I338898,I338981,I339295);
or I_19820 (I339326,I339247,I339216);
DFFARX1 I_19821  ( .D(I339326), .CLK(I2350), .RSTB(I338930), .Q(I338895) );
not I_19822 (I338901,I339247);
DFFARX1 I_19823  ( .D(I396659), .CLK(I2350), .RSTB(I338930), .Q(I339371) );
not I_19824 (I339388,I339371);
nor I_19825 (I339405,I339388,I338981);
DFFARX1 I_19826  ( .D(I339405), .CLK(I2350), .RSTB(I338930), .Q(I338907) );
nor I_19827 (I338922,I339247,I339388);
nor I_19828 (I338910,I339388,I339151);
not I_19829 (I339464,I339388);
and I_19830 (I339481,I339015,I339464);
nor I_19831 (I338916,I339151,I339481);
nand I_19832 (I338904,I339388,I339278);
not I_19833 (I339559,I2357);
not I_19834 (I339576,I238911);
nor I_19835 (I339593,I238884,I238902);
nand I_19836 (I339610,I339593,I238887);
nor I_19837 (I339627,I339576,I238884);
nand I_19838 (I339644,I339627,I238905);
not I_19839 (I339661,I238884);
not I_19840 (I339678,I339661);
not I_19841 (I339695,I238881);
nor I_19842 (I339712,I339695,I238908);
and I_19843 (I339729,I339712,I238899);
or I_19844 (I339746,I339729,I238890);
DFFARX1 I_19845  ( .D(I339746), .CLK(I2350), .RSTB(I339559), .Q(I339763) );
nand I_19846 (I339780,I339576,I238881);
or I_19847 (I339548,I339780,I339763);
not I_19848 (I339811,I339780);
nor I_19849 (I339828,I339763,I339811);
and I_19850 (I339845,I339661,I339828);
nand I_19851 (I339521,I339780,I339678);
DFFARX1 I_19852  ( .D(I238893), .CLK(I2350), .RSTB(I339559), .Q(I339876) );
or I_19853 (I339542,I339876,I339763);
nor I_19854 (I339907,I339876,I339644);
nor I_19855 (I339924,I339876,I339678);
nand I_19856 (I339527,I339610,I339924);
or I_19857 (I339955,I339876,I339845);
DFFARX1 I_19858  ( .D(I339955), .CLK(I2350), .RSTB(I339559), .Q(I339524) );
not I_19859 (I339530,I339876);
DFFARX1 I_19860  ( .D(I238896), .CLK(I2350), .RSTB(I339559), .Q(I340000) );
not I_19861 (I340017,I340000);
nor I_19862 (I340034,I340017,I339610);
DFFARX1 I_19863  ( .D(I340034), .CLK(I2350), .RSTB(I339559), .Q(I339536) );
nor I_19864 (I339551,I339876,I340017);
nor I_19865 (I339539,I340017,I339780);
not I_19866 (I340093,I340017);
and I_19867 (I340110,I339644,I340093);
nor I_19868 (I339545,I339780,I340110);
nand I_19869 (I339533,I340017,I339907);
not I_19870 (I340188,I2357);
not I_19871 (I340205,I197249);
nor I_19872 (I340222,I197258,I197261);
nand I_19873 (I340239,I340222,I197246);
nor I_19874 (I340256,I340205,I197258);
nand I_19875 (I340273,I340256,I197243);
not I_19876 (I340290,I197258);
not I_19877 (I340307,I340290);
not I_19878 (I340324,I197231);
nor I_19879 (I340341,I340324,I197237);
and I_19880 (I340358,I340341,I197234);
or I_19881 (I340375,I340358,I197255);
DFFARX1 I_19882  ( .D(I340375), .CLK(I2350), .RSTB(I340188), .Q(I340392) );
nand I_19883 (I340409,I340205,I197231);
or I_19884 (I340177,I340409,I340392);
not I_19885 (I340440,I340409);
nor I_19886 (I340457,I340392,I340440);
and I_19887 (I340474,I340290,I340457);
nand I_19888 (I340150,I340409,I340307);
DFFARX1 I_19889  ( .D(I197240), .CLK(I2350), .RSTB(I340188), .Q(I340505) );
or I_19890 (I340171,I340505,I340392);
nor I_19891 (I340536,I340505,I340273);
nor I_19892 (I340553,I340505,I340307);
nand I_19893 (I340156,I340239,I340553);
or I_19894 (I340584,I340505,I340474);
DFFARX1 I_19895  ( .D(I340584), .CLK(I2350), .RSTB(I340188), .Q(I340153) );
not I_19896 (I340159,I340505);
DFFARX1 I_19897  ( .D(I197252), .CLK(I2350), .RSTB(I340188), .Q(I340629) );
not I_19898 (I340646,I340629);
nor I_19899 (I340663,I340646,I340239);
DFFARX1 I_19900  ( .D(I340663), .CLK(I2350), .RSTB(I340188), .Q(I340165) );
nor I_19901 (I340180,I340505,I340646);
nor I_19902 (I340168,I340646,I340409);
not I_19903 (I340722,I340646);
and I_19904 (I340739,I340273,I340722);
nor I_19905 (I340174,I340409,I340739);
nand I_19906 (I340162,I340646,I340536);
not I_19907 (I340817,I2357);
not I_19908 (I340834,I59520);
nor I_19909 (I340851,I59538,I59517);
nand I_19910 (I340868,I340851,I59535);
nor I_19911 (I340885,I340834,I59538);
nand I_19912 (I340902,I340885,I59529);
not I_19913 (I340919,I59538);
not I_19914 (I340936,I340919);
not I_19915 (I340953,I59532);
nor I_19916 (I340970,I340953,I59526);
and I_19917 (I340987,I340970,I59523);
or I_19918 (I341004,I340987,I59514);
DFFARX1 I_19919  ( .D(I341004), .CLK(I2350), .RSTB(I340817), .Q(I341021) );
nand I_19920 (I341038,I340834,I59532);
or I_19921 (I340806,I341038,I341021);
not I_19922 (I341069,I341038);
nor I_19923 (I341086,I341021,I341069);
and I_19924 (I341103,I340919,I341086);
nand I_19925 (I340779,I341038,I340936);
DFFARX1 I_19926  ( .D(I59544), .CLK(I2350), .RSTB(I340817), .Q(I341134) );
or I_19927 (I340800,I341134,I341021);
nor I_19928 (I341165,I341134,I340902);
nor I_19929 (I341182,I341134,I340936);
nand I_19930 (I340785,I340868,I341182);
or I_19931 (I341213,I341134,I341103);
DFFARX1 I_19932  ( .D(I341213), .CLK(I2350), .RSTB(I340817), .Q(I340782) );
not I_19933 (I340788,I341134);
DFFARX1 I_19934  ( .D(I59541), .CLK(I2350), .RSTB(I340817), .Q(I341258) );
not I_19935 (I341275,I341258);
nor I_19936 (I341292,I341275,I340868);
DFFARX1 I_19937  ( .D(I341292), .CLK(I2350), .RSTB(I340817), .Q(I340794) );
nor I_19938 (I340809,I341134,I341275);
nor I_19939 (I340797,I341275,I341038);
not I_19940 (I341351,I341275);
and I_19941 (I341368,I340902,I341351);
nor I_19942 (I340803,I341038,I341368);
nand I_19943 (I340791,I341275,I341165);
not I_19944 (I341446,I2357);
not I_19945 (I341463,I11339);
nor I_19946 (I341480,I11342,I11351);
nand I_19947 (I341497,I341480,I11366);
nor I_19948 (I341514,I341463,I11342);
nand I_19949 (I341531,I341514,I11345);
not I_19950 (I341548,I11342);
not I_19951 (I341565,I341548);
not I_19952 (I341582,I11336);
nor I_19953 (I341599,I341582,I11360);
and I_19954 (I341616,I341599,I11348);
or I_19955 (I341633,I341616,I11354);
DFFARX1 I_19956  ( .D(I341633), .CLK(I2350), .RSTB(I341446), .Q(I341650) );
nand I_19957 (I341667,I341463,I11336);
or I_19958 (I341435,I341667,I341650);
not I_19959 (I341698,I341667);
nor I_19960 (I341715,I341650,I341698);
and I_19961 (I341732,I341548,I341715);
nand I_19962 (I341408,I341667,I341565);
DFFARX1 I_19963  ( .D(I11357), .CLK(I2350), .RSTB(I341446), .Q(I341763) );
or I_19964 (I341429,I341763,I341650);
nor I_19965 (I341794,I341763,I341531);
nor I_19966 (I341811,I341763,I341565);
nand I_19967 (I341414,I341497,I341811);
or I_19968 (I341842,I341763,I341732);
DFFARX1 I_19969  ( .D(I341842), .CLK(I2350), .RSTB(I341446), .Q(I341411) );
not I_19970 (I341417,I341763);
DFFARX1 I_19971  ( .D(I11363), .CLK(I2350), .RSTB(I341446), .Q(I341887) );
not I_19972 (I341904,I341887);
nor I_19973 (I341921,I341904,I341497);
DFFARX1 I_19974  ( .D(I341921), .CLK(I2350), .RSTB(I341446), .Q(I341423) );
nor I_19975 (I341438,I341763,I341904);
nor I_19976 (I341426,I341904,I341667);
not I_19977 (I341980,I341904);
and I_19978 (I341997,I341531,I341980);
nor I_19979 (I341432,I341667,I341997);
nand I_19980 (I341420,I341904,I341794);
not I_19981 (I342075,I2357);
not I_19982 (I342092,I56936);
nor I_19983 (I342109,I56954,I56933);
nand I_19984 (I342126,I342109,I56951);
nor I_19985 (I342143,I342092,I56954);
nand I_19986 (I342160,I342143,I56945);
not I_19987 (I342177,I56954);
not I_19988 (I342194,I342177);
not I_19989 (I342211,I56948);
nor I_19990 (I342228,I342211,I56942);
and I_19991 (I342245,I342228,I56939);
or I_19992 (I342262,I342245,I56930);
DFFARX1 I_19993  ( .D(I342262), .CLK(I2350), .RSTB(I342075), .Q(I342279) );
nand I_19994 (I342296,I342092,I56948);
or I_19995 (I342064,I342296,I342279);
not I_19996 (I342327,I342296);
nor I_19997 (I342344,I342279,I342327);
and I_19998 (I342361,I342177,I342344);
nand I_19999 (I342037,I342296,I342194);
DFFARX1 I_20000  ( .D(I56960), .CLK(I2350), .RSTB(I342075), .Q(I342392) );
or I_20001 (I342058,I342392,I342279);
nor I_20002 (I342423,I342392,I342160);
nor I_20003 (I342440,I342392,I342194);
nand I_20004 (I342043,I342126,I342440);
or I_20005 (I342471,I342392,I342361);
DFFARX1 I_20006  ( .D(I342471), .CLK(I2350), .RSTB(I342075), .Q(I342040) );
not I_20007 (I342046,I342392);
DFFARX1 I_20008  ( .D(I56957), .CLK(I2350), .RSTB(I342075), .Q(I342516) );
not I_20009 (I342533,I342516);
nor I_20010 (I342550,I342533,I342126);
DFFARX1 I_20011  ( .D(I342550), .CLK(I2350), .RSTB(I342075), .Q(I342052) );
nor I_20012 (I342067,I342392,I342533);
nor I_20013 (I342055,I342533,I342296);
not I_20014 (I342609,I342533);
and I_20015 (I342626,I342160,I342609);
nor I_20016 (I342061,I342296,I342626);
nand I_20017 (I342049,I342533,I342423);
not I_20018 (I342704,I2357);
not I_20019 (I342721,I69210);
nor I_20020 (I342738,I69228,I69207);
nand I_20021 (I342755,I342738,I69225);
nor I_20022 (I342772,I342721,I69228);
nand I_20023 (I342789,I342772,I69219);
not I_20024 (I342806,I69228);
not I_20025 (I342823,I342806);
not I_20026 (I342840,I69222);
nor I_20027 (I342857,I342840,I69216);
and I_20028 (I342874,I342857,I69213);
or I_20029 (I342891,I342874,I69204);
DFFARX1 I_20030  ( .D(I342891), .CLK(I2350), .RSTB(I342704), .Q(I342908) );
nand I_20031 (I342925,I342721,I69222);
or I_20032 (I342693,I342925,I342908);
not I_20033 (I342956,I342925);
nor I_20034 (I342973,I342908,I342956);
and I_20035 (I342990,I342806,I342973);
nand I_20036 (I342666,I342925,I342823);
DFFARX1 I_20037  ( .D(I69234), .CLK(I2350), .RSTB(I342704), .Q(I343021) );
or I_20038 (I342687,I343021,I342908);
nor I_20039 (I343052,I343021,I342789);
nor I_20040 (I343069,I343021,I342823);
nand I_20041 (I342672,I342755,I343069);
or I_20042 (I343100,I343021,I342990);
DFFARX1 I_20043  ( .D(I343100), .CLK(I2350), .RSTB(I342704), .Q(I342669) );
not I_20044 (I342675,I343021);
DFFARX1 I_20045  ( .D(I69231), .CLK(I2350), .RSTB(I342704), .Q(I343145) );
not I_20046 (I343162,I343145);
nor I_20047 (I343179,I343162,I342755);
DFFARX1 I_20048  ( .D(I343179), .CLK(I2350), .RSTB(I342704), .Q(I342681) );
nor I_20049 (I342696,I343021,I343162);
nor I_20050 (I342684,I343162,I342925);
not I_20051 (I343238,I343162);
and I_20052 (I343255,I342789,I343238);
nor I_20053 (I342690,I342925,I343255);
nand I_20054 (I342678,I343162,I343052);
not I_20055 (I343333,I2357);
not I_20056 (I343350,I23681);
nor I_20057 (I343367,I23684,I23693);
nand I_20058 (I343384,I343367,I23708);
nor I_20059 (I343401,I343350,I23684);
nand I_20060 (I343418,I343401,I23687);
not I_20061 (I343435,I23684);
not I_20062 (I343452,I343435);
not I_20063 (I343469,I23678);
nor I_20064 (I343486,I343469,I23702);
and I_20065 (I343503,I343486,I23690);
or I_20066 (I343520,I343503,I23696);
DFFARX1 I_20067  ( .D(I343520), .CLK(I2350), .RSTB(I343333), .Q(I343537) );
nand I_20068 (I343554,I343350,I23678);
or I_20069 (I343322,I343554,I343537);
not I_20070 (I343585,I343554);
nor I_20071 (I343602,I343537,I343585);
and I_20072 (I343619,I343435,I343602);
nand I_20073 (I343295,I343554,I343452);
DFFARX1 I_20074  ( .D(I23699), .CLK(I2350), .RSTB(I343333), .Q(I343650) );
or I_20075 (I343316,I343650,I343537);
nor I_20076 (I343681,I343650,I343418);
nor I_20077 (I343698,I343650,I343452);
nand I_20078 (I343301,I343384,I343698);
or I_20079 (I343729,I343650,I343619);
DFFARX1 I_20080  ( .D(I343729), .CLK(I2350), .RSTB(I343333), .Q(I343298) );
not I_20081 (I343304,I343650);
DFFARX1 I_20082  ( .D(I23705), .CLK(I2350), .RSTB(I343333), .Q(I343774) );
not I_20083 (I343791,I343774);
nor I_20084 (I343808,I343791,I343384);
DFFARX1 I_20085  ( .D(I343808), .CLK(I2350), .RSTB(I343333), .Q(I343310) );
nor I_20086 (I343325,I343650,I343791);
nor I_20087 (I343313,I343791,I343554);
not I_20088 (I343867,I343791);
and I_20089 (I343884,I343418,I343867);
nor I_20090 (I343319,I343554,I343884);
nand I_20091 (I343307,I343791,I343681);
not I_20092 (I343962,I2357);
not I_20093 (I343979,I332016);
nor I_20094 (I343996,I332019,I332028);
nand I_20095 (I344013,I343996,I332013);
nor I_20096 (I344030,I343979,I332019);
nand I_20097 (I344047,I344030,I332022);
not I_20098 (I344064,I332019);
not I_20099 (I344081,I344064);
not I_20100 (I344098,I332037);
nor I_20101 (I344115,I344098,I332025);
and I_20102 (I344132,I344115,I332010);
or I_20103 (I344149,I344132,I332007);
DFFARX1 I_20104  ( .D(I344149), .CLK(I2350), .RSTB(I343962), .Q(I344166) );
nand I_20105 (I344183,I343979,I332037);
or I_20106 (I343951,I344183,I344166);
not I_20107 (I344214,I344183);
nor I_20108 (I344231,I344166,I344214);
and I_20109 (I344248,I344064,I344231);
nand I_20110 (I343924,I344183,I344081);
DFFARX1 I_20111  ( .D(I332031), .CLK(I2350), .RSTB(I343962), .Q(I344279) );
or I_20112 (I343945,I344279,I344166);
nor I_20113 (I344310,I344279,I344047);
nor I_20114 (I344327,I344279,I344081);
nand I_20115 (I343930,I344013,I344327);
or I_20116 (I344358,I344279,I344248);
DFFARX1 I_20117  ( .D(I344358), .CLK(I2350), .RSTB(I343962), .Q(I343927) );
not I_20118 (I343933,I344279);
DFFARX1 I_20119  ( .D(I332034), .CLK(I2350), .RSTB(I343962), .Q(I344403) );
not I_20120 (I344420,I344403);
nor I_20121 (I344437,I344420,I344013);
DFFARX1 I_20122  ( .D(I344437), .CLK(I2350), .RSTB(I343962), .Q(I343939) );
nor I_20123 (I343954,I344279,I344420);
nor I_20124 (I343942,I344420,I344183);
not I_20125 (I344496,I344420);
and I_20126 (I344513,I344047,I344496);
nor I_20127 (I343948,I344183,I344513);
nand I_20128 (I343936,I344420,I344310);
not I_20129 (I344591,I2357);
not I_20130 (I344608,I151621);
nor I_20131 (I344625,I151627,I151606);
nand I_20132 (I344642,I344625,I151612);
nor I_20133 (I344659,I344608,I151627);
nand I_20134 (I344676,I344659,I151618);
not I_20135 (I344693,I151627);
not I_20136 (I344710,I344693);
not I_20137 (I344727,I151615);
nor I_20138 (I344744,I344727,I151633);
and I_20139 (I344761,I344744,I151624);
or I_20140 (I344778,I344761,I151603);
DFFARX1 I_20141  ( .D(I344778), .CLK(I2350), .RSTB(I344591), .Q(I344795) );
nand I_20142 (I344812,I344608,I151615);
or I_20143 (I344580,I344812,I344795);
not I_20144 (I344843,I344812);
nor I_20145 (I344860,I344795,I344843);
and I_20146 (I344877,I344693,I344860);
nand I_20147 (I344553,I344812,I344710);
DFFARX1 I_20148  ( .D(I151630), .CLK(I2350), .RSTB(I344591), .Q(I344908) );
or I_20149 (I344574,I344908,I344795);
nor I_20150 (I344939,I344908,I344676);
nor I_20151 (I344956,I344908,I344710);
nand I_20152 (I344559,I344642,I344956);
or I_20153 (I344987,I344908,I344877);
DFFARX1 I_20154  ( .D(I344987), .CLK(I2350), .RSTB(I344591), .Q(I344556) );
not I_20155 (I344562,I344908);
DFFARX1 I_20156  ( .D(I151609), .CLK(I2350), .RSTB(I344591), .Q(I345032) );
not I_20157 (I345049,I345032);
nor I_20158 (I345066,I345049,I344642);
DFFARX1 I_20159  ( .D(I345066), .CLK(I2350), .RSTB(I344591), .Q(I344568) );
nor I_20160 (I344583,I344908,I345049);
nor I_20161 (I344571,I345049,I344812);
not I_20162 (I345125,I345049);
and I_20163 (I345142,I344676,I345125);
nor I_20164 (I344577,I344812,I345142);
nand I_20165 (I344565,I345049,I344939);
not I_20166 (I345220,I2357);
not I_20167 (I345237,I381619);
nor I_20168 (I345254,I381643,I381628);
nand I_20169 (I345271,I345254,I381613);
nor I_20170 (I345288,I345237,I381643);
nand I_20171 (I345305,I345288,I381640);
not I_20172 (I345322,I381643);
not I_20173 (I345339,I345322);
not I_20174 (I345356,I381622);
nor I_20175 (I345373,I345356,I381616);
and I_20176 (I345390,I345373,I381637);
or I_20177 (I345407,I345390,I381625);
DFFARX1 I_20178  ( .D(I345407), .CLK(I2350), .RSTB(I345220), .Q(I345424) );
nand I_20179 (I345441,I345237,I381622);
or I_20180 (I345209,I345441,I345424);
not I_20181 (I345472,I345441);
nor I_20182 (I345489,I345424,I345472);
and I_20183 (I345506,I345322,I345489);
nand I_20184 (I345182,I345441,I345339);
DFFARX1 I_20185  ( .D(I381634), .CLK(I2350), .RSTB(I345220), .Q(I345537) );
or I_20186 (I345203,I345537,I345424);
nor I_20187 (I345568,I345537,I345305);
nor I_20188 (I345585,I345537,I345339);
nand I_20189 (I345188,I345271,I345585);
or I_20190 (I345616,I345537,I345506);
DFFARX1 I_20191  ( .D(I345616), .CLK(I2350), .RSTB(I345220), .Q(I345185) );
not I_20192 (I345191,I345537);
DFFARX1 I_20193  ( .D(I381631), .CLK(I2350), .RSTB(I345220), .Q(I345661) );
not I_20194 (I345678,I345661);
nor I_20195 (I345695,I345678,I345271);
DFFARX1 I_20196  ( .D(I345695), .CLK(I2350), .RSTB(I345220), .Q(I345197) );
nor I_20197 (I345212,I345537,I345678);
nor I_20198 (I345200,I345678,I345441);
not I_20199 (I345754,I345678);
and I_20200 (I345771,I345305,I345754);
nor I_20201 (I345206,I345441,I345771);
nand I_20202 (I345194,I345678,I345568);
not I_20203 (I345849,I2357);
not I_20204 (I345866,I186097);
nor I_20205 (I345883,I186103,I186082);
nand I_20206 (I345900,I345883,I186088);
nor I_20207 (I345917,I345866,I186103);
nand I_20208 (I345934,I345917,I186094);
not I_20209 (I345951,I186103);
not I_20210 (I345968,I345951);
not I_20211 (I345985,I186091);
nor I_20212 (I346002,I345985,I186109);
and I_20213 (I346019,I346002,I186100);
or I_20214 (I346036,I346019,I186079);
DFFARX1 I_20215  ( .D(I346036), .CLK(I2350), .RSTB(I345849), .Q(I346053) );
nand I_20216 (I346070,I345866,I186091);
or I_20217 (I345838,I346070,I346053);
not I_20218 (I346101,I346070);
nor I_20219 (I346118,I346053,I346101);
and I_20220 (I346135,I345951,I346118);
nand I_20221 (I345811,I346070,I345968);
DFFARX1 I_20222  ( .D(I186106), .CLK(I2350), .RSTB(I345849), .Q(I346166) );
or I_20223 (I345832,I346166,I346053);
nor I_20224 (I346197,I346166,I345934);
nor I_20225 (I346214,I346166,I345968);
nand I_20226 (I345817,I345900,I346214);
or I_20227 (I346245,I346166,I346135);
DFFARX1 I_20228  ( .D(I346245), .CLK(I2350), .RSTB(I345849), .Q(I345814) );
not I_20229 (I345820,I346166);
DFFARX1 I_20230  ( .D(I186085), .CLK(I2350), .RSTB(I345849), .Q(I346290) );
not I_20231 (I346307,I346290);
nor I_20232 (I346324,I346307,I345900);
DFFARX1 I_20233  ( .D(I346324), .CLK(I2350), .RSTB(I345849), .Q(I345826) );
nor I_20234 (I345841,I346166,I346307);
nor I_20235 (I345829,I346307,I346070);
not I_20236 (I346383,I346307);
and I_20237 (I346400,I345934,I346383);
nor I_20238 (I345835,I346070,I346400);
nand I_20239 (I345823,I346307,I346197);
not I_20240 (I346478,I2357);
not I_20241 (I346495,I62104);
nor I_20242 (I346512,I62122,I62101);
nand I_20243 (I346529,I346512,I62119);
nor I_20244 (I346546,I346495,I62122);
nand I_20245 (I346563,I346546,I62113);
not I_20246 (I346580,I62122);
not I_20247 (I346597,I346580);
not I_20248 (I346614,I62116);
nor I_20249 (I346631,I346614,I62110);
and I_20250 (I346648,I346631,I62107);
or I_20251 (I346665,I346648,I62098);
DFFARX1 I_20252  ( .D(I346665), .CLK(I2350), .RSTB(I346478), .Q(I346682) );
nand I_20253 (I346699,I346495,I62116);
or I_20254 (I346467,I346699,I346682);
not I_20255 (I346730,I346699);
nor I_20256 (I346747,I346682,I346730);
and I_20257 (I346764,I346580,I346747);
nand I_20258 (I346440,I346699,I346597);
DFFARX1 I_20259  ( .D(I62128), .CLK(I2350), .RSTB(I346478), .Q(I346795) );
or I_20260 (I346461,I346795,I346682);
nor I_20261 (I346826,I346795,I346563);
nor I_20262 (I346843,I346795,I346597);
nand I_20263 (I346446,I346529,I346843);
or I_20264 (I346874,I346795,I346764);
DFFARX1 I_20265  ( .D(I346874), .CLK(I2350), .RSTB(I346478), .Q(I346443) );
not I_20266 (I346449,I346795);
DFFARX1 I_20267  ( .D(I62125), .CLK(I2350), .RSTB(I346478), .Q(I346919) );
not I_20268 (I346936,I346919);
nor I_20269 (I346953,I346936,I346529);
DFFARX1 I_20270  ( .D(I346953), .CLK(I2350), .RSTB(I346478), .Q(I346455) );
nor I_20271 (I346470,I346795,I346936);
nor I_20272 (I346458,I346936,I346699);
not I_20273 (I347012,I346936);
and I_20274 (I347029,I346563,I347012);
nor I_20275 (I346464,I346699,I347029);
nand I_20276 (I346452,I346936,I346826);
not I_20277 (I347107,I2357);
not I_20278 (I347124,I155599);
nor I_20279 (I347141,I155605,I155584);
nand I_20280 (I347158,I347141,I155590);
nor I_20281 (I347175,I347124,I155605);
nand I_20282 (I347192,I347175,I155596);
not I_20283 (I347209,I155605);
not I_20284 (I347226,I347209);
not I_20285 (I347243,I155593);
nor I_20286 (I347260,I347243,I155611);
and I_20287 (I347277,I347260,I155602);
or I_20288 (I347294,I347277,I155581);
DFFARX1 I_20289  ( .D(I347294), .CLK(I2350), .RSTB(I347107), .Q(I347311) );
nand I_20290 (I347328,I347124,I155593);
or I_20291 (I347096,I347328,I347311);
not I_20292 (I347359,I347328);
nor I_20293 (I347376,I347311,I347359);
and I_20294 (I347393,I347209,I347376);
nand I_20295 (I347069,I347328,I347226);
DFFARX1 I_20296  ( .D(I155608), .CLK(I2350), .RSTB(I347107), .Q(I347424) );
or I_20297 (I347090,I347424,I347311);
nor I_20298 (I347455,I347424,I347192);
nor I_20299 (I347472,I347424,I347226);
nand I_20300 (I347075,I347158,I347472);
or I_20301 (I347503,I347424,I347393);
DFFARX1 I_20302  ( .D(I347503), .CLK(I2350), .RSTB(I347107), .Q(I347072) );
not I_20303 (I347078,I347424);
DFFARX1 I_20304  ( .D(I155587), .CLK(I2350), .RSTB(I347107), .Q(I347548) );
not I_20305 (I347565,I347548);
nor I_20306 (I347582,I347565,I347158);
DFFARX1 I_20307  ( .D(I347582), .CLK(I2350), .RSTB(I347107), .Q(I347084) );
nor I_20308 (I347099,I347424,I347565);
nor I_20309 (I347087,I347565,I347328);
not I_20310 (I347641,I347565);
and I_20311 (I347658,I347192,I347641);
nor I_20312 (I347093,I347328,I347658);
nand I_20313 (I347081,I347565,I347455);
not I_20314 (I347736,I2357);
not I_20315 (I347753,I168196);
nor I_20316 (I347770,I168202,I168181);
nand I_20317 (I347787,I347770,I168187);
nor I_20318 (I347804,I347753,I168202);
nand I_20319 (I347821,I347804,I168193);
not I_20320 (I347838,I168202);
not I_20321 (I347855,I347838);
not I_20322 (I347872,I168190);
nor I_20323 (I347889,I347872,I168208);
and I_20324 (I347906,I347889,I168199);
or I_20325 (I347923,I347906,I168178);
DFFARX1 I_20326  ( .D(I347923), .CLK(I2350), .RSTB(I347736), .Q(I347940) );
nand I_20327 (I347957,I347753,I168190);
or I_20328 (I347725,I347957,I347940);
not I_20329 (I347988,I347957);
nor I_20330 (I348005,I347940,I347988);
and I_20331 (I348022,I347838,I348005);
nand I_20332 (I347698,I347957,I347855);
DFFARX1 I_20333  ( .D(I168205), .CLK(I2350), .RSTB(I347736), .Q(I348053) );
or I_20334 (I347719,I348053,I347940);
nor I_20335 (I348084,I348053,I347821);
nor I_20336 (I348101,I348053,I347855);
nand I_20337 (I347704,I347787,I348101);
or I_20338 (I348132,I348053,I348022);
DFFARX1 I_20339  ( .D(I348132), .CLK(I2350), .RSTB(I347736), .Q(I347701) );
not I_20340 (I347707,I348053);
DFFARX1 I_20341  ( .D(I168184), .CLK(I2350), .RSTB(I347736), .Q(I348177) );
not I_20342 (I348194,I348177);
nor I_20343 (I348211,I348194,I347787);
DFFARX1 I_20344  ( .D(I348211), .CLK(I2350), .RSTB(I347736), .Q(I347713) );
nor I_20345 (I347728,I348053,I348194);
nor I_20346 (I347716,I348194,I347957);
not I_20347 (I348270,I348194);
and I_20348 (I348287,I347821,I348270);
nor I_20349 (I347722,I347957,I348287);
nand I_20350 (I347710,I348194,I348084);
not I_20351 (I348365,I2357);
not I_20352 (I348382,I33680);
nor I_20353 (I348399,I33698,I33677);
nand I_20354 (I348416,I348399,I33695);
nor I_20355 (I348433,I348382,I33698);
nand I_20356 (I348450,I348433,I33689);
not I_20357 (I348467,I33698);
not I_20358 (I348484,I348467);
not I_20359 (I348501,I33692);
nor I_20360 (I348518,I348501,I33686);
and I_20361 (I348535,I348518,I33683);
or I_20362 (I348552,I348535,I33674);
DFFARX1 I_20363  ( .D(I348552), .CLK(I2350), .RSTB(I348365), .Q(I348569) );
nand I_20364 (I348586,I348382,I33692);
or I_20365 (I348354,I348586,I348569);
not I_20366 (I348617,I348586);
nor I_20367 (I348634,I348569,I348617);
and I_20368 (I348651,I348467,I348634);
nand I_20369 (I348327,I348586,I348484);
DFFARX1 I_20370  ( .D(I33704), .CLK(I2350), .RSTB(I348365), .Q(I348682) );
or I_20371 (I348348,I348682,I348569);
nor I_20372 (I348713,I348682,I348450);
nor I_20373 (I348730,I348682,I348484);
nand I_20374 (I348333,I348416,I348730);
or I_20375 (I348761,I348682,I348651);
DFFARX1 I_20376  ( .D(I348761), .CLK(I2350), .RSTB(I348365), .Q(I348330) );
not I_20377 (I348336,I348682);
DFFARX1 I_20378  ( .D(I33701), .CLK(I2350), .RSTB(I348365), .Q(I348806) );
not I_20379 (I348823,I348806);
nor I_20380 (I348840,I348823,I348416);
DFFARX1 I_20381  ( .D(I348840), .CLK(I2350), .RSTB(I348365), .Q(I348342) );
nor I_20382 (I348357,I348682,I348823);
nor I_20383 (I348345,I348823,I348586);
not I_20384 (I348899,I348823);
and I_20385 (I348916,I348450,I348899);
nor I_20386 (I348351,I348586,I348916);
nand I_20387 (I348339,I348823,I348713);
not I_20388 (I348994,I2357);
not I_20389 (I349011,I156262);
nor I_20390 (I349028,I156268,I156247);
nand I_20391 (I349045,I349028,I156253);
nor I_20392 (I349062,I349011,I156268);
nand I_20393 (I349079,I349062,I156259);
not I_20394 (I349096,I156268);
not I_20395 (I349113,I349096);
not I_20396 (I349130,I156256);
nor I_20397 (I349147,I349130,I156274);
and I_20398 (I349164,I349147,I156265);
or I_20399 (I349181,I349164,I156244);
DFFARX1 I_20400  ( .D(I349181), .CLK(I2350), .RSTB(I348994), .Q(I349198) );
nand I_20401 (I349215,I349011,I156256);
or I_20402 (I348983,I349215,I349198);
not I_20403 (I349246,I349215);
nor I_20404 (I349263,I349198,I349246);
and I_20405 (I349280,I349096,I349263);
nand I_20406 (I348956,I349215,I349113);
DFFARX1 I_20407  ( .D(I156271), .CLK(I2350), .RSTB(I348994), .Q(I349311) );
or I_20408 (I348977,I349311,I349198);
nor I_20409 (I349342,I349311,I349079);
nor I_20410 (I349359,I349311,I349113);
nand I_20411 (I348962,I349045,I349359);
or I_20412 (I349390,I349311,I349280);
DFFARX1 I_20413  ( .D(I349390), .CLK(I2350), .RSTB(I348994), .Q(I348959) );
not I_20414 (I348965,I349311);
DFFARX1 I_20415  ( .D(I156250), .CLK(I2350), .RSTB(I348994), .Q(I349435) );
not I_20416 (I349452,I349435);
nor I_20417 (I349469,I349452,I349045);
DFFARX1 I_20418  ( .D(I349469), .CLK(I2350), .RSTB(I348994), .Q(I348971) );
nor I_20419 (I348986,I349311,I349452);
nor I_20420 (I348974,I349452,I349215);
not I_20421 (I349528,I349452);
and I_20422 (I349545,I349079,I349528);
nor I_20423 (I348980,I349215,I349545);
nand I_20424 (I348968,I349452,I349342);
not I_20425 (I349623,I2357);
not I_20426 (I349640,I171511);
nor I_20427 (I349657,I171517,I171496);
nand I_20428 (I349674,I349657,I171502);
nor I_20429 (I349691,I349640,I171517);
nand I_20430 (I349708,I349691,I171508);
not I_20431 (I349725,I171517);
not I_20432 (I349742,I349725);
not I_20433 (I349759,I171505);
nor I_20434 (I349776,I349759,I171523);
and I_20435 (I349793,I349776,I171514);
or I_20436 (I349810,I349793,I171493);
DFFARX1 I_20437  ( .D(I349810), .CLK(I2350), .RSTB(I349623), .Q(I349827) );
nand I_20438 (I349844,I349640,I171505);
or I_20439 (I349612,I349844,I349827);
not I_20440 (I349875,I349844);
nor I_20441 (I349892,I349827,I349875);
and I_20442 (I349909,I349725,I349892);
nand I_20443 (I349585,I349844,I349742);
DFFARX1 I_20444  ( .D(I171520), .CLK(I2350), .RSTB(I349623), .Q(I349940) );
or I_20445 (I349606,I349940,I349827);
nor I_20446 (I349971,I349940,I349708);
nor I_20447 (I349988,I349940,I349742);
nand I_20448 (I349591,I349674,I349988);
or I_20449 (I350019,I349940,I349909);
DFFARX1 I_20450  ( .D(I350019), .CLK(I2350), .RSTB(I349623), .Q(I349588) );
not I_20451 (I349594,I349940);
DFFARX1 I_20452  ( .D(I171499), .CLK(I2350), .RSTB(I349623), .Q(I350064) );
not I_20453 (I350081,I350064);
nor I_20454 (I350098,I350081,I349674);
DFFARX1 I_20455  ( .D(I350098), .CLK(I2350), .RSTB(I349623), .Q(I349600) );
nor I_20456 (I349615,I349940,I350081);
nor I_20457 (I349603,I350081,I349844);
not I_20458 (I350157,I350081);
and I_20459 (I350174,I349708,I350157);
nor I_20460 (I349609,I349844,I350174);
nand I_20461 (I349597,I350081,I349971);
not I_20462 (I350252,I2357);
not I_20463 (I350269,I6290);
nor I_20464 (I350286,I6293,I6302);
nand I_20465 (I350303,I350286,I6317);
nor I_20466 (I350320,I350269,I6293);
nand I_20467 (I350337,I350320,I6296);
not I_20468 (I350354,I6293);
not I_20469 (I350371,I350354);
not I_20470 (I350388,I6287);
nor I_20471 (I350405,I350388,I6311);
and I_20472 (I350422,I350405,I6299);
or I_20473 (I350439,I350422,I6305);
DFFARX1 I_20474  ( .D(I350439), .CLK(I2350), .RSTB(I350252), .Q(I350456) );
nand I_20475 (I350473,I350269,I6287);
or I_20476 (I350241,I350473,I350456);
not I_20477 (I350504,I350473);
nor I_20478 (I350521,I350456,I350504);
and I_20479 (I350538,I350354,I350521);
nand I_20480 (I350214,I350473,I350371);
DFFARX1 I_20481  ( .D(I6308), .CLK(I2350), .RSTB(I350252), .Q(I350569) );
or I_20482 (I350235,I350569,I350456);
nor I_20483 (I350600,I350569,I350337);
nor I_20484 (I350617,I350569,I350371);
nand I_20485 (I350220,I350303,I350617);
or I_20486 (I350648,I350569,I350538);
DFFARX1 I_20487  ( .D(I350648), .CLK(I2350), .RSTB(I350252), .Q(I350217) );
not I_20488 (I350223,I350569);
DFFARX1 I_20489  ( .D(I6314), .CLK(I2350), .RSTB(I350252), .Q(I350693) );
not I_20490 (I350710,I350693);
nor I_20491 (I350727,I350710,I350303);
DFFARX1 I_20492  ( .D(I350727), .CLK(I2350), .RSTB(I350252), .Q(I350229) );
nor I_20493 (I350244,I350569,I350710);
nor I_20494 (I350232,I350710,I350473);
not I_20495 (I350786,I350710);
and I_20496 (I350803,I350337,I350786);
nor I_20497 (I350238,I350473,I350803);
nand I_20498 (I350226,I350710,I350600);
not I_20499 (I350881,I2357);
not I_20500 (I350898,I162892);
nor I_20501 (I350915,I162898,I162877);
nand I_20502 (I350932,I350915,I162883);
nor I_20503 (I350949,I350898,I162898);
nand I_20504 (I350966,I350949,I162889);
not I_20505 (I350983,I162898);
not I_20506 (I351000,I350983);
not I_20507 (I351017,I162886);
nor I_20508 (I351034,I351017,I162904);
and I_20509 (I351051,I351034,I162895);
or I_20510 (I351068,I351051,I162874);
DFFARX1 I_20511  ( .D(I351068), .CLK(I2350), .RSTB(I350881), .Q(I351085) );
nand I_20512 (I351102,I350898,I162886);
or I_20513 (I350870,I351102,I351085);
not I_20514 (I351133,I351102);
nor I_20515 (I351150,I351085,I351133);
and I_20516 (I351167,I350983,I351150);
nand I_20517 (I350843,I351102,I351000);
DFFARX1 I_20518  ( .D(I162901), .CLK(I2350), .RSTB(I350881), .Q(I351198) );
or I_20519 (I350864,I351198,I351085);
nor I_20520 (I351229,I351198,I350966);
nor I_20521 (I351246,I351198,I351000);
nand I_20522 (I350849,I350932,I351246);
or I_20523 (I351277,I351198,I351167);
DFFARX1 I_20524  ( .D(I351277), .CLK(I2350), .RSTB(I350881), .Q(I350846) );
not I_20525 (I350852,I351198);
DFFARX1 I_20526  ( .D(I162880), .CLK(I2350), .RSTB(I350881), .Q(I351322) );
not I_20527 (I351339,I351322);
nor I_20528 (I351356,I351339,I350932);
DFFARX1 I_20529  ( .D(I351356), .CLK(I2350), .RSTB(I350881), .Q(I350858) );
nor I_20530 (I350873,I351198,I351339);
nor I_20531 (I350861,I351339,I351102);
not I_20532 (I351415,I351339);
and I_20533 (I351432,I350966,I351415);
nor I_20534 (I350867,I351102,I351432);
nand I_20535 (I350855,I351339,I351229);
not I_20536 (I351510,I2357);
not I_20537 (I351527,I142339);
nor I_20538 (I351544,I142345,I142324);
nand I_20539 (I351561,I351544,I142330);
nor I_20540 (I351578,I351527,I142345);
nand I_20541 (I351595,I351578,I142336);
not I_20542 (I351612,I142345);
not I_20543 (I351629,I351612);
not I_20544 (I351646,I142333);
nor I_20545 (I351663,I351646,I142351);
and I_20546 (I351680,I351663,I142342);
or I_20547 (I351697,I351680,I142321);
DFFARX1 I_20548  ( .D(I351697), .CLK(I2350), .RSTB(I351510), .Q(I351714) );
nand I_20549 (I351731,I351527,I142333);
or I_20550 (I351499,I351731,I351714);
not I_20551 (I351762,I351731);
nor I_20552 (I351779,I351714,I351762);
and I_20553 (I351796,I351612,I351779);
nand I_20554 (I351472,I351731,I351629);
DFFARX1 I_20555  ( .D(I142348), .CLK(I2350), .RSTB(I351510), .Q(I351827) );
or I_20556 (I351493,I351827,I351714);
nor I_20557 (I351858,I351827,I351595);
nor I_20558 (I351875,I351827,I351629);
nand I_20559 (I351478,I351561,I351875);
or I_20560 (I351906,I351827,I351796);
DFFARX1 I_20561  ( .D(I351906), .CLK(I2350), .RSTB(I351510), .Q(I351475) );
not I_20562 (I351481,I351827);
DFFARX1 I_20563  ( .D(I142327), .CLK(I2350), .RSTB(I351510), .Q(I351951) );
not I_20564 (I351968,I351951);
nor I_20565 (I351985,I351968,I351561);
DFFARX1 I_20566  ( .D(I351985), .CLK(I2350), .RSTB(I351510), .Q(I351487) );
nor I_20567 (I351502,I351827,I351968);
nor I_20568 (I351490,I351968,I351731);
not I_20569 (I352044,I351968);
and I_20570 (I352061,I351595,I352044);
nor I_20571 (I351496,I351731,I352061);
nand I_20572 (I351484,I351968,I351858);
not I_20573 (I352139,I2357);
not I_20574 (I352156,I223089);
nor I_20575 (I352173,I223098,I223101);
nand I_20576 (I352190,I352173,I223086);
nor I_20577 (I352207,I352156,I223098);
nand I_20578 (I352224,I352207,I223083);
not I_20579 (I352241,I223098);
not I_20580 (I352258,I352241);
not I_20581 (I352275,I223071);
nor I_20582 (I352292,I352275,I223077);
and I_20583 (I352309,I352292,I223074);
or I_20584 (I352326,I352309,I223095);
DFFARX1 I_20585  ( .D(I352326), .CLK(I2350), .RSTB(I352139), .Q(I352343) );
nand I_20586 (I352360,I352156,I223071);
or I_20587 (I352128,I352360,I352343);
not I_20588 (I352391,I352360);
nor I_20589 (I352408,I352343,I352391);
and I_20590 (I352425,I352241,I352408);
nand I_20591 (I352101,I352360,I352258);
DFFARX1 I_20592  ( .D(I223080), .CLK(I2350), .RSTB(I352139), .Q(I352456) );
or I_20593 (I352122,I352456,I352343);
nor I_20594 (I352487,I352456,I352224);
nor I_20595 (I352504,I352456,I352258);
nand I_20596 (I352107,I352190,I352504);
or I_20597 (I352535,I352456,I352425);
DFFARX1 I_20598  ( .D(I352535), .CLK(I2350), .RSTB(I352139), .Q(I352104) );
not I_20599 (I352110,I352456);
DFFARX1 I_20600  ( .D(I223092), .CLK(I2350), .RSTB(I352139), .Q(I352580) );
not I_20601 (I352597,I352580);
nor I_20602 (I352614,I352597,I352190);
DFFARX1 I_20603  ( .D(I352614), .CLK(I2350), .RSTB(I352139), .Q(I352116) );
nor I_20604 (I352131,I352456,I352597);
nor I_20605 (I352119,I352597,I352360);
not I_20606 (I352673,I352597);
and I_20607 (I352690,I352224,I352673);
nor I_20608 (I352125,I352360,I352690);
nand I_20609 (I352113,I352597,I352487);
not I_20610 (I352768,I2357);
not I_20611 (I352785,I238275);
nor I_20612 (I352802,I238299,I238278);
nand I_20613 (I352819,I352802,I238284);
nor I_20614 (I352836,I352785,I238299);
nand I_20615 (I352853,I352836,I238296);
not I_20616 (I352870,I238299);
not I_20617 (I352887,I352870);
not I_20618 (I352904,I238293);
nor I_20619 (I352921,I352904,I238272);
and I_20620 (I352938,I352921,I238269);
or I_20621 (I352955,I352938,I238281);
DFFARX1 I_20622  ( .D(I352955), .CLK(I2350), .RSTB(I352768), .Q(I352972) );
nand I_20623 (I352989,I352785,I238293);
or I_20624 (I352757,I352989,I352972);
not I_20625 (I353020,I352989);
nor I_20626 (I353037,I352972,I353020);
and I_20627 (I353054,I352870,I353037);
nand I_20628 (I352730,I352989,I352887);
DFFARX1 I_20629  ( .D(I238287), .CLK(I2350), .RSTB(I352768), .Q(I353085) );
or I_20630 (I352751,I353085,I352972);
nor I_20631 (I353116,I353085,I352853);
nor I_20632 (I353133,I353085,I352887);
nand I_20633 (I352736,I352819,I353133);
or I_20634 (I353164,I353085,I353054);
DFFARX1 I_20635  ( .D(I353164), .CLK(I2350), .RSTB(I352768), .Q(I352733) );
not I_20636 (I352739,I353085);
DFFARX1 I_20637  ( .D(I238290), .CLK(I2350), .RSTB(I352768), .Q(I353209) );
not I_20638 (I353226,I353209);
nor I_20639 (I353243,I353226,I352819);
DFFARX1 I_20640  ( .D(I353243), .CLK(I2350), .RSTB(I352768), .Q(I352745) );
nor I_20641 (I352760,I353085,I353226);
nor I_20642 (I352748,I353226,I352989);
not I_20643 (I353302,I353226);
and I_20644 (I353319,I352853,I353302);
nor I_20645 (I352754,I352989,I353319);
nand I_20646 (I352742,I353226,I353116);
not I_20647 (I353397,I2357);
not I_20648 (I353414,I309403);
nor I_20649 (I353431,I309421,I309400);
nand I_20650 (I353448,I353431,I309424);
nor I_20651 (I353465,I353414,I309421);
nand I_20652 (I353482,I353465,I309418);
not I_20653 (I353499,I309421);
not I_20654 (I353516,I353499);
not I_20655 (I353533,I309409);
nor I_20656 (I353550,I353533,I309397);
and I_20657 (I353567,I353550,I309415);
or I_20658 (I353584,I353567,I309427);
DFFARX1 I_20659  ( .D(I353584), .CLK(I2350), .RSTB(I353397), .Q(I353601) );
nand I_20660 (I353618,I353414,I309409);
or I_20661 (I353386,I353618,I353601);
not I_20662 (I353649,I353618);
nor I_20663 (I353666,I353601,I353649);
and I_20664 (I353683,I353499,I353666);
nand I_20665 (I353359,I353618,I353516);
DFFARX1 I_20666  ( .D(I309406), .CLK(I2350), .RSTB(I353397), .Q(I353714) );
or I_20667 (I353380,I353714,I353601);
nor I_20668 (I353745,I353714,I353482);
nor I_20669 (I353762,I353714,I353516);
nand I_20670 (I353365,I353448,I353762);
or I_20671 (I353793,I353714,I353683);
DFFARX1 I_20672  ( .D(I353793), .CLK(I2350), .RSTB(I353397), .Q(I353362) );
not I_20673 (I353368,I353714);
DFFARX1 I_20674  ( .D(I309412), .CLK(I2350), .RSTB(I353397), .Q(I353838) );
not I_20675 (I353855,I353838);
nor I_20676 (I353872,I353855,I353448);
DFFARX1 I_20677  ( .D(I353872), .CLK(I2350), .RSTB(I353397), .Q(I353374) );
nor I_20678 (I353389,I353714,I353855);
nor I_20679 (I353377,I353855,I353618);
not I_20680 (I353931,I353855);
and I_20681 (I353948,I353482,I353931);
nor I_20682 (I353383,I353618,I353948);
nand I_20683 (I353371,I353855,I353745);
not I_20684 (I354026,I2357);
not I_20685 (I354043,I1967);
nor I_20686 (I354060,I1719,I1351);
nand I_20687 (I354077,I354060,I1447);
nor I_20688 (I354094,I354043,I1719);
nand I_20689 (I354111,I354094,I2135);
not I_20690 (I354128,I1719);
not I_20691 (I354145,I354128);
not I_20692 (I354162,I2151);
nor I_20693 (I354179,I354162,I1407);
and I_20694 (I354196,I354179,I1703);
or I_20695 (I354213,I354196,I2087);
DFFARX1 I_20696  ( .D(I354213), .CLK(I2350), .RSTB(I354026), .Q(I354230) );
nand I_20697 (I354247,I354043,I2151);
or I_20698 (I354015,I354247,I354230);
not I_20699 (I354278,I354247);
nor I_20700 (I354295,I354230,I354278);
and I_20701 (I354312,I354128,I354295);
nand I_20702 (I353988,I354247,I354145);
DFFARX1 I_20703  ( .D(I1207), .CLK(I2350), .RSTB(I354026), .Q(I354343) );
or I_20704 (I354009,I354343,I354230);
nor I_20705 (I354374,I354343,I354111);
nor I_20706 (I354391,I354343,I354145);
nand I_20707 (I353994,I354077,I354391);
or I_20708 (I354422,I354343,I354312);
DFFARX1 I_20709  ( .D(I354422), .CLK(I2350), .RSTB(I354026), .Q(I353991) );
not I_20710 (I353997,I354343);
DFFARX1 I_20711  ( .D(I2215), .CLK(I2350), .RSTB(I354026), .Q(I354467) );
not I_20712 (I354484,I354467);
nor I_20713 (I354501,I354484,I354077);
DFFARX1 I_20714  ( .D(I354501), .CLK(I2350), .RSTB(I354026), .Q(I354003) );
nor I_20715 (I354018,I354343,I354484);
nor I_20716 (I354006,I354484,I354247);
not I_20717 (I354560,I354484);
and I_20718 (I354577,I354111,I354560);
nor I_20719 (I354012,I354247,I354577);
nand I_20720 (I354000,I354484,I354374);
not I_20721 (I354655,I2357);
not I_20722 (I354672,I286793);
nor I_20723 (I354689,I286811,I286790);
nand I_20724 (I354706,I354689,I286814);
nor I_20725 (I354723,I354672,I286811);
nand I_20726 (I354740,I354723,I286808);
not I_20727 (I354757,I286811);
not I_20728 (I354774,I354757);
not I_20729 (I354791,I286799);
nor I_20730 (I354808,I354791,I286787);
and I_20731 (I354825,I354808,I286805);
or I_20732 (I354842,I354825,I286817);
DFFARX1 I_20733  ( .D(I354842), .CLK(I2350), .RSTB(I354655), .Q(I354859) );
nand I_20734 (I354876,I354672,I286799);
or I_20735 (I354644,I354876,I354859);
not I_20736 (I354907,I354876);
nor I_20737 (I354924,I354859,I354907);
and I_20738 (I354941,I354757,I354924);
nand I_20739 (I354617,I354876,I354774);
DFFARX1 I_20740  ( .D(I286796), .CLK(I2350), .RSTB(I354655), .Q(I354972) );
or I_20741 (I354638,I354972,I354859);
nor I_20742 (I355003,I354972,I354740);
nor I_20743 (I355020,I354972,I354774);
nand I_20744 (I354623,I354706,I355020);
or I_20745 (I355051,I354972,I354941);
DFFARX1 I_20746  ( .D(I355051), .CLK(I2350), .RSTB(I354655), .Q(I354620) );
not I_20747 (I354626,I354972);
DFFARX1 I_20748  ( .D(I286802), .CLK(I2350), .RSTB(I354655), .Q(I355096) );
not I_20749 (I355113,I355096);
nor I_20750 (I355130,I355113,I354706);
DFFARX1 I_20751  ( .D(I355130), .CLK(I2350), .RSTB(I354655), .Q(I354632) );
nor I_20752 (I354647,I354972,I355113);
nor I_20753 (I354635,I355113,I354876);
not I_20754 (I355189,I355113);
and I_20755 (I355206,I354740,I355189);
nor I_20756 (I354641,I354876,I355206);
nand I_20757 (I354629,I355113,I355003);
not I_20758 (I355284,I2357);
not I_20759 (I355301,I221151);
nor I_20760 (I355318,I221160,I221163);
nand I_20761 (I355335,I355318,I221148);
nor I_20762 (I355352,I355301,I221160);
nand I_20763 (I355369,I355352,I221145);
not I_20764 (I355386,I221160);
not I_20765 (I355403,I355386);
not I_20766 (I355420,I221133);
nor I_20767 (I355437,I355420,I221139);
and I_20768 (I355454,I355437,I221136);
or I_20769 (I355471,I355454,I221157);
DFFARX1 I_20770  ( .D(I355471), .CLK(I2350), .RSTB(I355284), .Q(I355488) );
nand I_20771 (I355505,I355301,I221133);
or I_20772 (I355273,I355505,I355488);
not I_20773 (I355536,I355505);
nor I_20774 (I355553,I355488,I355536);
and I_20775 (I355570,I355386,I355553);
nand I_20776 (I355246,I355505,I355403);
DFFARX1 I_20777  ( .D(I221142), .CLK(I2350), .RSTB(I355284), .Q(I355601) );
or I_20778 (I355267,I355601,I355488);
nor I_20779 (I355632,I355601,I355369);
nor I_20780 (I355649,I355601,I355403);
nand I_20781 (I355252,I355335,I355649);
or I_20782 (I355680,I355601,I355570);
DFFARX1 I_20783  ( .D(I355680), .CLK(I2350), .RSTB(I355284), .Q(I355249) );
not I_20784 (I355255,I355601);
DFFARX1 I_20785  ( .D(I221154), .CLK(I2350), .RSTB(I355284), .Q(I355725) );
not I_20786 (I355742,I355725);
nor I_20787 (I355759,I355742,I355335);
DFFARX1 I_20788  ( .D(I355759), .CLK(I2350), .RSTB(I355284), .Q(I355261) );
nor I_20789 (I355276,I355601,I355742);
nor I_20790 (I355264,I355742,I355505);
not I_20791 (I355818,I355742);
and I_20792 (I355835,I355369,I355818);
nor I_20793 (I355270,I355505,I355835);
nand I_20794 (I355258,I355742,I355632);
not I_20795 (I355913,I2357);
not I_20796 (I355930,I1423);
nor I_20797 (I355947,I1639,I1647);
nand I_20798 (I355964,I355947,I2015);
nor I_20799 (I355981,I355930,I1639);
nand I_20800 (I355998,I355981,I1311);
not I_20801 (I356015,I1639);
not I_20802 (I356032,I356015);
not I_20803 (I356049,I1279);
nor I_20804 (I356066,I356049,I1271);
and I_20805 (I356083,I356066,I1471);
or I_20806 (I356100,I356083,I1231);
DFFARX1 I_20807  ( .D(I356100), .CLK(I2350), .RSTB(I355913), .Q(I356117) );
nand I_20808 (I356134,I355930,I1279);
or I_20809 (I355902,I356134,I356117);
not I_20810 (I356165,I356134);
nor I_20811 (I356182,I356117,I356165);
and I_20812 (I356199,I356015,I356182);
nand I_20813 (I355875,I356134,I356032);
DFFARX1 I_20814  ( .D(I1799), .CLK(I2350), .RSTB(I355913), .Q(I356230) );
or I_20815 (I355896,I356230,I356117);
nor I_20816 (I356261,I356230,I355998);
nor I_20817 (I356278,I356230,I356032);
nand I_20818 (I355881,I355964,I356278);
or I_20819 (I356309,I356230,I356199);
DFFARX1 I_20820  ( .D(I356309), .CLK(I2350), .RSTB(I355913), .Q(I355878) );
not I_20821 (I355884,I356230);
DFFARX1 I_20822  ( .D(I1399), .CLK(I2350), .RSTB(I355913), .Q(I356354) );
not I_20823 (I356371,I356354);
nor I_20824 (I356388,I356371,I355964);
DFFARX1 I_20825  ( .D(I356388), .CLK(I2350), .RSTB(I355913), .Q(I355890) );
nor I_20826 (I355905,I356230,I356371);
nor I_20827 (I355893,I356371,I356134);
not I_20828 (I356447,I356371);
and I_20829 (I356464,I355998,I356447);
nor I_20830 (I355899,I356134,I356464);
nand I_20831 (I355887,I356371,I356261);
not I_20832 (I356542,I2357);
not I_20833 (I356559,I104610);
nor I_20834 (I356576,I104601,I104625);
nand I_20835 (I356593,I356576,I104628);
nor I_20836 (I356610,I356559,I104601);
nand I_20837 (I356627,I356610,I104619);
not I_20838 (I356644,I104601);
not I_20839 (I356661,I356644);
not I_20840 (I356678,I104613);
nor I_20841 (I356695,I356678,I104607);
and I_20842 (I356712,I356695,I104616);
or I_20843 (I356729,I356712,I104604);
DFFARX1 I_20844  ( .D(I356729), .CLK(I2350), .RSTB(I356542), .Q(I356746) );
nand I_20845 (I356763,I356559,I104613);
or I_20846 (I356531,I356763,I356746);
not I_20847 (I356794,I356763);
nor I_20848 (I356811,I356746,I356794);
and I_20849 (I356828,I356644,I356811);
nand I_20850 (I356504,I356763,I356661);
DFFARX1 I_20851  ( .D(I104598), .CLK(I2350), .RSTB(I356542), .Q(I356859) );
or I_20852 (I356525,I356859,I356746);
nor I_20853 (I356890,I356859,I356627);
nor I_20854 (I356907,I356859,I356661);
nand I_20855 (I356510,I356593,I356907);
or I_20856 (I356938,I356859,I356828);
DFFARX1 I_20857  ( .D(I356938), .CLK(I2350), .RSTB(I356542), .Q(I356507) );
not I_20858 (I356513,I356859);
DFFARX1 I_20859  ( .D(I104622), .CLK(I2350), .RSTB(I356542), .Q(I356983) );
not I_20860 (I357000,I356983);
nor I_20861 (I357017,I357000,I356593);
DFFARX1 I_20862  ( .D(I357017), .CLK(I2350), .RSTB(I356542), .Q(I356519) );
nor I_20863 (I356534,I356859,I357000);
nor I_20864 (I356522,I357000,I356763);
not I_20865 (I357076,I357000);
and I_20866 (I357093,I356627,I357076);
nor I_20867 (I356528,I356763,I357093);
nand I_20868 (I356516,I357000,I356890);
not I_20869 (I357171,I2357);
not I_20870 (I357188,I28512);
nor I_20871 (I357205,I28530,I28509);
nand I_20872 (I357222,I357205,I28527);
nor I_20873 (I357239,I357188,I28530);
nand I_20874 (I357256,I357239,I28521);
not I_20875 (I357273,I28530);
not I_20876 (I357290,I357273);
not I_20877 (I357307,I28524);
nor I_20878 (I357324,I357307,I28518);
and I_20879 (I357341,I357324,I28515);
or I_20880 (I357358,I357341,I28506);
DFFARX1 I_20881  ( .D(I357358), .CLK(I2350), .RSTB(I357171), .Q(I357375) );
nand I_20882 (I357392,I357188,I28524);
or I_20883 (I357160,I357392,I357375);
not I_20884 (I357423,I357392);
nor I_20885 (I357440,I357375,I357423);
and I_20886 (I357457,I357273,I357440);
nand I_20887 (I357133,I357392,I357290);
DFFARX1 I_20888  ( .D(I28536), .CLK(I2350), .RSTB(I357171), .Q(I357488) );
or I_20889 (I357154,I357488,I357375);
nor I_20890 (I357519,I357488,I357256);
nor I_20891 (I357536,I357488,I357290);
nand I_20892 (I357139,I357222,I357536);
or I_20893 (I357567,I357488,I357457);
DFFARX1 I_20894  ( .D(I357567), .CLK(I2350), .RSTB(I357171), .Q(I357136) );
not I_20895 (I357142,I357488);
DFFARX1 I_20896  ( .D(I28533), .CLK(I2350), .RSTB(I357171), .Q(I357612) );
not I_20897 (I357629,I357612);
nor I_20898 (I357646,I357629,I357222);
DFFARX1 I_20899  ( .D(I357646), .CLK(I2350), .RSTB(I357171), .Q(I357148) );
nor I_20900 (I357163,I357488,I357629);
nor I_20901 (I357151,I357629,I357392);
not I_20902 (I357705,I357629);
and I_20903 (I357722,I357256,I357705);
nor I_20904 (I357157,I357392,I357722);
nand I_20905 (I357145,I357629,I357519);
not I_20906 (I357800,I2357);
not I_20907 (I357817,I97980);
nor I_20908 (I357834,I97971,I97995);
nand I_20909 (I357851,I357834,I97998);
nor I_20910 (I357868,I357817,I97971);
nand I_20911 (I357885,I357868,I97989);
not I_20912 (I357902,I97971);
not I_20913 (I357919,I357902);
not I_20914 (I357936,I97983);
nor I_20915 (I357953,I357936,I97977);
and I_20916 (I357970,I357953,I97986);
or I_20917 (I357987,I357970,I97974);
DFFARX1 I_20918  ( .D(I357987), .CLK(I2350), .RSTB(I357800), .Q(I358004) );
nand I_20919 (I358021,I357817,I97983);
or I_20920 (I357789,I358021,I358004);
not I_20921 (I358052,I358021);
nor I_20922 (I358069,I358004,I358052);
and I_20923 (I358086,I357902,I358069);
nand I_20924 (I357762,I358021,I357919);
DFFARX1 I_20925  ( .D(I97968), .CLK(I2350), .RSTB(I357800), .Q(I358117) );
or I_20926 (I357783,I358117,I358004);
nor I_20927 (I358148,I358117,I357885);
nor I_20928 (I358165,I358117,I357919);
nand I_20929 (I357768,I357851,I358165);
or I_20930 (I358196,I358117,I358086);
DFFARX1 I_20931  ( .D(I358196), .CLK(I2350), .RSTB(I357800), .Q(I357765) );
not I_20932 (I357771,I358117);
DFFARX1 I_20933  ( .D(I97992), .CLK(I2350), .RSTB(I357800), .Q(I358241) );
not I_20934 (I358258,I358241);
nor I_20935 (I358275,I358258,I357851);
DFFARX1 I_20936  ( .D(I358275), .CLK(I2350), .RSTB(I357800), .Q(I357777) );
nor I_20937 (I357792,I358117,I358258);
nor I_20938 (I357780,I358258,I358021);
not I_20939 (I358334,I358258);
and I_20940 (I358351,I357885,I358334);
nor I_20941 (I357786,I358021,I358351);
nand I_20942 (I357774,I358258,I358148);
not I_20943 (I358429,I2357);
not I_20944 (I358446,I282628);
nor I_20945 (I358463,I282646,I282625);
nand I_20946 (I358480,I358463,I282649);
nor I_20947 (I358497,I358446,I282646);
nand I_20948 (I358514,I358497,I282643);
not I_20949 (I358531,I282646);
not I_20950 (I358548,I358531);
not I_20951 (I358565,I282634);
nor I_20952 (I358582,I358565,I282622);
and I_20953 (I358599,I358582,I282640);
or I_20954 (I358616,I358599,I282652);
DFFARX1 I_20955  ( .D(I358616), .CLK(I2350), .RSTB(I358429), .Q(I358633) );
nand I_20956 (I358650,I358446,I282634);
or I_20957 (I358418,I358650,I358633);
not I_20958 (I358681,I358650);
nor I_20959 (I358698,I358633,I358681);
and I_20960 (I358715,I358531,I358698);
nand I_20961 (I358391,I358650,I358548);
DFFARX1 I_20962  ( .D(I282631), .CLK(I2350), .RSTB(I358429), .Q(I358746) );
or I_20963 (I358412,I358746,I358633);
nor I_20964 (I358777,I358746,I358514);
nor I_20965 (I358794,I358746,I358548);
nand I_20966 (I358397,I358480,I358794);
or I_20967 (I358825,I358746,I358715);
DFFARX1 I_20968  ( .D(I358825), .CLK(I2350), .RSTB(I358429), .Q(I358394) );
not I_20969 (I358400,I358746);
DFFARX1 I_20970  ( .D(I282637), .CLK(I2350), .RSTB(I358429), .Q(I358870) );
not I_20971 (I358887,I358870);
nor I_20972 (I358904,I358887,I358480);
DFFARX1 I_20973  ( .D(I358904), .CLK(I2350), .RSTB(I358429), .Q(I358406) );
nor I_20974 (I358421,I358746,I358887);
nor I_20975 (I358409,I358887,I358650);
not I_20976 (I358963,I358887);
and I_20977 (I358980,I358514,I358963);
nor I_20978 (I358415,I358650,I358980);
nand I_20979 (I358403,I358887,I358777);
not I_20980 (I359058,I2357);
not I_20981 (I359075,I105936);
nor I_20982 (I359092,I105927,I105951);
nand I_20983 (I359109,I359092,I105954);
nor I_20984 (I359126,I359075,I105927);
nand I_20985 (I359143,I359126,I105945);
not I_20986 (I359160,I105927);
not I_20987 (I359177,I359160);
not I_20988 (I359194,I105939);
nor I_20989 (I359211,I359194,I105933);
and I_20990 (I359228,I359211,I105942);
or I_20991 (I359245,I359228,I105930);
DFFARX1 I_20992  ( .D(I359245), .CLK(I2350), .RSTB(I359058), .Q(I359262) );
nand I_20993 (I359279,I359075,I105939);
or I_20994 (I359047,I359279,I359262);
not I_20995 (I359310,I359279);
nor I_20996 (I359327,I359262,I359310);
and I_20997 (I359344,I359160,I359327);
nand I_20998 (I359020,I359279,I359177);
DFFARX1 I_20999  ( .D(I105924), .CLK(I2350), .RSTB(I359058), .Q(I359375) );
or I_21000 (I359041,I359375,I359262);
nor I_21001 (I359406,I359375,I359143);
nor I_21002 (I359423,I359375,I359177);
nand I_21003 (I359026,I359109,I359423);
or I_21004 (I359454,I359375,I359344);
DFFARX1 I_21005  ( .D(I359454), .CLK(I2350), .RSTB(I359058), .Q(I359023) );
not I_21006 (I359029,I359375);
DFFARX1 I_21007  ( .D(I105948), .CLK(I2350), .RSTB(I359058), .Q(I359499) );
not I_21008 (I359516,I359499);
nor I_21009 (I359533,I359516,I359109);
DFFARX1 I_21010  ( .D(I359533), .CLK(I2350), .RSTB(I359058), .Q(I359035) );
nor I_21011 (I359050,I359375,I359516);
nor I_21012 (I359038,I359516,I359279);
not I_21013 (I359592,I359516);
and I_21014 (I359609,I359143,I359592);
nor I_21015 (I359044,I359279,I359609);
nand I_21016 (I359032,I359516,I359406);
not I_21017 (I359687,I2357);
not I_21018 (I359704,I34972);
nor I_21019 (I359721,I34990,I34969);
nand I_21020 (I359738,I359721,I34987);
nor I_21021 (I359755,I359704,I34990);
nand I_21022 (I359772,I359755,I34981);
not I_21023 (I359789,I34990);
not I_21024 (I359806,I359789);
not I_21025 (I359823,I34984);
nor I_21026 (I359840,I359823,I34978);
and I_21027 (I359857,I359840,I34975);
or I_21028 (I359874,I359857,I34966);
DFFARX1 I_21029  ( .D(I359874), .CLK(I2350), .RSTB(I359687), .Q(I359891) );
nand I_21030 (I359908,I359704,I34984);
or I_21031 (I359676,I359908,I359891);
not I_21032 (I359939,I359908);
nor I_21033 (I359956,I359891,I359939);
and I_21034 (I359973,I359789,I359956);
nand I_21035 (I359649,I359908,I359806);
DFFARX1 I_21036  ( .D(I34996), .CLK(I2350), .RSTB(I359687), .Q(I360004) );
or I_21037 (I359670,I360004,I359891);
nor I_21038 (I360035,I360004,I359772);
nor I_21039 (I360052,I360004,I359806);
nand I_21040 (I359655,I359738,I360052);
or I_21041 (I360083,I360004,I359973);
DFFARX1 I_21042  ( .D(I360083), .CLK(I2350), .RSTB(I359687), .Q(I359652) );
not I_21043 (I359658,I360004);
DFFARX1 I_21044  ( .D(I34993), .CLK(I2350), .RSTB(I359687), .Q(I360128) );
not I_21045 (I360145,I360128);
nor I_21046 (I360162,I360145,I359738);
DFFARX1 I_21047  ( .D(I360162), .CLK(I2350), .RSTB(I359687), .Q(I359664) );
nor I_21048 (I359679,I360004,I360145);
nor I_21049 (I359667,I360145,I359908);
not I_21050 (I360221,I360145);
and I_21051 (I360238,I359772,I360221);
nor I_21052 (I359673,I359908,I360238);
nand I_21053 (I359661,I360145,I360035);
not I_21054 (I360316,I2357);
not I_21055 (I360333,I274429);
nor I_21056 (I360350,I274414,I274435);
nand I_21057 (I360367,I360350,I274423);
nor I_21058 (I360384,I360333,I274414);
nand I_21059 (I360401,I360384,I274411);
not I_21060 (I360418,I274414);
not I_21061 (I360435,I360418);
not I_21062 (I360452,I274438);
nor I_21063 (I360469,I360452,I274426);
and I_21064 (I360486,I360469,I274420);
or I_21065 (I360503,I360486,I274417);
DFFARX1 I_21066  ( .D(I360503), .CLK(I2350), .RSTB(I360316), .Q(I360520) );
nand I_21067 (I360537,I360333,I274438);
or I_21068 (I360305,I360537,I360520);
not I_21069 (I360568,I360537);
nor I_21070 (I360585,I360520,I360568);
and I_21071 (I360602,I360418,I360585);
nand I_21072 (I360278,I360537,I360435);
DFFARX1 I_21073  ( .D(I274441), .CLK(I2350), .RSTB(I360316), .Q(I360633) );
or I_21074 (I360299,I360633,I360520);
nor I_21075 (I360664,I360633,I360401);
nor I_21076 (I360681,I360633,I360435);
nand I_21077 (I360284,I360367,I360681);
or I_21078 (I360712,I360633,I360602);
DFFARX1 I_21079  ( .D(I360712), .CLK(I2350), .RSTB(I360316), .Q(I360281) );
not I_21080 (I360287,I360633);
DFFARX1 I_21081  ( .D(I274432), .CLK(I2350), .RSTB(I360316), .Q(I360757) );
not I_21082 (I360774,I360757);
nor I_21083 (I360791,I360774,I360367);
DFFARX1 I_21084  ( .D(I360791), .CLK(I2350), .RSTB(I360316), .Q(I360293) );
nor I_21085 (I360308,I360633,I360774);
nor I_21086 (I360296,I360774,I360537);
not I_21087 (I360850,I360774);
and I_21088 (I360867,I360401,I360850);
nor I_21089 (I360302,I360537,I360867);
nand I_21090 (I360290,I360774,I360664);
not I_21091 (I360945,I2357);
not I_21092 (I360962,I279058);
nor I_21093 (I360979,I279076,I279055);
nand I_21094 (I360996,I360979,I279079);
nor I_21095 (I361013,I360962,I279076);
nand I_21096 (I361030,I361013,I279073);
not I_21097 (I361047,I279076);
not I_21098 (I361064,I361047);
not I_21099 (I361081,I279064);
nor I_21100 (I361098,I361081,I279052);
and I_21101 (I361115,I361098,I279070);
or I_21102 (I361132,I361115,I279082);
DFFARX1 I_21103  ( .D(I361132), .CLK(I2350), .RSTB(I360945), .Q(I361149) );
nand I_21104 (I361166,I360962,I279064);
or I_21105 (I360934,I361166,I361149);
not I_21106 (I361197,I361166);
nor I_21107 (I361214,I361149,I361197);
and I_21108 (I361231,I361047,I361214);
nand I_21109 (I360907,I361166,I361064);
DFFARX1 I_21110  ( .D(I279061), .CLK(I2350), .RSTB(I360945), .Q(I361262) );
or I_21111 (I360928,I361262,I361149);
nor I_21112 (I361293,I361262,I361030);
nor I_21113 (I361310,I361262,I361064);
nand I_21114 (I360913,I360996,I361310);
or I_21115 (I361341,I361262,I361231);
DFFARX1 I_21116  ( .D(I361341), .CLK(I2350), .RSTB(I360945), .Q(I360910) );
not I_21117 (I360916,I361262);
DFFARX1 I_21118  ( .D(I279067), .CLK(I2350), .RSTB(I360945), .Q(I361386) );
not I_21119 (I361403,I361386);
nor I_21120 (I361420,I361403,I360996);
DFFARX1 I_21121  ( .D(I361420), .CLK(I2350), .RSTB(I360945), .Q(I360922) );
nor I_21122 (I360937,I361262,I361403);
nor I_21123 (I360925,I361403,I361166);
not I_21124 (I361479,I361403);
and I_21125 (I361496,I361030,I361479);
nor I_21126 (I360931,I361166,I361496);
nand I_21127 (I360919,I361403,I361293);
not I_21128 (I361574,I2357);
not I_21129 (I361591,I15827);
nor I_21130 (I361608,I15830,I15839);
nand I_21131 (I361625,I361608,I15854);
nor I_21132 (I361642,I361591,I15830);
nand I_21133 (I361659,I361642,I15833);
not I_21134 (I361676,I15830);
not I_21135 (I361693,I361676);
not I_21136 (I361710,I15824);
nor I_21137 (I361727,I361710,I15848);
and I_21138 (I361744,I361727,I15836);
or I_21139 (I361761,I361744,I15842);
DFFARX1 I_21140  ( .D(I361761), .CLK(I2350), .RSTB(I361574), .Q(I361778) );
nand I_21141 (I361795,I361591,I15824);
or I_21142 (I361563,I361795,I361778);
not I_21143 (I361826,I361795);
nor I_21144 (I361843,I361778,I361826);
and I_21145 (I361860,I361676,I361843);
nand I_21146 (I361536,I361795,I361693);
DFFARX1 I_21147  ( .D(I15845), .CLK(I2350), .RSTB(I361574), .Q(I361891) );
or I_21148 (I361557,I361891,I361778);
nor I_21149 (I361922,I361891,I361659);
nor I_21150 (I361939,I361891,I361693);
nand I_21151 (I361542,I361625,I361939);
or I_21152 (I361970,I361891,I361860);
DFFARX1 I_21153  ( .D(I361970), .CLK(I2350), .RSTB(I361574), .Q(I361539) );
not I_21154 (I361545,I361891);
DFFARX1 I_21155  ( .D(I15851), .CLK(I2350), .RSTB(I361574), .Q(I362015) );
not I_21156 (I362032,I362015);
nor I_21157 (I362049,I362032,I361625);
DFFARX1 I_21158  ( .D(I362049), .CLK(I2350), .RSTB(I361574), .Q(I361551) );
nor I_21159 (I361566,I361891,I362032);
nor I_21160 (I361554,I362032,I361795);
not I_21161 (I362108,I362032);
and I_21162 (I362125,I361659,I362108);
nor I_21163 (I361560,I361795,I362125);
nand I_21164 (I361548,I362032,I361922);
not I_21165 (I362203,I2357);
not I_21166 (I362220,I243535);
nor I_21167 (I362237,I243508,I243526);
nand I_21168 (I362254,I362237,I243511);
nor I_21169 (I362271,I362220,I243508);
nand I_21170 (I362288,I362271,I243529);
not I_21171 (I362305,I243508);
not I_21172 (I362322,I362305);
not I_21173 (I362339,I243505);
nor I_21174 (I362356,I362339,I243532);
and I_21175 (I362373,I362356,I243523);
or I_21176 (I362390,I362373,I243514);
DFFARX1 I_21177  ( .D(I362390), .CLK(I2350), .RSTB(I362203), .Q(I362407) );
nand I_21178 (I362424,I362220,I243505);
or I_21179 (I362192,I362424,I362407);
not I_21180 (I362455,I362424);
nor I_21181 (I362472,I362407,I362455);
and I_21182 (I362489,I362305,I362472);
nand I_21183 (I362165,I362424,I362322);
DFFARX1 I_21184  ( .D(I243517), .CLK(I2350), .RSTB(I362203), .Q(I362520) );
or I_21185 (I362186,I362520,I362407);
nor I_21186 (I362551,I362520,I362288);
nor I_21187 (I362568,I362520,I362322);
nand I_21188 (I362171,I362254,I362568);
or I_21189 (I362599,I362520,I362489);
DFFARX1 I_21190  ( .D(I362599), .CLK(I2350), .RSTB(I362203), .Q(I362168) );
not I_21191 (I362174,I362520);
DFFARX1 I_21192  ( .D(I243520), .CLK(I2350), .RSTB(I362203), .Q(I362644) );
not I_21193 (I362661,I362644);
nor I_21194 (I362678,I362661,I362254);
DFFARX1 I_21195  ( .D(I362678), .CLK(I2350), .RSTB(I362203), .Q(I362180) );
nor I_21196 (I362195,I362520,I362661);
nor I_21197 (I362183,I362661,I362424);
not I_21198 (I362737,I362661);
and I_21199 (I362754,I362288,I362737);
nor I_21200 (I362189,I362424,I362754);
nand I_21201 (I362177,I362661,I362551);
not I_21202 (I362832,I2357);
not I_21203 (I362849,I24242);
nor I_21204 (I362866,I24245,I24254);
nand I_21205 (I362883,I362866,I24269);
nor I_21206 (I362900,I362849,I24245);
nand I_21207 (I362917,I362900,I24248);
not I_21208 (I362934,I24245);
not I_21209 (I362951,I362934);
not I_21210 (I362968,I24239);
nor I_21211 (I362985,I362968,I24263);
and I_21212 (I363002,I362985,I24251);
or I_21213 (I363019,I363002,I24257);
DFFARX1 I_21214  ( .D(I363019), .CLK(I2350), .RSTB(I362832), .Q(I363036) );
nand I_21215 (I363053,I362849,I24239);
or I_21216 (I362821,I363053,I363036);
not I_21217 (I363084,I363053);
nor I_21218 (I363101,I363036,I363084);
and I_21219 (I363118,I362934,I363101);
nand I_21220 (I362794,I363053,I362951);
DFFARX1 I_21221  ( .D(I24260), .CLK(I2350), .RSTB(I362832), .Q(I363149) );
or I_21222 (I362815,I363149,I363036);
nor I_21223 (I363180,I363149,I362917);
nor I_21224 (I363197,I363149,I362951);
nand I_21225 (I362800,I362883,I363197);
or I_21226 (I363228,I363149,I363118);
DFFARX1 I_21227  ( .D(I363228), .CLK(I2350), .RSTB(I362832), .Q(I362797) );
not I_21228 (I362803,I363149);
DFFARX1 I_21229  ( .D(I24266), .CLK(I2350), .RSTB(I362832), .Q(I363273) );
not I_21230 (I363290,I363273);
nor I_21231 (I363307,I363290,I362883);
DFFARX1 I_21232  ( .D(I363307), .CLK(I2350), .RSTB(I362832), .Q(I362809) );
nor I_21233 (I362824,I363149,I363290);
nor I_21234 (I362812,I363290,I363053);
not I_21235 (I363366,I363290);
and I_21236 (I363383,I362917,I363366);
nor I_21237 (I362818,I363053,I363383);
nand I_21238 (I362806,I363290,I363180);
not I_21239 (I363461,I2357);
not I_21240 (I363478,I27866);
nor I_21241 (I363495,I27884,I27863);
nand I_21242 (I363512,I363495,I27881);
nor I_21243 (I363529,I363478,I27884);
nand I_21244 (I363546,I363529,I27875);
not I_21245 (I363563,I27884);
not I_21246 (I363580,I363563);
not I_21247 (I363597,I27878);
nor I_21248 (I363614,I363597,I27872);
and I_21249 (I363631,I363614,I27869);
or I_21250 (I363648,I363631,I27860);
DFFARX1 I_21251  ( .D(I363648), .CLK(I2350), .RSTB(I363461), .Q(I363665) );
nand I_21252 (I363682,I363478,I27878);
or I_21253 (I363450,I363682,I363665);
not I_21254 (I363713,I363682);
nor I_21255 (I363730,I363665,I363713);
and I_21256 (I363747,I363563,I363730);
nand I_21257 (I363423,I363682,I363580);
DFFARX1 I_21258  ( .D(I27890), .CLK(I2350), .RSTB(I363461), .Q(I363778) );
or I_21259 (I363444,I363778,I363665);
nor I_21260 (I363809,I363778,I363546);
nor I_21261 (I363826,I363778,I363580);
nand I_21262 (I363429,I363512,I363826);
or I_21263 (I363857,I363778,I363747);
DFFARX1 I_21264  ( .D(I363857), .CLK(I2350), .RSTB(I363461), .Q(I363426) );
not I_21265 (I363432,I363778);
DFFARX1 I_21266  ( .D(I27887), .CLK(I2350), .RSTB(I363461), .Q(I363902) );
not I_21267 (I363919,I363902);
nor I_21268 (I363936,I363919,I363512);
DFFARX1 I_21269  ( .D(I363936), .CLK(I2350), .RSTB(I363461), .Q(I363438) );
nor I_21270 (I363453,I363778,I363919);
nor I_21271 (I363441,I363919,I363682);
not I_21272 (I363995,I363919);
and I_21273 (I364012,I363546,I363995);
nor I_21274 (I363447,I363682,I364012);
nand I_21275 (I363435,I363919,I363809);
not I_21276 (I364090,I2357);
not I_21277 (I364107,I395491);
nor I_21278 (I364124,I395515,I395500);
nand I_21279 (I364141,I364124,I395485);
nor I_21280 (I364158,I364107,I395515);
nand I_21281 (I364175,I364158,I395512);
not I_21282 (I364192,I395515);
not I_21283 (I364209,I364192);
not I_21284 (I364226,I395494);
nor I_21285 (I364243,I364226,I395488);
and I_21286 (I364260,I364243,I395509);
or I_21287 (I364277,I364260,I395497);
DFFARX1 I_21288  ( .D(I364277), .CLK(I2350), .RSTB(I364090), .Q(I364294) );
nand I_21289 (I364311,I364107,I395494);
or I_21290 (I364079,I364311,I364294);
not I_21291 (I364342,I364311);
nor I_21292 (I364359,I364294,I364342);
and I_21293 (I364376,I364192,I364359);
nand I_21294 (I364052,I364311,I364209);
DFFARX1 I_21295  ( .D(I395506), .CLK(I2350), .RSTB(I364090), .Q(I364407) );
or I_21296 (I364073,I364407,I364294);
nor I_21297 (I364438,I364407,I364175);
nor I_21298 (I364455,I364407,I364209);
nand I_21299 (I364058,I364141,I364455);
or I_21300 (I364486,I364407,I364376);
DFFARX1 I_21301  ( .D(I364486), .CLK(I2350), .RSTB(I364090), .Q(I364055) );
not I_21302 (I364061,I364407);
DFFARX1 I_21303  ( .D(I395503), .CLK(I2350), .RSTB(I364090), .Q(I364531) );
not I_21304 (I364548,I364531);
nor I_21305 (I364565,I364548,I364141);
DFFARX1 I_21306  ( .D(I364565), .CLK(I2350), .RSTB(I364090), .Q(I364067) );
nor I_21307 (I364082,I364407,I364548);
nor I_21308 (I364070,I364548,I364311);
not I_21309 (I364624,I364548);
and I_21310 (I364641,I364175,I364624);
nor I_21311 (I364076,I364311,I364641);
nand I_21312 (I364064,I364548,I364438);
not I_21313 (I364719,I2357);
not I_21314 (I364736,I53706);
nor I_21315 (I364753,I53724,I53703);
nand I_21316 (I364770,I364753,I53721);
nor I_21317 (I364787,I364736,I53724);
nand I_21318 (I364804,I364787,I53715);
not I_21319 (I364821,I53724);
not I_21320 (I364838,I364821);
not I_21321 (I364855,I53718);
nor I_21322 (I364872,I364855,I53712);
and I_21323 (I364889,I364872,I53709);
or I_21324 (I364906,I364889,I53700);
DFFARX1 I_21325  ( .D(I364906), .CLK(I2350), .RSTB(I364719), .Q(I364923) );
nand I_21326 (I364940,I364736,I53718);
or I_21327 (I364708,I364940,I364923);
not I_21328 (I364971,I364940);
nor I_21329 (I364988,I364923,I364971);
and I_21330 (I365005,I364821,I364988);
nand I_21331 (I364681,I364940,I364838);
DFFARX1 I_21332  ( .D(I53730), .CLK(I2350), .RSTB(I364719), .Q(I365036) );
or I_21333 (I364702,I365036,I364923);
nor I_21334 (I365067,I365036,I364804);
nor I_21335 (I365084,I365036,I364838);
nand I_21336 (I364687,I364770,I365084);
or I_21337 (I365115,I365036,I365005);
DFFARX1 I_21338  ( .D(I365115), .CLK(I2350), .RSTB(I364719), .Q(I364684) );
not I_21339 (I364690,I365036);
DFFARX1 I_21340  ( .D(I53727), .CLK(I2350), .RSTB(I364719), .Q(I365160) );
not I_21341 (I365177,I365160);
nor I_21342 (I365194,I365177,I364770);
DFFARX1 I_21343  ( .D(I365194), .CLK(I2350), .RSTB(I364719), .Q(I364696) );
nor I_21344 (I364711,I365036,I365177);
nor I_21345 (I364699,I365177,I364940);
not I_21346 (I365253,I365177);
and I_21347 (I365270,I364804,I365253);
nor I_21348 (I364705,I364940,I365270);
nand I_21349 (I364693,I365177,I365067);
not I_21350 (I365348,I2357);
not I_21351 (I365365,I242379);
nor I_21352 (I365382,I242352,I242370);
nand I_21353 (I365399,I365382,I242355);
nor I_21354 (I365416,I365365,I242352);
nand I_21355 (I365433,I365416,I242373);
not I_21356 (I365450,I242352);
not I_21357 (I365467,I365450);
not I_21358 (I365484,I242349);
nor I_21359 (I365501,I365484,I242376);
and I_21360 (I365518,I365501,I242367);
or I_21361 (I365535,I365518,I242358);
DFFARX1 I_21362  ( .D(I365535), .CLK(I2350), .RSTB(I365348), .Q(I365552) );
nand I_21363 (I365569,I365365,I242349);
or I_21364 (I365337,I365569,I365552);
not I_21365 (I365600,I365569);
nor I_21366 (I365617,I365552,I365600);
and I_21367 (I365634,I365450,I365617);
nand I_21368 (I365310,I365569,I365467);
DFFARX1 I_21369  ( .D(I242361), .CLK(I2350), .RSTB(I365348), .Q(I365665) );
or I_21370 (I365331,I365665,I365552);
nor I_21371 (I365696,I365665,I365433);
nor I_21372 (I365713,I365665,I365467);
nand I_21373 (I365316,I365399,I365713);
or I_21374 (I365744,I365665,I365634);
DFFARX1 I_21375  ( .D(I365744), .CLK(I2350), .RSTB(I365348), .Q(I365313) );
not I_21376 (I365319,I365665);
DFFARX1 I_21377  ( .D(I242364), .CLK(I2350), .RSTB(I365348), .Q(I365789) );
not I_21378 (I365806,I365789);
nor I_21379 (I365823,I365806,I365399);
DFFARX1 I_21380  ( .D(I365823), .CLK(I2350), .RSTB(I365348), .Q(I365325) );
nor I_21381 (I365340,I365665,I365806);
nor I_21382 (I365328,I365806,I365569);
not I_21383 (I365882,I365806);
and I_21384 (I365899,I365433,I365882);
nor I_21385 (I365334,I365569,I365899);
nand I_21386 (I365322,I365806,I365696);
not I_21387 (I365977,I2357);
not I_21388 (I365994,I64042);
nor I_21389 (I366011,I64060,I64039);
nand I_21390 (I366028,I366011,I64057);
nor I_21391 (I366045,I365994,I64060);
nand I_21392 (I366062,I366045,I64051);
not I_21393 (I366079,I64060);
not I_21394 (I366096,I366079);
not I_21395 (I366113,I64054);
nor I_21396 (I366130,I366113,I64048);
and I_21397 (I366147,I366130,I64045);
or I_21398 (I366164,I366147,I64036);
DFFARX1 I_21399  ( .D(I366164), .CLK(I2350), .RSTB(I365977), .Q(I366181) );
nand I_21400 (I366198,I365994,I64054);
or I_21401 (I365966,I366198,I366181);
not I_21402 (I366229,I366198);
nor I_21403 (I366246,I366181,I366229);
and I_21404 (I366263,I366079,I366246);
nand I_21405 (I365939,I366198,I366096);
DFFARX1 I_21406  ( .D(I64066), .CLK(I2350), .RSTB(I365977), .Q(I366294) );
or I_21407 (I365960,I366294,I366181);
nor I_21408 (I366325,I366294,I366062);
nor I_21409 (I366342,I366294,I366096);
nand I_21410 (I365945,I366028,I366342);
or I_21411 (I366373,I366294,I366263);
DFFARX1 I_21412  ( .D(I366373), .CLK(I2350), .RSTB(I365977), .Q(I365942) );
not I_21413 (I365948,I366294);
DFFARX1 I_21414  ( .D(I64063), .CLK(I2350), .RSTB(I365977), .Q(I366418) );
not I_21415 (I366435,I366418);
nor I_21416 (I366452,I366435,I366028);
DFFARX1 I_21417  ( .D(I366452), .CLK(I2350), .RSTB(I365977), .Q(I365954) );
nor I_21418 (I365969,I366294,I366435);
nor I_21419 (I365957,I366435,I366198);
not I_21420 (I366511,I366435);
and I_21421 (I366528,I366062,I366511);
nor I_21422 (I365963,I366198,I366528);
nand I_21423 (I365951,I366435,I366325);
not I_21424 (I366606,I2357);
not I_21425 (I366623,I101295);
nor I_21426 (I366640,I101286,I101310);
nand I_21427 (I366657,I366640,I101313);
nor I_21428 (I366674,I366623,I101286);
nand I_21429 (I366691,I366674,I101304);
not I_21430 (I366708,I101286);
not I_21431 (I366725,I366708);
not I_21432 (I366742,I101298);
nor I_21433 (I366759,I366742,I101292);
and I_21434 (I366776,I366759,I101301);
or I_21435 (I366793,I366776,I101289);
DFFARX1 I_21436  ( .D(I366793), .CLK(I2350), .RSTB(I366606), .Q(I366810) );
nand I_21437 (I366827,I366623,I101298);
or I_21438 (I366595,I366827,I366810);
not I_21439 (I366858,I366827);
nor I_21440 (I366875,I366810,I366858);
and I_21441 (I366892,I366708,I366875);
nand I_21442 (I366568,I366827,I366725);
DFFARX1 I_21443  ( .D(I101283), .CLK(I2350), .RSTB(I366606), .Q(I366923) );
or I_21444 (I366589,I366923,I366810);
nor I_21445 (I366954,I366923,I366691);
nor I_21446 (I366971,I366923,I366725);
nand I_21447 (I366574,I366657,I366971);
or I_21448 (I367002,I366923,I366892);
DFFARX1 I_21449  ( .D(I367002), .CLK(I2350), .RSTB(I366606), .Q(I366571) );
not I_21450 (I366577,I366923);
DFFARX1 I_21451  ( .D(I101307), .CLK(I2350), .RSTB(I366606), .Q(I367047) );
not I_21452 (I367064,I367047);
nor I_21453 (I367081,I367064,I366657);
DFFARX1 I_21454  ( .D(I367081), .CLK(I2350), .RSTB(I366606), .Q(I366583) );
nor I_21455 (I366598,I366923,I367064);
nor I_21456 (I366586,I367064,I366827);
not I_21457 (I367140,I367064);
and I_21458 (I367157,I366691,I367140);
nor I_21459 (I366592,I366827,I367157);
nand I_21460 (I366580,I367064,I366954);
not I_21461 (I367235,I2357);
not I_21462 (I367252,I203709);
nor I_21463 (I367269,I203718,I203721);
nand I_21464 (I367286,I367269,I203706);
nor I_21465 (I367303,I367252,I203718);
nand I_21466 (I367320,I367303,I203703);
not I_21467 (I367337,I203718);
not I_21468 (I367354,I367337);
not I_21469 (I367371,I203691);
nor I_21470 (I367388,I367371,I203697);
and I_21471 (I367405,I367388,I203694);
or I_21472 (I367422,I367405,I203715);
DFFARX1 I_21473  ( .D(I367422), .CLK(I2350), .RSTB(I367235), .Q(I367439) );
nand I_21474 (I367456,I367252,I203691);
or I_21475 (I367224,I367456,I367439);
not I_21476 (I367487,I367456);
nor I_21477 (I367504,I367439,I367487);
and I_21478 (I367521,I367337,I367504);
nand I_21479 (I367197,I367456,I367354);
DFFARX1 I_21480  ( .D(I203700), .CLK(I2350), .RSTB(I367235), .Q(I367552) );
or I_21481 (I367218,I367552,I367439);
nor I_21482 (I367583,I367552,I367320);
nor I_21483 (I367600,I367552,I367354);
nand I_21484 (I367203,I367286,I367600);
or I_21485 (I367631,I367552,I367521);
DFFARX1 I_21486  ( .D(I367631), .CLK(I2350), .RSTB(I367235), .Q(I367200) );
not I_21487 (I367206,I367552);
DFFARX1 I_21488  ( .D(I203712), .CLK(I2350), .RSTB(I367235), .Q(I367676) );
not I_21489 (I367693,I367676);
nor I_21490 (I367710,I367693,I367286);
DFFARX1 I_21491  ( .D(I367710), .CLK(I2350), .RSTB(I367235), .Q(I367212) );
nor I_21492 (I367227,I367552,I367693);
nor I_21493 (I367215,I367693,I367456);
not I_21494 (I367769,I367693);
and I_21495 (I367786,I367320,I367769);
nor I_21496 (I367221,I367456,I367786);
nand I_21497 (I367209,I367693,I367583);
not I_21498 (I367864,I2357);
not I_21499 (I367881,I314761);
nor I_21500 (I367898,I314764,I314773);
nand I_21501 (I367915,I367898,I314758);
nor I_21502 (I367932,I367881,I314764);
nand I_21503 (I367949,I367932,I314767);
not I_21504 (I367966,I314764);
not I_21505 (I367983,I367966);
not I_21506 (I368000,I314782);
nor I_21507 (I368017,I368000,I314770);
and I_21508 (I368034,I368017,I314755);
or I_21509 (I368051,I368034,I314752);
DFFARX1 I_21510  ( .D(I368051), .CLK(I2350), .RSTB(I367864), .Q(I368068) );
nand I_21511 (I368085,I367881,I314782);
or I_21512 (I367853,I368085,I368068);
not I_21513 (I368116,I368085);
nor I_21514 (I368133,I368068,I368116);
and I_21515 (I368150,I367966,I368133);
nand I_21516 (I367826,I368085,I367983);
DFFARX1 I_21517  ( .D(I314776), .CLK(I2350), .RSTB(I367864), .Q(I368181) );
or I_21518 (I367847,I368181,I368068);
nor I_21519 (I368212,I368181,I367949);
nor I_21520 (I368229,I368181,I367983);
nand I_21521 (I367832,I367915,I368229);
or I_21522 (I368260,I368181,I368150);
DFFARX1 I_21523  ( .D(I368260), .CLK(I2350), .RSTB(I367864), .Q(I367829) );
not I_21524 (I367835,I368181);
DFFARX1 I_21525  ( .D(I314779), .CLK(I2350), .RSTB(I367864), .Q(I368305) );
not I_21526 (I368322,I368305);
nor I_21527 (I368339,I368322,I367915);
DFFARX1 I_21528  ( .D(I368339), .CLK(I2350), .RSTB(I367864), .Q(I367841) );
nor I_21529 (I367856,I368181,I368322);
nor I_21530 (I367844,I368322,I368085);
not I_21531 (I368398,I368322);
and I_21532 (I368415,I367949,I368398);
nor I_21533 (I367850,I368085,I368415);
nand I_21534 (I367838,I368322,I368212);
not I_21535 (I368493,I2357);
not I_21536 (I368510,I178141);
nor I_21537 (I368527,I178147,I178126);
nand I_21538 (I368544,I368527,I178132);
nor I_21539 (I368561,I368510,I178147);
nand I_21540 (I368578,I368561,I178138);
not I_21541 (I368595,I178147);
not I_21542 (I368612,I368595);
not I_21543 (I368629,I178135);
nor I_21544 (I368646,I368629,I178153);
and I_21545 (I368663,I368646,I178144);
or I_21546 (I368680,I368663,I178123);
DFFARX1 I_21547  ( .D(I368680), .CLK(I2350), .RSTB(I368493), .Q(I368697) );
nand I_21548 (I368714,I368510,I178135);
or I_21549 (I368482,I368714,I368697);
not I_21550 (I368745,I368714);
nor I_21551 (I368762,I368697,I368745);
and I_21552 (I368779,I368595,I368762);
nand I_21553 (I368455,I368714,I368612);
DFFARX1 I_21554  ( .D(I178150), .CLK(I2350), .RSTB(I368493), .Q(I368810) );
or I_21555 (I368476,I368810,I368697);
nor I_21556 (I368841,I368810,I368578);
nor I_21557 (I368858,I368810,I368612);
nand I_21558 (I368461,I368544,I368858);
or I_21559 (I368889,I368810,I368779);
DFFARX1 I_21560  ( .D(I368889), .CLK(I2350), .RSTB(I368493), .Q(I368458) );
not I_21561 (I368464,I368810);
DFFARX1 I_21562  ( .D(I178129), .CLK(I2350), .RSTB(I368493), .Q(I368934) );
not I_21563 (I368951,I368934);
nor I_21564 (I368968,I368951,I368544);
DFFARX1 I_21565  ( .D(I368968), .CLK(I2350), .RSTB(I368493), .Q(I368470) );
nor I_21566 (I368485,I368810,I368951);
nor I_21567 (I368473,I368951,I368714);
not I_21568 (I369027,I368951);
and I_21569 (I369044,I368578,I369027);
nor I_21570 (I368479,I368714,I369044);
nand I_21571 (I368467,I368951,I368841);
not I_21572 (I369122,I2357);
not I_21573 (I369139,I282033);
nor I_21574 (I369156,I282051,I282030);
nand I_21575 (I369173,I369156,I282054);
nor I_21576 (I369190,I369139,I282051);
nand I_21577 (I369207,I369190,I282048);
not I_21578 (I369224,I282051);
not I_21579 (I369241,I369224);
not I_21580 (I369258,I282039);
nor I_21581 (I369275,I369258,I282027);
and I_21582 (I369292,I369275,I282045);
or I_21583 (I369309,I369292,I282057);
DFFARX1 I_21584  ( .D(I369309), .CLK(I2350), .RSTB(I369122), .Q(I369326) );
nand I_21585 (I369343,I369139,I282039);
or I_21586 (I369111,I369343,I369326);
not I_21587 (I369374,I369343);
nor I_21588 (I369391,I369326,I369374);
and I_21589 (I369408,I369224,I369391);
nand I_21590 (I369084,I369343,I369241);
DFFARX1 I_21591  ( .D(I282036), .CLK(I2350), .RSTB(I369122), .Q(I369439) );
or I_21592 (I369105,I369439,I369326);
nor I_21593 (I369470,I369439,I369207);
nor I_21594 (I369487,I369439,I369241);
nand I_21595 (I369090,I369173,I369487);
or I_21596 (I369518,I369439,I369408);
DFFARX1 I_21597  ( .D(I369518), .CLK(I2350), .RSTB(I369122), .Q(I369087) );
not I_21598 (I369093,I369439);
DFFARX1 I_21599  ( .D(I282042), .CLK(I2350), .RSTB(I369122), .Q(I369563) );
not I_21600 (I369580,I369563);
nor I_21601 (I369597,I369580,I369173);
DFFARX1 I_21602  ( .D(I369597), .CLK(I2350), .RSTB(I369122), .Q(I369099) );
nor I_21603 (I369114,I369439,I369580);
nor I_21604 (I369102,I369580,I369343);
not I_21605 (I369656,I369580);
and I_21606 (I369673,I369207,I369656);
nor I_21607 (I369108,I369343,I369673);
nand I_21608 (I369096,I369580,I369470);
not I_21609 (I369751,I2357);
not I_21610 (I369768,I26574);
nor I_21611 (I369785,I26592,I26571);
nand I_21612 (I369802,I369785,I26589);
nor I_21613 (I369819,I369768,I26592);
nand I_21614 (I369836,I369819,I26583);
not I_21615 (I369853,I26592);
not I_21616 (I369870,I369853);
not I_21617 (I369887,I26586);
nor I_21618 (I369904,I369887,I26580);
and I_21619 (I369921,I369904,I26577);
or I_21620 (I369938,I369921,I26568);
DFFARX1 I_21621  ( .D(I369938), .CLK(I2350), .RSTB(I369751), .Q(I369955) );
nand I_21622 (I369972,I369768,I26586);
or I_21623 (I369740,I369972,I369955);
not I_21624 (I370003,I369972);
nor I_21625 (I370020,I369955,I370003);
and I_21626 (I370037,I369853,I370020);
nand I_21627 (I369713,I369972,I369870);
DFFARX1 I_21628  ( .D(I26598), .CLK(I2350), .RSTB(I369751), .Q(I370068) );
or I_21629 (I369734,I370068,I369955);
nor I_21630 (I370099,I370068,I369836);
nor I_21631 (I370116,I370068,I369870);
nand I_21632 (I369719,I369802,I370116);
or I_21633 (I370147,I370068,I370037);
DFFARX1 I_21634  ( .D(I370147), .CLK(I2350), .RSTB(I369751), .Q(I369716) );
not I_21635 (I369722,I370068);
DFFARX1 I_21636  ( .D(I26595), .CLK(I2350), .RSTB(I369751), .Q(I370192) );
not I_21637 (I370209,I370192);
nor I_21638 (I370226,I370209,I369802);
DFFARX1 I_21639  ( .D(I370226), .CLK(I2350), .RSTB(I369751), .Q(I369728) );
nor I_21640 (I369743,I370068,I370209);
nor I_21641 (I369731,I370209,I369972);
not I_21642 (I370285,I370209);
and I_21643 (I370302,I369836,I370285);
nor I_21644 (I369737,I369972,I370302);
nand I_21645 (I369725,I370209,I370099);
not I_21646 (I370380,I2357);
not I_21647 (I370397,I281438);
nor I_21648 (I370414,I281456,I281435);
nand I_21649 (I370431,I370414,I281459);
nor I_21650 (I370448,I370397,I281456);
nand I_21651 (I370465,I370448,I281453);
not I_21652 (I370482,I281456);
not I_21653 (I370499,I370482);
not I_21654 (I370516,I281444);
nor I_21655 (I370533,I370516,I281432);
and I_21656 (I370550,I370533,I281450);
or I_21657 (I370567,I370550,I281462);
DFFARX1 I_21658  ( .D(I370567), .CLK(I2350), .RSTB(I370380), .Q(I370584) );
nand I_21659 (I370601,I370397,I281444);
or I_21660 (I370369,I370601,I370584);
not I_21661 (I370632,I370601);
nor I_21662 (I370649,I370584,I370632);
and I_21663 (I370666,I370482,I370649);
nand I_21664 (I370342,I370601,I370499);
DFFARX1 I_21665  ( .D(I281441), .CLK(I2350), .RSTB(I370380), .Q(I370697) );
or I_21666 (I370363,I370697,I370584);
nor I_21667 (I370728,I370697,I370465);
nor I_21668 (I370745,I370697,I370499);
nand I_21669 (I370348,I370431,I370745);
or I_21670 (I370776,I370697,I370666);
DFFARX1 I_21671  ( .D(I370776), .CLK(I2350), .RSTB(I370380), .Q(I370345) );
not I_21672 (I370351,I370697);
DFFARX1 I_21673  ( .D(I281447), .CLK(I2350), .RSTB(I370380), .Q(I370821) );
not I_21674 (I370838,I370821);
nor I_21675 (I370855,I370838,I370431);
DFFARX1 I_21676  ( .D(I370855), .CLK(I2350), .RSTB(I370380), .Q(I370357) );
nor I_21677 (I370372,I370697,I370838);
nor I_21678 (I370360,I370838,I370601);
not I_21679 (I370914,I370838);
and I_21680 (I370931,I370465,I370914);
nor I_21681 (I370366,I370601,I370931);
nand I_21682 (I370354,I370838,I370728);
not I_21683 (I371009,I2357);
not I_21684 (I371026,I285008);
nor I_21685 (I371043,I285026,I285005);
nand I_21686 (I371060,I371043,I285029);
nor I_21687 (I371077,I371026,I285026);
nand I_21688 (I371094,I371077,I285023);
not I_21689 (I371111,I285026);
not I_21690 (I371128,I371111);
not I_21691 (I371145,I285014);
nor I_21692 (I371162,I371145,I285002);
and I_21693 (I371179,I371162,I285020);
or I_21694 (I371196,I371179,I285032);
DFFARX1 I_21695  ( .D(I371196), .CLK(I2350), .RSTB(I371009), .Q(I371213) );
nand I_21696 (I371230,I371026,I285014);
or I_21697 (I370998,I371230,I371213);
not I_21698 (I371261,I371230);
nor I_21699 (I371278,I371213,I371261);
and I_21700 (I371295,I371111,I371278);
nand I_21701 (I370971,I371230,I371128);
DFFARX1 I_21702  ( .D(I285011), .CLK(I2350), .RSTB(I371009), .Q(I371326) );
or I_21703 (I370992,I371326,I371213);
nor I_21704 (I371357,I371326,I371094);
nor I_21705 (I371374,I371326,I371128);
nand I_21706 (I370977,I371060,I371374);
or I_21707 (I371405,I371326,I371295);
DFFARX1 I_21708  ( .D(I371405), .CLK(I2350), .RSTB(I371009), .Q(I370974) );
not I_21709 (I370980,I371326);
DFFARX1 I_21710  ( .D(I285017), .CLK(I2350), .RSTB(I371009), .Q(I371450) );
not I_21711 (I371467,I371450);
nor I_21712 (I371484,I371467,I371060);
DFFARX1 I_21713  ( .D(I371484), .CLK(I2350), .RSTB(I371009), .Q(I370986) );
nor I_21714 (I371001,I371326,I371467);
nor I_21715 (I370989,I371467,I371230);
not I_21716 (I371543,I371467);
and I_21717 (I371560,I371094,I371543);
nor I_21718 (I370995,I371230,I371560);
nand I_21719 (I370983,I371467,I371357);
not I_21720 (I371638,I2357);
not I_21721 (I371655,I298098);
nor I_21722 (I371672,I298116,I298095);
nand I_21723 (I371689,I371672,I298119);
nor I_21724 (I371706,I371655,I298116);
nand I_21725 (I371723,I371706,I298113);
not I_21726 (I371740,I298116);
not I_21727 (I371757,I371740);
not I_21728 (I371774,I298104);
nor I_21729 (I371791,I371774,I298092);
and I_21730 (I371808,I371791,I298110);
or I_21731 (I371825,I371808,I298122);
DFFARX1 I_21732  ( .D(I371825), .CLK(I2350), .RSTB(I371638), .Q(I371842) );
nand I_21733 (I371859,I371655,I298104);
or I_21734 (I371627,I371859,I371842);
not I_21735 (I371890,I371859);
nor I_21736 (I371907,I371842,I371890);
and I_21737 (I371924,I371740,I371907);
nand I_21738 (I371600,I371859,I371757);
DFFARX1 I_21739  ( .D(I298101), .CLK(I2350), .RSTB(I371638), .Q(I371955) );
or I_21740 (I371621,I371955,I371842);
nor I_21741 (I371986,I371955,I371723);
nor I_21742 (I372003,I371955,I371757);
nand I_21743 (I371606,I371689,I372003);
or I_21744 (I372034,I371955,I371924);
DFFARX1 I_21745  ( .D(I372034), .CLK(I2350), .RSTB(I371638), .Q(I371603) );
not I_21746 (I371609,I371955);
DFFARX1 I_21747  ( .D(I298107), .CLK(I2350), .RSTB(I371638), .Q(I372079) );
not I_21748 (I372096,I372079);
nor I_21749 (I372113,I372096,I371689);
DFFARX1 I_21750  ( .D(I372113), .CLK(I2350), .RSTB(I371638), .Q(I371615) );
nor I_21751 (I371630,I371955,I372096);
nor I_21752 (I371618,I372096,I371859);
not I_21753 (I372172,I372096);
and I_21754 (I372189,I371723,I372172);
nor I_21755 (I371624,I371859,I372189);
nand I_21756 (I371612,I372096,I371986);
not I_21757 (I372267,I2357);
not I_21758 (I372284,I70502);
nor I_21759 (I372301,I70520,I70499);
nand I_21760 (I372318,I372301,I70517);
nor I_21761 (I372335,I372284,I70520);
nand I_21762 (I372352,I372335,I70511);
not I_21763 (I372369,I70520);
not I_21764 (I372386,I372369);
not I_21765 (I372403,I70514);
nor I_21766 (I372420,I372403,I70508);
and I_21767 (I372437,I372420,I70505);
or I_21768 (I372454,I372437,I70496);
DFFARX1 I_21769  ( .D(I372454), .CLK(I2350), .RSTB(I372267), .Q(I372471) );
nand I_21770 (I372488,I372284,I70514);
or I_21771 (I372256,I372488,I372471);
not I_21772 (I372519,I372488);
nor I_21773 (I372536,I372471,I372519);
and I_21774 (I372553,I372369,I372536);
nand I_21775 (I372229,I372488,I372386);
DFFARX1 I_21776  ( .D(I70526), .CLK(I2350), .RSTB(I372267), .Q(I372584) );
or I_21777 (I372250,I372584,I372471);
nor I_21778 (I372615,I372584,I372352);
nor I_21779 (I372632,I372584,I372386);
nand I_21780 (I372235,I372318,I372632);
or I_21781 (I372663,I372584,I372553);
DFFARX1 I_21782  ( .D(I372663), .CLK(I2350), .RSTB(I372267), .Q(I372232) );
not I_21783 (I372238,I372584);
DFFARX1 I_21784  ( .D(I70523), .CLK(I2350), .RSTB(I372267), .Q(I372708) );
not I_21785 (I372725,I372708);
nor I_21786 (I372742,I372725,I372318);
DFFARX1 I_21787  ( .D(I372742), .CLK(I2350), .RSTB(I372267), .Q(I372244) );
nor I_21788 (I372259,I372584,I372725);
nor I_21789 (I372247,I372725,I372488);
not I_21790 (I372801,I372725);
and I_21791 (I372818,I372352,I372801);
nor I_21792 (I372253,I372488,I372818);
nand I_21793 (I372241,I372725,I372615);
not I_21794 (I372896,I2357);
not I_21795 (I372913,I90024);
nor I_21796 (I372930,I90015,I90039);
nand I_21797 (I372947,I372930,I90042);
nor I_21798 (I372964,I372913,I90015);
nand I_21799 (I372981,I372964,I90033);
not I_21800 (I372998,I90015);
not I_21801 (I373015,I372998);
not I_21802 (I373032,I90027);
nor I_21803 (I373049,I373032,I90021);
and I_21804 (I373066,I373049,I90030);
or I_21805 (I373083,I373066,I90018);
DFFARX1 I_21806  ( .D(I373083), .CLK(I2350), .RSTB(I372896), .Q(I373100) );
nand I_21807 (I373117,I372913,I90027);
or I_21808 (I372885,I373117,I373100);
not I_21809 (I373148,I373117);
nor I_21810 (I373165,I373100,I373148);
and I_21811 (I373182,I372998,I373165);
nand I_21812 (I372858,I373117,I373015);
DFFARX1 I_21813  ( .D(I90012), .CLK(I2350), .RSTB(I372896), .Q(I373213) );
or I_21814 (I372879,I373213,I373100);
nor I_21815 (I373244,I373213,I372981);
nor I_21816 (I373261,I373213,I373015);
nand I_21817 (I372864,I372947,I373261);
or I_21818 (I373292,I373213,I373182);
DFFARX1 I_21819  ( .D(I373292), .CLK(I2350), .RSTB(I372896), .Q(I372861) );
not I_21820 (I372867,I373213);
DFFARX1 I_21821  ( .D(I90036), .CLK(I2350), .RSTB(I372896), .Q(I373337) );
not I_21822 (I373354,I373337);
nor I_21823 (I373371,I373354,I372947);
DFFARX1 I_21824  ( .D(I373371), .CLK(I2350), .RSTB(I372896), .Q(I372873) );
nor I_21825 (I372888,I373213,I373354);
nor I_21826 (I372876,I373354,I373117);
not I_21827 (I373430,I373354);
and I_21828 (I373447,I372981,I373430);
nor I_21829 (I372882,I373117,I373447);
nand I_21830 (I372870,I373354,I373244);
not I_21831 (I373525,I2357);
not I_21832 (I373542,I218567);
nor I_21833 (I373559,I218576,I218579);
nand I_21834 (I373576,I373559,I218564);
nor I_21835 (I373593,I373542,I218576);
nand I_21836 (I373610,I373593,I218561);
not I_21837 (I373627,I218576);
not I_21838 (I373644,I373627);
not I_21839 (I373661,I218549);
nor I_21840 (I373678,I373661,I218555);
and I_21841 (I373695,I373678,I218552);
or I_21842 (I373712,I373695,I218573);
DFFARX1 I_21843  ( .D(I373712), .CLK(I2350), .RSTB(I373525), .Q(I373729) );
nand I_21844 (I373746,I373542,I218549);
or I_21845 (I373514,I373746,I373729);
not I_21846 (I373777,I373746);
nor I_21847 (I373794,I373729,I373777);
and I_21848 (I373811,I373627,I373794);
nand I_21849 (I373487,I373746,I373644);
DFFARX1 I_21850  ( .D(I218558), .CLK(I2350), .RSTB(I373525), .Q(I373842) );
or I_21851 (I373508,I373842,I373729);
nor I_21852 (I373873,I373842,I373610);
nor I_21853 (I373890,I373842,I373644);
nand I_21854 (I373493,I373576,I373890);
or I_21855 (I373921,I373842,I373811);
DFFARX1 I_21856  ( .D(I373921), .CLK(I2350), .RSTB(I373525), .Q(I373490) );
not I_21857 (I373496,I373842);
DFFARX1 I_21858  ( .D(I218570), .CLK(I2350), .RSTB(I373525), .Q(I373966) );
not I_21859 (I373983,I373966);
nor I_21860 (I374000,I373983,I373576);
DFFARX1 I_21861  ( .D(I374000), .CLK(I2350), .RSTB(I373525), .Q(I373502) );
nor I_21862 (I373517,I373842,I373983);
nor I_21863 (I373505,I373983,I373746);
not I_21864 (I374059,I373983);
and I_21865 (I374076,I373610,I374059);
nor I_21866 (I373511,I373746,I374076);
nand I_21867 (I373499,I373983,I373873);
not I_21868 (I374154,I2357);
not I_21869 (I374171,I198541);
nor I_21870 (I374188,I198550,I198553);
nand I_21871 (I374205,I374188,I198538);
nor I_21872 (I374222,I374171,I198550);
nand I_21873 (I374239,I374222,I198535);
not I_21874 (I374256,I198550);
not I_21875 (I374273,I374256);
not I_21876 (I374290,I198523);
nor I_21877 (I374307,I374290,I198529);
and I_21878 (I374324,I374307,I198526);
or I_21879 (I374341,I374324,I198547);
DFFARX1 I_21880  ( .D(I374341), .CLK(I2350), .RSTB(I374154), .Q(I374358) );
nand I_21881 (I374375,I374171,I198523);
or I_21882 (I374143,I374375,I374358);
not I_21883 (I374406,I374375);
nor I_21884 (I374423,I374358,I374406);
and I_21885 (I374440,I374256,I374423);
nand I_21886 (I374116,I374375,I374273);
DFFARX1 I_21887  ( .D(I198532), .CLK(I2350), .RSTB(I374154), .Q(I374471) );
or I_21888 (I374137,I374471,I374358);
nor I_21889 (I374502,I374471,I374239);
nor I_21890 (I374519,I374471,I374273);
nand I_21891 (I374122,I374205,I374519);
or I_21892 (I374550,I374471,I374440);
DFFARX1 I_21893  ( .D(I374550), .CLK(I2350), .RSTB(I374154), .Q(I374119) );
not I_21894 (I374125,I374471);
DFFARX1 I_21895  ( .D(I198544), .CLK(I2350), .RSTB(I374154), .Q(I374595) );
not I_21896 (I374612,I374595);
nor I_21897 (I374629,I374612,I374205);
DFFARX1 I_21898  ( .D(I374629), .CLK(I2350), .RSTB(I374154), .Q(I374131) );
nor I_21899 (I374146,I374471,I374612);
nor I_21900 (I374134,I374612,I374375);
not I_21901 (I374688,I374612);
and I_21902 (I374705,I374239,I374688);
nor I_21903 (I374140,I374375,I374705);
nand I_21904 (I374128,I374612,I374502);
not I_21905 (I374783,I2357);
not I_21906 (I374800,I17510);
nor I_21907 (I374817,I17513,I17522);
nand I_21908 (I374834,I374817,I17537);
nor I_21909 (I374851,I374800,I17513);
nand I_21910 (I374868,I374851,I17516);
not I_21911 (I374885,I17513);
not I_21912 (I374902,I374885);
not I_21913 (I374919,I17507);
nor I_21914 (I374936,I374919,I17531);
and I_21915 (I374953,I374936,I17519);
or I_21916 (I374970,I374953,I17525);
DFFARX1 I_21917  ( .D(I374970), .CLK(I2350), .RSTB(I374783), .Q(I374987) );
nand I_21918 (I375004,I374800,I17507);
or I_21919 (I374772,I375004,I374987);
not I_21920 (I375035,I375004);
nor I_21921 (I375052,I374987,I375035);
and I_21922 (I375069,I374885,I375052);
nand I_21923 (I374745,I375004,I374902);
DFFARX1 I_21924  ( .D(I17528), .CLK(I2350), .RSTB(I374783), .Q(I375100) );
or I_21925 (I374766,I375100,I374987);
nor I_21926 (I375131,I375100,I374868);
nor I_21927 (I375148,I375100,I374902);
nand I_21928 (I374751,I374834,I375148);
or I_21929 (I375179,I375100,I375069);
DFFARX1 I_21930  ( .D(I375179), .CLK(I2350), .RSTB(I374783), .Q(I374748) );
not I_21931 (I374754,I375100);
DFFARX1 I_21932  ( .D(I17534), .CLK(I2350), .RSTB(I374783), .Q(I375224) );
not I_21933 (I375241,I375224);
nor I_21934 (I375258,I375241,I374834);
DFFARX1 I_21935  ( .D(I375258), .CLK(I2350), .RSTB(I374783), .Q(I374760) );
nor I_21936 (I374775,I375100,I375241);
nor I_21937 (I374763,I375241,I375004);
not I_21938 (I375317,I375241);
and I_21939 (I375334,I374868,I375317);
nor I_21940 (I374769,I375004,I375334);
nand I_21941 (I374757,I375241,I375131);
not I_21942 (I375412,I2357);
not I_21943 (I375429,I2363);
nor I_21944 (I375446,I2366,I2375);
nand I_21945 (I375463,I375446,I2390);
nor I_21946 (I375480,I375429,I2366);
nand I_21947 (I375497,I375480,I2369);
not I_21948 (I375514,I2366);
not I_21949 (I375531,I375514);
not I_21950 (I375548,I2360);
nor I_21951 (I375565,I375548,I2384);
and I_21952 (I375582,I375565,I2372);
or I_21953 (I375599,I375582,I2378);
DFFARX1 I_21954  ( .D(I375599), .CLK(I2350), .RSTB(I375412), .Q(I375616) );
nand I_21955 (I375633,I375429,I2360);
or I_21956 (I375401,I375633,I375616);
not I_21957 (I375664,I375633);
nor I_21958 (I375681,I375616,I375664);
and I_21959 (I375698,I375514,I375681);
nand I_21960 (I375374,I375633,I375531);
DFFARX1 I_21961  ( .D(I2381), .CLK(I2350), .RSTB(I375412), .Q(I375729) );
or I_21962 (I375395,I375729,I375616);
nor I_21963 (I375760,I375729,I375497);
nor I_21964 (I375777,I375729,I375531);
nand I_21965 (I375380,I375463,I375777);
or I_21966 (I375808,I375729,I375698);
DFFARX1 I_21967  ( .D(I375808), .CLK(I2350), .RSTB(I375412), .Q(I375377) );
not I_21968 (I375383,I375729);
DFFARX1 I_21969  ( .D(I2387), .CLK(I2350), .RSTB(I375412), .Q(I375853) );
not I_21970 (I375870,I375853);
nor I_21971 (I375887,I375870,I375463);
DFFARX1 I_21972  ( .D(I375887), .CLK(I2350), .RSTB(I375412), .Q(I375389) );
nor I_21973 (I375404,I375729,I375870);
nor I_21974 (I375392,I375870,I375633);
not I_21975 (I375946,I375870);
and I_21976 (I375963,I375497,I375946);
nor I_21977 (I375398,I375633,I375963);
nand I_21978 (I375386,I375870,I375760);
not I_21979 (I376041,I2357);
not I_21980 (I376058,I140350);
nor I_21981 (I376075,I140356,I140335);
nand I_21982 (I376092,I376075,I140341);
nor I_21983 (I376109,I376058,I140356);
nand I_21984 (I376126,I376109,I140347);
not I_21985 (I376143,I140356);
not I_21986 (I376160,I376143);
not I_21987 (I376177,I140344);
nor I_21988 (I376194,I376177,I140362);
and I_21989 (I376211,I376194,I140353);
or I_21990 (I376228,I376211,I140332);
DFFARX1 I_21991  ( .D(I376228), .CLK(I2350), .RSTB(I376041), .Q(I376245) );
nand I_21992 (I376262,I376058,I140344);
or I_21993 (I376030,I376262,I376245);
not I_21994 (I376293,I376262);
nor I_21995 (I376310,I376245,I376293);
and I_21996 (I376327,I376143,I376310);
nand I_21997 (I376003,I376262,I376160);
DFFARX1 I_21998  ( .D(I140359), .CLK(I2350), .RSTB(I376041), .Q(I376358) );
or I_21999 (I376024,I376358,I376245);
nor I_22000 (I376389,I376358,I376126);
nor I_22001 (I376406,I376358,I376160);
nand I_22002 (I376009,I376092,I376406);
or I_22003 (I376437,I376358,I376327);
DFFARX1 I_22004  ( .D(I376437), .CLK(I2350), .RSTB(I376041), .Q(I376006) );
not I_22005 (I376012,I376358);
DFFARX1 I_22006  ( .D(I140338), .CLK(I2350), .RSTB(I376041), .Q(I376482) );
not I_22007 (I376499,I376482);
nor I_22008 (I376516,I376499,I376092);
DFFARX1 I_22009  ( .D(I376516), .CLK(I2350), .RSTB(I376041), .Q(I376018) );
nor I_22010 (I376033,I376358,I376499);
nor I_22011 (I376021,I376499,I376262);
not I_22012 (I376575,I376499);
and I_22013 (I376592,I376126,I376575);
nor I_22014 (I376027,I376262,I376592);
nand I_22015 (I376015,I376499,I376389);
not I_22016 (I376670,I2357);
not I_22017 (I376687,I5729);
nor I_22018 (I376704,I5732,I5741);
nand I_22019 (I376721,I376704,I5756);
nor I_22020 (I376738,I376687,I5732);
nand I_22021 (I376755,I376738,I5735);
not I_22022 (I376772,I5732);
not I_22023 (I376789,I376772);
not I_22024 (I376806,I5726);
nor I_22025 (I376823,I376806,I5750);
and I_22026 (I376840,I376823,I5738);
or I_22027 (I376857,I376840,I5744);
DFFARX1 I_22028  ( .D(I376857), .CLK(I2350), .RSTB(I376670), .Q(I376874) );
nand I_22029 (I376891,I376687,I5726);
or I_22030 (I376659,I376891,I376874);
not I_22031 (I376922,I376891);
nor I_22032 (I376939,I376874,I376922);
and I_22033 (I376956,I376772,I376939);
nand I_22034 (I376632,I376891,I376789);
DFFARX1 I_22035  ( .D(I5747), .CLK(I2350), .RSTB(I376670), .Q(I376987) );
or I_22036 (I376653,I376987,I376874);
nor I_22037 (I377018,I376987,I376755);
nor I_22038 (I377035,I376987,I376789);
nand I_22039 (I376638,I376721,I377035);
or I_22040 (I377066,I376987,I376956);
DFFARX1 I_22041  ( .D(I377066), .CLK(I2350), .RSTB(I376670), .Q(I376635) );
not I_22042 (I376641,I376987);
DFFARX1 I_22043  ( .D(I5753), .CLK(I2350), .RSTB(I376670), .Q(I377111) );
not I_22044 (I377128,I377111);
nor I_22045 (I377145,I377128,I376721);
DFFARX1 I_22046  ( .D(I377145), .CLK(I2350), .RSTB(I376670), .Q(I376647) );
nor I_22047 (I376662,I376987,I377128);
nor I_22048 (I376650,I377128,I376891);
not I_22049 (I377204,I377128);
and I_22050 (I377221,I376755,I377204);
nor I_22051 (I376656,I376891,I377221);
nand I_22052 (I376644,I377128,I377018);
not I_22053 (I377299,I2357);
not I_22054 (I377316,I107925);
nor I_22055 (I377333,I107916,I107940);
nand I_22056 (I377350,I377333,I107943);
nor I_22057 (I377367,I377316,I107916);
nand I_22058 (I377384,I377367,I107934);
not I_22059 (I377401,I107916);
not I_22060 (I377418,I377401);
not I_22061 (I377435,I107928);
nor I_22062 (I377452,I377435,I107922);
and I_22063 (I377469,I377452,I107931);
or I_22064 (I377486,I377469,I107919);
DFFARX1 I_22065  ( .D(I377486), .CLK(I2350), .RSTB(I377299), .Q(I377503) );
nand I_22066 (I377520,I377316,I107928);
or I_22067 (I377288,I377520,I377503);
not I_22068 (I377551,I377520);
nor I_22069 (I377568,I377503,I377551);
and I_22070 (I377585,I377401,I377568);
nand I_22071 (I377261,I377520,I377418);
DFFARX1 I_22072  ( .D(I107913), .CLK(I2350), .RSTB(I377299), .Q(I377616) );
or I_22073 (I377282,I377616,I377503);
nor I_22074 (I377647,I377616,I377384);
nor I_22075 (I377664,I377616,I377418);
nand I_22076 (I377267,I377350,I377664);
or I_22077 (I377695,I377616,I377585);
DFFARX1 I_22078  ( .D(I377695), .CLK(I2350), .RSTB(I377299), .Q(I377264) );
not I_22079 (I377270,I377616);
DFFARX1 I_22080  ( .D(I107937), .CLK(I2350), .RSTB(I377299), .Q(I377740) );
not I_22081 (I377757,I377740);
nor I_22082 (I377774,I377757,I377350);
DFFARX1 I_22083  ( .D(I377774), .CLK(I2350), .RSTB(I377299), .Q(I377276) );
nor I_22084 (I377291,I377616,I377757);
nor I_22085 (I377279,I377757,I377520);
not I_22086 (I377833,I377757);
and I_22087 (I377850,I377384,I377833);
nor I_22088 (I377285,I377520,I377850);
nand I_22089 (I377273,I377757,I377647);
not I_22090 (I377928,I2357);
not I_22091 (I377945,I299883);
nor I_22092 (I377962,I299901,I299880);
nand I_22093 (I377979,I377962,I299904);
nor I_22094 (I377996,I377945,I299901);
nand I_22095 (I378013,I377996,I299898);
not I_22096 (I378030,I299901);
not I_22097 (I378047,I378030);
not I_22098 (I378064,I299889);
nor I_22099 (I378081,I378064,I299877);
and I_22100 (I378098,I378081,I299895);
or I_22101 (I378115,I378098,I299907);
DFFARX1 I_22102  ( .D(I378115), .CLK(I2350), .RSTB(I377928), .Q(I378132) );
nand I_22103 (I378149,I377945,I299889);
or I_22104 (I377917,I378149,I378132);
not I_22105 (I378180,I378149);
nor I_22106 (I378197,I378132,I378180);
and I_22107 (I378214,I378030,I378197);
nand I_22108 (I377890,I378149,I378047);
DFFARX1 I_22109  ( .D(I299886), .CLK(I2350), .RSTB(I377928), .Q(I378245) );
or I_22110 (I377911,I378245,I378132);
nor I_22111 (I378276,I378245,I378013);
nor I_22112 (I378293,I378245,I378047);
nand I_22113 (I377896,I377979,I378293);
or I_22114 (I378324,I378245,I378214);
DFFARX1 I_22115  ( .D(I378324), .CLK(I2350), .RSTB(I377928), .Q(I377893) );
not I_22116 (I377899,I378245);
DFFARX1 I_22117  ( .D(I299892), .CLK(I2350), .RSTB(I377928), .Q(I378369) );
not I_22118 (I378386,I378369);
nor I_22119 (I378403,I378386,I377979);
DFFARX1 I_22120  ( .D(I378403), .CLK(I2350), .RSTB(I377928), .Q(I377905) );
nor I_22121 (I377920,I378245,I378386);
nor I_22122 (I377908,I378386,I378149);
not I_22123 (I378462,I378386);
and I_22124 (I378479,I378013,I378462);
nor I_22125 (I377914,I378149,I378479);
nand I_22126 (I377902,I378386,I378276);
not I_22127 (I378557,I2357);
not I_22128 (I378574,I232133);
nor I_22129 (I378591,I232142,I232145);
nand I_22130 (I378608,I378591,I232130);
nor I_22131 (I378625,I378574,I232142);
nand I_22132 (I378642,I378625,I232127);
not I_22133 (I378659,I232142);
not I_22134 (I378676,I378659);
not I_22135 (I378693,I232115);
nor I_22136 (I378710,I378693,I232121);
and I_22137 (I378727,I378710,I232118);
or I_22138 (I378744,I378727,I232139);
DFFARX1 I_22139  ( .D(I378744), .CLK(I2350), .RSTB(I378557), .Q(I378761) );
nand I_22140 (I378778,I378574,I232115);
or I_22141 (I378546,I378778,I378761);
not I_22142 (I378809,I378778);
nor I_22143 (I378826,I378761,I378809);
and I_22144 (I378843,I378659,I378826);
nand I_22145 (I378519,I378778,I378676);
DFFARX1 I_22146  ( .D(I232124), .CLK(I2350), .RSTB(I378557), .Q(I378874) );
or I_22147 (I378540,I378874,I378761);
nor I_22148 (I378905,I378874,I378642);
nor I_22149 (I378922,I378874,I378676);
nand I_22150 (I378525,I378608,I378922);
or I_22151 (I378953,I378874,I378843);
DFFARX1 I_22152  ( .D(I378953), .CLK(I2350), .RSTB(I378557), .Q(I378522) );
not I_22153 (I378528,I378874);
DFFARX1 I_22154  ( .D(I232136), .CLK(I2350), .RSTB(I378557), .Q(I378998) );
not I_22155 (I379015,I378998);
nor I_22156 (I379032,I379015,I378608);
DFFARX1 I_22157  ( .D(I379032), .CLK(I2350), .RSTB(I378557), .Q(I378534) );
nor I_22158 (I378549,I378874,I379015);
nor I_22159 (I378537,I379015,I378778);
not I_22160 (I379091,I379015);
and I_22161 (I379108,I378642,I379091);
nor I_22162 (I378543,I378778,I379108);
nand I_22163 (I378531,I379015,I378905);
not I_22164 (I379186,I2357);
not I_22165 (I379203,I27220);
nor I_22166 (I379220,I27238,I27217);
nand I_22167 (I379237,I379220,I27235);
nor I_22168 (I379254,I379203,I27238);
nand I_22169 (I379271,I379254,I27229);
not I_22170 (I379288,I27238);
not I_22171 (I379305,I379288);
not I_22172 (I379322,I27232);
nor I_22173 (I379339,I379322,I27226);
and I_22174 (I379356,I379339,I27223);
or I_22175 (I379373,I379356,I27214);
DFFARX1 I_22176  ( .D(I379373), .CLK(I2350), .RSTB(I379186), .Q(I379390) );
nand I_22177 (I379407,I379203,I27232);
or I_22178 (I379175,I379407,I379390);
not I_22179 (I379438,I379407);
nor I_22180 (I379455,I379390,I379438);
and I_22181 (I379472,I379288,I379455);
nand I_22182 (I379148,I379407,I379305);
DFFARX1 I_22183  ( .D(I27244), .CLK(I2350), .RSTB(I379186), .Q(I379503) );
or I_22184 (I379169,I379503,I379390);
nor I_22185 (I379534,I379503,I379271);
nor I_22186 (I379551,I379503,I379305);
nand I_22187 (I379154,I379237,I379551);
or I_22188 (I379582,I379503,I379472);
DFFARX1 I_22189  ( .D(I379582), .CLK(I2350), .RSTB(I379186), .Q(I379151) );
not I_22190 (I379157,I379503);
DFFARX1 I_22191  ( .D(I27241), .CLK(I2350), .RSTB(I379186), .Q(I379627) );
not I_22192 (I379644,I379627);
nor I_22193 (I379661,I379644,I379237);
DFFARX1 I_22194  ( .D(I379661), .CLK(I2350), .RSTB(I379186), .Q(I379163) );
nor I_22195 (I379178,I379503,I379644);
nor I_22196 (I379166,I379644,I379407);
not I_22197 (I379720,I379644);
and I_22198 (I379737,I379271,I379720);
nor I_22199 (I379172,I379407,I379737);
nand I_22200 (I379160,I379644,I379534);
not I_22201 (I379815,I2357);
not I_22202 (I379832,I49830);
nor I_22203 (I379849,I49848,I49827);
nand I_22204 (I379866,I379849,I49845);
nor I_22205 (I379883,I379832,I49848);
nand I_22206 (I379900,I379883,I49839);
not I_22207 (I379917,I49848);
not I_22208 (I379934,I379917);
not I_22209 (I379951,I49842);
nor I_22210 (I379968,I379951,I49836);
and I_22211 (I379985,I379968,I49833);
or I_22212 (I380002,I379985,I49824);
DFFARX1 I_22213  ( .D(I380002), .CLK(I2350), .RSTB(I379815), .Q(I380019) );
nand I_22214 (I380036,I379832,I49842);
or I_22215 (I379804,I380036,I380019);
not I_22216 (I380067,I380036);
nor I_22217 (I380084,I380019,I380067);
and I_22218 (I380101,I379917,I380084);
nand I_22219 (I379777,I380036,I379934);
DFFARX1 I_22220  ( .D(I49854), .CLK(I2350), .RSTB(I379815), .Q(I380132) );
or I_22221 (I379798,I380132,I380019);
nor I_22222 (I380163,I380132,I379900);
nor I_22223 (I380180,I380132,I379934);
nand I_22224 (I379783,I379866,I380180);
or I_22225 (I380211,I380132,I380101);
DFFARX1 I_22226  ( .D(I380211), .CLK(I2350), .RSTB(I379815), .Q(I379780) );
not I_22227 (I379786,I380132);
DFFARX1 I_22228  ( .D(I49851), .CLK(I2350), .RSTB(I379815), .Q(I380256) );
not I_22229 (I380273,I380256);
nor I_22230 (I380290,I380273,I379866);
DFFARX1 I_22231  ( .D(I380290), .CLK(I2350), .RSTB(I379815), .Q(I379792) );
nor I_22232 (I379807,I380132,I380273);
nor I_22233 (I379795,I380273,I380036);
not I_22234 (I380349,I380273);
and I_22235 (I380366,I379900,I380349);
nor I_22236 (I379801,I380036,I380366);
nand I_22237 (I379789,I380273,I380163);
not I_22238 (I380444,I2357);
not I_22239 (I380461,I129380);
nor I_22240 (I380478,I129356,I129371);
nand I_22241 (I380495,I380478,I129353);
nor I_22242 (I380512,I380461,I129356);
nand I_22243 (I380529,I380512,I129368);
not I_22244 (I380546,I129356);
not I_22245 (I380563,I380546);
not I_22246 (I380580,I129359);
nor I_22247 (I380597,I380580,I129374);
and I_22248 (I380614,I380597,I129365);
or I_22249 (I380631,I380614,I129350);
DFFARX1 I_22250  ( .D(I380631), .CLK(I2350), .RSTB(I380444), .Q(I380648) );
nand I_22251 (I380665,I380461,I129359);
or I_22252 (I380433,I380665,I380648);
not I_22253 (I380696,I380665);
nor I_22254 (I380713,I380648,I380696);
and I_22255 (I380730,I380546,I380713);
nand I_22256 (I380406,I380665,I380563);
DFFARX1 I_22257  ( .D(I129362), .CLK(I2350), .RSTB(I380444), .Q(I380761) );
or I_22258 (I380427,I380761,I380648);
nor I_22259 (I380792,I380761,I380529);
nor I_22260 (I380809,I380761,I380563);
nand I_22261 (I380412,I380495,I380809);
or I_22262 (I380840,I380761,I380730);
DFFARX1 I_22263  ( .D(I380840), .CLK(I2350), .RSTB(I380444), .Q(I380409) );
not I_22264 (I380415,I380761);
DFFARX1 I_22265  ( .D(I129377), .CLK(I2350), .RSTB(I380444), .Q(I380885) );
not I_22266 (I380902,I380885);
nor I_22267 (I380919,I380902,I380495);
DFFARX1 I_22268  ( .D(I380919), .CLK(I2350), .RSTB(I380444), .Q(I380421) );
nor I_22269 (I380436,I380761,I380902);
nor I_22270 (I380424,I380902,I380665);
not I_22271 (I380978,I380902);
and I_22272 (I380995,I380529,I380978);
nor I_22273 (I380430,I380665,I380995);
nand I_22274 (I380418,I380902,I380792);
not I_22275 (I381073,I2357);
nand I_22276 (I381090,I132340,I132328);
and I_22277 (I381107,I381090,I132352);
DFFARX1 I_22278  ( .D(I381107), .CLK(I2350), .RSTB(I381073), .Q(I381124) );
not I_22279 (I381062,I381124);
DFFARX1 I_22280  ( .D(I381124), .CLK(I2350), .RSTB(I381073), .Q(I381155) );
not I_22281 (I381050,I381155);
nor I_22282 (I381186,I132346,I132328);
not I_22283 (I381203,I381186);
nor I_22284 (I381220,I381124,I381203);
DFFARX1 I_22285  ( .D(I132325), .CLK(I2350), .RSTB(I381073), .Q(I381237) );
not I_22286 (I381254,I381237);
nand I_22287 (I381053,I381237,I381203);
DFFARX1 I_22288  ( .D(I381237), .CLK(I2350), .RSTB(I381073), .Q(I381285) );
and I_22289 (I381038,I381124,I381285);
nand I_22290 (I381316,I132355,I132337);
and I_22291 (I381333,I381316,I132343);
DFFARX1 I_22292  ( .D(I381333), .CLK(I2350), .RSTB(I381073), .Q(I381350) );
nor I_22293 (I381367,I381350,I381254);
and I_22294 (I381384,I381186,I381367);
nor I_22295 (I381401,I381350,I381124);
DFFARX1 I_22296  ( .D(I381350), .CLK(I2350), .RSTB(I381073), .Q(I381044) );
DFFARX1 I_22297  ( .D(I132331), .CLK(I2350), .RSTB(I381073), .Q(I381432) );
and I_22298 (I381449,I381432,I132349);
or I_22299 (I381466,I381449,I381384);
DFFARX1 I_22300  ( .D(I381466), .CLK(I2350), .RSTB(I381073), .Q(I381056) );
nand I_22301 (I381065,I381449,I381401);
DFFARX1 I_22302  ( .D(I381449), .CLK(I2350), .RSTB(I381073), .Q(I381035) );
DFFARX1 I_22303  ( .D(I132334), .CLK(I2350), .RSTB(I381073), .Q(I381525) );
nand I_22304 (I381059,I381525,I381220);
DFFARX1 I_22305  ( .D(I381525), .CLK(I2350), .RSTB(I381073), .Q(I381047) );
nand I_22306 (I381570,I381525,I381186);
and I_22307 (I381587,I381237,I381570);
DFFARX1 I_22308  ( .D(I381587), .CLK(I2350), .RSTB(I381073), .Q(I381041) );
not I_22309 (I381651,I2357);
nand I_22310 (I381668,I47261,I47246);
and I_22311 (I381685,I381668,I47240);
DFFARX1 I_22312  ( .D(I381685), .CLK(I2350), .RSTB(I381651), .Q(I381702) );
not I_22313 (I381640,I381702);
DFFARX1 I_22314  ( .D(I381702), .CLK(I2350), .RSTB(I381651), .Q(I381733) );
not I_22315 (I381628,I381733);
nor I_22316 (I381764,I47267,I47246);
not I_22317 (I381781,I381764);
nor I_22318 (I381798,I381702,I381781);
DFFARX1 I_22319  ( .D(I47270), .CLK(I2350), .RSTB(I381651), .Q(I381815) );
not I_22320 (I381832,I381815);
nand I_22321 (I381631,I381815,I381781);
DFFARX1 I_22322  ( .D(I381815), .CLK(I2350), .RSTB(I381651), .Q(I381863) );
and I_22323 (I381616,I381702,I381863);
nand I_22324 (I381894,I47252,I47255);
and I_22325 (I381911,I381894,I47258);
DFFARX1 I_22326  ( .D(I381911), .CLK(I2350), .RSTB(I381651), .Q(I381928) );
nor I_22327 (I381945,I381928,I381832);
and I_22328 (I381962,I381764,I381945);
nor I_22329 (I381979,I381928,I381702);
DFFARX1 I_22330  ( .D(I381928), .CLK(I2350), .RSTB(I381651), .Q(I381622) );
DFFARX1 I_22331  ( .D(I47264), .CLK(I2350), .RSTB(I381651), .Q(I382010) );
and I_22332 (I382027,I382010,I47249);
or I_22333 (I382044,I382027,I381962);
DFFARX1 I_22334  ( .D(I382044), .CLK(I2350), .RSTB(I381651), .Q(I381634) );
nand I_22335 (I381643,I382027,I381979);
DFFARX1 I_22336  ( .D(I382027), .CLK(I2350), .RSTB(I381651), .Q(I381613) );
DFFARX1 I_22337  ( .D(I47243), .CLK(I2350), .RSTB(I381651), .Q(I382103) );
nand I_22338 (I381637,I382103,I381798);
DFFARX1 I_22339  ( .D(I382103), .CLK(I2350), .RSTB(I381651), .Q(I381625) );
nand I_22340 (I382148,I382103,I381764);
and I_22341 (I382165,I381815,I382148);
DFFARX1 I_22342  ( .D(I382165), .CLK(I2350), .RSTB(I381651), .Q(I381619) );
not I_22343 (I382229,I2357);
nand I_22344 (I382246,I14726,I14711);
and I_22345 (I382263,I382246,I14720);
DFFARX1 I_22346  ( .D(I382263), .CLK(I2350), .RSTB(I382229), .Q(I382280) );
not I_22347 (I382218,I382280);
DFFARX1 I_22348  ( .D(I382280), .CLK(I2350), .RSTB(I382229), .Q(I382311) );
not I_22349 (I382206,I382311);
nor I_22350 (I382342,I14732,I14711);
not I_22351 (I382359,I382342);
nor I_22352 (I382376,I382280,I382359);
DFFARX1 I_22353  ( .D(I14723), .CLK(I2350), .RSTB(I382229), .Q(I382393) );
not I_22354 (I382410,I382393);
nand I_22355 (I382209,I382393,I382359);
DFFARX1 I_22356  ( .D(I382393), .CLK(I2350), .RSTB(I382229), .Q(I382441) );
and I_22357 (I382194,I382280,I382441);
nand I_22358 (I382472,I14708,I14702);
and I_22359 (I382489,I382472,I14717);
DFFARX1 I_22360  ( .D(I382489), .CLK(I2350), .RSTB(I382229), .Q(I382506) );
nor I_22361 (I382523,I382506,I382410);
and I_22362 (I382540,I382342,I382523);
nor I_22363 (I382557,I382506,I382280);
DFFARX1 I_22364  ( .D(I382506), .CLK(I2350), .RSTB(I382229), .Q(I382200) );
DFFARX1 I_22365  ( .D(I14705), .CLK(I2350), .RSTB(I382229), .Q(I382588) );
and I_22366 (I382605,I382588,I14729);
or I_22367 (I382622,I382605,I382540);
DFFARX1 I_22368  ( .D(I382622), .CLK(I2350), .RSTB(I382229), .Q(I382212) );
nand I_22369 (I382221,I382605,I382557);
DFFARX1 I_22370  ( .D(I382605), .CLK(I2350), .RSTB(I382229), .Q(I382191) );
DFFARX1 I_22371  ( .D(I14714), .CLK(I2350), .RSTB(I382229), .Q(I382681) );
nand I_22372 (I382215,I382681,I382376);
DFFARX1 I_22373  ( .D(I382681), .CLK(I2350), .RSTB(I382229), .Q(I382203) );
nand I_22374 (I382726,I382681,I382342);
and I_22375 (I382743,I382393,I382726);
DFFARX1 I_22376  ( .D(I382743), .CLK(I2350), .RSTB(I382229), .Q(I382197) );
not I_22377 (I382807,I2357);
nand I_22378 (I382824,I193373,I193376);
and I_22379 (I382841,I382824,I193355);
DFFARX1 I_22380  ( .D(I382841), .CLK(I2350), .RSTB(I382807), .Q(I382858) );
not I_22381 (I382796,I382858);
DFFARX1 I_22382  ( .D(I382858), .CLK(I2350), .RSTB(I382807), .Q(I382889) );
not I_22383 (I382784,I382889);
nor I_22384 (I382920,I193370,I193376);
not I_22385 (I382937,I382920);
nor I_22386 (I382954,I382858,I382937);
DFFARX1 I_22387  ( .D(I193379), .CLK(I2350), .RSTB(I382807), .Q(I382971) );
not I_22388 (I382988,I382971);
nand I_22389 (I382787,I382971,I382937);
DFFARX1 I_22390  ( .D(I382971), .CLK(I2350), .RSTB(I382807), .Q(I383019) );
and I_22391 (I382772,I382858,I383019);
nand I_22392 (I383050,I193367,I193385);
and I_22393 (I383067,I383050,I193361);
DFFARX1 I_22394  ( .D(I383067), .CLK(I2350), .RSTB(I382807), .Q(I383084) );
nor I_22395 (I383101,I383084,I382988);
and I_22396 (I383118,I382920,I383101);
nor I_22397 (I383135,I383084,I382858);
DFFARX1 I_22398  ( .D(I383084), .CLK(I2350), .RSTB(I382807), .Q(I382778) );
DFFARX1 I_22399  ( .D(I193358), .CLK(I2350), .RSTB(I382807), .Q(I383166) );
and I_22400 (I383183,I383166,I193364);
or I_22401 (I383200,I383183,I383118);
DFFARX1 I_22402  ( .D(I383200), .CLK(I2350), .RSTB(I382807), .Q(I382790) );
nand I_22403 (I382799,I383183,I383135);
DFFARX1 I_22404  ( .D(I383183), .CLK(I2350), .RSTB(I382807), .Q(I382769) );
DFFARX1 I_22405  ( .D(I193382), .CLK(I2350), .RSTB(I382807), .Q(I383259) );
nand I_22406 (I382793,I383259,I382954);
DFFARX1 I_22407  ( .D(I383259), .CLK(I2350), .RSTB(I382807), .Q(I382781) );
nand I_22408 (I383304,I383259,I382920);
and I_22409 (I383321,I382971,I383304);
DFFARX1 I_22410  ( .D(I383321), .CLK(I2350), .RSTB(I382807), .Q(I382775) );
not I_22411 (I383385,I2357);
nand I_22412 (I383402,I96642,I96672);
and I_22413 (I383419,I383402,I96654);
DFFARX1 I_22414  ( .D(I383419), .CLK(I2350), .RSTB(I383385), .Q(I383436) );
not I_22415 (I383374,I383436);
DFFARX1 I_22416  ( .D(I383436), .CLK(I2350), .RSTB(I383385), .Q(I383467) );
not I_22417 (I383362,I383467);
nor I_22418 (I383498,I96651,I96672);
not I_22419 (I383515,I383498);
nor I_22420 (I383532,I383436,I383515);
DFFARX1 I_22421  ( .D(I96645), .CLK(I2350), .RSTB(I383385), .Q(I383549) );
not I_22422 (I383566,I383549);
nand I_22423 (I383365,I383549,I383515);
DFFARX1 I_22424  ( .D(I383549), .CLK(I2350), .RSTB(I383385), .Q(I383597) );
and I_22425 (I383350,I383436,I383597);
nand I_22426 (I383628,I96648,I96663);
and I_22427 (I383645,I383628,I96660);
DFFARX1 I_22428  ( .D(I383645), .CLK(I2350), .RSTB(I383385), .Q(I383662) );
nor I_22429 (I383679,I383662,I383566);
and I_22430 (I383696,I383498,I383679);
nor I_22431 (I383713,I383662,I383436);
DFFARX1 I_22432  ( .D(I383662), .CLK(I2350), .RSTB(I383385), .Q(I383356) );
DFFARX1 I_22433  ( .D(I96657), .CLK(I2350), .RSTB(I383385), .Q(I383744) );
and I_22434 (I383761,I383744,I96669);
or I_22435 (I383778,I383761,I383696);
DFFARX1 I_22436  ( .D(I383778), .CLK(I2350), .RSTB(I383385), .Q(I383368) );
nand I_22437 (I383377,I383761,I383713);
DFFARX1 I_22438  ( .D(I383761), .CLK(I2350), .RSTB(I383385), .Q(I383347) );
DFFARX1 I_22439  ( .D(I96666), .CLK(I2350), .RSTB(I383385), .Q(I383837) );
nand I_22440 (I383371,I383837,I383532);
DFFARX1 I_22441  ( .D(I383837), .CLK(I2350), .RSTB(I383385), .Q(I383359) );
nand I_22442 (I383882,I383837,I383498);
and I_22443 (I383899,I383549,I383882);
DFFARX1 I_22444  ( .D(I383899), .CLK(I2350), .RSTB(I383385), .Q(I383353) );
not I_22445 (I383963,I2357);
nand I_22446 (I383980,I304063,I304045);
and I_22447 (I383997,I383980,I304060);
DFFARX1 I_22448  ( .D(I383997), .CLK(I2350), .RSTB(I383963), .Q(I384014) );
not I_22449 (I383952,I384014);
DFFARX1 I_22450  ( .D(I384014), .CLK(I2350), .RSTB(I383963), .Q(I384045) );
not I_22451 (I383940,I384045);
nor I_22452 (I384076,I304051,I304045);
not I_22453 (I384093,I384076);
nor I_22454 (I384110,I384014,I384093);
DFFARX1 I_22455  ( .D(I304066), .CLK(I2350), .RSTB(I383963), .Q(I384127) );
not I_22456 (I384144,I384127);
nand I_22457 (I383943,I384127,I384093);
DFFARX1 I_22458  ( .D(I384127), .CLK(I2350), .RSTB(I383963), .Q(I384175) );
and I_22459 (I383928,I384014,I384175);
nand I_22460 (I384206,I304042,I304048);
and I_22461 (I384223,I384206,I304054);
DFFARX1 I_22462  ( .D(I384223), .CLK(I2350), .RSTB(I383963), .Q(I384240) );
nor I_22463 (I384257,I384240,I384144);
and I_22464 (I384274,I384076,I384257);
nor I_22465 (I384291,I384240,I384014);
DFFARX1 I_22466  ( .D(I384240), .CLK(I2350), .RSTB(I383963), .Q(I383934) );
DFFARX1 I_22467  ( .D(I304069), .CLK(I2350), .RSTB(I383963), .Q(I384322) );
and I_22468 (I384339,I384322,I304057);
or I_22469 (I384356,I384339,I384274);
DFFARX1 I_22470  ( .D(I384356), .CLK(I2350), .RSTB(I383963), .Q(I383946) );
nand I_22471 (I383955,I384339,I384291);
DFFARX1 I_22472  ( .D(I384339), .CLK(I2350), .RSTB(I383963), .Q(I383925) );
DFFARX1 I_22473  ( .D(I304072), .CLK(I2350), .RSTB(I383963), .Q(I384415) );
nand I_22474 (I383949,I384415,I384110);
DFFARX1 I_22475  ( .D(I384415), .CLK(I2350), .RSTB(I383963), .Q(I383937) );
nand I_22476 (I384460,I384415,I384076);
and I_22477 (I384477,I384127,I384460);
DFFARX1 I_22478  ( .D(I384477), .CLK(I2350), .RSTB(I383963), .Q(I383931) );
not I_22479 (I384541,I2357);
nand I_22480 (I384558,I189403,I189400);
and I_22481 (I384575,I384558,I189424);
DFFARX1 I_22482  ( .D(I384575), .CLK(I2350), .RSTB(I384541), .Q(I384592) );
not I_22483 (I384530,I384592);
DFFARX1 I_22484  ( .D(I384592), .CLK(I2350), .RSTB(I384541), .Q(I384623) );
not I_22485 (I384518,I384623);
nor I_22486 (I384654,I189406,I189400);
not I_22487 (I384671,I384654);
nor I_22488 (I384688,I384592,I384671);
DFFARX1 I_22489  ( .D(I189421), .CLK(I2350), .RSTB(I384541), .Q(I384705) );
not I_22490 (I384722,I384705);
nand I_22491 (I384521,I384705,I384671);
DFFARX1 I_22492  ( .D(I384705), .CLK(I2350), .RSTB(I384541), .Q(I384753) );
and I_22493 (I384506,I384592,I384753);
nand I_22494 (I384784,I189409,I189394);
and I_22495 (I384801,I384784,I189412);
DFFARX1 I_22496  ( .D(I384801), .CLK(I2350), .RSTB(I384541), .Q(I384818) );
nor I_22497 (I384835,I384818,I384722);
and I_22498 (I384852,I384654,I384835);
nor I_22499 (I384869,I384818,I384592);
DFFARX1 I_22500  ( .D(I384818), .CLK(I2350), .RSTB(I384541), .Q(I384512) );
DFFARX1 I_22501  ( .D(I189415), .CLK(I2350), .RSTB(I384541), .Q(I384900) );
and I_22502 (I384917,I384900,I189418);
or I_22503 (I384934,I384917,I384852);
DFFARX1 I_22504  ( .D(I384934), .CLK(I2350), .RSTB(I384541), .Q(I384524) );
nand I_22505 (I384533,I384917,I384869);
DFFARX1 I_22506  ( .D(I384917), .CLK(I2350), .RSTB(I384541), .Q(I384503) );
DFFARX1 I_22507  ( .D(I189397), .CLK(I2350), .RSTB(I384541), .Q(I384993) );
nand I_22508 (I384527,I384993,I384688);
DFFARX1 I_22509  ( .D(I384993), .CLK(I2350), .RSTB(I384541), .Q(I384515) );
nand I_22510 (I385038,I384993,I384654);
and I_22511 (I385055,I384705,I385038);
DFFARX1 I_22512  ( .D(I385055), .CLK(I2350), .RSTB(I384541), .Q(I384509) );
not I_22513 (I385119,I2357);
nand I_22514 (I385136,I164209,I164206);
and I_22515 (I385153,I385136,I164230);
DFFARX1 I_22516  ( .D(I385153), .CLK(I2350), .RSTB(I385119), .Q(I385170) );
not I_22517 (I385108,I385170);
DFFARX1 I_22518  ( .D(I385170), .CLK(I2350), .RSTB(I385119), .Q(I385201) );
not I_22519 (I385096,I385201);
nor I_22520 (I385232,I164212,I164206);
not I_22521 (I385249,I385232);
nor I_22522 (I385266,I385170,I385249);
DFFARX1 I_22523  ( .D(I164227), .CLK(I2350), .RSTB(I385119), .Q(I385283) );
not I_22524 (I385300,I385283);
nand I_22525 (I385099,I385283,I385249);
DFFARX1 I_22526  ( .D(I385283), .CLK(I2350), .RSTB(I385119), .Q(I385331) );
and I_22527 (I385084,I385170,I385331);
nand I_22528 (I385362,I164215,I164200);
and I_22529 (I385379,I385362,I164218);
DFFARX1 I_22530  ( .D(I385379), .CLK(I2350), .RSTB(I385119), .Q(I385396) );
nor I_22531 (I385413,I385396,I385300);
and I_22532 (I385430,I385232,I385413);
nor I_22533 (I385447,I385396,I385170);
DFFARX1 I_22534  ( .D(I385396), .CLK(I2350), .RSTB(I385119), .Q(I385090) );
DFFARX1 I_22535  ( .D(I164221), .CLK(I2350), .RSTB(I385119), .Q(I385478) );
and I_22536 (I385495,I385478,I164224);
or I_22537 (I385512,I385495,I385430);
DFFARX1 I_22538  ( .D(I385512), .CLK(I2350), .RSTB(I385119), .Q(I385102) );
nand I_22539 (I385111,I385495,I385447);
DFFARX1 I_22540  ( .D(I385495), .CLK(I2350), .RSTB(I385119), .Q(I385081) );
DFFARX1 I_22541  ( .D(I164203), .CLK(I2350), .RSTB(I385119), .Q(I385571) );
nand I_22542 (I385105,I385571,I385266);
DFFARX1 I_22543  ( .D(I385571), .CLK(I2350), .RSTB(I385119), .Q(I385093) );
nand I_22544 (I385616,I385571,I385232);
and I_22545 (I385633,I385283,I385616);
DFFARX1 I_22546  ( .D(I385633), .CLK(I2350), .RSTB(I385119), .Q(I385087) );
not I_22547 (I385697,I2357);
nand I_22548 (I385714,I190066,I190063);
and I_22549 (I385731,I385714,I190087);
DFFARX1 I_22550  ( .D(I385731), .CLK(I2350), .RSTB(I385697), .Q(I385748) );
not I_22551 (I385686,I385748);
DFFARX1 I_22552  ( .D(I385748), .CLK(I2350), .RSTB(I385697), .Q(I385779) );
not I_22553 (I385674,I385779);
nor I_22554 (I385810,I190069,I190063);
not I_22555 (I385827,I385810);
nor I_22556 (I385844,I385748,I385827);
DFFARX1 I_22557  ( .D(I190084), .CLK(I2350), .RSTB(I385697), .Q(I385861) );
not I_22558 (I385878,I385861);
nand I_22559 (I385677,I385861,I385827);
DFFARX1 I_22560  ( .D(I385861), .CLK(I2350), .RSTB(I385697), .Q(I385909) );
and I_22561 (I385662,I385748,I385909);
nand I_22562 (I385940,I190072,I190057);
and I_22563 (I385957,I385940,I190075);
DFFARX1 I_22564  ( .D(I385957), .CLK(I2350), .RSTB(I385697), .Q(I385974) );
nor I_22565 (I385991,I385974,I385878);
and I_22566 (I386008,I385810,I385991);
nor I_22567 (I386025,I385974,I385748);
DFFARX1 I_22568  ( .D(I385974), .CLK(I2350), .RSTB(I385697), .Q(I385668) );
DFFARX1 I_22569  ( .D(I190078), .CLK(I2350), .RSTB(I385697), .Q(I386056) );
and I_22570 (I386073,I386056,I190081);
or I_22571 (I386090,I386073,I386008);
DFFARX1 I_22572  ( .D(I386090), .CLK(I2350), .RSTB(I385697), .Q(I385680) );
nand I_22573 (I385689,I386073,I386025);
DFFARX1 I_22574  ( .D(I386073), .CLK(I2350), .RSTB(I385697), .Q(I385659) );
DFFARX1 I_22575  ( .D(I190060), .CLK(I2350), .RSTB(I385697), .Q(I386149) );
nand I_22576 (I385683,I386149,I385844);
DFFARX1 I_22577  ( .D(I386149), .CLK(I2350), .RSTB(I385697), .Q(I385671) );
nand I_22578 (I386194,I386149,I385810);
and I_22579 (I386211,I385861,I386194);
DFFARX1 I_22580  ( .D(I386211), .CLK(I2350), .RSTB(I385697), .Q(I385665) );
not I_22581 (I386275,I2357);
nand I_22582 (I386292,I106587,I106617);
and I_22583 (I386309,I386292,I106599);
DFFARX1 I_22584  ( .D(I386309), .CLK(I2350), .RSTB(I386275), .Q(I386326) );
not I_22585 (I386264,I386326);
DFFARX1 I_22586  ( .D(I386326), .CLK(I2350), .RSTB(I386275), .Q(I386357) );
not I_22587 (I386252,I386357);
nor I_22588 (I386388,I106596,I106617);
not I_22589 (I386405,I386388);
nor I_22590 (I386422,I386326,I386405);
DFFARX1 I_22591  ( .D(I106590), .CLK(I2350), .RSTB(I386275), .Q(I386439) );
not I_22592 (I386456,I386439);
nand I_22593 (I386255,I386439,I386405);
DFFARX1 I_22594  ( .D(I386439), .CLK(I2350), .RSTB(I386275), .Q(I386487) );
and I_22595 (I386240,I386326,I386487);
nand I_22596 (I386518,I106593,I106608);
and I_22597 (I386535,I386518,I106605);
DFFARX1 I_22598  ( .D(I386535), .CLK(I2350), .RSTB(I386275), .Q(I386552) );
nor I_22599 (I386569,I386552,I386456);
and I_22600 (I386586,I386388,I386569);
nor I_22601 (I386603,I386552,I386326);
DFFARX1 I_22602  ( .D(I386552), .CLK(I2350), .RSTB(I386275), .Q(I386246) );
DFFARX1 I_22603  ( .D(I106602), .CLK(I2350), .RSTB(I386275), .Q(I386634) );
and I_22604 (I386651,I386634,I106614);
or I_22605 (I386668,I386651,I386586);
DFFARX1 I_22606  ( .D(I386668), .CLK(I2350), .RSTB(I386275), .Q(I386258) );
nand I_22607 (I386267,I386651,I386603);
DFFARX1 I_22608  ( .D(I386651), .CLK(I2350), .RSTB(I386275), .Q(I386237) );
DFFARX1 I_22609  ( .D(I106611), .CLK(I2350), .RSTB(I386275), .Q(I386727) );
nand I_22610 (I386261,I386727,I386422);
DFFARX1 I_22611  ( .D(I386727), .CLK(I2350), .RSTB(I386275), .Q(I386249) );
nand I_22612 (I386772,I386727,I386388);
and I_22613 (I386789,I386439,I386772);
DFFARX1 I_22614  ( .D(I386789), .CLK(I2350), .RSTB(I386275), .Q(I386243) );
not I_22615 (I386853,I2357);
nand I_22616 (I386870,I268473,I268491);
and I_22617 (I386887,I386870,I268467);
DFFARX1 I_22618  ( .D(I386887), .CLK(I2350), .RSTB(I386853), .Q(I386904) );
not I_22619 (I386842,I386904);
DFFARX1 I_22620  ( .D(I386904), .CLK(I2350), .RSTB(I386853), .Q(I386935) );
not I_22621 (I386830,I386935);
nor I_22622 (I386966,I268479,I268491);
not I_22623 (I386983,I386966);
nor I_22624 (I387000,I386904,I386983);
DFFARX1 I_22625  ( .D(I268470), .CLK(I2350), .RSTB(I386853), .Q(I387017) );
not I_22626 (I387034,I387017);
nand I_22627 (I386833,I387017,I386983);
DFFARX1 I_22628  ( .D(I387017), .CLK(I2350), .RSTB(I386853), .Q(I387065) );
and I_22629 (I386818,I386904,I387065);
nand I_22630 (I387096,I268485,I268464);
and I_22631 (I387113,I387096,I268482);
DFFARX1 I_22632  ( .D(I387113), .CLK(I2350), .RSTB(I386853), .Q(I387130) );
nor I_22633 (I387147,I387130,I387034);
and I_22634 (I387164,I386966,I387147);
nor I_22635 (I387181,I387130,I386904);
DFFARX1 I_22636  ( .D(I387130), .CLK(I2350), .RSTB(I386853), .Q(I386824) );
DFFARX1 I_22637  ( .D(I268488), .CLK(I2350), .RSTB(I386853), .Q(I387212) );
and I_22638 (I387229,I387212,I268476);
or I_22639 (I387246,I387229,I387164);
DFFARX1 I_22640  ( .D(I387246), .CLK(I2350), .RSTB(I386853), .Q(I386836) );
nand I_22641 (I386845,I387229,I387181);
DFFARX1 I_22642  ( .D(I387229), .CLK(I2350), .RSTB(I386853), .Q(I386815) );
DFFARX1 I_22643  ( .D(I268461), .CLK(I2350), .RSTB(I386853), .Q(I387305) );
nand I_22644 (I386839,I387305,I387000);
DFFARX1 I_22645  ( .D(I387305), .CLK(I2350), .RSTB(I386853), .Q(I386827) );
nand I_22646 (I387350,I387305,I386966);
and I_22647 (I387367,I387017,I387350);
DFFARX1 I_22648  ( .D(I387367), .CLK(I2350), .RSTB(I386853), .Q(I386821) );
not I_22649 (I387431,I2357);
nand I_22650 (I387448,I22019,I22004);
and I_22651 (I387465,I387448,I22013);
DFFARX1 I_22652  ( .D(I387465), .CLK(I2350), .RSTB(I387431), .Q(I387482) );
not I_22653 (I387420,I387482);
DFFARX1 I_22654  ( .D(I387482), .CLK(I2350), .RSTB(I387431), .Q(I387513) );
not I_22655 (I387408,I387513);
nor I_22656 (I387544,I22025,I22004);
not I_22657 (I387561,I387544);
nor I_22658 (I387578,I387482,I387561);
DFFARX1 I_22659  ( .D(I22016), .CLK(I2350), .RSTB(I387431), .Q(I387595) );
not I_22660 (I387612,I387595);
nand I_22661 (I387411,I387595,I387561);
DFFARX1 I_22662  ( .D(I387595), .CLK(I2350), .RSTB(I387431), .Q(I387643) );
and I_22663 (I387396,I387482,I387643);
nand I_22664 (I387674,I22001,I21995);
and I_22665 (I387691,I387674,I22010);
DFFARX1 I_22666  ( .D(I387691), .CLK(I2350), .RSTB(I387431), .Q(I387708) );
nor I_22667 (I387725,I387708,I387612);
and I_22668 (I387742,I387544,I387725);
nor I_22669 (I387759,I387708,I387482);
DFFARX1 I_22670  ( .D(I387708), .CLK(I2350), .RSTB(I387431), .Q(I387402) );
DFFARX1 I_22671  ( .D(I21998), .CLK(I2350), .RSTB(I387431), .Q(I387790) );
and I_22672 (I387807,I387790,I22022);
or I_22673 (I387824,I387807,I387742);
DFFARX1 I_22674  ( .D(I387824), .CLK(I2350), .RSTB(I387431), .Q(I387414) );
nand I_22675 (I387423,I387807,I387759);
DFFARX1 I_22676  ( .D(I387807), .CLK(I2350), .RSTB(I387431), .Q(I387393) );
DFFARX1 I_22677  ( .D(I22007), .CLK(I2350), .RSTB(I387431), .Q(I387883) );
nand I_22678 (I387417,I387883,I387578);
DFFARX1 I_22679  ( .D(I387883), .CLK(I2350), .RSTB(I387431), .Q(I387405) );
nand I_22680 (I387928,I387883,I387544);
and I_22681 (I387945,I387595,I387928);
DFFARX1 I_22682  ( .D(I387945), .CLK(I2350), .RSTB(I387431), .Q(I387399) );
not I_22683 (I388009,I2357);
nand I_22684 (I388026,I196603,I196606);
and I_22685 (I388043,I388026,I196585);
DFFARX1 I_22686  ( .D(I388043), .CLK(I2350), .RSTB(I388009), .Q(I388060) );
not I_22687 (I387998,I388060);
DFFARX1 I_22688  ( .D(I388060), .CLK(I2350), .RSTB(I388009), .Q(I388091) );
not I_22689 (I387986,I388091);
nor I_22690 (I388122,I196600,I196606);
not I_22691 (I388139,I388122);
nor I_22692 (I388156,I388060,I388139);
DFFARX1 I_22693  ( .D(I196609), .CLK(I2350), .RSTB(I388009), .Q(I388173) );
not I_22694 (I388190,I388173);
nand I_22695 (I387989,I388173,I388139);
DFFARX1 I_22696  ( .D(I388173), .CLK(I2350), .RSTB(I388009), .Q(I388221) );
and I_22697 (I387974,I388060,I388221);
nand I_22698 (I388252,I196597,I196615);
and I_22699 (I388269,I388252,I196591);
DFFARX1 I_22700  ( .D(I388269), .CLK(I2350), .RSTB(I388009), .Q(I388286) );
nor I_22701 (I388303,I388286,I388190);
and I_22702 (I388320,I388122,I388303);
nor I_22703 (I388337,I388286,I388060);
DFFARX1 I_22704  ( .D(I388286), .CLK(I2350), .RSTB(I388009), .Q(I387980) );
DFFARX1 I_22705  ( .D(I196588), .CLK(I2350), .RSTB(I388009), .Q(I388368) );
and I_22706 (I388385,I388368,I196594);
or I_22707 (I388402,I388385,I388320);
DFFARX1 I_22708  ( .D(I388402), .CLK(I2350), .RSTB(I388009), .Q(I387992) );
nand I_22709 (I388001,I388385,I388337);
DFFARX1 I_22710  ( .D(I388385), .CLK(I2350), .RSTB(I388009), .Q(I387971) );
DFFARX1 I_22711  ( .D(I196612), .CLK(I2350), .RSTB(I388009), .Q(I388461) );
nand I_22712 (I387995,I388461,I388156);
DFFARX1 I_22713  ( .D(I388461), .CLK(I2350), .RSTB(I388009), .Q(I387983) );
nand I_22714 (I388506,I388461,I388122);
and I_22715 (I388523,I388173,I388506);
DFFARX1 I_22716  ( .D(I388523), .CLK(I2350), .RSTB(I388009), .Q(I387977) );
not I_22717 (I388587,I2357);
nand I_22718 (I388604,I67287,I67272);
and I_22719 (I388621,I388604,I67266);
DFFARX1 I_22720  ( .D(I388621), .CLK(I2350), .RSTB(I388587), .Q(I388638) );
not I_22721 (I388576,I388638);
DFFARX1 I_22722  ( .D(I388638), .CLK(I2350), .RSTB(I388587), .Q(I388669) );
not I_22723 (I388564,I388669);
nor I_22724 (I388700,I67293,I67272);
not I_22725 (I388717,I388700);
nor I_22726 (I388734,I388638,I388717);
DFFARX1 I_22727  ( .D(I67296), .CLK(I2350), .RSTB(I388587), .Q(I388751) );
not I_22728 (I388768,I388751);
nand I_22729 (I388567,I388751,I388717);
DFFARX1 I_22730  ( .D(I388751), .CLK(I2350), .RSTB(I388587), .Q(I388799) );
and I_22731 (I388552,I388638,I388799);
nand I_22732 (I388830,I67278,I67281);
and I_22733 (I388847,I388830,I67284);
DFFARX1 I_22734  ( .D(I388847), .CLK(I2350), .RSTB(I388587), .Q(I388864) );
nor I_22735 (I388881,I388864,I388768);
and I_22736 (I388898,I388700,I388881);
nor I_22737 (I388915,I388864,I388638);
DFFARX1 I_22738  ( .D(I388864), .CLK(I2350), .RSTB(I388587), .Q(I388558) );
DFFARX1 I_22739  ( .D(I67290), .CLK(I2350), .RSTB(I388587), .Q(I388946) );
and I_22740 (I388963,I388946,I67275);
or I_22741 (I388980,I388963,I388898);
DFFARX1 I_22742  ( .D(I388980), .CLK(I2350), .RSTB(I388587), .Q(I388570) );
nand I_22743 (I388579,I388963,I388915);
DFFARX1 I_22744  ( .D(I388963), .CLK(I2350), .RSTB(I388587), .Q(I388549) );
DFFARX1 I_22745  ( .D(I67269), .CLK(I2350), .RSTB(I388587), .Q(I389039) );
nand I_22746 (I388573,I389039,I388734);
DFFARX1 I_22747  ( .D(I389039), .CLK(I2350), .RSTB(I388587), .Q(I388561) );
nand I_22748 (I389084,I389039,I388700);
and I_22749 (I389101,I388751,I389084);
DFFARX1 I_22750  ( .D(I389101), .CLK(I2350), .RSTB(I388587), .Q(I388555) );
not I_22751 (I389165,I2357);
nand I_22752 (I389182,I84083,I84068);
and I_22753 (I389199,I389182,I84062);
DFFARX1 I_22754  ( .D(I389199), .CLK(I2350), .RSTB(I389165), .Q(I389216) );
not I_22755 (I389154,I389216);
DFFARX1 I_22756  ( .D(I389216), .CLK(I2350), .RSTB(I389165), .Q(I389247) );
not I_22757 (I389142,I389247);
nor I_22758 (I389278,I84089,I84068);
not I_22759 (I389295,I389278);
nor I_22760 (I389312,I389216,I389295);
DFFARX1 I_22761  ( .D(I84092), .CLK(I2350), .RSTB(I389165), .Q(I389329) );
not I_22762 (I389346,I389329);
nand I_22763 (I389145,I389329,I389295);
DFFARX1 I_22764  ( .D(I389329), .CLK(I2350), .RSTB(I389165), .Q(I389377) );
and I_22765 (I389130,I389216,I389377);
nand I_22766 (I389408,I84074,I84077);
and I_22767 (I389425,I389408,I84080);
DFFARX1 I_22768  ( .D(I389425), .CLK(I2350), .RSTB(I389165), .Q(I389442) );
nor I_22769 (I389459,I389442,I389346);
and I_22770 (I389476,I389278,I389459);
nor I_22771 (I389493,I389442,I389216);
DFFARX1 I_22772  ( .D(I389442), .CLK(I2350), .RSTB(I389165), .Q(I389136) );
DFFARX1 I_22773  ( .D(I84086), .CLK(I2350), .RSTB(I389165), .Q(I389524) );
and I_22774 (I389541,I389524,I84071);
or I_22775 (I389558,I389541,I389476);
DFFARX1 I_22776  ( .D(I389558), .CLK(I2350), .RSTB(I389165), .Q(I389148) );
nand I_22777 (I389157,I389541,I389493);
DFFARX1 I_22778  ( .D(I389541), .CLK(I2350), .RSTB(I389165), .Q(I389127) );
DFFARX1 I_22779  ( .D(I84065), .CLK(I2350), .RSTB(I389165), .Q(I389617) );
nand I_22780 (I389151,I389617,I389312);
DFFARX1 I_22781  ( .D(I389617), .CLK(I2350), .RSTB(I389165), .Q(I389139) );
nand I_22782 (I389662,I389617,I389278);
and I_22783 (I389679,I389329,I389662);
DFFARX1 I_22784  ( .D(I389679), .CLK(I2350), .RSTB(I389165), .Q(I389133) );
not I_22785 (I389743,I2357);
nand I_22786 (I389760,I200479,I200482);
and I_22787 (I389777,I389760,I200461);
DFFARX1 I_22788  ( .D(I389777), .CLK(I2350), .RSTB(I389743), .Q(I389794) );
not I_22789 (I389732,I389794);
DFFARX1 I_22790  ( .D(I389794), .CLK(I2350), .RSTB(I389743), .Q(I389825) );
not I_22791 (I389720,I389825);
nor I_22792 (I389856,I200476,I200482);
not I_22793 (I389873,I389856);
nor I_22794 (I389890,I389794,I389873);
DFFARX1 I_22795  ( .D(I200485), .CLK(I2350), .RSTB(I389743), .Q(I389907) );
not I_22796 (I389924,I389907);
nand I_22797 (I389723,I389907,I389873);
DFFARX1 I_22798  ( .D(I389907), .CLK(I2350), .RSTB(I389743), .Q(I389955) );
and I_22799 (I389708,I389794,I389955);
nand I_22800 (I389986,I200473,I200491);
and I_22801 (I390003,I389986,I200467);
DFFARX1 I_22802  ( .D(I390003), .CLK(I2350), .RSTB(I389743), .Q(I390020) );
nor I_22803 (I390037,I390020,I389924);
and I_22804 (I390054,I389856,I390037);
nor I_22805 (I390071,I390020,I389794);
DFFARX1 I_22806  ( .D(I390020), .CLK(I2350), .RSTB(I389743), .Q(I389714) );
DFFARX1 I_22807  ( .D(I200464), .CLK(I2350), .RSTB(I389743), .Q(I390102) );
and I_22808 (I390119,I390102,I200470);
or I_22809 (I390136,I390119,I390054);
DFFARX1 I_22810  ( .D(I390136), .CLK(I2350), .RSTB(I389743), .Q(I389726) );
nand I_22811 (I389735,I390119,I390071);
DFFARX1 I_22812  ( .D(I390119), .CLK(I2350), .RSTB(I389743), .Q(I389705) );
DFFARX1 I_22813  ( .D(I200488), .CLK(I2350), .RSTB(I389743), .Q(I390195) );
nand I_22814 (I389729,I390195,I389890);
DFFARX1 I_22815  ( .D(I390195), .CLK(I2350), .RSTB(I389743), .Q(I389717) );
nand I_22816 (I390240,I390195,I389856);
and I_22817 (I390257,I389907,I390240);
DFFARX1 I_22818  ( .D(I390257), .CLK(I2350), .RSTB(I389743), .Q(I389711) );
not I_22819 (I390321,I2357);
nand I_22820 (I390338,I315963,I315942);
and I_22821 (I390355,I390338,I315960);
DFFARX1 I_22822  ( .D(I390355), .CLK(I2350), .RSTB(I390321), .Q(I390372) );
not I_22823 (I390310,I390372);
DFFARX1 I_22824  ( .D(I390372), .CLK(I2350), .RSTB(I390321), .Q(I390403) );
not I_22825 (I390298,I390403);
nor I_22826 (I390434,I315972,I315942);
not I_22827 (I390451,I390434);
nor I_22828 (I390468,I390372,I390451);
DFFARX1 I_22829  ( .D(I315948), .CLK(I2350), .RSTB(I390321), .Q(I390485) );
not I_22830 (I390502,I390485);
nand I_22831 (I390301,I390485,I390451);
DFFARX1 I_22832  ( .D(I390485), .CLK(I2350), .RSTB(I390321), .Q(I390533) );
and I_22833 (I390286,I390372,I390533);
nand I_22834 (I390564,I315957,I315945);
and I_22835 (I390581,I390564,I315969);
DFFARX1 I_22836  ( .D(I390581), .CLK(I2350), .RSTB(I390321), .Q(I390598) );
nor I_22837 (I390615,I390598,I390502);
and I_22838 (I390632,I390434,I390615);
nor I_22839 (I390649,I390598,I390372);
DFFARX1 I_22840  ( .D(I390598), .CLK(I2350), .RSTB(I390321), .Q(I390292) );
DFFARX1 I_22841  ( .D(I315954), .CLK(I2350), .RSTB(I390321), .Q(I390680) );
and I_22842 (I390697,I390680,I315966);
or I_22843 (I390714,I390697,I390632);
DFFARX1 I_22844  ( .D(I390714), .CLK(I2350), .RSTB(I390321), .Q(I390304) );
nand I_22845 (I390313,I390697,I390649);
DFFARX1 I_22846  ( .D(I390697), .CLK(I2350), .RSTB(I390321), .Q(I390283) );
DFFARX1 I_22847  ( .D(I315951), .CLK(I2350), .RSTB(I390321), .Q(I390773) );
nand I_22848 (I390307,I390773,I390468);
DFFARX1 I_22849  ( .D(I390773), .CLK(I2350), .RSTB(I390321), .Q(I390295) );
nand I_22850 (I390818,I390773,I390434);
and I_22851 (I390835,I390485,I390818);
DFFARX1 I_22852  ( .D(I390835), .CLK(I2350), .RSTB(I390321), .Q(I390289) );
not I_22853 (I390899,I2357);
nand I_22854 (I390916,I64703,I64688);
and I_22855 (I390933,I390916,I64682);
DFFARX1 I_22856  ( .D(I390933), .CLK(I2350), .RSTB(I390899), .Q(I390950) );
not I_22857 (I390888,I390950);
DFFARX1 I_22858  ( .D(I390950), .CLK(I2350), .RSTB(I390899), .Q(I390981) );
not I_22859 (I390876,I390981);
nor I_22860 (I391012,I64709,I64688);
not I_22861 (I391029,I391012);
nor I_22862 (I391046,I390950,I391029);
DFFARX1 I_22863  ( .D(I64712), .CLK(I2350), .RSTB(I390899), .Q(I391063) );
not I_22864 (I391080,I391063);
nand I_22865 (I390879,I391063,I391029);
DFFARX1 I_22866  ( .D(I391063), .CLK(I2350), .RSTB(I390899), .Q(I391111) );
and I_22867 (I390864,I390950,I391111);
nand I_22868 (I391142,I64694,I64697);
and I_22869 (I391159,I391142,I64700);
DFFARX1 I_22870  ( .D(I391159), .CLK(I2350), .RSTB(I390899), .Q(I391176) );
nor I_22871 (I391193,I391176,I391080);
and I_22872 (I391210,I391012,I391193);
nor I_22873 (I391227,I391176,I390950);
DFFARX1 I_22874  ( .D(I391176), .CLK(I2350), .RSTB(I390899), .Q(I390870) );
DFFARX1 I_22875  ( .D(I64706), .CLK(I2350), .RSTB(I390899), .Q(I391258) );
and I_22876 (I391275,I391258,I64691);
or I_22877 (I391292,I391275,I391210);
DFFARX1 I_22878  ( .D(I391292), .CLK(I2350), .RSTB(I390899), .Q(I390882) );
nand I_22879 (I390891,I391275,I391227);
DFFARX1 I_22880  ( .D(I391275), .CLK(I2350), .RSTB(I390899), .Q(I390861) );
DFFARX1 I_22881  ( .D(I64685), .CLK(I2350), .RSTB(I390899), .Q(I391351) );
nand I_22882 (I390885,I391351,I391046);
DFFARX1 I_22883  ( .D(I391351), .CLK(I2350), .RSTB(I390899), .Q(I390873) );
nand I_22884 (I391396,I391351,I391012);
and I_22885 (I391413,I391063,I391396);
DFFARX1 I_22886  ( .D(I391413), .CLK(I2350), .RSTB(I390899), .Q(I390867) );
not I_22887 (I391477,I2357);
nand I_22888 (I391494,I260848,I260866);
and I_22889 (I391511,I391494,I260857);
DFFARX1 I_22890  ( .D(I391511), .CLK(I2350), .RSTB(I391477), .Q(I391528) );
not I_22891 (I391466,I391528);
DFFARX1 I_22892  ( .D(I391528), .CLK(I2350), .RSTB(I391477), .Q(I391559) );
not I_22893 (I391454,I391559);
nor I_22894 (I391590,I260854,I260866);
not I_22895 (I391607,I391590);
nor I_22896 (I391624,I391528,I391607);
DFFARX1 I_22897  ( .D(I260845), .CLK(I2350), .RSTB(I391477), .Q(I391641) );
not I_22898 (I391658,I391641);
nand I_22899 (I391457,I391641,I391607);
DFFARX1 I_22900  ( .D(I391641), .CLK(I2350), .RSTB(I391477), .Q(I391689) );
and I_22901 (I391442,I391528,I391689);
nand I_22902 (I391720,I260863,I260875);
and I_22903 (I391737,I391720,I260869);
DFFARX1 I_22904  ( .D(I391737), .CLK(I2350), .RSTB(I391477), .Q(I391754) );
nor I_22905 (I391771,I391754,I391658);
and I_22906 (I391788,I391590,I391771);
nor I_22907 (I391805,I391754,I391528);
DFFARX1 I_22908  ( .D(I391754), .CLK(I2350), .RSTB(I391477), .Q(I391448) );
DFFARX1 I_22909  ( .D(I260851), .CLK(I2350), .RSTB(I391477), .Q(I391836) );
and I_22910 (I391853,I391836,I260860);
or I_22911 (I391870,I391853,I391788);
DFFARX1 I_22912  ( .D(I391870), .CLK(I2350), .RSTB(I391477), .Q(I391460) );
nand I_22913 (I391469,I391853,I391805);
DFFARX1 I_22914  ( .D(I391853), .CLK(I2350), .RSTB(I391477), .Q(I391439) );
DFFARX1 I_22915  ( .D(I260872), .CLK(I2350), .RSTB(I391477), .Q(I391929) );
nand I_22916 (I391463,I391929,I391624);
DFFARX1 I_22917  ( .D(I391929), .CLK(I2350), .RSTB(I391477), .Q(I391451) );
nand I_22918 (I391974,I391929,I391590);
and I_22919 (I391991,I391641,I391974);
DFFARX1 I_22920  ( .D(I391991), .CLK(I2350), .RSTB(I391477), .Q(I391445) );
not I_22921 (I392055,I2357);
nand I_22922 (I392072,I65349,I65334);
and I_22923 (I392089,I392072,I65328);
DFFARX1 I_22924  ( .D(I392089), .CLK(I2350), .RSTB(I392055), .Q(I392106) );
not I_22925 (I392044,I392106);
DFFARX1 I_22926  ( .D(I392106), .CLK(I2350), .RSTB(I392055), .Q(I392137) );
not I_22927 (I392032,I392137);
nor I_22928 (I392168,I65355,I65334);
not I_22929 (I392185,I392168);
nor I_22930 (I392202,I392106,I392185);
DFFARX1 I_22931  ( .D(I65358), .CLK(I2350), .RSTB(I392055), .Q(I392219) );
not I_22932 (I392236,I392219);
nand I_22933 (I392035,I392219,I392185);
DFFARX1 I_22934  ( .D(I392219), .CLK(I2350), .RSTB(I392055), .Q(I392267) );
and I_22935 (I392020,I392106,I392267);
nand I_22936 (I392298,I65340,I65343);
and I_22937 (I392315,I392298,I65346);
DFFARX1 I_22938  ( .D(I392315), .CLK(I2350), .RSTB(I392055), .Q(I392332) );
nor I_22939 (I392349,I392332,I392236);
and I_22940 (I392366,I392168,I392349);
nor I_22941 (I392383,I392332,I392106);
DFFARX1 I_22942  ( .D(I392332), .CLK(I2350), .RSTB(I392055), .Q(I392026) );
DFFARX1 I_22943  ( .D(I65352), .CLK(I2350), .RSTB(I392055), .Q(I392414) );
and I_22944 (I392431,I392414,I65337);
or I_22945 (I392448,I392431,I392366);
DFFARX1 I_22946  ( .D(I392448), .CLK(I2350), .RSTB(I392055), .Q(I392038) );
nand I_22947 (I392047,I392431,I392383);
DFFARX1 I_22948  ( .D(I392431), .CLK(I2350), .RSTB(I392055), .Q(I392017) );
DFFARX1 I_22949  ( .D(I65331), .CLK(I2350), .RSTB(I392055), .Q(I392507) );
nand I_22950 (I392041,I392507,I392202);
DFFARX1 I_22951  ( .D(I392507), .CLK(I2350), .RSTB(I392055), .Q(I392029) );
nand I_22952 (I392552,I392507,I392168);
and I_22953 (I392569,I392219,I392552);
DFFARX1 I_22954  ( .D(I392569), .CLK(I2350), .RSTB(I392055), .Q(I392023) );
not I_22955 (I392633,I2357);
nand I_22956 (I392650,I307633,I307615);
and I_22957 (I392667,I392650,I307630);
DFFARX1 I_22958  ( .D(I392667), .CLK(I2350), .RSTB(I392633), .Q(I392684) );
not I_22959 (I392622,I392684);
DFFARX1 I_22960  ( .D(I392684), .CLK(I2350), .RSTB(I392633), .Q(I392715) );
not I_22961 (I392610,I392715);
nor I_22962 (I392746,I307621,I307615);
not I_22963 (I392763,I392746);
nor I_22964 (I392780,I392684,I392763);
DFFARX1 I_22965  ( .D(I307636), .CLK(I2350), .RSTB(I392633), .Q(I392797) );
not I_22966 (I392814,I392797);
nand I_22967 (I392613,I392797,I392763);
DFFARX1 I_22968  ( .D(I392797), .CLK(I2350), .RSTB(I392633), .Q(I392845) );
and I_22969 (I392598,I392684,I392845);
nand I_22970 (I392876,I307612,I307618);
and I_22971 (I392893,I392876,I307624);
DFFARX1 I_22972  ( .D(I392893), .CLK(I2350), .RSTB(I392633), .Q(I392910) );
nor I_22973 (I392927,I392910,I392814);
and I_22974 (I392944,I392746,I392927);
nor I_22975 (I392961,I392910,I392684);
DFFARX1 I_22976  ( .D(I392910), .CLK(I2350), .RSTB(I392633), .Q(I392604) );
DFFARX1 I_22977  ( .D(I307639), .CLK(I2350), .RSTB(I392633), .Q(I392992) );
and I_22978 (I393009,I392992,I307627);
or I_22979 (I393026,I393009,I392944);
DFFARX1 I_22980  ( .D(I393026), .CLK(I2350), .RSTB(I392633), .Q(I392616) );
nand I_22981 (I392625,I393009,I392961);
DFFARX1 I_22982  ( .D(I393009), .CLK(I2350), .RSTB(I392633), .Q(I392595) );
DFFARX1 I_22983  ( .D(I307642), .CLK(I2350), .RSTB(I392633), .Q(I393085) );
nand I_22984 (I392619,I393085,I392780);
DFFARX1 I_22985  ( .D(I393085), .CLK(I2350), .RSTB(I392633), .Q(I392607) );
nand I_22986 (I393130,I393085,I392746);
and I_22987 (I393147,I392797,I393130);
DFFARX1 I_22988  ( .D(I393147), .CLK(I2350), .RSTB(I392633), .Q(I392601) );
not I_22989 (I393211,I2357);
nand I_22990 (I393228,I307038,I307020);
and I_22991 (I393245,I393228,I307035);
DFFARX1 I_22992  ( .D(I393245), .CLK(I2350), .RSTB(I393211), .Q(I393262) );
not I_22993 (I393200,I393262);
DFFARX1 I_22994  ( .D(I393262), .CLK(I2350), .RSTB(I393211), .Q(I393293) );
not I_22995 (I393188,I393293);
nor I_22996 (I393324,I307026,I307020);
not I_22997 (I393341,I393324);
nor I_22998 (I393358,I393262,I393341);
DFFARX1 I_22999  ( .D(I307041), .CLK(I2350), .RSTB(I393211), .Q(I393375) );
not I_23000 (I393392,I393375);
nand I_23001 (I393191,I393375,I393341);
DFFARX1 I_23002  ( .D(I393375), .CLK(I2350), .RSTB(I393211), .Q(I393423) );
and I_23003 (I393176,I393262,I393423);
nand I_23004 (I393454,I307017,I307023);
and I_23005 (I393471,I393454,I307029);
DFFARX1 I_23006  ( .D(I393471), .CLK(I2350), .RSTB(I393211), .Q(I393488) );
nor I_23007 (I393505,I393488,I393392);
and I_23008 (I393522,I393324,I393505);
nor I_23009 (I393539,I393488,I393262);
DFFARX1 I_23010  ( .D(I393488), .CLK(I2350), .RSTB(I393211), .Q(I393182) );
DFFARX1 I_23011  ( .D(I307044), .CLK(I2350), .RSTB(I393211), .Q(I393570) );
and I_23012 (I393587,I393570,I307032);
or I_23013 (I393604,I393587,I393522);
DFFARX1 I_23014  ( .D(I393604), .CLK(I2350), .RSTB(I393211), .Q(I393194) );
nand I_23015 (I393203,I393587,I393539);
DFFARX1 I_23016  ( .D(I393587), .CLK(I2350), .RSTB(I393211), .Q(I393173) );
DFFARX1 I_23017  ( .D(I307047), .CLK(I2350), .RSTB(I393211), .Q(I393663) );
nand I_23018 (I393197,I393663,I393358);
DFFARX1 I_23019  ( .D(I393663), .CLK(I2350), .RSTB(I393211), .Q(I393185) );
nand I_23020 (I393708,I393663,I393324);
and I_23021 (I393725,I393375,I393708);
DFFARX1 I_23022  ( .D(I393725), .CLK(I2350), .RSTB(I393211), .Q(I393179) );
not I_23023 (I393789,I2357);
nand I_23024 (I393806,I270309,I270327);
and I_23025 (I393823,I393806,I270303);
DFFARX1 I_23026  ( .D(I393823), .CLK(I2350), .RSTB(I393789), .Q(I393840) );
not I_23027 (I393778,I393840);
DFFARX1 I_23028  ( .D(I393840), .CLK(I2350), .RSTB(I393789), .Q(I393871) );
not I_23029 (I393766,I393871);
nor I_23030 (I393902,I270315,I270327);
not I_23031 (I393919,I393902);
nor I_23032 (I393936,I393840,I393919);
DFFARX1 I_23033  ( .D(I270306), .CLK(I2350), .RSTB(I393789), .Q(I393953) );
not I_23034 (I393970,I393953);
nand I_23035 (I393769,I393953,I393919);
DFFARX1 I_23036  ( .D(I393953), .CLK(I2350), .RSTB(I393789), .Q(I394001) );
and I_23037 (I393754,I393840,I394001);
nand I_23038 (I394032,I270321,I270300);
and I_23039 (I394049,I394032,I270318);
DFFARX1 I_23040  ( .D(I394049), .CLK(I2350), .RSTB(I393789), .Q(I394066) );
nor I_23041 (I394083,I394066,I393970);
and I_23042 (I394100,I393902,I394083);
nor I_23043 (I394117,I394066,I393840);
DFFARX1 I_23044  ( .D(I394066), .CLK(I2350), .RSTB(I393789), .Q(I393760) );
DFFARX1 I_23045  ( .D(I270324), .CLK(I2350), .RSTB(I393789), .Q(I394148) );
and I_23046 (I394165,I394148,I270312);
or I_23047 (I394182,I394165,I394100);
DFFARX1 I_23048  ( .D(I394182), .CLK(I2350), .RSTB(I393789), .Q(I393772) );
nand I_23049 (I393781,I394165,I394117);
DFFARX1 I_23050  ( .D(I394165), .CLK(I2350), .RSTB(I393789), .Q(I393751) );
DFFARX1 I_23051  ( .D(I270297), .CLK(I2350), .RSTB(I393789), .Q(I394241) );
nand I_23052 (I393775,I394241,I393936);
DFFARX1 I_23053  ( .D(I394241), .CLK(I2350), .RSTB(I393789), .Q(I393763) );
nand I_23054 (I394286,I394241,I393902);
and I_23055 (I394303,I393953,I394286);
DFFARX1 I_23056  ( .D(I394303), .CLK(I2350), .RSTB(I393789), .Q(I393757) );
not I_23057 (I394367,I2357);
nand I_23058 (I394384,I206939,I206942);
and I_23059 (I394401,I394384,I206921);
DFFARX1 I_23060  ( .D(I394401), .CLK(I2350), .RSTB(I394367), .Q(I394418) );
not I_23061 (I394356,I394418);
DFFARX1 I_23062  ( .D(I394418), .CLK(I2350), .RSTB(I394367), .Q(I394449) );
not I_23063 (I394344,I394449);
nor I_23064 (I394480,I206936,I206942);
not I_23065 (I394497,I394480);
nor I_23066 (I394514,I394418,I394497);
DFFARX1 I_23067  ( .D(I206945), .CLK(I2350), .RSTB(I394367), .Q(I394531) );
not I_23068 (I394548,I394531);
nand I_23069 (I394347,I394531,I394497);
DFFARX1 I_23070  ( .D(I394531), .CLK(I2350), .RSTB(I394367), .Q(I394579) );
and I_23071 (I394332,I394418,I394579);
nand I_23072 (I394610,I206933,I206951);
and I_23073 (I394627,I394610,I206927);
DFFARX1 I_23074  ( .D(I394627), .CLK(I2350), .RSTB(I394367), .Q(I394644) );
nor I_23075 (I394661,I394644,I394548);
and I_23076 (I394678,I394480,I394661);
nor I_23077 (I394695,I394644,I394418);
DFFARX1 I_23078  ( .D(I394644), .CLK(I2350), .RSTB(I394367), .Q(I394338) );
DFFARX1 I_23079  ( .D(I206924), .CLK(I2350), .RSTB(I394367), .Q(I394726) );
and I_23080 (I394743,I394726,I206930);
or I_23081 (I394760,I394743,I394678);
DFFARX1 I_23082  ( .D(I394760), .CLK(I2350), .RSTB(I394367), .Q(I394350) );
nand I_23083 (I394359,I394743,I394695);
DFFARX1 I_23084  ( .D(I394743), .CLK(I2350), .RSTB(I394367), .Q(I394329) );
DFFARX1 I_23085  ( .D(I206948), .CLK(I2350), .RSTB(I394367), .Q(I394819) );
nand I_23086 (I394353,I394819,I394514);
DFFARX1 I_23087  ( .D(I394819), .CLK(I2350), .RSTB(I394367), .Q(I394341) );
nand I_23088 (I394864,I394819,I394480);
and I_23089 (I394881,I394531,I394864);
DFFARX1 I_23090  ( .D(I394881), .CLK(I2350), .RSTB(I394367), .Q(I394335) );
not I_23091 (I394945,I2357);
nand I_23092 (I394962,I168850,I168847);
and I_23093 (I394979,I394962,I168871);
DFFARX1 I_23094  ( .D(I394979), .CLK(I2350), .RSTB(I394945), .Q(I394996) );
not I_23095 (I394934,I394996);
DFFARX1 I_23096  ( .D(I394996), .CLK(I2350), .RSTB(I394945), .Q(I395027) );
not I_23097 (I394922,I395027);
nor I_23098 (I395058,I168853,I168847);
not I_23099 (I395075,I395058);
nor I_23100 (I395092,I394996,I395075);
DFFARX1 I_23101  ( .D(I168868), .CLK(I2350), .RSTB(I394945), .Q(I395109) );
not I_23102 (I395126,I395109);
nand I_23103 (I394925,I395109,I395075);
DFFARX1 I_23104  ( .D(I395109), .CLK(I2350), .RSTB(I394945), .Q(I395157) );
and I_23105 (I394910,I394996,I395157);
nand I_23106 (I395188,I168856,I168841);
and I_23107 (I395205,I395188,I168859);
DFFARX1 I_23108  ( .D(I395205), .CLK(I2350), .RSTB(I394945), .Q(I395222) );
nor I_23109 (I395239,I395222,I395126);
and I_23110 (I395256,I395058,I395239);
nor I_23111 (I395273,I395222,I394996);
DFFARX1 I_23112  ( .D(I395222), .CLK(I2350), .RSTB(I394945), .Q(I394916) );
DFFARX1 I_23113  ( .D(I168862), .CLK(I2350), .RSTB(I394945), .Q(I395304) );
and I_23114 (I395321,I395304,I168865);
or I_23115 (I395338,I395321,I395256);
DFFARX1 I_23116  ( .D(I395338), .CLK(I2350), .RSTB(I394945), .Q(I394928) );
nand I_23117 (I394937,I395321,I395273);
DFFARX1 I_23118  ( .D(I395321), .CLK(I2350), .RSTB(I394945), .Q(I394907) );
DFFARX1 I_23119  ( .D(I168844), .CLK(I2350), .RSTB(I394945), .Q(I395397) );
nand I_23120 (I394931,I395397,I395092);
DFFARX1 I_23121  ( .D(I395397), .CLK(I2350), .RSTB(I394945), .Q(I394919) );
nand I_23122 (I395442,I395397,I395058);
and I_23123 (I395459,I395109,I395442);
DFFARX1 I_23124  ( .D(I395459), .CLK(I2350), .RSTB(I394945), .Q(I394913) );
not I_23125 (I395523,I2357);
nand I_23126 (I395540,I153601,I153598);
and I_23127 (I395557,I395540,I153622);
DFFARX1 I_23128  ( .D(I395557), .CLK(I2350), .RSTB(I395523), .Q(I395574) );
not I_23129 (I395512,I395574);
DFFARX1 I_23130  ( .D(I395574), .CLK(I2350), .RSTB(I395523), .Q(I395605) );
not I_23131 (I395500,I395605);
nor I_23132 (I395636,I153604,I153598);
not I_23133 (I395653,I395636);
nor I_23134 (I395670,I395574,I395653);
DFFARX1 I_23135  ( .D(I153619), .CLK(I2350), .RSTB(I395523), .Q(I395687) );
not I_23136 (I395704,I395687);
nand I_23137 (I395503,I395687,I395653);
DFFARX1 I_23138  ( .D(I395687), .CLK(I2350), .RSTB(I395523), .Q(I395735) );
and I_23139 (I395488,I395574,I395735);
nand I_23140 (I395766,I153607,I153592);
and I_23141 (I395783,I395766,I153610);
DFFARX1 I_23142  ( .D(I395783), .CLK(I2350), .RSTB(I395523), .Q(I395800) );
nor I_23143 (I395817,I395800,I395704);
and I_23144 (I395834,I395636,I395817);
nor I_23145 (I395851,I395800,I395574);
DFFARX1 I_23146  ( .D(I395800), .CLK(I2350), .RSTB(I395523), .Q(I395494) );
DFFARX1 I_23147  ( .D(I153613), .CLK(I2350), .RSTB(I395523), .Q(I395882) );
and I_23148 (I395899,I395882,I153616);
or I_23149 (I395916,I395899,I395834);
DFFARX1 I_23150  ( .D(I395916), .CLK(I2350), .RSTB(I395523), .Q(I395506) );
nand I_23151 (I395515,I395899,I395851);
DFFARX1 I_23152  ( .D(I395899), .CLK(I2350), .RSTB(I395523), .Q(I395485) );
DFFARX1 I_23153  ( .D(I153595), .CLK(I2350), .RSTB(I395523), .Q(I395975) );
nand I_23154 (I395509,I395975,I395670);
DFFARX1 I_23155  ( .D(I395975), .CLK(I2350), .RSTB(I395523), .Q(I395497) );
nand I_23156 (I396020,I395975,I395636);
and I_23157 (I396037,I395687,I396020);
DFFARX1 I_23158  ( .D(I396037), .CLK(I2350), .RSTB(I395523), .Q(I395491) );
not I_23159 (I396101,I2357);
nand I_23160 (I396118,I7433,I7418);
and I_23161 (I396135,I396118,I7427);
DFFARX1 I_23162  ( .D(I396135), .CLK(I2350), .RSTB(I396101), .Q(I396152) );
not I_23163 (I396090,I396152);
DFFARX1 I_23164  ( .D(I396152), .CLK(I2350), .RSTB(I396101), .Q(I396183) );
not I_23165 (I396078,I396183);
nor I_23166 (I396214,I7439,I7418);
not I_23167 (I396231,I396214);
nor I_23168 (I396248,I396152,I396231);
DFFARX1 I_23169  ( .D(I7430), .CLK(I2350), .RSTB(I396101), .Q(I396265) );
not I_23170 (I396282,I396265);
nand I_23171 (I396081,I396265,I396231);
DFFARX1 I_23172  ( .D(I396265), .CLK(I2350), .RSTB(I396101), .Q(I396313) );
and I_23173 (I396066,I396152,I396313);
nand I_23174 (I396344,I7415,I7409);
and I_23175 (I396361,I396344,I7424);
DFFARX1 I_23176  ( .D(I396361), .CLK(I2350), .RSTB(I396101), .Q(I396378) );
nor I_23177 (I396395,I396378,I396282);
and I_23178 (I396412,I396214,I396395);
nor I_23179 (I396429,I396378,I396152);
DFFARX1 I_23180  ( .D(I396378), .CLK(I2350), .RSTB(I396101), .Q(I396072) );
DFFARX1 I_23181  ( .D(I7412), .CLK(I2350), .RSTB(I396101), .Q(I396460) );
and I_23182 (I396477,I396460,I7436);
or I_23183 (I396494,I396477,I396412);
DFFARX1 I_23184  ( .D(I396494), .CLK(I2350), .RSTB(I396101), .Q(I396084) );
nand I_23185 (I396093,I396477,I396429);
DFFARX1 I_23186  ( .D(I396477), .CLK(I2350), .RSTB(I396101), .Q(I396063) );
DFFARX1 I_23187  ( .D(I7421), .CLK(I2350), .RSTB(I396101), .Q(I396553) );
nand I_23188 (I396087,I396553,I396248);
DFFARX1 I_23189  ( .D(I396553), .CLK(I2350), .RSTB(I396101), .Q(I396075) );
nand I_23190 (I396598,I396553,I396214);
and I_23191 (I396615,I396265,I396598);
DFFARX1 I_23192  ( .D(I396615), .CLK(I2350), .RSTB(I396101), .Q(I396069) );
not I_23193 (I396679,I2357);
nand I_23194 (I396696,I246398,I246416);
and I_23195 (I396713,I396696,I246407);
DFFARX1 I_23196  ( .D(I396713), .CLK(I2350), .RSTB(I396679), .Q(I396730) );
not I_23197 (I396668,I396730);
DFFARX1 I_23198  ( .D(I396730), .CLK(I2350), .RSTB(I396679), .Q(I396761) );
not I_23199 (I396656,I396761);
nor I_23200 (I396792,I246404,I246416);
not I_23201 (I396809,I396792);
nor I_23202 (I396826,I396730,I396809);
DFFARX1 I_23203  ( .D(I246395), .CLK(I2350), .RSTB(I396679), .Q(I396843) );
not I_23204 (I396860,I396843);
nand I_23205 (I396659,I396843,I396809);
DFFARX1 I_23206  ( .D(I396843), .CLK(I2350), .RSTB(I396679), .Q(I396891) );
and I_23207 (I396644,I396730,I396891);
nand I_23208 (I396922,I246413,I246425);
and I_23209 (I396939,I396922,I246419);
DFFARX1 I_23210  ( .D(I396939), .CLK(I2350), .RSTB(I396679), .Q(I396956) );
nor I_23211 (I396973,I396956,I396860);
and I_23212 (I396990,I396792,I396973);
nor I_23213 (I397007,I396956,I396730);
DFFARX1 I_23214  ( .D(I396956), .CLK(I2350), .RSTB(I396679), .Q(I396650) );
DFFARX1 I_23215  ( .D(I246401), .CLK(I2350), .RSTB(I396679), .Q(I397038) );
and I_23216 (I397055,I397038,I246410);
or I_23217 (I397072,I397055,I396990);
DFFARX1 I_23218  ( .D(I397072), .CLK(I2350), .RSTB(I396679), .Q(I396662) );
nand I_23219 (I396671,I397055,I397007);
DFFARX1 I_23220  ( .D(I397055), .CLK(I2350), .RSTB(I396679), .Q(I396641) );
DFFARX1 I_23221  ( .D(I246422), .CLK(I2350), .RSTB(I396679), .Q(I397131) );
nand I_23222 (I396665,I397131,I396826);
DFFARX1 I_23223  ( .D(I397131), .CLK(I2350), .RSTB(I396679), .Q(I396653) );
nand I_23224 (I397176,I397131,I396792);
and I_23225 (I397193,I396843,I397176);
DFFARX1 I_23226  ( .D(I397193), .CLK(I2350), .RSTB(I396679), .Q(I396647) );
not I_23227 (I397257,I2357);
nand I_23228 (I397274,I80853,I80838);
and I_23229 (I397291,I397274,I80832);
DFFARX1 I_23230  ( .D(I397291), .CLK(I2350), .RSTB(I397257), .Q(I397308) );
not I_23231 (I397246,I397308);
DFFARX1 I_23232  ( .D(I397308), .CLK(I2350), .RSTB(I397257), .Q(I397339) );
not I_23233 (I397234,I397339);
nor I_23234 (I397370,I80859,I80838);
not I_23235 (I397387,I397370);
nor I_23236 (I397404,I397308,I397387);
DFFARX1 I_23237  ( .D(I80862), .CLK(I2350), .RSTB(I397257), .Q(I397421) );
not I_23238 (I397438,I397421);
nand I_23239 (I397237,I397421,I397387);
DFFARX1 I_23240  ( .D(I397421), .CLK(I2350), .RSTB(I397257), .Q(I397469) );
and I_23241 (I397222,I397308,I397469);
nand I_23242 (I397500,I80844,I80847);
and I_23243 (I397517,I397500,I80850);
DFFARX1 I_23244  ( .D(I397517), .CLK(I2350), .RSTB(I397257), .Q(I397534) );
nor I_23245 (I397551,I397534,I397438);
and I_23246 (I397568,I397370,I397551);
nor I_23247 (I397585,I397534,I397308);
DFFARX1 I_23248  ( .D(I397534), .CLK(I2350), .RSTB(I397257), .Q(I397228) );
DFFARX1 I_23249  ( .D(I80856), .CLK(I2350), .RSTB(I397257), .Q(I397616) );
and I_23250 (I397633,I397616,I80841);
or I_23251 (I397650,I397633,I397568);
DFFARX1 I_23252  ( .D(I397650), .CLK(I2350), .RSTB(I397257), .Q(I397240) );
nand I_23253 (I397249,I397633,I397585);
DFFARX1 I_23254  ( .D(I397633), .CLK(I2350), .RSTB(I397257), .Q(I397219) );
DFFARX1 I_23255  ( .D(I80835), .CLK(I2350), .RSTB(I397257), .Q(I397709) );
nand I_23256 (I397243,I397709,I397404);
DFFARX1 I_23257  ( .D(I397709), .CLK(I2350), .RSTB(I397257), .Q(I397231) );
nand I_23258 (I397754,I397709,I397370);
and I_23259 (I397771,I397421,I397754);
DFFARX1 I_23260  ( .D(I397771), .CLK(I2350), .RSTB(I397257), .Q(I397225) );
endmodule


