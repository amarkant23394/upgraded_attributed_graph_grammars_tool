module test_final(IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_4_2_l_6,IN_5_2_l_6,IN_1_6_l_6,IN_2_6_l_6,IN_3_6_l_6,IN_4_6_l_6,IN_5_6_l_6,IN_1_9_l_6,IN_2_9_l_6,IN_3_9_l_6,IN_4_9_l_6,IN_5_9_l_6,blif_clk_net_5_r_13,blif_reset_net_5_r_13,N1371_0_r_13,N1508_0_r_13,n_429_or_0_5_r_13,G78_5_r_13,n_576_5_r_13,n_547_5_r_13,G42_7_r_13,n_572_7_r_13,n_573_7_r_13,n_549_7_r_13,n_569_7_r_13,n_452_7_r_13);
input IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_4_2_l_6,IN_5_2_l_6,IN_1_6_l_6,IN_2_6_l_6,IN_3_6_l_6,IN_4_6_l_6,IN_5_6_l_6,IN_1_9_l_6,IN_2_9_l_6,IN_3_9_l_6,IN_4_9_l_6,IN_5_9_l_6,blif_clk_net_5_r_13,blif_reset_net_5_r_13;
output N1371_0_r_13,N1508_0_r_13,n_429_or_0_5_r_13,G78_5_r_13,n_576_5_r_13,n_547_5_r_13,G42_7_r_13,n_572_7_r_13,n_573_7_r_13,n_549_7_r_13,n_569_7_r_13,n_452_7_r_13;
wire N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,I_BUFF_1_9_r_6,N1372_10_r_6,N1508_10_r_6,N3_8_r_6,n30_6,n31_6,n32_6,n33_6,n34_6,n35_6,n36_6,n37_6,n38_6,n39_6,n40_6,n41_6,n42_6,n43_6,n44_6,n45_6,n46_6,n47_6,n48_6,n49_6,n50_6,n51_6,n52_6,n53_6,n54_6,n_102_5_r_13,n4_7_l_13,n9_13,n62_13,n33_13,n_431_5_r_13,n1_13,n34_13,n35_13,n36_13,n37_13,n38_13,n39_13,n40_13,n41_13,n42_13,n43_13,n44_13,n45_13,n46_13,n47_13,n48_13,n49_13,n50_13,n51_13,n52_13,n53_13,n54_13,n55_13,n56_13,n57_13,n58_13,n59_13,n60_13,n61_13;
nor I_0(N1371_0_r_6,n30_6,n33_6);
nor I_1(N1508_0_r_6,n33_6,n44_6);
not I_2(N1372_1_r_6,n41_6);
nor I_3(N1508_1_r_6,n40_6,n41_6);
nor I_4(N1507_6_r_6,n39_6,n45_6);
nor I_5(N1508_6_r_6,n37_6,n38_6);
nor I_6(n_42_8_r_6,n30_6,n31_6);
DFFARX1 I_7(N3_8_r_6,blif_clk_net_5_r_13,n9_13,G199_8_r_6,);
nor I_8(N6147_9_r_6,n32_6,n33_6);
nor I_9(N6134_9_r_6,I_BUFF_1_9_r_6,n35_6);
not I_10(I_BUFF_1_9_r_6,n37_6);
not I_11(N1372_10_r_6,n43_6);
nor I_12(N1508_10_r_6,n42_6,n43_6);
nor I_13(N3_8_r_6,IN_1_9_l_6,n36_6);
nor I_14(n30_6,IN_5_9_l_6,n53_6);
not I_15(n31_6,n36_6);
nor I_16(n32_6,I_BUFF_1_9_r_6,n34_6);
not I_17(n33_6,IN_1_9_l_6);
not I_18(n34_6,n35_6);
nand I_19(n35_6,IN_2_6_l_6,n49_6);
nand I_20(n36_6,IN_5_6_l_6,n51_6);
nand I_21(n37_6,IN_2_9_l_6,n54_6);
or I_22(n38_6,n35_6,n39_6);
nor I_23(n39_6,n40_6,n45_6);
and I_24(n40_6,n46_6,n47_6);
nand I_25(n41_6,n30_6,n31_6);
nor I_26(n42_6,n34_6,n40_6);
nand I_27(n43_6,IN_1_9_l_6,n30_6);
nor I_28(n44_6,n31_6,n40_6);
nor I_29(n45_6,n35_6,n36_6);
nor I_30(n46_6,IN_1_2_l_6,IN_2_2_l_6);
or I_31(n47_6,IN_5_2_l_6,n48_6);
nor I_32(n48_6,IN_3_2_l_6,IN_4_2_l_6);
and I_33(n49_6,IN_1_6_l_6,n50_6);
nand I_34(n50_6,n51_6,n52_6);
nand I_35(n51_6,IN_3_6_l_6,IN_4_6_l_6);
not I_36(n52_6,IN_5_6_l_6);
nor I_37(n53_6,IN_3_9_l_6,IN_4_9_l_6);
or I_38(n54_6,IN_3_9_l_6,IN_4_9_l_6);
nor I_39(N1371_0_r_13,n59_13,n61_13);
nor I_40(N1508_0_r_13,n59_13,n60_13);
not I_41(n_429_or_0_5_r_13,n46_13);
DFFARX1 I_42(n_431_5_r_13,blif_clk_net_5_r_13,n9_13,G78_5_r_13,);
nand I_43(n_576_5_r_13,n_102_5_r_13,n34_13);
nor I_44(n_102_5_r_13,N1508_1_r_6,N6134_9_r_6);
nand I_45(n_547_5_r_13,n48_13,n49_13);
DFFARX1 I_46(n1_13,blif_clk_net_5_r_13,n9_13,G42_7_r_13,);
nor I_47(n_572_7_r_13,n40_13,n41_13);
nand I_48(n_573_7_r_13,n37_13,n38_13);
nor I_49(n_549_7_r_13,n46_13,n47_13);
nand I_50(n_569_7_r_13,n37_13,n43_13);
nand I_51(n_452_7_r_13,n52_13,n53_13);
nor I_52(n4_7_l_13,N1508_10_r_6,N1508_0_r_6);
not I_53(n9_13,blif_reset_net_5_r_13);
DFFARX1 I_54(n4_7_l_13,blif_clk_net_5_r_13,n9_13,n62_13,);
not I_55(n33_13,n62_13);
nand I_56(n_431_5_r_13,n54_13,n55_13);
not I_57(n1_13,n52_13);
nor I_58(n34_13,n35_13,n36_13);
nor I_59(n35_13,n42_13,N1371_0_r_6);
nand I_60(n36_13,n50_13,n58_13);
nand I_61(n37_13,n44_13,n45_13);
or I_62(n38_13,n39_13,N1372_1_r_6);
nand I_63(n39_13,N1508_6_r_6,G199_8_r_6);
not I_64(n40_13,n36_13);
nor I_65(n41_13,n35_13,N1508_1_r_6);
not I_66(n42_13,N1372_10_r_6);
or I_67(n43_13,N1508_10_r_6,N1372_1_r_6);
not I_68(n44_13,N1371_0_r_6);
not I_69(n45_13,N6147_9_r_6);
nor I_70(n46_13,n39_13,n40_13);
nor I_71(n47_13,N1508_10_r_6,N1372_1_r_6);
nor I_72(n48_13,n50_13,n51_13);
nor I_73(n49_13,N1371_0_r_6,N6147_9_r_6);
not I_74(n50_13,n59_13);
not I_75(n51_13,n_102_5_r_13);
nand I_76(n52_13,n33_13,n39_13);
nand I_77(n53_13,n33_13,N1372_1_r_6);
nor I_78(n54_13,N6134_9_r_6,N1372_1_r_6);
nand I_79(n55_13,n62_13,n56_13);
nor I_80(n56_13,n39_13,n57_13);
not I_81(n57_13,N1508_10_r_6);
or I_82(n58_13,N1507_6_r_6,n_42_8_r_6);
nand I_83(n59_13,N1508_0_r_6,N1371_0_r_6);
nor I_84(n60_13,n51_13,N1372_1_r_6);
nor I_85(n61_13,n39_13,N1372_1_r_6);
endmodule


