module test_final(IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_4_2_l_6,IN_5_2_l_6,IN_1_6_l_6,IN_2_6_l_6,IN_3_6_l_6,IN_4_6_l_6,IN_5_6_l_6,IN_1_9_l_6,IN_2_9_l_6,IN_3_9_l_6,IN_4_9_l_6,IN_5_9_l_6,blif_clk_net_5_r_15,blif_reset_net_5_r_15,N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15);
input IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_4_2_l_6,IN_5_2_l_6,IN_1_6_l_6,IN_2_6_l_6,IN_3_6_l_6,IN_4_6_l_6,IN_5_6_l_6,IN_1_9_l_6,IN_2_9_l_6,IN_3_9_l_6,IN_4_9_l_6,IN_5_9_l_6,blif_clk_net_5_r_15,blif_reset_net_5_r_15;
output N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15;
wire N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,I_BUFF_1_9_r_6,N1372_10_r_6,N1508_10_r_6,N3_8_r_6,n30_6,n31_6,n32_6,n33_6,n34_6,n35_6,n36_6,n37_6,n38_6,n39_6,n40_6,n41_6,n42_6,n43_6,n44_6,n45_6,n46_6,n47_6,n48_6,n49_6,n50_6,n51_6,n52_6,n53_6,n54_6,N1371_0_r_15,N1508_0_r_15,N1372_1_r_15,n_102_5_r_15,n_431_5_r_15,n9_15,n31_15,n32_15,n33_15,n34_15,n35_15,n36_15,n37_15,n38_15,n39_15,n40_15,n41_15,n42_15,n43_15,n44_15,n45_15,n46_15,n47_15,n48_15,n49_15,n50_15,n51_15,n52_15,n53_15,n54_15,n55_15;
nor I_0(N1371_0_r_6,n30_6,n33_6);
nor I_1(N1508_0_r_6,n33_6,n44_6);
not I_2(N1372_1_r_6,n41_6);
nor I_3(N1508_1_r_6,n40_6,n41_6);
nor I_4(N1507_6_r_6,n39_6,n45_6);
nor I_5(N1508_6_r_6,n37_6,n38_6);
nor I_6(n_42_8_r_6,n30_6,n31_6);
DFFARX1 I_7(N3_8_r_6,blif_clk_net_5_r_15,n9_15,G199_8_r_6,);
nor I_8(N6147_9_r_6,n32_6,n33_6);
nor I_9(N6134_9_r_6,I_BUFF_1_9_r_6,n35_6);
not I_10(I_BUFF_1_9_r_6,n37_6);
not I_11(N1372_10_r_6,n43_6);
nor I_12(N1508_10_r_6,n42_6,n43_6);
nor I_13(N3_8_r_6,IN_1_9_l_6,n36_6);
nor I_14(n30_6,IN_5_9_l_6,n53_6);
not I_15(n31_6,n36_6);
nor I_16(n32_6,I_BUFF_1_9_r_6,n34_6);
not I_17(n33_6,IN_1_9_l_6);
not I_18(n34_6,n35_6);
nand I_19(n35_6,IN_2_6_l_6,n49_6);
nand I_20(n36_6,IN_5_6_l_6,n51_6);
nand I_21(n37_6,IN_2_9_l_6,n54_6);
or I_22(n38_6,n35_6,n39_6);
nor I_23(n39_6,n40_6,n45_6);
and I_24(n40_6,n46_6,n47_6);
nand I_25(n41_6,n30_6,n31_6);
nor I_26(n42_6,n34_6,n40_6);
nand I_27(n43_6,IN_1_9_l_6,n30_6);
nor I_28(n44_6,n31_6,n40_6);
nor I_29(n45_6,n35_6,n36_6);
nor I_30(n46_6,IN_1_2_l_6,IN_2_2_l_6);
or I_31(n47_6,IN_5_2_l_6,n48_6);
nor I_32(n48_6,IN_3_2_l_6,IN_4_2_l_6);
and I_33(n49_6,IN_1_6_l_6,n50_6);
nand I_34(n50_6,n51_6,n52_6);
nand I_35(n51_6,IN_3_6_l_6,IN_4_6_l_6);
not I_36(n52_6,IN_5_6_l_6);
nor I_37(n53_6,IN_3_9_l_6,IN_4_9_l_6);
or I_38(n54_6,IN_3_9_l_6,IN_4_9_l_6);
and I_39(N1371_0_r_15,N1508_0_r_15,n_102_5_r_15);
nor I_40(N1508_0_r_15,n55_15,N1371_0_r_6);
nor I_41(N1372_1_r_15,n_102_5_r_15,n46_15);
nor I_42(N1508_1_r_15,N1508_0_r_15,n45_15);
not I_43(N1372_4_r_15,n39_15);
nor I_44(N1508_4_r_15,n39_15,n43_15);
nand I_45(n_429_or_0_5_r_15,n36_15,n38_15);
DFFARX1 I_46(n_431_5_r_15,blif_clk_net_5_r_15,n9_15,G78_5_r_15,);
nand I_47(n_576_5_r_15,n31_15,n32_15);
not I_48(n_102_5_r_15,n33_15);
nand I_49(n_547_5_r_15,N1371_0_r_15,n35_15);
nor I_50(N1507_6_r_15,n42_15,n46_15);
nand I_51(N1508_6_r_15,n39_15,n40_15);
nand I_52(n_431_5_r_15,n36_15,n37_15);
not I_53(n9_15,blif_reset_net_5_r_15);
nor I_54(n31_15,n33_15,n34_15);
nor I_55(n32_15,n44_15,N1508_1_r_6);
nor I_56(n33_15,n54_15,n55_15);
nand I_57(n34_15,n49_15,N1508_0_r_6);
nand I_58(n35_15,N1508_6_r_6,N1371_0_r_6);
not I_59(n36_15,n32_15);
nand I_60(n37_15,n34_15,n38_15);
not I_61(n38_15,n46_15);
nand I_62(n39_15,n38_15,n41_15);
nand I_63(n40_15,n41_15,n42_15);
and I_64(n41_15,n51_15,N1508_10_r_6);
and I_65(n42_15,n47_15,N1508_6_r_6);
and I_66(n43_15,n34_15,n36_15);
or I_67(n44_15,n_42_8_r_6,N6134_9_r_6);
not I_68(n45_15,N1372_1_r_15);
nand I_69(n46_15,n53_15,N1508_6_r_6);
nor I_70(n47_15,n34_15,n48_15);
not I_71(n48_15,N1371_0_r_6);
and I_72(n49_15,n50_15,N1372_1_r_6);
nand I_73(n50_15,n51_15,n52_15);
nand I_74(n51_15,N1508_0_r_6,N1507_6_r_6);
not I_75(n52_15,N1508_10_r_6);
nor I_76(n53_15,n48_15,N1372_1_r_6);
nor I_77(n54_15,G199_8_r_6,N1372_10_r_6);
not I_78(n55_15,N6147_9_r_6);
endmodule


