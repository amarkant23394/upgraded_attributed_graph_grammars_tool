module test_I5802(I4629,I1477,I4824,I4886,I1470,I4725,I4578,I5802);
input I4629,I1477,I4824,I4886,I1470,I4725,I4578;
output I5802;
wire I5751,I4515,I4595,I4524,I4544,I5785,I4742,I5768,I4530;
not I_0(I5751,I1477);
not I_1(I4515,I4629);
DFFARX1 I_2(I4578,I1470,I4544,,,I4595,);
nor I_3(I4524,I4742,I4595);
not I_4(I4544,I1477);
and I_5(I5785,I5768,I4524);
DFFARX1 I_6(I4725,I1470,I4544,,,I4742,);
DFFARX1 I_7(I5785,I1470,I5751,,,I5802,);
nand I_8(I5768,I4530,I4515);
nor I_9(I4530,I4824,I4886);
endmodule


