module test_I6459(I2742,I4017,I2727,I1470,I3983,I6459);
input I2742,I4017,I2727,I1470,I3983;
output I6459;
wire I3975,I3954,I6442,I4308,I4068,I4034,I2724;
nor I_0(I3975,I4308,I4034);
not I_1(I3954,I4068);
nor I_2(I6442,I3975,I3954);
DFFARX1 I_3(I2727,I1470,I3983,,,I4308,);
nor I_4(I4068,I2742,I2724);
DFFARX1 I_5(I4017,I1470,I3983,,,I4034,);
not I_6(I6459,I6442);
DFFARX1 I_7(I1470,,,I2724,);
endmodule


