module test_I2181_rst(I1477_rst,I2181_rst);
,I2181_rst);
input I1477_rst;
output I2181_rst;
wire ;
not I_0(I2181_rst,I1477_rst);
endmodule


