module test_I1914(I1322,I2087,I1294,I1331,I2406,I1301,I1914);
input I1322,I2087,I1294,I1331,I2406,I1301;
output I1914;
wire I2440,I2313,I1937,I1342,I2234,I2423,I2457,I1509,I1304,I1954;
and I_0(I2440,I2313,I2423);
DFFARX1 I_1(I2457,I1294,I1937,,,I1914,);
DFFARX1 I_2(I1331,I1294,I1937,,,I2313,);
not I_3(I1937,I1301);
not I_4(I1342,I1301);
nand I_5(I2234,I1954,I1304);
nor I_6(I2423,I2406,I2087);
or I_7(I2457,I2234,I2440);
DFFARX1 I_8(I1294,I1342,,,I1509,);
DFFARX1 I_9(I1509,I1294,I1342,,,I1304,);
not I_10(I1954,I1322);
endmodule


