module test_I15928(I11956,I1477,I1470,I15928);
input I11956,I1477,I1470;
output I15928;
wire I14083,I13746,I14066,I13775,I15611,I14049;
DFFARX1 I_0(I14066,I1470,I13775,,,I14083,);
not I_1(I13746,I14083);
and I_2(I14066,I14049,I11956);
not I_3(I13775,I1477);
not I_4(I15611,I1477);
DFFARX1 I_5(I1470,I13775,,,I14049,);
DFFARX1 I_6(I13746,I1470,I15611,,,I15928,);
endmodule


