module test_I10086(I1477,I6294,I6476,I7881,I6318,I1470,I10086);
input I1477,I6294,I6476,I7881,I6318,I1470;
output I10086;
wire I6781,I6315,I6297,I7621,I7652,I7669,I7714,I7946,I7535,I10069,I7570,I7559,I7604,I7544;
DFFARX1 I_0(I1470,,,I6781,);
nand I_1(I6315,I6781,I6476);
DFFARX1 I_2(I1470,,,I6297,);
nand I_3(I7621,I7604,I6315);
nor I_4(I7652,I6297);
nand I_5(I7669,I7652,I6318);
not I_6(I7714,I6297);
DFFARX1 I_7(I7881,I1470,I7570,,,I7946,);
and I_8(I7535,I7714,I7946);
nand I_9(I10069,I7559,I7535);
and I_10(I10086,I10069,I7544);
not I_11(I7570,I1477);
not I_12(I7559,I7669);
nor I_13(I7604,I6297,I6294);
DFFARX1 I_14(I7621,I1470,I7570,,,I7544,);
endmodule


