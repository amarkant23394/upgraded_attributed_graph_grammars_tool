module test_I5067(I1477,I1470,I5067);
input I1477,I1470;
output I5067;
wire I5625,I3377,I3747,I5105,I5642;
DFFARX1 I_0(I3377,I1470,I5105,,,I5625,);
DFFARX1 I_1(I5642,I1470,I5105,,,I5067,);
not I_2(I3377,I3747);
DFFARX1 I_3(I1470,,,I3747,);
not I_4(I5105,I1477);
not I_5(I5642,I5625);
endmodule


