module test_I11813(I6992,I1477,I7026,I1470,I11813);
input I6992,I1477,I7026,I1470;
output I11813;
wire I9320,I6875,I8854,I9303,I9179,I8862,I11310,I6896;
not I_0(I9320,I9303);
DFFARX1 I_1(I1470,,,I6875,);
nor I_2(I8854,I9179,I9320);
DFFARX1 I_3(I8854,I1470,I11310,,,I11813,);
DFFARX1 I_4(I6875,I1470,I8862,,,I9303,);
DFFARX1 I_5(I6896,I1470,I8862,,,I9179,);
not I_6(I8862,I1477);
not I_7(I11310,I1477);
nor I_8(I6896,I6992,I7026);
endmodule


