module test_I14344(I13697,I13180,I1477,I13168,I1470,I13635,I14344);
input I13697,I13180,I1477,I13168,I1470,I13635;
output I14344;
wire I14667,I13189,I13197,I14503,I14520,I13174,I14370,I14650,I13165,I14537,I14715;
and I_0(I14667,I14650,I13189);
DFFARX1 I_1(I13635,I1470,I13197,,,I13189,);
not I_2(I13197,I1477);
nand I_3(I14344,I14537,I14715);
nand I_4(I14503,I13180,I13168);
and I_5(I14520,I14503,I13174);
DFFARX1 I_6(I13697,I1470,I13197,,,I13174,);
not I_7(I14370,I1477);
DFFARX1 I_8(I13165,I1470,I14370,,,I14650,);
DFFARX1 I_9(I1470,I13197,,,I13165,);
DFFARX1 I_10(I14520,I1470,I14370,,,I14537,);
not I_11(I14715,I14667);
endmodule


