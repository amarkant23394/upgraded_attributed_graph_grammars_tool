module test_I15628(I1477,I1470,I15628);
input I1477,I1470;
output I15628;
wire I13743,I13891,I13775,I12075,I11944;
DFFARX1 I_0(I13891,I1470,I13775,,,I13743,);
not I_1(I15628,I13743);
DFFARX1 I_2(I11944,I1470,I13775,,,I13891,);
not I_3(I13775,I1477);
DFFARX1 I_4(I1470,,,I12075,);
not I_5(I11944,I12075);
endmodule


