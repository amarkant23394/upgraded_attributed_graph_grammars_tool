module test_I11460(I9396,I6881,I8879,I8947,I11460);
input I9396,I6881,I8879,I8947;
output I11460;
wire I11429,I8848,I9083,I9413;
not I_0(I11429,I8848);
not I_1(I11460,I11429);
nor I_2(I8848,I9083,I9413);
nand I_3(I9083,I8879,I6881);
and I_4(I9413,I8947,I9396);
endmodule


