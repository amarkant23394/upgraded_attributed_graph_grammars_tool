module test_I3464(I2668,I2733,I2600,I3103,I1923,I1294,I2566,I1301,I3464);
input I2668,I2733,I2600,I3103,I1923,I1294,I2566,I1301;
output I3464;
wire I3120,I3137,I2897,I2551,I2575,I2583,I2557,I3413,I3430,I3447;
or I_0(I3464,I3447,I2575);
nand I_1(I3120,I3103,I2668);
and I_2(I3137,I2897,I3120);
nand I_3(I2897,I2600,I1923);
DFFARX1 I_4(I2897,I1294,I2583,,,I2551,);
DFFARX1 I_5(I3137,I1294,I2583,,,I2575,);
not I_6(I2583,I1301);
nand I_7(I2557,I2668,I2733);
not I_8(I3413,I2566);
nor I_9(I3430,I3413,I2557);
and I_10(I3447,I3430,I2551);
endmodule


