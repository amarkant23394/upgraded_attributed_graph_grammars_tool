module test_I3422(I1383,I1477,I1215,I1470,I1569,I3422);
input I1383,I1477,I1215,I1470,I1569;
output I3422;
wire I1518,I1637,I1480,I1976,I1880,I1483,I1959;
not I_0(I1518,I1477);
not I_1(I1637,I1215);
or I_2(I3422,I1483,I1480);
DFFARX1 I_3(I1976,I1470,I1518,,,I1480,);
and I_4(I1976,I1637,I1959);
DFFARX1 I_5(I1383,I1470,I1518,,,I1880,);
DFFARX1 I_6(I1880,I1470,I1518,,,I1483,);
nand I_7(I1959,I1880,I1569);
endmodule


