module test_I5013(I1477,I1303,I1470,I4725,I5013);
input I1477,I1303,I1470,I4725;
output I5013;
wire I2167,I4629,I4979,I4996,I4544,I2328,I4869,I4962,I2633,I2540,I2143,I4807,I2173,I2181,I2170,I2557,I2232,I2509,I4742,I4824;
nand I_0(I2167,I2633,I2328);
nor I_1(I4629,I2167,I2173);
nor I_2(I4979,I4742,I4962);
and I_3(I4996,I4629,I4979);
not I_4(I4544,I1477);
nor I_5(I2328,I2232);
DFFARX1 I_6(I1470,I4544,,,I4869,);
not I_7(I4962,I4869);
DFFARX1 I_8(I1470,I2181,,,I2633,);
DFFARX1 I_9(I1470,I2181,,,I2540,);
DFFARX1 I_10(I2557,I1470,I2181,,,I2143,);
or I_11(I5013,I4824,I4996);
DFFARX1 I_12(I2170,I1470,I4544,,,I4807,);
nand I_13(I2173,I2557,I2509);
not I_14(I2181,I1477);
not I_15(I2170,I2232);
and I_16(I2557,I2540,I1303);
DFFARX1 I_17(I1470,I2181,,,I2232,);
nor I_18(I2509,I2232);
DFFARX1 I_19(I4725,I1470,I4544,,,I4742,);
and I_20(I4824,I4807,I2143);
endmodule


