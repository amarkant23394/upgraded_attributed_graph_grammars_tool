module test_I10120(I1477,I7587,I6843,I1470,I10120);
input I1477,I7587,I6843,I1470;
output I10120;
wire I7898,I6297,I7538,I7714,I7946,I7570,I7881,I7816,I6329,I7535,I7915,I6291;
nand I_0(I7898,I7881,I7816);
DFFARX1 I_1(I6843,I1470,I6329,,,I6297,);
DFFARX1 I_2(I7915,I1470,I7570,,,I7538,);
not I_3(I7714,I6297);
DFFARX1 I_4(I7881,I1470,I7570,,,I7946,);
not I_5(I7570,I1477);
nand I_6(I7881,I7587,I6291);
DFFARX1 I_7(I1470,I7570,,,I7816,);
not I_8(I6329,I1477);
and I_9(I7535,I7714,I7946);
and I_10(I7915,I7881,I7898);
DFFARX1 I_11(I1470,I6329,,,I6291,);
nor I_12(I10120,I7538,I7535);
endmodule


