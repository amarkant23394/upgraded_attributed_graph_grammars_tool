module test_I4524(I2173,I1477,I1470,I2311,I2146,I4524);
input I2173,I1477,I1470,I2311,I2146;
output I4524;
wire I4595,I4544,I4561,I2164,I4708,I2152,I2345,I4742,I4725,I4578,I2161,I2263,I2158;
DFFARX1 I_0(I4578,I1470,I4544,,,I4595,);
not I_1(I4544,I1477);
nor I_2(I4524,I4742,I4595);
nand I_3(I4561,I2152,I2173);
DFFARX1 I_4(I1470,,,I2164,);
nand I_5(I4708,I2146,I2164);
DFFARX1 I_6(I1470,,,I2152,);
DFFARX1 I_7(I1470,,,I2345,);
DFFARX1 I_8(I4725,I1470,I4544,,,I4742,);
and I_9(I4725,I4708,I2158);
and I_10(I4578,I4561,I2161);
nand I_11(I2161,I2345,I2311);
DFFARX1 I_12(I1470,,,I2263,);
not I_13(I2158,I2263);
endmodule


