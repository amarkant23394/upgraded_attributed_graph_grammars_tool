module test_final(IN_1_2_l_2,IN_2_2_l_2,IN_3_2_l_2,IN_6_2_l_2,IN_1_3_l_2,IN_2_3_l_2,IN_4_3_l_2,IN_1_4_l_2,IN_2_4_l_2,IN_3_4_l_2,IN_6_4_l_2,blif_clk_net_1_r_7,blif_reset_net_1_r_7,G42_1_r_7,n_572_1_r_7,n_573_1_r_7,n_549_1_r_7,n_569_1_r_7,G199_4_r_7,G214_4_r_7,ACVQN1_5_r_7,P6_5_r_7);
input IN_1_2_l_2,IN_2_2_l_2,IN_3_2_l_2,IN_6_2_l_2,IN_1_3_l_2,IN_2_3_l_2,IN_4_3_l_2,IN_1_4_l_2,IN_2_4_l_2,IN_3_4_l_2,IN_6_4_l_2,blif_clk_net_1_r_7,blif_reset_net_1_r_7;
output G42_1_r_7,n_572_1_r_7,n_573_1_r_7,n_549_1_r_7,n_569_1_r_7,G199_4_r_7,G214_4_r_7,ACVQN1_5_r_7,P6_5_r_7;
wire G42_1_r_2,n_572_1_r_2,n_573_1_r_2,n_549_1_r_2,n_569_1_r_2,n_452_1_r_2,n_42_2_r_2,G199_2_r_2,ACVQN1_5_r_2,P6_5_r_2,N3_2_l_2,G199_2_l_2,n13_2,ACVQN2_3_l_2,n16_2,N1_4_l_2,n26_2,n17_internal_2,n17_2,n4_1_r_2,N3_2_r_2,P6_5_r_internal_2,n18_2,n19_2,n20_2,n21_2,n22_2,n23_2,n24_2,n25_2,n_431_0_l_7,n8_7,n43_7,n27_7,ACVQN1_5_l_7,n44_7,n4_1_r_7,N1_4_r_7,n26_7,n5_7,P6_5_r_internal_7,n28_7,n29_7,n30_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7;
DFFARX1 I_0(n4_1_r_2,blif_clk_net_1_r_7,n8_7,G42_1_r_2,);
nor I_1(n_572_1_r_2,n26_2,n18_2);
nand I_2(n_573_1_r_2,n17_2,n19_2);
nor I_3(n_549_1_r_2,G199_2_l_2,n20_2);
nand I_4(n_569_1_r_2,n13_2,n19_2);
not I_5(n_452_1_r_2,n_573_1_r_2);
nor I_6(n_42_2_r_2,ACVQN2_3_l_2,n18_2);
DFFARX1 I_7(N3_2_r_2,blif_clk_net_1_r_7,n8_7,G199_2_r_2,);
DFFARX1 I_8(ACVQN2_3_l_2,blif_clk_net_1_r_7,n8_7,ACVQN1_5_r_2,);
not I_9(P6_5_r_2,P6_5_r_internal_2);
and I_10(N3_2_l_2,IN_6_2_l_2,n24_2);
DFFARX1 I_11(N3_2_l_2,blif_clk_net_1_r_7,n8_7,G199_2_l_2,);
not I_12(n13_2,G199_2_l_2);
DFFARX1 I_13(IN_1_3_l_2,blif_clk_net_1_r_7,n8_7,ACVQN2_3_l_2,);
DFFARX1 I_14(IN_2_3_l_2,blif_clk_net_1_r_7,n8_7,n16_2,);
and I_15(N1_4_l_2,IN_6_4_l_2,n25_2);
DFFARX1 I_16(N1_4_l_2,blif_clk_net_1_r_7,n8_7,n26_2,);
DFFARX1 I_17(IN_3_4_l_2,blif_clk_net_1_r_7,n8_7,n17_internal_2,);
not I_18(n17_2,n17_internal_2);
nor I_19(n4_1_r_2,n26_2,n22_2);
nor I_20(N3_2_r_2,n17_2,n23_2);
DFFARX1 I_21(G199_2_l_2,blif_clk_net_1_r_7,n8_7,P6_5_r_internal_2,);
nor I_22(n18_2,IN_1_2_l_2,IN_3_2_l_2);
nand I_23(n19_2,IN_4_3_l_2,n16_2);
nor I_24(n20_2,n26_2,n21_2);
not I_25(n21_2,n18_2);
and I_26(n22_2,IN_4_3_l_2,n16_2);
nor I_27(n23_2,n13_2,n21_2);
nand I_28(n24_2,IN_2_2_l_2,IN_3_2_l_2);
nand I_29(n25_2,IN_1_4_l_2,IN_2_4_l_2);
DFFARX1 I_30(n4_1_r_7,blif_clk_net_1_r_7,n8_7,G42_1_r_7,);
nor I_31(n_572_1_r_7,n30_7,n31_7);
nand I_32(n_573_1_r_7,n28_7,G42_1_r_2);
nor I_33(n_549_1_r_7,ACVQN1_5_l_7,n35_7);
nand I_34(n_569_1_r_7,n32_7,n33_7);
DFFARX1 I_35(N1_4_r_7,blif_clk_net_1_r_7,n8_7,G199_4_r_7,);
DFFARX1 I_36(n26_7,blif_clk_net_1_r_7,n8_7,G214_4_r_7,);
DFFARX1 I_37(n5_7,blif_clk_net_1_r_7,n8_7,ACVQN1_5_r_7,);
not I_38(P6_5_r_7,P6_5_r_internal_7);
or I_39(n_431_0_l_7,n36_7,n_42_2_r_2);
not I_40(n8_7,blif_reset_net_1_r_7);
DFFARX1 I_41(n_431_0_l_7,blif_clk_net_1_r_7,n8_7,n43_7,);
not I_42(n27_7,n43_7);
DFFARX1 I_43(P6_5_r_2,blif_clk_net_1_r_7,n8_7,ACVQN1_5_l_7,);
DFFARX1 I_44(G199_2_r_2,blif_clk_net_1_r_7,n8_7,n44_7,);
nor I_45(n4_1_r_7,n30_7,n38_7);
nor I_46(N1_4_r_7,n27_7,n40_7);
nand I_47(n26_7,n39_7,G42_1_r_2);
not I_48(n5_7,n_572_1_r_2);
DFFARX1 I_49(ACVQN1_5_l_7,blif_clk_net_1_r_7,n8_7,P6_5_r_internal_7,);
nor I_50(n28_7,n26_7,n29_7);
not I_51(n29_7,n_452_1_r_2);
not I_52(n30_7,n_549_1_r_2);
nand I_53(n31_7,n27_7,n29_7);
nor I_54(n32_7,ACVQN1_5_l_7,n34_7);
nor I_55(n33_7,n29_7,n_572_1_r_2);
not I_56(n34_7,G42_1_r_2);
nor I_57(n35_7,n43_7,n44_7);
and I_58(n36_7,n37_7,ACVQN1_5_r_2);
nor I_59(n37_7,n30_7,n_572_1_r_2);
nand I_60(n38_7,n29_7,n_572_1_r_2);
nor I_61(n39_7,n_569_1_r_2,n_572_1_r_2);
nor I_62(n40_7,n44_7,n41_7);
nor I_63(n41_7,n34_7,n42_7);
nand I_64(n42_7,n5_7,n_452_1_r_2);
endmodule


