module Benchmark_testing100(I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1451,I1458,I2059,I2083,I2065,I2068,I2056,I2074,I2077,I2062,I2071,I2080);
input I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1451,I1458;
output I2059,I2083,I2065,I2068,I2056,I2074,I2077,I2062,I2071,I2080;
wire I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1451,I1458,I1493,I2595,I1519,I1536,I1485,I1558,I2592,I1584,I1592,I1609,I2598,I1626,I2583,I1643,I1660,I2586,I1677,I2607,I1694,I2604,I1711,I1461,I1742,I1759,I1776,I1793,I1473,I1467,I1838,I1482,I1476,I1883,I1900,I2589,I1917,I2601,I1934,I1960,I1968,I1470,I1464,I2022,I2030,I1479,I2091,I3161,I2117,I2125,I3176,I2142,I3179,I2168,I2190,I3185,I2216,I2224,I3167,I2241,I2267,I2289,I3164,I2329,I2346,I2354,I2371,I2402,I3170,I2419,I3182,I2445,I2453,I2498,I3173,I2515,I2615,I2641,I2649,I2666,I2683,I2709,I2717,I2743,I2751,I2768,I2785,I2802,I2842,I2850,I2867,I2884,I2901,I2932,I2949,I2975,I2983,I3014,I3045,I3062,I3093,I3193,I3219,I3227,I3267,I3275,I3292,I3309,I3349,I3371,I3388,I3414,I3422,I3439,I3456,I3473,I3490,I3535,I3566,I3583,I3609,I3617,I3648,I3665,I3682,I3699;
not I_0 (I1493,I1458);
DFFARX1 I_1 (I2595,I1451,I1493,I1519,);
DFFARX1 I_2 (I1519,I1451,I1493,I1536,);
not I_3 (I1485,I1536);
not I_4 (I1558,I1519);
DFFARX1 I_5 (I2592,I1451,I1493,I1584,);
not I_6 (I1592,I1584);
and I_7 (I1609,I1558,I2598);
not I_8 (I1626,I2583);
nand I_9 (I1643,I1626,I2598);
not I_10 (I1660,I2586);
nor I_11 (I1677,I1660,I2607);
nand I_12 (I1694,I1677,I2604);
nor I_13 (I1711,I1694,I1643);
DFFARX1 I_14 (I1711,I1451,I1493,I1461,);
not I_15 (I1742,I1694);
not I_16 (I1759,I2607);
nand I_17 (I1776,I1759,I2598);
nor I_18 (I1793,I2607,I2583);
nand I_19 (I1473,I1609,I1793);
nand I_20 (I1467,I1558,I2607);
nand I_21 (I1838,I1660,I2583);
DFFARX1 I_22 (I1838,I1451,I1493,I1482,);
DFFARX1 I_23 (I1838,I1451,I1493,I1476,);
not I_24 (I1883,I2583);
nor I_25 (I1900,I1883,I2589);
and I_26 (I1917,I1900,I2601);
or I_27 (I1934,I1917,I2586);
DFFARX1 I_28 (I1934,I1451,I1493,I1960,);
nand I_29 (I1968,I1960,I1626);
nor I_30 (I1470,I1968,I1776);
nor I_31 (I1464,I1960,I1592);
DFFARX1 I_32 (I1960,I1451,I1493,I2022,);
not I_33 (I2030,I2022);
nor I_34 (I1479,I2030,I1742);
not I_35 (I2091,I1458);
DFFARX1 I_36 (I3161,I1451,I2091,I2117,);
nand I_37 (I2125,I3176,I3161);
and I_38 (I2142,I2125,I3179);
DFFARX1 I_39 (I2142,I1451,I2091,I2168,);
nor I_40 (I2059,I2168,I2117);
not I_41 (I2190,I2168);
DFFARX1 I_42 (I3185,I1451,I2091,I2216,);
nand I_43 (I2224,I2216,I3167);
not I_44 (I2241,I2224);
DFFARX1 I_45 (I2241,I1451,I2091,I2267,);
not I_46 (I2083,I2267);
nor I_47 (I2289,I2117,I2224);
nor I_48 (I2065,I2168,I2289);
DFFARX1 I_49 (I3164,I1451,I2091,I2329,);
DFFARX1 I_50 (I2329,I1451,I2091,I2346,);
not I_51 (I2354,I2346);
not I_52 (I2371,I2329);
nand I_53 (I2068,I2371,I2190);
nand I_54 (I2402,I3164,I3170);
and I_55 (I2419,I2402,I3182);
DFFARX1 I_56 (I2419,I1451,I2091,I2445,);
nor I_57 (I2453,I2445,I2117);
DFFARX1 I_58 (I2453,I1451,I2091,I2056,);
DFFARX1 I_59 (I2445,I1451,I2091,I2074,);
nor I_60 (I2498,I3173,I3170);
not I_61 (I2515,I2498);
nor I_62 (I2077,I2354,I2515);
nand I_63 (I2062,I2371,I2515);
nor I_64 (I2071,I2117,I2498);
DFFARX1 I_65 (I2498,I1451,I2091,I2080,);
not I_66 (I2615,I1458);
DFFARX1 I_67 (I1412,I1451,I2615,I2641,);
not I_68 (I2649,I2641);
nand I_69 (I2666,I1404,I1364);
and I_70 (I2683,I2666,I1420);
DFFARX1 I_71 (I2683,I1451,I2615,I2709,);
not I_72 (I2717,I1372);
DFFARX1 I_73 (I1388,I1451,I2615,I2743,);
not I_74 (I2751,I2743);
nor I_75 (I2768,I2751,I2649);
and I_76 (I2785,I2768,I1372);
nor I_77 (I2802,I2751,I2717);
nor I_78 (I2598,I2709,I2802);
DFFARX1 I_79 (I1436,I1451,I2615,I2842,);
nor I_80 (I2850,I2842,I2709);
not I_81 (I2867,I2850);
not I_82 (I2884,I2842);
nor I_83 (I2901,I2884,I2785);
DFFARX1 I_84 (I2901,I1451,I2615,I2601,);
nand I_85 (I2932,I1380,I1428);
and I_86 (I2949,I2932,I1396);
DFFARX1 I_87 (I2949,I1451,I2615,I2975,);
nor I_88 (I2983,I2975,I2842);
DFFARX1 I_89 (I2983,I1451,I2615,I2583,);
nand I_90 (I3014,I2975,I2884);
nand I_91 (I2592,I2867,I3014);
not I_92 (I3045,I2975);
nor I_93 (I3062,I3045,I2785);
DFFARX1 I_94 (I3062,I1451,I2615,I2604,);
nor I_95 (I3093,I1444,I1428);
or I_96 (I2595,I2842,I3093);
nor I_97 (I2586,I2975,I3093);
or I_98 (I2589,I2709,I3093);
DFFARX1 I_99 (I3093,I1451,I2615,I2607,);
not I_100 (I3193,I1458);
DFFARX1 I_101 (I1461,I1451,I3193,I3219,);
and I_102 (I3227,I3219,I1464);
DFFARX1 I_103 (I3227,I1451,I3193,I3176,);
DFFARX1 I_104 (I1464,I1451,I3193,I3267,);
not I_105 (I3275,I1479);
not I_106 (I3292,I1485);
nand I_107 (I3309,I3292,I3275);
nor I_108 (I3164,I3267,I3309);
DFFARX1 I_109 (I3309,I1451,I3193,I3349,);
not I_110 (I3185,I3349);
not I_111 (I3371,I1473);
nand I_112 (I3388,I3292,I3371);
DFFARX1 I_113 (I3388,I1451,I3193,I3414,);
not I_114 (I3422,I3414);
not I_115 (I3439,I1470);
nand I_116 (I3456,I3439,I1467);
and I_117 (I3473,I3275,I3456);
nor I_118 (I3490,I3388,I3473);
DFFARX1 I_119 (I3490,I1451,I3193,I3161,);
DFFARX1 I_120 (I3473,I1451,I3193,I3182,);
nor I_121 (I3535,I1470,I1461);
nor I_122 (I3173,I3388,I3535);
or I_123 (I3566,I1470,I1461);
nor I_124 (I3583,I1476,I1482);
DFFARX1 I_125 (I3583,I1451,I3193,I3609,);
not I_126 (I3617,I3609);
nor I_127 (I3179,I3617,I3422);
nand I_128 (I3648,I3617,I3267);
not I_129 (I3665,I1476);
nand I_130 (I3682,I3665,I3371);
nand I_131 (I3699,I3617,I3682);
nand I_132 (I3170,I3699,I3648);
nand I_133 (I3167,I3682,I3566);
endmodule


