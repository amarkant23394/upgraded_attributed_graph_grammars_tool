module test_I5070(I1477,I1470,I3504,I5070);
input I1477,I1470,I3504;
output I5070;
wire I5416,I3388,I3350,I3521,I3380,I3846,I5122,I1495,I3555,I3589,I5249,I3747,I3356,I5105,I5481;
nand I_0(I5416,I5122,I3356);
not I_1(I3388,I1477);
DFFARX1 I_2(I1470,I3388,,,I3350,);
nor I_3(I3521,I3504,I1495);
nand I_4(I3380,I3521,I3846);
and I_5(I5070,I5249,I5481);
nor I_6(I3846,I3747,I3555);
not I_7(I5122,I3350);
DFFARX1 I_8(I1470,,,I1495,);
DFFARX1 I_9(I1470,I3388,,,I3555,);
and I_10(I3589,I3521);
not I_11(I5249,I3380);
DFFARX1 I_12(I1470,I3388,,,I3747,);
DFFARX1 I_13(I3589,I1470,I3388,,,I3356,);
not I_14(I5105,I1477);
DFFARX1 I_15(I5416,I1470,I5105,,,I5481,);
endmodule


