module test_I1458(I1287,I1215,I1247,I1223,I1263,I1458);
input I1287,I1215,I1247,I1223,I1263;
output I1458;
wire I1376,I1393,I1441,I1359,I1424;
nor I_0(I1376,I1215,I1223);
nand I_1(I1393,I1376,I1287);
nand I_2(I1441,I1424,I1247);
nand I_3(I1458,I1441,I1393);
not I_4(I1359,I1263);
nor I_5(I1424,I1359,I1215);
endmodule


