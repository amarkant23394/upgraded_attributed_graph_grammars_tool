module test_I8527(I4629,I1477,I6011,I1470,I4824,I8527);
input I4629,I1477,I6011,I1470,I4824;
output I8527;
wire I8233,I5751,I5713,I6028,I6110,I6127,I4533,I4509,I5722;
nand I_0(I8527,I8233,I5713);
not I_1(I8233,I5722);
not I_2(I5751,I1477);
DFFARX1 I_3(I6127,I1470,I5751,,,I5713,);
DFFARX1 I_4(I6011,I1470,I5751,,,I6028,);
DFFARX1 I_5(I4509,I1470,I5751,,,I6110,);
and I_6(I6127,I6110,I4533);
or I_7(I4533,I4824,I4629);
DFFARX1 I_8(I1470,,,I4509,);
DFFARX1 I_9(I6028,I1470,I5751,,,I5722,);
endmodule


