module test_final(G18_1_l_14,G15_1_l_14,IN_1_1_l_14,IN_4_1_l_14,IN_5_1_l_14,IN_7_1_l_14,IN_9_1_l_14,IN_10_1_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_4_3_l_14,blif_clk_net_1_r_12,blif_reset_net_1_r_12,G42_1_r_12,n_572_1_r_12,n_573_1_r_12,n_549_1_r_12,n_42_2_r_12,G199_2_r_12,ACVQN1_5_r_12,P6_5_r_12);
input G18_1_l_14,G15_1_l_14,IN_1_1_l_14,IN_4_1_l_14,IN_5_1_l_14,IN_7_1_l_14,IN_9_1_l_14,IN_10_1_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_4_3_l_14,blif_clk_net_1_r_12,blif_reset_net_1_r_12;
output G42_1_r_12,n_572_1_r_12,n_573_1_r_12,n_549_1_r_12,n_42_2_r_12,G199_2_r_12,ACVQN1_5_r_12,P6_5_r_12;
wire G42_1_r_14,n_572_1_r_14,n_573_1_r_14,n_549_1_r_14,n_569_1_r_14,n_452_1_r_14,n_42_2_r_14,G199_2_r_14,ACVQN1_5_r_14,P6_5_r_14,n4_1_l_14,n15_internal_14,n15_14,ACVQN2_3_l_14,ACVQN1_3_l_14,N3_2_r_14,n_572_1_l_14,P6_5_r_internal_14,n16_14,n17_14,n18_14,n19_14,n20_14,n21_14,n22_14,n23_14,n24_14,n25_14,n26_14,n27_14,n28_14,n_431_0_l_12,n8_12,n41_12,ACVQN1_5_l_12,n22_12,n42_12,n4_1_r_12,N3_2_r_12,n3_12,P6_5_r_internal_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12;
DFFARX1 I_0(n_452_1_r_14,blif_clk_net_1_r_12,n8_12,G42_1_r_14,);
and I_1(n_572_1_r_14,n18_14,n19_14);
nand I_2(n_573_1_r_14,n16_14,n17_14);
nor I_3(n_549_1_r_14,n20_14,n21_14);
or I_4(n_569_1_r_14,n_572_1_l_14,n20_14);
nor I_5(n_452_1_r_14,IN_10_1_l_14,n23_14);
nor I_6(n_42_2_r_14,n20_14,n22_14);
DFFARX1 I_7(N3_2_r_14,blif_clk_net_1_r_12,n8_12,G199_2_r_14,);
DFFARX1 I_8(n_572_1_l_14,blif_clk_net_1_r_12,n8_12,ACVQN1_5_r_14,);
not I_9(P6_5_r_14,P6_5_r_internal_14);
nor I_10(n4_1_l_14,G18_1_l_14,IN_1_1_l_14);
DFFARX1 I_11(n4_1_l_14,blif_clk_net_1_r_12,n8_12,n15_internal_14,);
not I_12(n15_14,n15_internal_14);
DFFARX1 I_13(IN_1_3_l_14,blif_clk_net_1_r_12,n8_12,ACVQN2_3_l_14,);
DFFARX1 I_14(IN_2_3_l_14,blif_clk_net_1_r_12,n8_12,ACVQN1_3_l_14,);
and I_15(N3_2_r_14,n26_14,n27_14);
nor I_16(n_572_1_l_14,G15_1_l_14,IN_7_1_l_14);
DFFARX1 I_17(ACVQN2_3_l_14,blif_clk_net_1_r_12,n8_12,P6_5_r_internal_14,);
nor I_18(n16_14,IN_9_1_l_14,IN_10_1_l_14);
not I_19(n17_14,n_572_1_l_14);
nor I_20(n18_14,IN_5_1_l_14,IN_9_1_l_14);
nand I_21(n19_14,IN_4_3_l_14,ACVQN1_3_l_14);
nor I_22(n20_14,G18_1_l_14,IN_5_1_l_14);
nor I_23(n21_14,n15_14,n22_14);
nand I_24(n22_14,n24_14,n25_14);
nand I_25(n23_14,n15_14,n24_14);
not I_26(n24_14,IN_9_1_l_14);
not I_27(n25_14,IN_5_1_l_14);
nor I_28(n26_14,IN_10_1_l_14,n20_14);
nand I_29(n27_14,IN_4_1_l_14,n28_14);
not I_30(n28_14,G15_1_l_14);
DFFARX1 I_31(n4_1_r_12,blif_clk_net_1_r_12,n8_12,G42_1_r_12,);
nor I_32(n_572_1_r_12,n29_12,n30_12);
nand I_33(n_573_1_r_12,n26_12,n27_12);
nor I_34(n_549_1_r_12,n33_12,n34_12);
and I_35(n_42_2_r_12,n42_12,n39_12);
DFFARX1 I_36(N3_2_r_12,blif_clk_net_1_r_12,n8_12,G199_2_r_12,);
DFFARX1 I_37(n3_12,blif_clk_net_1_r_12,n8_12,ACVQN1_5_r_12,);
not I_38(P6_5_r_12,P6_5_r_internal_12);
or I_39(n_431_0_l_12,n36_12,ACVQN1_5_r_14);
not I_40(n8_12,blif_reset_net_1_r_12);
DFFARX1 I_41(n_431_0_l_12,blif_clk_net_1_r_12,n8_12,n41_12,);
DFFARX1 I_42(G42_1_r_14,blif_clk_net_1_r_12,n8_12,ACVQN1_5_l_12,);
not I_43(n22_12,ACVQN1_5_l_12);
DFFARX1 I_44(n_569_1_r_14,blif_clk_net_1_r_12,n8_12,n42_12,);
nor I_45(n4_1_r_12,n41_12,n31_12);
nor I_46(N3_2_r_12,n22_12,n40_12);
not I_47(n3_12,n39_12);
DFFARX1 I_48(ACVQN1_5_l_12,blif_clk_net_1_r_12,n8_12,P6_5_r_internal_12,);
and I_49(n26_12,n_573_1_r_14,n_549_1_r_14);
nor I_50(n27_12,n28_12,n29_12);
not I_51(n28_12,n_572_1_r_14);
nand I_52(n29_12,n31_12,n32_12);
nand I_53(n30_12,n42_12,n_572_1_r_14);
not I_54(n31_12,P6_5_r_14);
not I_55(n32_12,G199_2_r_14);
nand I_56(n33_12,n31_12,n35_12);
nand I_57(n34_12,n_573_1_r_14,n_549_1_r_14);
nand I_58(n35_12,n41_12,n42_12);
and I_59(n36_12,n37_12,n_42_2_r_14);
nor I_60(n37_12,n38_12,n_572_1_r_14);
not I_61(n38_12,G42_1_r_14);
nor I_62(n39_12,n38_12,n_573_1_r_14);
nor I_63(n40_12,n39_12,P6_5_r_14);
endmodule


