module test_final(IN_1_0_l_5,IN_2_0_l_5,IN_3_0_l_5,IN_4_0_l_5,IN_1_1_l_5,IN_2_1_l_5,IN_3_1_l_5,IN_1_10_l_5,IN_2_10_l_5,IN_3_10_l_5,IN_4_10_l_5,blif_clk_net_5_r_4,blif_reset_net_5_r_4,N1508_0_r_4,N6147_2_r_4,n_429_or_0_5_r_4,G78_5_r_4,n_576_5_r_4,n_547_5_r_4,N1507_6_r_4,N1508_6_r_4);
input IN_1_0_l_5,IN_2_0_l_5,IN_3_0_l_5,IN_4_0_l_5,IN_1_1_l_5,IN_2_1_l_5,IN_3_1_l_5,IN_1_10_l_5,IN_2_10_l_5,IN_3_10_l_5,IN_4_10_l_5,blif_clk_net_5_r_4,blif_reset_net_5_r_4;
output N1508_0_r_4,N6147_2_r_4,n_429_or_0_5_r_4,G78_5_r_4,n_576_5_r_4,n_547_5_r_4,N1507_6_r_4,N1508_6_r_4;
wire N1371_0_r_5,N1508_0_r_5,N6147_2_r_5,n_429_or_0_5_r_5,G78_5_r_5,n_576_5_r_5,n_102_5_r_5,n_547_5_r_5,N1507_6_r_5,N1508_6_r_5,n_431_5_r_5,n26_5,n27_5,n28_5,n29_5,n30_5,n31_5,n32_5,n33_5,n34_5,n35_5,n36_5,n37_5,n38_5,n39_5,n40_5,n41_5,n42_5,n43_5,n44_5,N1371_0_r_4,n_102_5_r_4,n_431_5_r_4,n4_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4;
nor I_0(N1371_0_r_5,n28_5,n39_5);
not I_1(N1508_0_r_5,n39_5);
nor I_2(N6147_2_r_5,n28_5,n37_5);
nand I_3(n_429_or_0_5_r_5,n30_5,n32_5);
DFFARX1 I_4(n_431_5_r_5,blif_clk_net_5_r_4,n4_4,G78_5_r_5,);
nand I_5(n_576_5_r_5,n26_5,n27_5);
not I_6(n_102_5_r_5,n28_5);
nand I_7(n_547_5_r_5,n31_5,n32_5);
nor I_8(N1507_6_r_5,n30_5,n32_5);
nor I_9(N1508_6_r_5,n39_5,n41_5);
nand I_10(n_431_5_r_5,n34_5,n35_5);
nor I_11(n26_5,n29_5,n30_5);
nor I_12(n27_5,IN_2_0_l_5,n28_5);
nor I_13(n28_5,n29_5,n44_5);
not I_14(n29_5,IN_1_0_l_5);
nand I_15(n30_5,N1508_0_r_5,n43_5);
nor I_16(n31_5,n28_5,n33_5);
nor I_17(n32_5,IN_3_1_l_5,n40_5);
nor I_18(n33_5,IN_2_0_l_5,n29_5);
or I_19(n34_5,IN_2_0_l_5,n29_5);
nand I_20(n35_5,n32_5,n36_5);
not I_21(n36_5,n30_5);
nor I_22(n37_5,N1507_6_r_5,n38_5);
and I_23(n38_5,n39_5,n40_5);
nand I_24(n39_5,IN_1_10_l_5,IN_2_10_l_5);
nand I_25(n40_5,IN_1_1_l_5,IN_2_1_l_5);
nand I_26(n41_5,n28_5,n42_5);
or I_27(n42_5,n32_5,n36_5);
or I_28(n43_5,IN_3_10_l_5,IN_4_10_l_5);
nor I_29(n44_5,IN_3_0_l_5,IN_4_0_l_5);
nor I_30(N1371_0_r_4,n25_4,n29_4);
nor I_31(N1508_0_r_4,n25_4,n32_4);
nor I_32(N6147_2_r_4,n24_4,n31_4);
or I_33(n_429_or_0_5_r_4,n23_4,n30_4);
DFFARX1 I_34(n_431_5_r_4,blif_clk_net_5_r_4,n4_4,G78_5_r_4,);
nand I_35(n_576_5_r_4,n22_4,n23_4);
nand I_36(n_102_5_r_4,n34_4,n35_4);
nand I_37(n_547_5_r_4,n26_4,n27_4);
nor I_38(N1507_6_r_4,n27_4,n30_4);
nor I_39(N1508_6_r_4,n30_4,n33_4);
nand I_40(n_431_5_r_4,n_102_5_r_4,n28_4);
not I_41(n4_4,blif_reset_net_5_r_4);
nor I_42(n22_4,n24_4,n25_4);
nor I_43(n23_4,n37_4,G78_5_r_5);
not I_44(n24_4,n_102_5_r_4);
nand I_45(n25_4,n_429_or_0_5_r_5,n_547_5_r_5);
nor I_46(n26_4,n23_4,n24_4);
not I_47(n27_4,n25_4);
nand I_48(n28_4,n23_4,n29_4);
nor I_49(n29_4,n25_4,n_102_5_r_5);
not I_50(n30_4,n29_4);
nor I_51(n31_4,N1371_0_r_4,n32_4);
nor I_52(n32_4,n23_4,n29_4);
nand I_53(n33_4,n23_4,n24_4);
nor I_54(n34_4,N6147_2_r_5,n_576_5_r_5);
or I_55(n35_4,n36_4,N1371_0_r_5);
nor I_56(n36_4,N1508_6_r_5,n_429_or_0_5_r_5);
or I_57(n37_4,N1371_0_r_5,N6147_2_r_5);
endmodule


