module test_I17594(I15713,I1477,I13746,I15880,I1470,I17594);
input I15713,I1477,I13746,I15880,I1470;
output I17594;
wire I15897,I15928,I15576,I15611,I16007;
and I_0(I15897,I15713,I15880);
DFFARX1 I_1(I13746,I1470,I15611,,,I15928,);
DFFARX1 I_2(I16007,I1470,I15611,,,I15576,);
not I_3(I15611,I1477);
not I_4(I17594,I15576);
or I_5(I16007,I15928,I15897);
endmodule


