module test_I2155(I1477,I1470,I1239,I2155);
input I1477,I1470,I1239;
output I2155;
wire I2181,I2633;
not I_0(I2181,I1477);
DFFARX1 I_1(I2633,I1470,I2181,,,I2155,);
DFFARX1 I_2(I1239,I1470,I2181,,,I2633,);
endmodule


