module test_I2600_rst(I1301_rst,I2600_rst);
,I2600_rst);
input I1301_rst;
output I2600_rst;
wire ;
not I_0(I2600_rst,I1301_rst);
endmodule


