module test_I13197_rst(I1477_rst,I13197_rst);
,I13197_rst);
input I1477_rst;
output I13197_rst;
wire ;
not I_0(I13197_rst,I1477_rst);
endmodule


