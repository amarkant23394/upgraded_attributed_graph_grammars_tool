module test_I16503(I14350,I1477,I1470,I14825,I14359,I16503);
input I14350,I1477,I1470,I14825,I14359;
output I16503;
wire I14362,I16452,I16469,I16240,I16435,I14370;
DFFARX1 I_0(I14825,I1470,I14370,,,I14362,);
and I_1(I16452,I16435,I14362);
DFFARX1 I_2(I16452,I1470,I16240,,,I16469,);
not I_3(I16240,I1477);
nand I_4(I16435,I14359,I14350);
not I_5(I16503,I16469);
not I_6(I14370,I1477);
endmodule


