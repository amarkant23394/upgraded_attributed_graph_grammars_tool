module test_I1410(I1239,I1223,I1410);
input I1239,I1223;
output I1410;
wire ;
nor I_0(I1410,I1223,I1239);
endmodule


