module test_final(IN_1_1_l_2,IN_2_1_l_2,IN_3_1_l_2,G18_7_l_2,G15_7_l_2,IN_1_7_l_2,IN_4_7_l_2,IN_5_7_l_2,IN_7_7_l_2,IN_9_7_l_2,IN_10_7_l_2,IN_1_8_l_2,IN_2_8_l_2,IN_3_8_l_2,IN_6_8_l_2,blif_clk_net_5_r_9,blif_reset_net_5_r_9,N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,G78_5_r_9,n_576_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9);
input IN_1_1_l_2,IN_2_1_l_2,IN_3_1_l_2,G18_7_l_2,G15_7_l_2,IN_1_7_l_2,IN_4_7_l_2,IN_5_7_l_2,IN_7_7_l_2,IN_9_7_l_2,IN_10_7_l_2,IN_1_8_l_2,IN_2_8_l_2,IN_3_8_l_2,IN_6_8_l_2,blif_clk_net_5_r_9,blif_reset_net_5_r_9;
output N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,G78_5_r_9,n_576_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9;
wire N1371_0_r_2,N1508_0_r_2,N1372_1_r_2,N1508_1_r_2,N6147_2_r_2,N1507_6_r_2,N1508_6_r_2,G42_7_r_2,n_572_7_r_2,n_573_7_r_2,n_549_7_r_2,n_569_7_r_2,n_452_7_r_2,n4_7_l_2,n59_2,n33_2,N3_8_l_2,n32_internal_2,n32_2,n4_7_r_2,n34_2,n35_2,n36_2,n37_2,n38_2,n39_2,n40_2,n41_2,n42_2,n43_2,n44_2,n45_2,n46_2,n47_2,n48_2,n49_2,n50_2,n51_2,n52_2,n53_2,n54_2,n55_2,n56_2,n57_2,n58_2,n_429_or_0_5_r_9,n_102_5_r_9,I_BUFF_1_9_r_9,n4_7_l_9,n10_9,n62_9,N3_8_l_9,n63_9,n38_9,n_431_5_r_9,N3_8_r_9,n39_9,n40_9,n41_9,n42_9,n43_9,n44_9,n45_9,n46_9,n47_9,n48_9,n49_9,n50_9,n51_9,n52_9,n53_9,n54_9,n55_9,n56_9,n57_9,n58_9,n59_9,n60_9,n61_9;
nor I_0(N1371_0_r_2,n32_2,n35_2);
nor I_1(N1508_0_r_2,n32_2,n55_2);
not I_2(N1372_1_r_2,n54_2);
nor I_3(N1508_1_r_2,n59_2,n54_2);
nor I_4(N6147_2_r_2,n42_2,n43_2);
nor I_5(N1507_6_r_2,n40_2,n53_2);
nor I_6(N1508_6_r_2,n33_2,n50_2);
DFFARX1 I_7(n4_7_r_2,blif_clk_net_5_r_9,n10_9,G42_7_r_2,);
nor I_8(n_572_7_r_2,n36_2,n37_2);
or I_9(n_573_7_r_2,n34_2,n35_2);
nor I_10(n_549_7_r_2,n40_2,n41_2);
nand I_11(n_569_7_r_2,n38_2,n39_2);
nor I_12(n_452_7_r_2,n59_2,n35_2);
nor I_13(n4_7_l_2,G18_7_l_2,IN_1_7_l_2);
DFFARX1 I_14(n4_7_l_2,blif_clk_net_5_r_9,n10_9,n59_2,);
not I_15(n33_2,n59_2);
and I_16(N3_8_l_2,IN_6_8_l_2,n49_2);
DFFARX1 I_17(N3_8_l_2,blif_clk_net_5_r_9,n10_9,n32_internal_2,);
not I_18(n32_2,n32_internal_2);
nor I_19(n4_7_r_2,n59_2,n36_2);
not I_20(n34_2,n39_2);
nor I_21(n35_2,IN_1_8_l_2,IN_3_8_l_2);
nor I_22(n36_2,G18_7_l_2,IN_5_7_l_2);
or I_23(n37_2,IN_9_7_l_2,IN_10_7_l_2);
not I_24(n38_2,n40_2);
nand I_25(n39_2,n45_2,n57_2);
nor I_26(n40_2,IN_3_1_l_2,n47_2);
nor I_27(n41_2,n32_2,n36_2);
not I_28(n42_2,n53_2);
nand I_29(n43_2,n44_2,n45_2);
nand I_30(n44_2,n38_2,n46_2);
not I_31(n45_2,IN_10_7_l_2);
nand I_32(n46_2,n47_2,n48_2);
nand I_33(n47_2,IN_1_1_l_2,IN_2_1_l_2);
or I_34(n48_2,G15_7_l_2,IN_7_7_l_2);
nand I_35(n49_2,IN_2_8_l_2,IN_3_8_l_2);
nand I_36(n50_2,n51_2,n52_2);
not I_37(n51_2,n47_2);
nand I_38(n52_2,n38_2,n53_2);
nor I_39(n53_2,IN_5_7_l_2,IN_9_7_l_2);
nand I_40(n54_2,n42_2,n56_2);
nor I_41(n55_2,n34_2,n56_2);
nor I_42(n56_2,G15_7_l_2,IN_7_7_l_2);
nand I_43(n57_2,IN_4_7_l_2,n58_2);
not I_44(n58_2,G15_7_l_2);
nor I_45(N6147_2_r_9,n62_9,n46_9);
not I_46(N1372_4_r_9,n59_9);
nor I_47(N1508_4_r_9,n58_9,n59_9);
nand I_48(n_429_or_0_5_r_9,n_431_5_r_9,n42_9);
DFFARX1 I_49(n_431_5_r_9,blif_clk_net_5_r_9,n10_9,G78_5_r_9,);
nand I_50(n_576_5_r_9,n39_9,n40_9);
not I_51(n_102_5_r_9,I_BUFF_1_9_r_9);
nand I_52(n_547_5_r_9,n43_9,N1507_6_r_2);
and I_53(n_42_8_r_9,n44_9,n_572_7_r_2);
DFFARX1 I_54(N3_8_r_9,blif_clk_net_5_r_9,n10_9,G199_8_r_9,);
nor I_55(N6147_9_r_9,n41_9,n45_9);
nor I_56(N6134_9_r_9,n45_9,n51_9);
nor I_57(I_BUFF_1_9_r_9,n41_9,N1507_6_r_2);
nor I_58(n4_7_l_9,N1508_6_r_2,n_572_7_r_2);
not I_59(n10_9,blif_reset_net_5_r_9);
DFFARX1 I_60(n4_7_l_9,blif_clk_net_5_r_9,n10_9,n62_9,);
and I_61(N3_8_l_9,n57_9,n_569_7_r_2);
DFFARX1 I_62(N3_8_l_9,blif_clk_net_5_r_9,n10_9,n63_9,);
not I_63(n38_9,n63_9);
nor I_64(n_431_5_r_9,N1372_1_r_2,n_549_7_r_2);
nor I_65(N3_8_r_9,n_102_5_r_9,n53_9);
nor I_66(n39_9,I_BUFF_1_9_r_9,n42_9);
not I_67(n40_9,n41_9);
nand I_68(n41_9,N1371_0_r_2,n_452_7_r_2);
nor I_69(n42_9,N6147_2_r_2,N1371_0_r_2);
nor I_70(n43_9,n63_9,n41_9);
nor I_71(n44_9,n_573_7_r_2,N1371_0_r_2);
and I_72(n45_9,n52_9,N1508_1_r_2);
nor I_73(n46_9,n47_9,n48_9);
nor I_74(n47_9,n49_9,n50_9);
not I_75(n48_9,n_429_or_0_5_r_9);
not I_76(n49_9,n42_9);
or I_77(n50_9,n63_9,n51_9);
nor I_78(n51_9,N1508_0_r_2,N1372_1_r_2);
nor I_79(n52_9,n49_9,n_549_7_r_2);
nor I_80(n53_9,n54_9,n55_9);
nor I_81(n54_9,n56_9,n_549_7_r_2);
or I_82(n55_9,n44_9,N6147_2_r_2);
not I_83(n56_9,N1508_1_r_2);
nand I_84(n57_9,G42_7_r_2,N1508_0_r_2);
nor I_85(n58_9,n62_9,n60_9);
nand I_86(n59_9,n51_9,n61_9);
nor I_87(n60_9,n38_9,n44_9);
nor I_88(n61_9,n_572_7_r_2,n_573_7_r_2);
endmodule


