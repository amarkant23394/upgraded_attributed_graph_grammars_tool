module test_I6640(I1477,I6572,I2742,I4017,I2727,I1470,I6640);
input I1477,I6572,I2742,I4017,I2727,I1470;
output I6640;
wire I6442,I3983,I6510,I3954,I6329,I4068,I2724,I3975,I3966,I6493,I4308,I4034,I6606,I3960,I6589,I6623;
and I_0(I6640,I6442,I6623);
nor I_1(I6442,I3975,I3954);
not I_2(I3983,I1477);
not I_3(I6510,I6493);
not I_4(I3954,I4068);
not I_5(I6329,I1477);
nor I_6(I4068,I2742,I2724);
DFFARX1 I_7(I1470,,,I2724,);
nor I_8(I3975,I4308,I4034);
or I_9(I3966,I4068,I4034);
DFFARX1 I_10(I3966,I1470,I6329,,,I6493,);
DFFARX1 I_11(I2727,I1470,I3983,,,I4308,);
DFFARX1 I_12(I4017,I1470,I3983,,,I4034,);
DFFARX1 I_13(I6589,I1470,I6329,,,I6606,);
DFFARX1 I_14(I1470,I3983,,,I3960,);
and I_15(I6589,I6572,I3960);
nor I_16(I6623,I6606,I6510);
endmodule


