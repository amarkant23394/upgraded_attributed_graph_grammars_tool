module test_I3359(I1750,I1477,I1603,I1470,I3359);
input I1750,I1477,I1603,I1470;
output I3359;
wire I1518,I3388,I1504,I1880,I3747,I1897,I1767;
not I_0(I1518,I1477);
not I_1(I3388,I1477);
nand I_2(I1504,I1767,I1897);
DFFARX1 I_3(I1470,I1518,,,I1880,);
DFFARX1 I_4(I1504,I1470,I3388,,,I3747,);
DFFARX1 I_5(I3747,I1470,I3388,,,I3359,);
nor I_6(I1897,I1880,I1603);
DFFARX1 I_7(I1750,I1470,I1518,,,I1767,);
endmodule


