module test_final(IN_1_2_l_3,IN_2_2_l_3,IN_3_2_l_3,IN_4_2_l_3,IN_5_2_l_3,IN_1_6_l_3,IN_2_6_l_3,IN_3_6_l_3,IN_4_6_l_3,IN_5_6_l_3,IN_1_9_l_3,IN_2_9_l_3,IN_3_9_l_3,IN_4_9_l_3,IN_5_9_l_3,blif_clk_net_7_r_4,blif_reset_net_7_r_4,N1371_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6134_9_r_4);
input IN_1_2_l_3,IN_2_2_l_3,IN_3_2_l_3,IN_4_2_l_3,IN_5_2_l_3,IN_1_6_l_3,IN_2_6_l_3,IN_3_6_l_3,IN_4_6_l_3,IN_5_6_l_3,IN_1_9_l_3,IN_2_9_l_3,IN_3_9_l_3,IN_4_9_l_3,IN_5_9_l_3,blif_clk_net_7_r_4,blif_reset_net_7_r_4;
output N1371_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6134_9_r_4;
wire N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_572_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6147_9_r_3,N6134_9_r_3,I_BUFF_1_9_r_3,n4_7_r_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3,n40_3,n41_3,n42_3,n43_3,n44_3,n45_3,n46_3,n47_3,n48_3,n49_3,n50_3,n51_3,N1508_0_r_4,n_573_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4,n4_7_r_4,n6_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4,n38_4,n39_4,n40_4,n41_4;
not I_0(N1372_1_r_3,n40_3);
nor I_1(N1508_1_r_3,N6147_9_r_3,n40_3);
nor I_2(N1507_6_r_3,n31_3,n42_3);
nor I_3(N1508_6_r_3,n30_3,n38_3);
DFFARX1 I_4(n4_7_r_3,blif_clk_net_7_r_4,n6_4,G42_7_r_3,);
nor I_5(n_572_7_r_3,I_BUFF_1_9_r_3,n35_3);
nand I_6(n_573_7_r_3,n30_3,n31_3);
nor I_7(n_549_7_r_3,N6147_9_r_3,n33_3);
nand I_8(n_569_7_r_3,n30_3,n32_3);
nor I_9(n_452_7_r_3,IN_1_9_l_3,n35_3);
not I_10(N6147_9_r_3,n32_3);
nor I_11(N6134_9_r_3,n36_3,n37_3);
not I_12(I_BUFF_1_9_r_3,n45_3);
nor I_13(n4_7_r_3,IN_1_9_l_3,I_BUFF_1_9_r_3);
not I_14(n30_3,n39_3);
not I_15(n31_3,n35_3);
nand I_16(n32_3,IN_5_6_l_3,n41_3);
nor I_17(n33_3,I_BUFF_1_9_r_3,n34_3);
nand I_18(n34_3,IN_2_6_l_3,n46_3);
nor I_19(n35_3,n43_3,n44_3);
not I_20(n36_3,n34_3);
nor I_21(n37_3,IN_1_9_l_3,N6147_9_r_3);
or I_22(n38_3,n_572_7_r_3,n34_3);
nor I_23(n39_3,IN_5_9_l_3,n44_3);
nand I_24(n40_3,IN_1_9_l_3,n39_3);
nand I_25(n41_3,IN_3_6_l_3,IN_4_6_l_3);
nor I_26(n42_3,n34_3,n45_3);
not I_27(n43_3,IN_2_9_l_3);
nor I_28(n44_3,IN_3_9_l_3,IN_4_9_l_3);
nand I_29(n45_3,n49_3,n50_3);
and I_30(n46_3,IN_1_6_l_3,n47_3);
nand I_31(n47_3,n41_3,n48_3);
not I_32(n48_3,IN_5_6_l_3);
nor I_33(n49_3,IN_1_2_l_3,IN_2_2_l_3);
or I_34(n50_3,IN_5_2_l_3,n51_3);
nor I_35(n51_3,IN_3_2_l_3,IN_4_2_l_3);
nor I_36(N1371_0_r_4,n25_4,n_452_7_r_3);
not I_37(N1508_0_r_4,n25_4);
nor I_38(N1507_6_r_4,n32_4,n33_4);
nor I_39(N1508_6_r_4,n22_4,n29_4);
DFFARX1 I_40(n4_7_r_4,blif_clk_net_7_r_4,n6_4,G42_7_r_4,);
not I_41(n_572_7_r_4,n_573_7_r_4);
nand I_42(n_573_7_r_4,n21_4,n22_4);
nor I_43(n_549_7_r_4,n24_4,n_452_7_r_3);
nand I_44(n_569_7_r_4,n22_4,n23_4);
nor I_45(n_452_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4);
not I_46(N6147_9_r_4,n28_4);
nor I_47(N6134_9_r_4,N1508_0_r_4,n28_4);
not I_48(I_BUFF_1_9_r_4,n21_4);
nor I_49(n4_7_r_4,N6147_9_r_4,n_452_7_r_3);
not I_50(n6_4,blif_reset_net_7_r_4);
nand I_51(n21_4,n39_4,n40_4);
or I_52(n22_4,n31_4,N1372_1_r_3);
not I_53(n23_4,n_452_7_r_3);
nor I_54(n24_4,n25_4,n26_4);
nand I_55(n25_4,n_549_7_r_3,N1508_1_r_3);
nand I_56(n26_4,n21_4,n27_4);
nand I_57(n27_4,n36_4,n37_4);
nand I_58(n28_4,n38_4,N1508_6_r_3);
nand I_59(n29_4,N1508_0_r_4,n30_4);
nand I_60(n30_4,n34_4,n35_4);
nor I_61(n31_4,N1507_6_r_3,n_573_7_r_3);
not I_62(n32_4,n30_4);
nor I_63(n33_4,n21_4,n28_4);
nand I_64(n34_4,N6147_9_r_4,I_BUFF_1_9_r_4);
nand I_65(n35_4,N1508_0_r_4,n27_4);
not I_66(n36_4,N1372_1_r_3);
nand I_67(n37_4,N1508_6_r_3,N1507_6_r_3);
or I_68(n38_4,N1507_6_r_3,n_573_7_r_3);
nor I_69(n39_4,N6134_9_r_3,G42_7_r_3);
or I_70(n40_4,n41_4,n_569_7_r_3);
nor I_71(n41_4,N1508_1_r_3,G42_7_r_3);
endmodule


