module test_I17563(I13749,I15696,I16145,I15628,I17563);
input I13749,I15696,I16145,I15628;
output I17563;
wire I17532,I15832,I16162,I15597;
not I_0(I17563,I17532);
not I_1(I17532,I15597);
nand I_2(I15832,I15628,I13749);
and I_3(I16162,I15696,I16145);
nor I_4(I15597,I15832,I16162);
endmodule


