module test_final(G18_1_l_14,G15_1_l_14,IN_1_1_l_14,IN_4_1_l_14,IN_5_1_l_14,IN_7_1_l_14,IN_9_1_l_14,IN_10_1_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_4_3_l_14,blif_clk_net_1_r_4,blif_reset_net_1_r_4,G42_1_r_4,n_572_1_r_4,n_573_1_r_4,n_549_1_r_4,n_569_1_r_4,ACVQN2_3_r_4,n_266_and_0_3_r_4,ACVQN1_5_r_4,P6_5_r_4);
input G18_1_l_14,G15_1_l_14,IN_1_1_l_14,IN_4_1_l_14,IN_5_1_l_14,IN_7_1_l_14,IN_9_1_l_14,IN_10_1_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_4_3_l_14,blif_clk_net_1_r_4,blif_reset_net_1_r_4;
output G42_1_r_4,n_572_1_r_4,n_573_1_r_4,n_549_1_r_4,n_569_1_r_4,ACVQN2_3_r_4,n_266_and_0_3_r_4,ACVQN1_5_r_4,P6_5_r_4;
wire G42_1_r_14,n_572_1_r_14,n_573_1_r_14,n_549_1_r_14,n_569_1_r_14,n_452_1_r_14,n_42_2_r_14,G199_2_r_14,ACVQN1_5_r_14,P6_5_r_14,n4_1_l_14,n15_internal_14,n15_14,ACVQN2_3_l_14,ACVQN1_3_l_14,N3_2_r_14,n_572_1_l_14,P6_5_r_internal_14,n16_14,n17_14,n18_14,n19_14,n20_14,n21_14,n22_14,n23_14,n24_14,n25_14,n26_14,n27_14,n28_14,n_431_0_l_4,n6_4,G78_0_l_4,ACVQN1_5_l_4,n16_4,n17_internal_4,n17_4,n4_1_r_4,n19_4,n15_internal_4,n15_4,P6_5_r_internal_4,n20_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4;
DFFARX1 I_0(n_452_1_r_14,blif_clk_net_1_r_4,n6_4,G42_1_r_14,);
and I_1(n_572_1_r_14,n18_14,n19_14);
nand I_2(n_573_1_r_14,n16_14,n17_14);
nor I_3(n_549_1_r_14,n20_14,n21_14);
or I_4(n_569_1_r_14,n_572_1_l_14,n20_14);
nor I_5(n_452_1_r_14,IN_10_1_l_14,n23_14);
nor I_6(n_42_2_r_14,n20_14,n22_14);
DFFARX1 I_7(N3_2_r_14,blif_clk_net_1_r_4,n6_4,G199_2_r_14,);
DFFARX1 I_8(n_572_1_l_14,blif_clk_net_1_r_4,n6_4,ACVQN1_5_r_14,);
not I_9(P6_5_r_14,P6_5_r_internal_14);
nor I_10(n4_1_l_14,G18_1_l_14,IN_1_1_l_14);
DFFARX1 I_11(n4_1_l_14,blif_clk_net_1_r_4,n6_4,n15_internal_14,);
not I_12(n15_14,n15_internal_14);
DFFARX1 I_13(IN_1_3_l_14,blif_clk_net_1_r_4,n6_4,ACVQN2_3_l_14,);
DFFARX1 I_14(IN_2_3_l_14,blif_clk_net_1_r_4,n6_4,ACVQN1_3_l_14,);
and I_15(N3_2_r_14,n26_14,n27_14);
nor I_16(n_572_1_l_14,G15_1_l_14,IN_7_1_l_14);
DFFARX1 I_17(ACVQN2_3_l_14,blif_clk_net_1_r_4,n6_4,P6_5_r_internal_14,);
nor I_18(n16_14,IN_9_1_l_14,IN_10_1_l_14);
not I_19(n17_14,n_572_1_l_14);
nor I_20(n18_14,IN_5_1_l_14,IN_9_1_l_14);
nand I_21(n19_14,IN_4_3_l_14,ACVQN1_3_l_14);
nor I_22(n20_14,G18_1_l_14,IN_5_1_l_14);
nor I_23(n21_14,n15_14,n22_14);
nand I_24(n22_14,n24_14,n25_14);
nand I_25(n23_14,n15_14,n24_14);
not I_26(n24_14,IN_9_1_l_14);
not I_27(n25_14,IN_5_1_l_14);
nor I_28(n26_14,IN_10_1_l_14,n20_14);
nand I_29(n27_14,IN_4_1_l_14,n28_14);
not I_30(n28_14,G15_1_l_14);
DFFARX1 I_31(n4_1_r_4,blif_clk_net_1_r_4,n6_4,G42_1_r_4,);
nor I_32(n_572_1_r_4,G78_0_l_4,n17_4);
nand I_33(n_573_1_r_4,n16_4,n_572_1_r_14);
nor I_34(n_549_1_r_4,n22_4,n23_4);
nand I_35(n_569_1_r_4,n20_4,n21_4);
DFFARX1 I_36(n19_4,blif_clk_net_1_r_4,n6_4,ACVQN2_3_r_4,);
nor I_37(n_266_and_0_3_r_4,n15_4,n29_4);
DFFARX1 I_38(n19_4,blif_clk_net_1_r_4,n6_4,ACVQN1_5_r_4,);
not I_39(P6_5_r_4,P6_5_r_internal_4);
or I_40(n_431_0_l_4,n26_4,n_572_1_r_14);
not I_41(n6_4,blif_reset_net_1_r_4);
DFFARX1 I_42(n_431_0_l_4,blif_clk_net_1_r_4,n6_4,G78_0_l_4,);
DFFARX1 I_43(n_573_1_r_14,blif_clk_net_1_r_4,n6_4,ACVQN1_5_l_4,);
not I_44(n16_4,ACVQN1_5_l_4);
DFFARX1 I_45(P6_5_r_14,blif_clk_net_1_r_4,n6_4,n17_internal_4,);
not I_46(n17_4,n17_internal_4);
nor I_47(n4_1_r_4,n30_4,n31_4);
nand I_48(n19_4,n33_4,G42_1_r_14);
DFFARX1 I_49(G78_0_l_4,blif_clk_net_1_r_4,n6_4,n15_internal_4,);
not I_50(n15_4,n15_internal_4);
DFFARX1 I_51(ACVQN1_5_l_4,blif_clk_net_1_r_4,n6_4,P6_5_r_internal_4,);
and I_52(n20_4,n16_4,n_549_1_r_14);
nor I_53(n21_4,n_569_1_r_14,n_572_1_r_14);
nand I_54(n22_4,G78_0_l_4,n25_4);
nand I_55(n23_4,n24_4,n_549_1_r_14);
not I_56(n24_4,n_572_1_r_14);
not I_57(n25_4,n_569_1_r_14);
and I_58(n26_4,n27_4,ACVQN1_5_r_14);
nor I_59(n27_4,n28_4,n_42_2_r_14);
not I_60(n28_4,G42_1_r_14);
not I_61(n29_4,n30_4);
nand I_62(n30_4,n32_4,G199_2_r_14);
nand I_63(n31_4,n25_4,n_549_1_r_14);
nor I_64(n32_4,n33_4,n_572_1_r_14);
not I_65(n33_4,G42_1_r_14);
endmodule


