module test_I8674(I8233,I1477,I4533,I1470,I8674);
input I8233,I1477,I4533,I1470;
output I8674;
wire I8640,I8216,I6110,I8623,I5743,I8657,I6028,I6127,I6079,I5802,I8298,I5719,I5740,I8315;
and I_0(I8674,I8623,I8657);
not I_1(I8640,I8623);
not I_2(I8216,I1477);
DFFARX1 I_3(I1470,,,I6110,);
DFFARX1 I_4(I5743,I1470,I8216,,,I8623,);
nand I_5(I5743,I6127,I6079);
nor I_6(I8657,I8315,I8640);
DFFARX1 I_7(I1470,,,I6028,);
and I_8(I6127,I6110,I4533);
nor I_9(I6079,I6028,I5802);
DFFARX1 I_10(I1470,,,I5802,);
nor I_11(I8298,I8233,I5719);
DFFARX1 I_12(I1470,,,I5719,);
not I_13(I5740,I5802);
nand I_14(I8315,I8298,I5740);
endmodule


