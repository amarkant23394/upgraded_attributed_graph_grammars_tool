module test_I11299(I8830,I9396,I9049,I1470,I6881,I8879,I8862,I8947,I11299);
input I8830,I9396,I9049,I1470,I6881,I8879,I8862,I8947;
output I11299;
wire I11378,I11429,I9066,I11395,I8848,I11327,I9083,I8851,I9413;
nor I_0(I11378,I11327,I8848);
not I_1(I11429,I8848);
DFFARX1 I_2(I9049,I1470,I8862,,,I9066,);
nor I_3(I11299,I11395,I11429);
nand I_4(I11395,I11378,I8851);
nor I_5(I8848,I9083,I9413);
not I_6(I11327,I8830);
nand I_7(I9083,I8879,I6881);
or I_8(I8851,I9083,I9066);
and I_9(I9413,I8947,I9396);
endmodule


