module test_I11895(I9320,I8830,I1477,I11395,I11542,I1470,I11895);
input I9320,I8830,I1477,I11395,I11542,I1470;
output I11895;
wire I9179,I11559,I11641,I11412,I8854,I8827,I11830,I11624,I11576,I8862,I9258,I11813,I11327,I11310;
DFFARX1 I_0(I1470,I8862,,,I9179,);
DFFARX1 I_1(I11542,I1470,I11310,,,I11559,);
and I_2(I11641,I11624,I11576);
not I_3(I11412,I11395);
nor I_4(I8854,I9179,I9320);
DFFARX1 I_5(I9258,I1470,I8862,,,I8827,);
not I_6(I11830,I11813);
nand I_7(I11624,I11327,I8827);
nor I_8(I11576,I11559,I11412);
or I_9(I11895,I11830,I11641);
not I_10(I8862,I1477);
or I_11(I9258,I9179);
DFFARX1 I_12(I8854,I1470,I11310,,,I11813,);
not I_13(I11327,I8830);
not I_14(I11310,I1477);
endmodule


