module test_I11720(I1477,I1470,I9083,I8947,I11720);
input I1477,I1470,I9083,I8947;
output I11720;
wire I9320,I11672,I11429,I8836,I9303,I9210,I9179,I11460,I8848,I11310,I9413;
not I_0(I9320,I9303);
DFFARX1 I_1(I8836,I1470,I11310,,,I11672,);
not I_2(I11429,I8848);
nor I_3(I11720,I11672,I11460);
nand I_4(I8836,I9320,I9210);
DFFARX1 I_5(I1470,,,I9303,);
nor I_6(I9210,I9179,I8947);
DFFARX1 I_7(I1470,,,I9179,);
not I_8(I11460,I11429);
nor I_9(I8848,I9083,I9413);
not I_10(I11310,I1477);
and I_11(I9413,I8947);
endmodule


