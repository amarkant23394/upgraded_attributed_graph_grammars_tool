module test_I5481(I1477,I3521,I1470,I3572,I3685,I5481);
input I1477,I3521,I1470,I3572,I3685;
output I5481;
wire I5416,I3388,I3350,I5122,I3589,I3356,I5105;
nand I_0(I5416,I5122,I3356);
not I_1(I3388,I1477);
DFFARX1 I_2(I3685,I1470,I3388,,,I3350,);
not I_3(I5122,I3350);
and I_4(I3589,I3521,I3572);
DFFARX1 I_5(I3589,I1470,I3388,,,I3356,);
not I_6(I5105,I1477);
DFFARX1 I_7(I5416,I1470,I5105,,,I5481,);
endmodule


