module test_final(IN_1_0_l_1,IN_2_0_l_1,IN_3_0_l_1,IN_4_0_l_1,IN_1_1_l_1,IN_2_1_l_1,IN_3_1_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_3_3_l_1,IN_1_6_l_1,IN_2_6_l_1,IN_3_6_l_1,IN_4_6_l_1,IN_5_6_l_1,blif_clk_net_7_r_14,blif_reset_net_7_r_14,N1371_0_r_14,N1508_0_r_14,N1507_6_r_14,N1508_6_r_14,G42_7_r_14,n_572_7_r_14,n_573_7_r_14,n_549_7_r_14,n_569_7_r_14,n_452_7_r_14,N6147_9_r_14,N6134_9_r_14);
input IN_1_0_l_1,IN_2_0_l_1,IN_3_0_l_1,IN_4_0_l_1,IN_1_1_l_1,IN_2_1_l_1,IN_3_1_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_3_3_l_1,IN_1_6_l_1,IN_2_6_l_1,IN_3_6_l_1,IN_4_6_l_1,IN_5_6_l_1,blif_clk_net_7_r_14,blif_reset_net_7_r_14;
output N1371_0_r_14,N1508_0_r_14,N1507_6_r_14,N1508_6_r_14,G42_7_r_14,n_572_7_r_14,n_573_7_r_14,n_549_7_r_14,n_569_7_r_14,n_452_7_r_14,N6147_9_r_14,N6134_9_r_14;
wire N1371_0_r_1,N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,n_452_7_r_1,N6147_9_r_1,N6134_9_r_1,I_BUFF_1_9_r_1,n4_7_r_1,n29_1,n30_1,n31_1,n32_1,n33_1,n34_1,n35_1,n36_1,n37_1,n38_1,n39_1,n40_1,n41_1,n42_1,n43_1,n44_1,n45_1,n46_1,n47_1,n48_1,n49_1,n50_1,n51_1,n52_1,n53_1,n54_1,n55_1,I_BUFF_1_9_r_14,N3_8_l_14,n8_14,n47_14,n4_7_r_14,n26_14,n27_14,n28_14,n29_14,n30_14,n31_14,n32_14,n33_14,n34_14,n35_14,n36_14,n37_14,n38_14,n39_14,n40_14,n41_14,n42_14,n43_14,n44_14,n45_14,n46_14;
and I_0(N1371_0_r_1,I_BUFF_1_9_r_1,n55_1);
nor I_1(N1508_0_r_1,n40_1,n44_1);
nor I_2(N1507_6_r_1,n43_1,n49_1);
nor I_3(N1508_6_r_1,n41_1,n42_1);
DFFARX1 I_4(n4_7_r_1,blif_clk_net_7_r_14,n8_14,G42_7_r_1,);
nor I_5(n_572_7_r_1,n29_1,n30_1);
not I_6(n_573_7_r_1,n_452_7_r_1);
nor I_7(n_549_7_r_1,N1371_0_r_1,n31_1);
or I_8(n_569_7_r_1,n30_1,n31_1);
nor I_9(n_452_7_r_1,n30_1,n32_1);
nor I_10(N6147_9_r_1,n35_1,n36_1);
nand I_11(N6134_9_r_1,n38_1,n39_1);
not I_12(I_BUFF_1_9_r_1,n40_1);
nor I_13(n4_7_r_1,I_BUFF_1_9_r_1,n30_1);
nor I_14(n29_1,IN_2_0_l_1,n34_1);
nor I_15(n30_1,n33_1,n34_1);
nor I_16(n31_1,IN_1_3_l_1,n54_1);
not I_17(n32_1,n48_1);
nor I_18(n33_1,IN_3_0_l_1,IN_4_0_l_1);
not I_19(n34_1,IN_1_0_l_1);
nor I_20(n35_1,I_BUFF_1_9_r_1,n37_1);
not I_21(n36_1,n29_1);
not I_22(n37_1,n41_1);
nand I_23(n38_1,IN_3_1_l_1,I_BUFF_1_9_r_1);
nand I_24(n39_1,n37_1,n40_1);
nand I_25(n40_1,IN_1_1_l_1,IN_2_1_l_1);
nand I_26(n41_1,IN_5_6_l_1,n52_1);
or I_27(n42_1,n36_1,n43_1);
nor I_28(n43_1,n32_1,n49_1);
nand I_29(n44_1,n45_1,n46_1);
nand I_30(n45_1,n47_1,n48_1);
not I_31(n46_1,IN_3_1_l_1);
not I_32(n47_1,n31_1);
nand I_33(n48_1,IN_2_6_l_1,n50_1);
nor I_34(n49_1,n41_1,n47_1);
and I_35(n50_1,IN_1_6_l_1,n51_1);
nand I_36(n51_1,n52_1,n53_1);
nand I_37(n52_1,IN_3_6_l_1,IN_4_6_l_1);
not I_38(n53_1,IN_5_6_l_1);
or I_39(n54_1,IN_2_3_l_1,IN_3_3_l_1);
nor I_40(n55_1,IN_3_1_l_1,n29_1);
nor I_41(N1371_0_r_14,n47_14,n30_14);
nor I_42(N1508_0_r_14,n30_14,n41_14);
nor I_43(N1507_6_r_14,n37_14,n44_14);
nor I_44(N1508_6_r_14,n30_14,n39_14);
DFFARX1 I_45(n4_7_r_14,blif_clk_net_7_r_14,n8_14,G42_7_r_14,);
nor I_46(n_572_7_r_14,n28_14,n29_14);
nand I_47(n_573_7_r_14,n26_14,n27_14);
nor I_48(n_549_7_r_14,n31_14,n32_14);
nand I_49(n_569_7_r_14,n26_14,n30_14);
nor I_50(n_452_7_r_14,n47_14,n28_14);
nor I_51(N6147_9_r_14,n36_14,n37_14);
nor I_52(N6134_9_r_14,n28_14,n36_14);
not I_53(I_BUFF_1_9_r_14,n26_14);
and I_54(N3_8_l_14,n38_14,n_569_7_r_1);
not I_55(n8_14,blif_reset_net_7_r_14);
DFFARX1 I_56(N3_8_l_14,blif_clk_net_7_r_14,n8_14,n47_14,);
nor I_57(n4_7_r_14,n47_14,n35_14);
nand I_58(n26_14,n_573_7_r_1,N6147_9_r_1);
not I_59(n27_14,n28_14);
nor I_60(n28_14,n43_14,N1508_6_r_1);
not I_61(n29_14,n33_14);
not I_62(n30_14,n31_14);
nor I_63(n31_14,n46_14,n_549_7_r_1);
and I_64(n32_14,n33_14,n34_14);
nand I_65(n33_14,I_BUFF_1_9_r_14,n45_14);
nor I_66(n34_14,n42_14,n43_14);
nor I_67(n35_14,N1508_6_r_1,n_572_7_r_1);
nor I_68(n36_14,n47_14,n34_14);
not I_69(n37_14,n35_14);
nand I_70(n38_14,N1507_6_r_1,n_572_7_r_1);
nand I_71(n39_14,n29_14,n40_14);
nand I_72(n40_14,n27_14,n37_14);
nor I_73(n41_14,I_BUFF_1_9_r_14,n34_14);
nor I_74(n42_14,N6134_9_r_1,G42_7_r_1);
not I_75(n43_14,G42_7_r_1);
nor I_76(n44_14,n27_14,n33_14);
or I_77(n45_14,n_572_7_r_1,N1508_0_r_1);
or I_78(n46_14,N1508_0_r_1,N1507_6_r_1);
endmodule


