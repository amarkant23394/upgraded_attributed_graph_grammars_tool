module test_I3137(I2005,I2583,I1316,I1908,I1294,I2488,I2070,I1937,I2457,I1988,I3137);
input I2005,I2583,I1316,I1908,I1294,I2488,I2070,I1937,I2457,I1988;
output I3137;
wire I2668,I1911,I1914,I2313,I2022,I2897,I2600,I2344,I2651,I1920,I3120,I1923,I3086,I3103;
nand I_0(I2668,I2651,I1914);
nand I_1(I1911,I2070,I2488);
DFFARX1 I_2(I2457,I1294,I1937,,,I1914,);
DFFARX1 I_3(I1294,I1937,,,I2313,);
nand I_4(I2022,I2005,I1316);
nand I_5(I2897,I2600,I1923);
and I_6(I3137,I2897,I3120);
not I_7(I2600,I1911);
nor I_8(I2344,I2313,I1988);
nor I_9(I2651,I2600,I1908);
not I_10(I1920,I2313);
nand I_11(I3120,I3103,I2668);
nand I_12(I1923,I2022,I2344);
DFFARX1 I_13(I1920,I1294,I2583,,,I3086,);
not I_14(I3103,I3086);
endmodule


