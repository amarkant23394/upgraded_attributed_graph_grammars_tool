module test_I4509(I2167,I2170,I1477,I2557,I4962,I1470,I4509);
input I2167,I2170,I1477,I2557,I4962,I1470;
output I4509;
wire I4629,I4996,I4979,I2143,I2173,I2181,I4544,I5013,I4742,I4807,I4824;
nor I_0(I4629,I2167,I2173);
and I_1(I4996,I4629,I4979);
nor I_2(I4979,I4742,I4962);
DFFARX1 I_3(I2557,I1470,I2181,,,I2143,);
nand I_4(I2173,I2557);
not I_5(I2181,I1477);
not I_6(I4544,I1477);
or I_7(I5013,I4824,I4996);
DFFARX1 I_8(I1470,I4544,,,I4742,);
DFFARX1 I_9(I2170,I1470,I4544,,,I4807,);
and I_10(I4824,I4807,I2143);
DFFARX1 I_11(I5013,I1470,I4544,,,I4509,);
endmodule


