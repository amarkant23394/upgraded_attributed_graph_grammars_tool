module test_final(IN_1_2_l_2,IN_2_2_l_2,IN_3_2_l_2,IN_6_2_l_2,IN_1_3_l_2,IN_2_3_l_2,IN_4_3_l_2,IN_1_4_l_2,IN_2_4_l_2,IN_3_4_l_2,IN_6_4_l_2,blif_clk_net_1_r_9,blif_reset_net_1_r_9,G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9);
input IN_1_2_l_2,IN_2_2_l_2,IN_3_2_l_2,IN_6_2_l_2,IN_1_3_l_2,IN_2_3_l_2,IN_4_3_l_2,IN_1_4_l_2,IN_2_4_l_2,IN_3_4_l_2,IN_6_4_l_2,blif_clk_net_1_r_9,blif_reset_net_1_r_9;
output G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9;
wire G42_1_r_2,n_572_1_r_2,n_573_1_r_2,n_549_1_r_2,n_569_1_r_2,n_452_1_r_2,n_42_2_r_2,G199_2_r_2,ACVQN1_5_r_2,P6_5_r_2,N3_2_l_2,G199_2_l_2,n13_2,ACVQN2_3_l_2,n16_2,N1_4_l_2,n26_2,n17_internal_2,n17_2,n4_1_r_2,N3_2_r_2,P6_5_r_internal_2,n18_2,n19_2,n20_2,n21_2,n22_2,n23_2,n24_2,n25_2,n_452_1_r_9,N3_2_l_9,n5_9,n27_9,n16_9,n26_9,n15_9,n29_internal_9,n29_9,N1_4_l_9,n25_9,n28_internal_9,n28_9,n4_1_r_9,N3_2_r_9,N1_4_r_9,n_42_2_l_9,n17_9,n18_9,n19_9,n20_9,n21_9,n22_9,n23_9,n24_9;
DFFARX1 I_0(n4_1_r_2,blif_clk_net_1_r_9,n5_9,G42_1_r_2,);
nor I_1(n_572_1_r_2,n26_2,n18_2);
nand I_2(n_573_1_r_2,n17_2,n19_2);
nor I_3(n_549_1_r_2,G199_2_l_2,n20_2);
nand I_4(n_569_1_r_2,n13_2,n19_2);
not I_5(n_452_1_r_2,n_573_1_r_2);
nor I_6(n_42_2_r_2,ACVQN2_3_l_2,n18_2);
DFFARX1 I_7(N3_2_r_2,blif_clk_net_1_r_9,n5_9,G199_2_r_2,);
DFFARX1 I_8(ACVQN2_3_l_2,blif_clk_net_1_r_9,n5_9,ACVQN1_5_r_2,);
not I_9(P6_5_r_2,P6_5_r_internal_2);
and I_10(N3_2_l_2,IN_6_2_l_2,n24_2);
DFFARX1 I_11(N3_2_l_2,blif_clk_net_1_r_9,n5_9,G199_2_l_2,);
not I_12(n13_2,G199_2_l_2);
DFFARX1 I_13(IN_1_3_l_2,blif_clk_net_1_r_9,n5_9,ACVQN2_3_l_2,);
DFFARX1 I_14(IN_2_3_l_2,blif_clk_net_1_r_9,n5_9,n16_2,);
and I_15(N1_4_l_2,IN_6_4_l_2,n25_2);
DFFARX1 I_16(N1_4_l_2,blif_clk_net_1_r_9,n5_9,n26_2,);
DFFARX1 I_17(IN_3_4_l_2,blif_clk_net_1_r_9,n5_9,n17_internal_2,);
not I_18(n17_2,n17_internal_2);
nor I_19(n4_1_r_2,n26_2,n22_2);
nor I_20(N3_2_r_2,n17_2,n23_2);
DFFARX1 I_21(G199_2_l_2,blif_clk_net_1_r_9,n5_9,P6_5_r_internal_2,);
nor I_22(n18_2,IN_1_2_l_2,IN_3_2_l_2);
nand I_23(n19_2,IN_4_3_l_2,n16_2);
nor I_24(n20_2,n26_2,n21_2);
not I_25(n21_2,n18_2);
and I_26(n22_2,IN_4_3_l_2,n16_2);
nor I_27(n23_2,n13_2,n21_2);
nand I_28(n24_2,IN_2_2_l_2,IN_3_2_l_2);
nand I_29(n25_2,IN_1_4_l_2,IN_2_4_l_2);
DFFARX1 I_30(n4_1_r_9,blif_clk_net_1_r_9,n5_9,G42_1_r_9,);
nor I_31(n_572_1_r_9,n27_9,n_42_2_l_9);
or I_32(n_573_1_r_9,n25_9,n_42_2_l_9);
nand I_33(n_549_1_r_9,n17_9,n18_9);
or I_34(n_569_1_r_9,n26_9,n_42_2_l_9);
nor I_35(n_452_1_r_9,n26_9,n25_9);
nor I_36(n_42_2_r_9,n25_9,n19_9);
DFFARX1 I_37(N3_2_r_9,blif_clk_net_1_r_9,n5_9,G199_2_r_9,);
DFFARX1 I_38(N1_4_r_9,blif_clk_net_1_r_9,n5_9,G199_4_r_9,);
DFFARX1 I_39(n_42_2_l_9,blif_clk_net_1_r_9,n5_9,G214_4_r_9,);
and I_40(N3_2_l_9,n22_9,n_549_1_r_2);
not I_41(n5_9,blif_reset_net_1_r_9);
DFFARX1 I_42(N3_2_l_9,blif_clk_net_1_r_9,n5_9,n27_9,);
not I_43(n16_9,n27_9);
DFFARX1 I_44(n_569_1_r_2,blif_clk_net_1_r_9,n5_9,n26_9,);
not I_45(n15_9,n26_9);
DFFARX1 I_46(G199_2_r_2,blif_clk_net_1_r_9,n5_9,n29_internal_9,);
not I_47(n29_9,n29_internal_9);
and I_48(N1_4_l_9,n24_9,G42_1_r_2);
DFFARX1 I_49(N1_4_l_9,blif_clk_net_1_r_9,n5_9,n25_9,);
DFFARX1 I_50(n_572_1_r_2,blif_clk_net_1_r_9,n5_9,n28_internal_9,);
not I_51(n28_9,n28_internal_9);
nor I_52(n4_1_r_9,n27_9,n26_9);
nor I_53(N3_2_r_9,n15_9,n21_9);
nor I_54(N1_4_r_9,n16_9,n21_9);
nor I_55(n_42_2_l_9,n_42_2_r_2,G42_1_r_2);
not I_56(n17_9,n_452_1_r_9);
nand I_57(n18_9,n27_9,n15_9);
nor I_58(n19_9,n29_9,n20_9);
not I_59(n20_9,n_572_1_r_2);
and I_60(n21_9,n23_9,n_572_1_r_2);
nand I_61(n22_9,P6_5_r_2,G42_1_r_2);
nor I_62(n23_9,n29_9,n28_9);
nand I_63(n24_9,n_452_1_r_2,ACVQN1_5_r_2);
endmodule


