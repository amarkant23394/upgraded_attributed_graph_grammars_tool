module test_final(IN_1_0_l_14,IN_2_0_l_14,IN_4_0_l_14,IN_1_1_l_14,IN_2_1_l_14,IN_3_1_l_14,IN_6_1_l_14,IN_1_5_l_14,IN_2_5_l_14,IN_3_5_l_14,IN_6_5_l_14,blif_reset_net_0_r_6,blif_clk_net_0_r_6,ACVQN2_0_r_6,n_266_and_0_0_r_6,ACVQN1_2_r_6,P6_2_r_6,n_429_or_0_3_r_6,G78_3_r_6,n_576_3_r_6,n_102_3_r_6,n_547_3_r_6,n_42_5_r_6,G199_5_r_6);
input IN_1_0_l_14,IN_2_0_l_14,IN_4_0_l_14,IN_1_1_l_14,IN_2_1_l_14,IN_3_1_l_14,IN_6_1_l_14,IN_1_5_l_14,IN_2_5_l_14,IN_3_5_l_14,IN_6_5_l_14,blif_reset_net_0_r_6,blif_clk_net_0_r_6;
output ACVQN2_0_r_6,n_266_and_0_0_r_6,ACVQN1_2_r_6,P6_2_r_6,n_429_or_0_3_r_6,G78_3_r_6,n_576_3_r_6,n_102_3_r_6,n_547_3_r_6,n_42_5_r_6,G199_5_r_6;
wire ACVQN2_0_r_14,n_266_and_0_0_r_14,G199_1_r_14,G214_1_r_14,ACVQN1_2_r_14,P6_2_r_14,n_429_or_0_3_r_14,G78_3_r_14,n_576_3_r_14,n_102_3_r_14,n_547_3_r_14,ACVQN2_0_l_14,n_266_and_0_0_l_14,ACVQN1_0_l_14,N1_1_l_14,G199_1_l_14,G214_1_l_14,n3_1_l_14,n_42_5_l_14,N3_5_l_14,G199_5_l_14,n3_5_l_14,ACVQN1_0_r_14,N1_1_r_14,n3_1_r_14,P6_internal_2_r_14,n12_3_r_14,n_431_3_r_14,n11_3_r_14,n13_3_r_14,n14_3_r_14,n15_3_r_14,n16_3_r_14,n1_0_r_6,ACVQN1_2_l_6,P6_2_l_6,P6_internal_2_l_6,n_429_or_0_3_l_6,n12_3_l_6,n_431_3_l_6,G78_3_l_6,n_576_3_l_6,n11_3_l_6,n_102_3_l_6,n_547_3_l_6,n13_3_l_6,n14_3_l_6,n15_3_l_6,n16_3_l_6,ACVQN1_0_r_6,P6_internal_2_r_6,n12_3_r_6,n_431_3_r_6,n11_3_r_6,n13_3_r_6,n14_3_r_6,n15_3_r_6,n16_3_r_6,N3_5_r_6,n3_5_r_6;
DFFARX1 I_0(n_266_and_0_0_l_14,blif_clk_net_0_r_6,n1_0_r_6,ACVQN2_0_r_14,);
and I_1(n_266_and_0_0_r_14,G199_5_l_14,ACVQN1_0_r_14);
DFFARX1 I_2(N1_1_r_14,blif_clk_net_0_r_6,n1_0_r_6,G199_1_r_14,);
DFFARX1 I_3(G199_1_l_14,blif_clk_net_0_r_6,n1_0_r_6,G214_1_r_14,);
DFFARX1 I_4(ACVQN2_0_l_14,blif_clk_net_0_r_6,n1_0_r_6,ACVQN1_2_r_14,);
not I_5(P6_2_r_14,P6_internal_2_r_14);
nand I_6(n_429_or_0_3_r_14,G214_1_l_14,n12_3_r_14);
DFFARX1 I_7(n_431_3_r_14,blif_clk_net_0_r_6,n1_0_r_6,G78_3_r_14,);
nand I_8(n_576_3_r_14,ACVQN2_0_l_14,n11_3_r_14);
not I_9(n_102_3_r_14,G199_5_l_14);
nand I_10(n_547_3_r_14,n_266_and_0_0_l_14,n13_3_r_14);
DFFARX1 I_11(IN_1_0_l_14,blif_clk_net_0_r_6,n1_0_r_6,ACVQN2_0_l_14,);
and I_12(n_266_and_0_0_l_14,IN_4_0_l_14,ACVQN1_0_l_14);
DFFARX1 I_13(IN_2_0_l_14,blif_clk_net_0_r_6,n1_0_r_6,ACVQN1_0_l_14,);
and I_14(N1_1_l_14,IN_6_1_l_14,n3_1_l_14);
DFFARX1 I_15(N1_1_l_14,blif_clk_net_0_r_6,n1_0_r_6,G199_1_l_14,);
DFFARX1 I_16(IN_3_1_l_14,blif_clk_net_0_r_6,n1_0_r_6,G214_1_l_14,);
nand I_17(n3_1_l_14,IN_1_1_l_14,IN_2_1_l_14);
nor I_18(n_42_5_l_14,IN_1_5_l_14,IN_3_5_l_14);
and I_19(N3_5_l_14,IN_6_5_l_14,n3_5_l_14);
DFFARX1 I_20(N3_5_l_14,blif_clk_net_0_r_6,n1_0_r_6,G199_5_l_14,);
nand I_21(n3_5_l_14,IN_2_5_l_14,IN_3_5_l_14);
DFFARX1 I_22(G214_1_l_14,blif_clk_net_0_r_6,n1_0_r_6,ACVQN1_0_r_14,);
and I_23(N1_1_r_14,G214_1_l_14,n3_1_r_14);
nand I_24(n3_1_r_14,ACVQN2_0_l_14,n_42_5_l_14);
DFFARX1 I_25(G199_5_l_14,blif_clk_net_0_r_6,n1_0_r_6,P6_internal_2_r_14,);
not I_26(n12_3_r_14,n_42_5_l_14);
or I_27(n_431_3_r_14,n_266_and_0_0_l_14,n14_3_r_14);
nor I_28(n11_3_r_14,G199_5_l_14,n12_3_r_14);
nor I_29(n13_3_r_14,G199_1_l_14,G199_5_l_14);
and I_30(n14_3_r_14,n_42_5_l_14,n15_3_r_14);
nor I_31(n15_3_r_14,G199_1_l_14,n16_3_r_14);
not I_32(n16_3_r_14,G214_1_l_14);
DFFARX1 I_33(G78_3_l_6,blif_clk_net_0_r_6,n1_0_r_6,ACVQN2_0_r_6,);
and I_34(n_266_and_0_0_r_6,n_429_or_0_3_l_6,ACVQN1_0_r_6);
DFFARX1 I_35(G78_3_l_6,blif_clk_net_0_r_6,n1_0_r_6,ACVQN1_2_r_6,);
not I_36(P6_2_r_6,P6_internal_2_r_6);
nand I_37(n_429_or_0_3_r_6,n_102_3_l_6,n12_3_r_6);
DFFARX1 I_38(n_431_3_r_6,blif_clk_net_0_r_6,n1_0_r_6,G78_3_r_6,);
nand I_39(n_576_3_r_6,P6_2_l_6,n11_3_r_6);
not I_40(n_102_3_r_6,ACVQN1_2_l_6);
nand I_41(n_547_3_r_6,n_576_3_l_6,n13_3_r_6);
nor I_42(n_42_5_r_6,ACVQN1_2_l_6,n_429_or_0_3_l_6);
DFFARX1 I_43(N3_5_r_6,blif_clk_net_0_r_6,n1_0_r_6,G199_5_r_6,);
not I_44(n1_0_r_6,blif_reset_net_0_r_6);
DFFARX1 I_45(n_102_3_r_14,blif_clk_net_0_r_6,n1_0_r_6,ACVQN1_2_l_6,);
not I_46(P6_2_l_6,P6_internal_2_l_6);
DFFARX1 I_47(ACVQN1_2_r_14,blif_clk_net_0_r_6,n1_0_r_6,P6_internal_2_l_6,);
nand I_48(n_429_or_0_3_l_6,n12_3_l_6,n_547_3_r_14);
not I_49(n12_3_l_6,n_429_or_0_3_r_14);
or I_50(n_431_3_l_6,n14_3_l_6,ACVQN2_0_r_14);
DFFARX1 I_51(n_431_3_l_6,blif_clk_net_0_r_6,n1_0_r_6,G78_3_l_6,);
nand I_52(n_576_3_l_6,n11_3_l_6,P6_2_r_14);
nor I_53(n11_3_l_6,n12_3_l_6,n_266_and_0_0_r_14);
not I_54(n_102_3_l_6,n_266_and_0_0_r_14);
nand I_55(n_547_3_l_6,n13_3_l_6,G199_1_r_14);
nor I_56(n13_3_l_6,n_266_and_0_0_r_14,G214_1_r_14);
and I_57(n14_3_l_6,n15_3_l_6,G78_3_r_14);
nor I_58(n15_3_l_6,n16_3_l_6,n_576_3_r_14);
not I_59(n16_3_l_6,n_547_3_r_14);
DFFARX1 I_60(G78_3_l_6,blif_clk_net_0_r_6,n1_0_r_6,ACVQN1_0_r_6,);
DFFARX1 I_61(n_576_3_l_6,blif_clk_net_0_r_6,n1_0_r_6,P6_internal_2_r_6,);
not I_62(n12_3_r_6,P6_2_l_6);
or I_63(n_431_3_r_6,n_429_or_0_3_l_6,n14_3_r_6);
nor I_64(n11_3_r_6,ACVQN1_2_l_6,n12_3_r_6);
nor I_65(n13_3_r_6,ACVQN1_2_l_6,n_547_3_l_6);
and I_66(n14_3_r_6,ACVQN1_2_l_6,n15_3_r_6);
nor I_67(n15_3_r_6,P6_2_l_6,n16_3_r_6);
not I_68(n16_3_r_6,n_102_3_l_6);
and I_69(N3_5_r_6,n_102_3_l_6,n3_5_r_6);
nand I_70(n3_5_r_6,n_429_or_0_3_l_6,n_547_3_l_6);
endmodule


