module test_I14356(I13183,I1477,I14387,I13296,I13618,I1470,I14356);
input I13183,I1477,I14387,I13296,I13618,I1470;
output I14356;
wire I14667,I14856,I14421,I14650,I13165,I14808,I14370,I13162,I13197,I13635,I13248,I13361,I13189,I14404;
and I_0(I14667,I14650,I13189);
nor I_1(I14856,I14808,I14421);
DFFARX1 I_2(I14404,I1470,I14370,,,I14421,);
DFFARX1 I_3(I13165,I1470,I14370,,,I14650,);
DFFARX1 I_4(I13248,I1470,I13197,,,I13165,);
nand I_5(I14356,I14667,I14856);
DFFARX1 I_6(I13162,I1470,I14370,,,I14808,);
not I_7(I14370,I1477);
and I_8(I13162,I13248,I13361);
not I_9(I13197,I1477);
and I_10(I13635,I13296,I13618);
DFFARX1 I_11(I1470,I13197,,,I13248,);
DFFARX1 I_12(I1470,I13197,,,I13361,);
DFFARX1 I_13(I13635,I1470,I13197,,,I13189,);
and I_14(I14404,I14387,I13183);
endmodule


