module test_I2121(I1215,I1294,I1492,I1301,I2121);
input I1215,I1294,I1492,I1301;
output I2121;
wire I1325,I2104,I1342,I1509,I1304,I1780;
not I_0(I1325,I1780);
not I_1(I2104,I1304);
nor I_2(I2121,I2104,I1325);
not I_3(I1342,I1301);
DFFARX1 I_4(I1492,I1294,I1342,,,I1509,);
DFFARX1 I_5(I1509,I1294,I1342,,,I1304,);
DFFARX1 I_6(I1215,I1294,I1342,,,I1780,);
endmodule


