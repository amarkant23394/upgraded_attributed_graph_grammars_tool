module test_I1342(I1301,I1342);
input I1301;
output I1342;
wire ;
not I_0(I1342,I1301);
endmodule


