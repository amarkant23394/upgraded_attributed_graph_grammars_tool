module test_I11973_rst(I1477_rst,I11973_rst);
,I11973_rst);
input I1477_rst;
output I11973_rst;
wire ;
not I_0(I11973_rst,I1477_rst);
endmodule


