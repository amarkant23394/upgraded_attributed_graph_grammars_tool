module test_final(IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_4_l_4,IN_2_4_l_4,IN_3_4_l_4,IN_4_4_l_4,IN_5_4_l_4,IN_1_9_l_4,IN_2_9_l_4,IN_3_9_l_4,IN_4_9_l_4,IN_5_9_l_4,blif_clk_net_5_r_13,blif_reset_net_5_r_13,N1371_0_r_13,N1508_0_r_13,n_429_or_0_5_r_13,G78_5_r_13,n_576_5_r_13,n_547_5_r_13,G42_7_r_13,n_572_7_r_13,n_573_7_r_13,n_549_7_r_13,n_569_7_r_13,n_452_7_r_13);
input IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_4_l_4,IN_2_4_l_4,IN_3_4_l_4,IN_4_4_l_4,IN_5_4_l_4,IN_1_9_l_4,IN_2_9_l_4,IN_3_9_l_4,IN_4_9_l_4,IN_5_9_l_4,blif_clk_net_5_r_13,blif_reset_net_5_r_13;
output N1371_0_r_13,N1508_0_r_13,n_429_or_0_5_r_13,G78_5_r_13,n_576_5_r_13,n_547_5_r_13,G42_7_r_13,n_572_7_r_13,n_573_7_r_13,n_549_7_r_13,n_569_7_r_13,n_452_7_r_13;
wire N1371_0_r_4,N1508_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_573_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6147_9_r_4,N6134_9_r_4,I_BUFF_1_9_r_4,n4_7_r_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4,n38_4,n39_4,n40_4,n41_4,n_102_5_r_13,n4_7_l_13,n9_13,n62_13,n33_13,n_431_5_r_13,n1_13,n34_13,n35_13,n36_13,n37_13,n38_13,n39_13,n40_13,n41_13,n42_13,n43_13,n44_13,n45_13,n46_13,n47_13,n48_13,n49_13,n50_13,n51_13,n52_13,n53_13,n54_13,n55_13,n56_13,n57_13,n58_13,n59_13,n60_13,n61_13;
nor I_0(N1371_0_r_4,IN_1_9_l_4,n25_4);
not I_1(N1508_0_r_4,n25_4);
nor I_2(N1507_6_r_4,n32_4,n33_4);
nor I_3(N1508_6_r_4,n22_4,n29_4);
DFFARX1 I_4(n4_7_r_4,blif_clk_net_5_r_13,n9_13,G42_7_r_4,);
not I_5(n_572_7_r_4,n_573_7_r_4);
nand I_6(n_573_7_r_4,n21_4,n22_4);
nor I_7(n_549_7_r_4,IN_1_9_l_4,n24_4);
nand I_8(n_569_7_r_4,n22_4,n23_4);
nor I_9(n_452_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4);
not I_10(N6147_9_r_4,n28_4);
nor I_11(N6134_9_r_4,N1508_0_r_4,n28_4);
not I_12(I_BUFF_1_9_r_4,n21_4);
nor I_13(n4_7_r_4,IN_1_9_l_4,N6147_9_r_4);
nand I_14(n21_4,n39_4,n40_4);
or I_15(n22_4,IN_5_9_l_4,n31_4);
not I_16(n23_4,IN_1_9_l_4);
nor I_17(n24_4,n25_4,n26_4);
nand I_18(n25_4,IN_1_4_l_4,IN_2_4_l_4);
nand I_19(n26_4,n21_4,n27_4);
nand I_20(n27_4,n36_4,n37_4);
nand I_21(n28_4,IN_2_9_l_4,n38_4);
nand I_22(n29_4,N1508_0_r_4,n30_4);
nand I_23(n30_4,n34_4,n35_4);
nor I_24(n31_4,IN_3_9_l_4,IN_4_9_l_4);
not I_25(n32_4,n30_4);
nor I_26(n33_4,n21_4,n28_4);
nand I_27(n34_4,N6147_9_r_4,I_BUFF_1_9_r_4);
nand I_28(n35_4,N1508_0_r_4,n27_4);
not I_29(n36_4,IN_5_4_l_4);
nand I_30(n37_4,IN_3_4_l_4,IN_4_4_l_4);
or I_31(n38_4,IN_3_9_l_4,IN_4_9_l_4);
nor I_32(n39_4,IN_1_2_l_4,IN_2_2_l_4);
or I_33(n40_4,IN_5_2_l_4,n41_4);
nor I_34(n41_4,IN_3_2_l_4,IN_4_2_l_4);
nor I_35(N1371_0_r_13,n59_13,n61_13);
nor I_36(N1508_0_r_13,n59_13,n60_13);
not I_37(n_429_or_0_5_r_13,n46_13);
DFFARX1 I_38(n_431_5_r_13,blif_clk_net_5_r_13,n9_13,G78_5_r_13,);
nand I_39(n_576_5_r_13,n_102_5_r_13,n34_13);
nor I_40(n_102_5_r_13,N1371_0_r_4,n_572_7_r_4);
nand I_41(n_547_5_r_13,n48_13,n49_13);
DFFARX1 I_42(n1_13,blif_clk_net_5_r_13,n9_13,G42_7_r_13,);
nor I_43(n_572_7_r_13,n40_13,n41_13);
nand I_44(n_573_7_r_13,n37_13,n38_13);
nor I_45(n_549_7_r_13,n46_13,n47_13);
nand I_46(n_569_7_r_13,n37_13,n43_13);
nand I_47(n_452_7_r_13,n52_13,n53_13);
nor I_48(n4_7_l_13,n_549_7_r_4,n_569_7_r_4);
not I_49(n9_13,blif_reset_net_5_r_13);
DFFARX1 I_50(n4_7_l_13,blif_clk_net_5_r_13,n9_13,n62_13,);
not I_51(n33_13,n62_13);
nand I_52(n_431_5_r_13,n54_13,n55_13);
not I_53(n1_13,n52_13);
nor I_54(n34_13,n35_13,n36_13);
nor I_55(n35_13,n42_13,n_572_7_r_4);
nand I_56(n36_13,n50_13,n58_13);
nand I_57(n37_13,n44_13,n45_13);
or I_58(n38_13,n39_13,N1507_6_r_4);
nand I_59(n39_13,G42_7_r_4,n_569_7_r_4);
not I_60(n40_13,n36_13);
nor I_61(n41_13,n35_13,n_572_7_r_4);
not I_62(n42_13,n_452_7_r_4);
or I_63(n43_13,N1507_6_r_4,n_549_7_r_4);
not I_64(n44_13,n_572_7_r_4);
not I_65(n45_13,n_549_7_r_4);
nor I_66(n46_13,n39_13,n40_13);
nor I_67(n47_13,N1507_6_r_4,n_549_7_r_4);
nor I_68(n48_13,n50_13,n51_13);
nor I_69(n49_13,n_572_7_r_4,n_549_7_r_4);
not I_70(n50_13,n59_13);
not I_71(n51_13,n_102_5_r_13);
nand I_72(n52_13,n33_13,n39_13);
nand I_73(n53_13,n33_13,N1507_6_r_4);
nor I_74(n54_13,N1371_0_r_4,N1507_6_r_4);
nand I_75(n55_13,n62_13,n56_13);
nor I_76(n56_13,n39_13,n57_13);
not I_77(n57_13,n_549_7_r_4);
or I_78(n58_13,N6134_9_r_4,N1371_0_r_4);
nand I_79(n59_13,N1508_6_r_4,G42_7_r_4);
nor I_80(n60_13,n51_13,N1507_6_r_4);
nor I_81(n61_13,n39_13,N1507_6_r_4);
endmodule


