module test_I13183(I11296,I1477,I11281,I8848,I13392,I8851,I1470,I13183);
input I11296,I1477,I11281,I8848,I13392,I8851,I1470;
output I13183;
wire I11768,I13525,I13601,I11395,I13197,I11299,I11378,I11429,I13426,I11272,I13508,I13491,I11310,I13409;
nand I_0(I13183,I13601,I13525);
and I_1(I11768,I11429);
nor I_2(I13525,I13508,I13426);
DFFARX1 I_3(I11299,I1470,I13197,,,I13601,);
nand I_4(I11395,I11378,I8851);
not I_5(I13197,I1477);
nor I_6(I11299,I11395,I11429);
nor I_7(I11378,I8848);
not I_8(I11429,I8848);
DFFARX1 I_9(I13409,I1470,I13197,,,I13426,);
DFFARX1 I_10(I11768,I1470,I11310,,,I11272,);
and I_11(I13508,I13491,I11272);
DFFARX1 I_12(I11296,I1470,I13197,,,I13491,);
not I_13(I11310,I1477);
and I_14(I13409,I13392,I11281);
endmodule


