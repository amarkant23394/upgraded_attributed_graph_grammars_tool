module test_final(IN_1_1_l_0,IN_2_1_l_0,IN_3_1_l_0,IN_1_8_l_0,IN_2_8_l_0,IN_3_8_l_0,IN_6_8_l_0,IN_1_10_l_0,IN_2_10_l_0,IN_3_10_l_0,IN_4_10_l_0,blif_clk_net_5_r_6,blif_reset_net_5_r_6,N1371_0_r_6,N1508_0_r_6,N6147_3_r_6,G78_5_r_6,n_576_5_r_6,n_547_5_r_6,N1372_10_r_6,N1508_10_r_6);
input IN_1_1_l_0,IN_2_1_l_0,IN_3_1_l_0,IN_1_8_l_0,IN_2_8_l_0,IN_3_8_l_0,IN_6_8_l_0,IN_1_10_l_0,IN_2_10_l_0,IN_3_10_l_0,IN_4_10_l_0,blif_clk_net_5_r_6,blif_reset_net_5_r_6;
output N1371_0_r_6,N1508_0_r_6,N6147_3_r_6,G78_5_r_6,n_576_5_r_6,n_547_5_r_6,N1372_10_r_6,N1508_10_r_6;
wire N1371_0_r_0,N1508_0_r_0,N6147_2_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_102_5_r_0,n_547_5_r_0,N1507_6_r_0,N1508_6_r_0,N3_8_l_0,n40_0,n4_0,n23_0,n24_0,n25_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0,n37_0,n38_0,n39_0,n_429_or_0_5_r_6,n_102_5_r_6,n_431_5_r_6,n6_6,n24_6,n25_6,n26_6,n27_6,n28_6,n29_6,n30_6,n31_6,n32_6,n33_6,n34_6,n35_6,n36_6,n37_6,n38_6,n39_6,n40_6,n41_6,n42_6;
nor I_0(N1371_0_r_0,n24_0,n25_0);
not I_1(N1508_0_r_0,n25_0);
nor I_2(N6147_2_r_0,n28_0,n29_0);
nand I_3(n_429_or_0_5_r_0,n4_0,n25_0);
DFFARX1 I_4(n4_0,blif_clk_net_5_r_6,n6_6,G78_5_r_0,);
nand I_5(n_576_5_r_0,n23_0,n24_0);
not I_6(n_102_5_r_0,n40_0);
nand I_7(n_547_5_r_0,n26_0,n27_0);
nor I_8(N1507_6_r_0,n_102_5_r_0,n37_0);
nor I_9(N1508_6_r_0,n25_0,n33_0);
and I_10(N3_8_l_0,IN_6_8_l_0,n32_0);
DFFARX1 I_11(N3_8_l_0,blif_clk_net_5_r_6,n6_6,n40_0,);
not I_12(n4_0,n31_0);
nor I_13(n23_0,n40_0,n25_0);
and I_14(n24_0,n4_0,n39_0);
nand I_15(n25_0,IN_1_1_l_0,IN_2_1_l_0);
nor I_16(n26_0,n40_0,n24_0);
nor I_17(n27_0,IN_1_8_l_0,IN_3_8_l_0);
nor I_18(n28_0,IN_3_1_l_0,n25_0);
nand I_19(n29_0,n_102_5_r_0,n30_0);
nand I_20(n30_0,n27_0,n31_0);
nand I_21(n31_0,IN_1_10_l_0,IN_2_10_l_0);
nand I_22(n32_0,IN_2_8_l_0,IN_3_8_l_0);
nand I_23(n33_0,n34_0,n35_0);
nand I_24(n34_0,n_102_5_r_0,n36_0);
not I_25(n35_0,IN_3_1_l_0);
not I_26(n36_0,n27_0);
nor I_27(n37_0,n36_0,n38_0);
nand I_28(n38_0,N1508_0_r_0,n35_0);
or I_29(n39_0,IN_3_10_l_0,IN_4_10_l_0);
nor I_30(N1371_0_r_6,n26_6,n38_6);
not I_31(N1508_0_r_6,n38_6);
nor I_32(N6147_3_r_6,n30_6,n35_6);
nand I_33(n_429_or_0_5_r_6,n30_6,n32_6);
DFFARX1 I_34(n_431_5_r_6,blif_clk_net_5_r_6,n6_6,G78_5_r_6,);
nand I_35(n_576_5_r_6,n24_6,n25_6);
not I_36(n_102_5_r_6,n26_6);
or I_37(n_547_5_r_6,n_429_or_0_5_r_6,n26_6);
not I_38(N1372_10_r_6,n37_6);
nor I_39(N1508_10_r_6,n36_6,n37_6);
nand I_40(n_431_5_r_6,n_102_5_r_6,n28_6);
not I_41(n6_6,blif_reset_net_5_r_6);
nor I_42(n24_6,n33_6,n34_6);
nor I_43(n25_6,n26_6,n27_6);
nor I_44(n26_6,n40_6,N1371_0_r_0);
nand I_45(n27_6,G78_5_r_0,n_429_or_0_5_r_0);
nand I_46(n28_6,n29_6,n30_6);
nor I_47(n29_6,n31_6,N6147_2_r_0);
not I_48(n30_6,n27_6);
nor I_49(n31_6,n39_6,n40_6);
nor I_50(n32_6,n24_6,N6147_2_r_0);
not I_51(n33_6,n_429_or_0_5_r_0);
not I_52(n34_6,n_547_5_r_0);
or I_53(n35_6,n26_6,n31_6);
and I_54(n36_6,n38_6,N6147_2_r_0);
nand I_55(n37_6,n30_6,n31_6);
nand I_56(n38_6,n41_6,n_547_5_r_0);
nor I_57(n39_6,N1507_6_r_0,N1508_6_r_0);
not I_58(n40_6,n_576_5_r_0);
nor I_59(n41_6,n33_6,n42_6);
nor I_60(n42_6,N6147_2_r_0,N1371_0_r_0);
endmodule


