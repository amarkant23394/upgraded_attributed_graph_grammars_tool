module test_I9720(I8479,I8753,I1477,I8196,I1470,I9720);
input I8479,I8753,I1477,I8196,I1470;
output I9720;
wire I9491,I9655,I9689,I8190,I9672,I8208;
not I_0(I9491,I1477);
not I_1(I9720,I9689);
nand I_2(I9655,I8190,I8196);
DFFARX1 I_3(I9672,I1470,I9491,,,I9689,);
DFFARX1 I_4(I1470,,,I8190,);
and I_5(I9672,I9655,I8208);
nand I_6(I8208,I8753,I8479);
endmodule


