module test_I17321(I14951,I15064,I1477,I15276,I1470,I15502,I17321);
input I14951,I15064,I1477,I15276,I1470,I15502;
output I17321;
wire I14927,I14948,I14954,I15310,I14965,I17304,I14933,I17205,I17092,I16818,I17109,I17287,I15293,I17270,I16886;
DFFARX1 I_0(I15502,I1470,I14965,,,I14927,);
or I_1(I17321,I17109,I17304);
DFFARX1 I_2(I1470,I14965,,,I14948,);
not I_3(I14954,I15064);
and I_4(I15310,I15276,I15293);
not I_5(I14965,I1477);
and I_6(I17304,I17205,I17287);
DFFARX1 I_7(I15310,I1470,I14965,,,I14933,);
DFFARX1 I_8(I14927,I1470,I16818,,,I17205,);
DFFARX1 I_9(I14954,I1470,I16818,,,I17092,);
not I_10(I16818,I1477);
and I_11(I17109,I17092,I14933);
nor I_12(I17287,I16886,I17270);
nand I_13(I15293,I15276);
not I_14(I17270,I17205);
nor I_15(I16886,I14951,I14948);
endmodule


