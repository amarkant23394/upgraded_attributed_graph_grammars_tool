module Benchmark_rules100(I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1294,I1301,I3186,I3201,I3183,I3198,I3180,I3177,I3192,I3189,I3195,I3204,I3174);
input I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1294,I1301;
output I3186,I3201,I3183,I3198,I3180,I3177,I3192,I3189,I3195,I3204,I3174;
wire I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1294,I1301,I1342,I1359,I1376,I1393,I1410,I1427,I1444,I1461,I1478,I1495,I1512,I1529,I1546,I1563,I1331,I1594,I1611,I1628,I1304,I1659,I1325,I1690,I1707,I1310,I1738,I1307,I1313,I1783,I1800,I1817,I1319,I1334,I1322,I1876,I1893,I1328,I1316,I1971,I1988,I2005,I2022,I1960,I2053,I1948,I2084,I2101,I2118,I2135,I2152,I1951,I2183,I1936,I2214,I2231,I2248,I2265,I2282,I2299,I1942,I2330,I2347,I2364,I1954,I1963,I1933,I2423,I1957,I1945,I2468,I2485,I1939,I2549,I2566,I2583,I2600,I2520,I2631,I2648,I2665,I2682,I2699,I2716,I2733,I2750,I2767,I2784,I2535,I2532,I2829,I2517,I2860,I2514,I2891,I2908,I2925,I2942,I2959,I2976,I2541,I3007,I2529,I2523,I3052,I3069,I2538,I3100,I3117,I3134,I2526,I2511,I3212,I3229,I3246,I3263,I3294,I3311,I3356,I3373,I3390,I3407,I3424,I3441,I3458,I3475,I3492,I3523,I3540,I3557,I3588,I3619,I3636,I3653,I3670,I3701,I3732,I3749,I3766;
not I_0 (I1342,I1301);
not I_1 (I1359,I1247);
nor I_2 (I1376,I1207,I1239);
nand I_3 (I1393,I1376,I1223);
nor I_4 (I1410,I1359,I1207);
nand I_5 (I1427,I1410,I1279);
not I_6 (I1444,I1207);
not I_7 (I1461,I1444);
not I_8 (I1478,I1215);
nor I_9 (I1495,I1478,I1255);
and I_10 (I1512,I1495,I1263);
or I_11 (I1529,I1512,I1287);
dffarx1 I_12 (I1546,I1529,I1294,I1342);
nand I_13 (I1563,I1359,I1215);
or I_14 (I1331,I1563,I1546);
not I_15 (I1594,I1563);
nor I_16 (I1611,I1546,I1594);
and I_17 (I1628,I1444,I1611);
nand I_18 (I1304,I1563,I1461);
dffarx1 I_19 (I1659,I1231,I1294,I1342);
or I_20 (I1325,I1659,I1546);
nor I_21 (I1690,I1659,I1427);
nor I_22 (I1707,I1659,I1461);
nand I_23 (I1310,I1393,I1707);
or I_24 (I1738,I1659,I1628);
dffarx1 I_25 (I1307,I1738,I1294,I1342);
not I_26 (I1313,I1659);
dffarx1 I_27 (I1783,I1271,I1294,I1342);
not I_28 (I1800,I1783);
nor I_29 (I1817,I1800,I1393);
dffarx1 I_30 (I1319,I1817,I1294,I1342);
nor I_31 (I1334,I1659,I1800);
nor I_32 (I1322,I1800,I1563);
not I_33 (I1876,I1800);
and I_34 (I1893,I1427,I1876);
nor I_35 (I1328,I1563,I1893);
nand I_36 (I1316,I1800,I1690);
not I_37 (I1971,I1301);
nand I_38 (I1988,I1307,I1325);
and I_39 (I2005,I1988,I1322);
dffarx1 I_40 (I2022,I2005,I1294,I1971);
not I_41 (I1960,I2022);
dffarx1 I_42 (I2053,I2022,I1294,I1971);
not I_43 (I1948,I2053);
nor I_44 (I2084,I1328,I1325);
not I_45 (I2101,I2084);
nor I_46 (I2118,I2022,I2101);
dffarx1 I_47 (I2135,I1331,I1294,I1971);
not I_48 (I2152,I2135);
nand I_49 (I1951,I2135,I2101);
dffarx1 I_50 (I2183,I2135,I1294,I1971);
and I_51 (I1936,I2022,I2183);
nand I_52 (I2214,I1316,I1310);
and I_53 (I2231,I2214,I1313);
dffarx1 I_54 (I2248,I2231,I1294,I1971);
nor I_55 (I2265,I2248,I2152);
and I_56 (I2282,I2084,I2265);
nor I_57 (I2299,I2248,I2022);
dffarx1 I_58 (I1942,I2248,I1294,I1971);
dffarx1 I_59 (I2330,I1319,I1294,I1971);
and I_60 (I2347,I2330,I1304);
or I_61 (I2364,I2347,I2282);
dffarx1 I_62 (I1954,I2364,I1294,I1971);
nand I_63 (I1963,I2347,I2299);
dffarx1 I_64 (I1933,I2347,I1294,I1971);
dffarx1 I_65 (I2423,I1334,I1294,I1971);
nand I_66 (I1957,I2423,I2118);
dffarx1 I_67 (I1945,I2423,I1294,I1971);
nand I_68 (I2468,I2423,I2084);
and I_69 (I2485,I2135,I2468);
dffarx1 I_70 (I1939,I2485,I1294,I1971);
not I_71 (I2549,I1301);
not I_72 (I2566,I1957);
nor I_73 (I2583,I1936,I1948);
nand I_74 (I2600,I2583,I1942);
dffarx1 I_75 (I2520,I2600,I1294,I2549);
nor I_76 (I2631,I2566,I1936);
nand I_77 (I2648,I2631,I1963);
nand I_78 (I2665,I2648,I2600);
not I_79 (I2682,I1936);
not I_80 (I2699,I1939);
nor I_81 (I2716,I2699,I1951);
and I_82 (I2733,I2716,I1954);
or I_83 (I2750,I2733,I1960);
dffarx1 I_84 (I2767,I2750,I1294,I2549);
nor I_85 (I2784,I2767,I2648);
nand I_86 (I2535,I2682,I2784);
not I_87 (I2532,I2767);
and I_88 (I2829,I2767,I2665);
dffarx1 I_89 (I2517,I2829,I1294,I2549);
dffarx1 I_90 (I2860,I2767,I1294,I2549);
and I_91 (I2514,I2682,I2860);
nand I_92 (I2891,I2566,I1939);
not I_93 (I2908,I2891);
nor I_94 (I2925,I2767,I2908);
dffarx1 I_95 (I2942,I1933,I1294,I2549);
nand I_96 (I2959,I2942,I2891);
and I_97 (I2976,I2682,I2959);
dffarx1 I_98 (I2541,I2976,I1294,I2549);
not I_99 (I3007,I2942);
nand I_100 (I2529,I2942,I2925);
nand I_101 (I2523,I2942,I2908);
dffarx1 I_102 (I3052,I1945,I1294,I2549);
not I_103 (I3069,I3052);
nor I_104 (I2538,I2942,I3069);
nor I_105 (I3100,I3069,I3007);
and I_106 (I3117,I2648,I3100);
or I_107 (I3134,I2891,I3117);
dffarx1 I_108 (I2526,I3134,I1294,I2549);
dffarx1 I_109 (I2511,I3069,I1294,I2549);
not I_110 (I3212,I1301);
not I_111 (I3229,I2529);
nor I_112 (I3246,I2517,I2523);
nand I_113 (I3263,I3246,I2532);
dffarx1 I_114 (I3186,I3263,I1294,I3212);
nor I_115 (I3294,I3229,I2517);
nand I_116 (I3311,I3294,I2520);
not I_117 (I3201,I3311);
dffarx1 I_118 (I3183,I3311,I1294,I3212);
not I_119 (I3356,I2517);
not I_120 (I3373,I3356);
not I_121 (I3390,I2541);
nor I_122 (I3407,I3390,I2514);
and I_123 (I3424,I3407,I2535);
or I_124 (I3441,I3424,I2526);
dffarx1 I_125 (I3458,I3441,I1294,I3212);
nor I_126 (I3475,I3458,I3311);
nor I_127 (I3492,I3458,I3373);
nand I_128 (I3198,I3263,I3492);
nand I_129 (I3523,I3229,I2541);
nand I_130 (I3540,I3523,I3458);
and I_131 (I3557,I3523,I3540);
dffarx1 I_132 (I3180,I3557,I1294,I3212);
dffarx1 I_133 (I3588,I3523,I1294,I3212);
and I_134 (I3177,I3356,I3588);
dffarx1 I_135 (I3619,I2511,I1294,I3212);
not I_136 (I3636,I3619);
nor I_137 (I3653,I3311,I3636);
and I_138 (I3670,I3619,I3653);
nand I_139 (I3192,I3619,I3373);
dffarx1 I_140 (I3701,I3619,I1294,I3212);
not I_141 (I3189,I3701);
dffarx1 I_142 (I3732,I2538,I1294,I3212);
not I_143 (I3749,I3732);
or I_144 (I3766,I3749,I3670);
dffarx1 I_145 (I3195,I3766,I1294,I3212);
nand I_146 (I3204,I3749,I3475);
dffarx1 I_147 (I3174,I3749,I1294,I3212);
endmodule


