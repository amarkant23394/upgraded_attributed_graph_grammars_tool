module test_final(G18_1_l_13,G15_1_l_13,IN_1_1_l_13,IN_4_1_l_13,IN_5_1_l_13,IN_7_1_l_13,IN_9_1_l_13,IN_10_1_l_13,IN_1_3_l_13,IN_2_3_l_13,IN_4_3_l_13,blif_clk_net_1_r_2,blif_reset_net_1_r_2,G42_1_r_2,n_572_1_r_2,n_549_1_r_2,n_569_1_r_2,n_452_1_r_2,n_42_2_r_2,G199_2_r_2,ACVQN1_5_r_2,P6_5_r_2);
input G18_1_l_13,G15_1_l_13,IN_1_1_l_13,IN_4_1_l_13,IN_5_1_l_13,IN_7_1_l_13,IN_9_1_l_13,IN_10_1_l_13,IN_1_3_l_13,IN_2_3_l_13,IN_4_3_l_13,blif_clk_net_1_r_2,blif_reset_net_1_r_2;
output G42_1_r_2,n_572_1_r_2,n_549_1_r_2,n_569_1_r_2,n_452_1_r_2,n_42_2_r_2,G199_2_r_2,ACVQN1_5_r_2,P6_5_r_2;
wire G42_1_r_13,n_572_1_r_13,n_573_1_r_13,n_549_1_r_13,n_569_1_r_13,n_452_1_r_13,ACVQN2_3_r_13,n_266_and_0_3_r_13,ACVQN1_5_r_13,P6_5_r_13,n4_1_l_13,n17_internal_13,n17_13,n28_13,ACVQN1_3_l_13,n4_1_r_13,n_266_and_0_3_l_13,n_573_1_l_13,n14_internal_13,n14_13,n_549_1_l_13,n_569_1_l_13,P6_5_r_internal_13,n18_13,n19_13,n20_13,n21_13,n22_13,n23_13,n24_13,n25_13,n26_13,n27_13,n_573_1_r_2,N3_2_l_2,n5_2,G199_2_l_2,n13_2,ACVQN2_3_l_2,n16_2,N1_4_l_2,n26_2,n17_internal_2,n17_2,n4_1_r_2,N3_2_r_2,P6_5_r_internal_2,n18_2,n19_2,n20_2,n21_2,n22_2,n23_2,n24_2,n25_2;
DFFARX1 I_0(n4_1_r_13,blif_clk_net_1_r_2,n5_2,G42_1_r_13,);
nor I_1(n_572_1_r_13,n28_13,n_569_1_l_13);
nand I_2(n_573_1_r_13,n18_13,n19_13);
nand I_3(n_549_1_r_13,n_569_1_r_13,n22_13);
nand I_4(n_569_1_r_13,n17_13,n18_13);
nor I_5(n_452_1_r_13,n_573_1_l_13,n25_13);
DFFARX1 I_6(n_266_and_0_3_l_13,blif_clk_net_1_r_2,n5_2,ACVQN2_3_r_13,);
nor I_7(n_266_and_0_3_r_13,n17_13,n14_13);
DFFARX1 I_8(n_549_1_l_13,blif_clk_net_1_r_2,n5_2,ACVQN1_5_r_13,);
not I_9(P6_5_r_13,P6_5_r_internal_13);
nor I_10(n4_1_l_13,G18_1_l_13,IN_1_1_l_13);
DFFARX1 I_11(n4_1_l_13,blif_clk_net_1_r_2,n5_2,n17_internal_13,);
not I_12(n17_13,n17_internal_13);
DFFARX1 I_13(IN_1_3_l_13,blif_clk_net_1_r_2,n5_2,n28_13,);
DFFARX1 I_14(IN_2_3_l_13,blif_clk_net_1_r_2,n5_2,ACVQN1_3_l_13,);
nor I_15(n4_1_r_13,n_573_1_l_13,n_549_1_l_13);
and I_16(n_266_and_0_3_l_13,IN_4_3_l_13,ACVQN1_3_l_13);
nand I_17(n_573_1_l_13,n20_13,n24_13);
DFFARX1 I_18(n_573_1_l_13,blif_clk_net_1_r_2,n5_2,n14_internal_13,);
not I_19(n14_13,n14_internal_13);
and I_20(n_549_1_l_13,n21_13,n26_13);
nand I_21(n_569_1_l_13,n20_13,n21_13);
DFFARX1 I_22(n_569_1_l_13,blif_clk_net_1_r_2,n5_2,P6_5_r_internal_13,);
nand I_23(n18_13,n23_13,n24_13);
or I_24(n19_13,G15_1_l_13,IN_7_1_l_13);
not I_25(n20_13,IN_9_1_l_13);
not I_26(n21_13,IN_10_1_l_13);
nand I_27(n22_13,n17_13,n28_13);
not I_28(n23_13,G18_1_l_13);
not I_29(n24_13,IN_5_1_l_13);
nor I_30(n25_13,G15_1_l_13,IN_7_1_l_13);
nand I_31(n26_13,IN_4_1_l_13,n27_13);
not I_32(n27_13,G15_1_l_13);
DFFARX1 I_33(n4_1_r_2,blif_clk_net_1_r_2,n5_2,G42_1_r_2,);
nor I_34(n_572_1_r_2,n26_2,n18_2);
nand I_35(n_573_1_r_2,n17_2,n19_2);
nor I_36(n_549_1_r_2,G199_2_l_2,n20_2);
nand I_37(n_569_1_r_2,n13_2,n19_2);
not I_38(n_452_1_r_2,n_573_1_r_2);
nor I_39(n_42_2_r_2,ACVQN2_3_l_2,n18_2);
DFFARX1 I_40(N3_2_r_2,blif_clk_net_1_r_2,n5_2,G199_2_r_2,);
DFFARX1 I_41(ACVQN2_3_l_2,blif_clk_net_1_r_2,n5_2,ACVQN1_5_r_2,);
not I_42(P6_5_r_2,P6_5_r_internal_2);
and I_43(N3_2_l_2,n24_2,ACVQN2_3_r_13);
not I_44(n5_2,blif_reset_net_1_r_2);
DFFARX1 I_45(N3_2_l_2,blif_clk_net_1_r_2,n5_2,G199_2_l_2,);
not I_46(n13_2,G199_2_l_2);
DFFARX1 I_47(G42_1_r_13,blif_clk_net_1_r_2,n5_2,ACVQN2_3_l_2,);
DFFARX1 I_48(P6_5_r_13,blif_clk_net_1_r_2,n5_2,n16_2,);
and I_49(N1_4_l_2,n25_2,n_572_1_r_13);
DFFARX1 I_50(N1_4_l_2,blif_clk_net_1_r_2,n5_2,n26_2,);
DFFARX1 I_51(n_573_1_r_13,blif_clk_net_1_r_2,n5_2,n17_internal_2,);
not I_52(n17_2,n17_internal_2);
nor I_53(n4_1_r_2,n26_2,n22_2);
nor I_54(N3_2_r_2,n17_2,n23_2);
DFFARX1 I_55(G199_2_l_2,blif_clk_net_1_r_2,n5_2,P6_5_r_internal_2,);
nor I_56(n18_2,n_549_1_r_13,n_266_and_0_3_r_13);
nand I_57(n19_2,n16_2,n_572_1_r_13);
nor I_58(n20_2,n26_2,n21_2);
not I_59(n21_2,n18_2);
and I_60(n22_2,n16_2,n_572_1_r_13);
nor I_61(n23_2,n13_2,n21_2);
nand I_62(n24_2,n_549_1_r_13,n_452_1_r_13);
nand I_63(n25_2,G42_1_r_13,ACVQN1_5_r_13);
endmodule


