module test_final(IN_1_2_l_2,IN_2_2_l_2,IN_3_2_l_2,IN_6_2_l_2,IN_1_3_l_2,IN_2_3_l_2,IN_4_3_l_2,IN_1_4_l_2,IN_2_4_l_2,IN_3_4_l_2,IN_6_4_l_2,blif_clk_net_1_r_17,blif_reset_net_1_r_17,G42_1_r_17,n_572_1_r_17,n_573_1_r_17,n_549_1_r_17,n_569_1_r_17,n_452_1_r_17,ACVQN2_3_r_17,n_266_and_0_3_r_17,G199_4_r_17,G214_4_r_17);
input IN_1_2_l_2,IN_2_2_l_2,IN_3_2_l_2,IN_6_2_l_2,IN_1_3_l_2,IN_2_3_l_2,IN_4_3_l_2,IN_1_4_l_2,IN_2_4_l_2,IN_3_4_l_2,IN_6_4_l_2,blif_clk_net_1_r_17,blif_reset_net_1_r_17;
output G42_1_r_17,n_572_1_r_17,n_573_1_r_17,n_549_1_r_17,n_569_1_r_17,n_452_1_r_17,ACVQN2_3_r_17,n_266_and_0_3_r_17,G199_4_r_17,G214_4_r_17;
wire G42_1_r_2,n_572_1_r_2,n_573_1_r_2,n_549_1_r_2,n_569_1_r_2,n_452_1_r_2,n_42_2_r_2,G199_2_r_2,ACVQN1_5_r_2,P6_5_r_2,N3_2_l_2,G199_2_l_2,n13_2,ACVQN2_3_l_2,n16_2,N1_4_l_2,n26_2,n17_internal_2,n17_2,n4_1_r_2,N3_2_r_2,P6_5_r_internal_2,n18_2,n19_2,n20_2,n21_2,n22_2,n23_2,n24_2,n25_2,n_431_0_l_17,n6_17,n20_internal_17,n20_17,ACVQN1_5_l_17,n19_internal_17,n19_17,n4_1_r_17,n2_17,n17_internal_17,n17_17,N1_4_r_17,n5_17,n21_17,n22_17,n23_17,n24_17,n25_17,n26_17,n27_17,n28_17,n29_17,n30_17,n31_17,n32_17;
DFFARX1 I_0(n4_1_r_2,blif_clk_net_1_r_17,n6_17,G42_1_r_2,);
nor I_1(n_572_1_r_2,n26_2,n18_2);
nand I_2(n_573_1_r_2,n17_2,n19_2);
nor I_3(n_549_1_r_2,G199_2_l_2,n20_2);
nand I_4(n_569_1_r_2,n13_2,n19_2);
not I_5(n_452_1_r_2,n_573_1_r_2);
nor I_6(n_42_2_r_2,ACVQN2_3_l_2,n18_2);
DFFARX1 I_7(N3_2_r_2,blif_clk_net_1_r_17,n6_17,G199_2_r_2,);
DFFARX1 I_8(ACVQN2_3_l_2,blif_clk_net_1_r_17,n6_17,ACVQN1_5_r_2,);
not I_9(P6_5_r_2,P6_5_r_internal_2);
and I_10(N3_2_l_2,IN_6_2_l_2,n24_2);
DFFARX1 I_11(N3_2_l_2,blif_clk_net_1_r_17,n6_17,G199_2_l_2,);
not I_12(n13_2,G199_2_l_2);
DFFARX1 I_13(IN_1_3_l_2,blif_clk_net_1_r_17,n6_17,ACVQN2_3_l_2,);
DFFARX1 I_14(IN_2_3_l_2,blif_clk_net_1_r_17,n6_17,n16_2,);
and I_15(N1_4_l_2,IN_6_4_l_2,n25_2);
DFFARX1 I_16(N1_4_l_2,blif_clk_net_1_r_17,n6_17,n26_2,);
DFFARX1 I_17(IN_3_4_l_2,blif_clk_net_1_r_17,n6_17,n17_internal_2,);
not I_18(n17_2,n17_internal_2);
nor I_19(n4_1_r_2,n26_2,n22_2);
nor I_20(N3_2_r_2,n17_2,n23_2);
DFFARX1 I_21(G199_2_l_2,blif_clk_net_1_r_17,n6_17,P6_5_r_internal_2,);
nor I_22(n18_2,IN_1_2_l_2,IN_3_2_l_2);
nand I_23(n19_2,IN_4_3_l_2,n16_2);
nor I_24(n20_2,n26_2,n21_2);
not I_25(n21_2,n18_2);
and I_26(n22_2,IN_4_3_l_2,n16_2);
nor I_27(n23_2,n13_2,n21_2);
nand I_28(n24_2,IN_2_2_l_2,IN_3_2_l_2);
nand I_29(n25_2,IN_1_4_l_2,IN_2_4_l_2);
DFFARX1 I_30(n4_1_r_17,blif_clk_net_1_r_17,n6_17,G42_1_r_17,);
nor I_31(n_572_1_r_17,ACVQN1_5_l_17,n19_17);
nand I_32(n_573_1_r_17,n20_17,n21_17);
nand I_33(n_549_1_r_17,n23_17,n24_17);
nand I_34(n_569_1_r_17,n21_17,n22_17);
not I_35(n_452_1_r_17,n23_17);
DFFARX1 I_36(n19_17,blif_clk_net_1_r_17,n6_17,ACVQN2_3_r_17,);
nor I_37(n_266_and_0_3_r_17,n17_17,n29_17);
DFFARX1 I_38(N1_4_r_17,blif_clk_net_1_r_17,n6_17,G199_4_r_17,);
DFFARX1 I_39(n5_17,blif_clk_net_1_r_17,n6_17,G214_4_r_17,);
or I_40(n_431_0_l_17,n26_17,n_569_1_r_2);
not I_41(n6_17,blif_reset_net_1_r_17);
DFFARX1 I_42(n_431_0_l_17,blif_clk_net_1_r_17,n6_17,n20_internal_17,);
not I_43(n20_17,n20_internal_17);
DFFARX1 I_44(n_452_1_r_2,blif_clk_net_1_r_17,n6_17,ACVQN1_5_l_17,);
DFFARX1 I_45(G42_1_r_2,blif_clk_net_1_r_17,n6_17,n19_internal_17,);
not I_46(n19_17,n19_internal_17);
nor I_47(n4_1_r_17,n5_17,n25_17);
not I_48(n2_17,n29_17);
DFFARX1 I_49(n2_17,blif_clk_net_1_r_17,n6_17,n17_internal_17,);
not I_50(n17_17,n17_internal_17);
nor I_51(N1_4_r_17,n29_17,n31_17);
not I_52(n5_17,n_572_1_r_2);
and I_53(n21_17,n32_17,n_42_2_r_2);
not I_54(n22_17,n25_17);
nand I_55(n23_17,n20_17,n22_17);
nand I_56(n24_17,n19_17,n22_17);
nand I_57(n25_17,n30_17,G199_2_r_2);
and I_58(n26_17,n27_17,ACVQN1_5_r_2);
nor I_59(n27_17,n28_17,G42_1_r_2);
not I_60(n28_17,P6_5_r_2);
nor I_61(n29_17,n28_17,n_549_1_r_2);
and I_62(n30_17,n5_17,n_549_1_r_2);
nor I_63(n31_17,n21_17,n_572_1_r_2);
nor I_64(n32_17,n_572_1_r_2,n_549_1_r_2);
endmodule


