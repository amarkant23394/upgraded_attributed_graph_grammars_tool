module test_I13443(I13214,I11290,I1477,I1470,I11284,I13443);
input I13214,I11290,I1477,I1470,I11284;
output I13443;
wire I11287,I13231,I13392,I11281,I13197,I13265,I13426,I11593,I13248,I13409;
DFFARX1 I_0(I1470,,,I11287,);
and I_1(I13231,I13214,I11290);
nand I_2(I13392,I11287,I11284);
not I_3(I11281,I11593);
not I_4(I13197,I1477);
not I_5(I13265,I13248);
DFFARX1 I_6(I13409,I1470,I13197,,,I13426,);
DFFARX1 I_7(I1470,,,I11593,);
DFFARX1 I_8(I13231,I1470,I13197,,,I13248,);
nor I_9(I13443,I13426,I13265);
and I_10(I13409,I13392,I11281);
endmodule


