module test_final(IN_1_0_l_14,IN_2_0_l_14,IN_3_0_l_14,IN_4_0_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_3_3_l_14,IN_1_8_l_14,IN_2_8_l_14,IN_3_8_l_14,IN_6_8_l_14,IN_1_10_l_14,IN_2_10_l_14,IN_3_10_l_14,IN_4_10_l_14,blif_clk_net_8_r_8,blif_reset_net_8_r_8,N1371_0_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,N1508_10_r_8);
input IN_1_0_l_14,IN_2_0_l_14,IN_3_0_l_14,IN_4_0_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_3_3_l_14,IN_1_8_l_14,IN_2_8_l_14,IN_3_8_l_14,IN_6_8_l_14,IN_1_10_l_14,IN_2_10_l_14,IN_3_10_l_14,IN_4_10_l_14,blif_clk_net_8_r_8,blif_reset_net_8_r_8;
output N1371_0_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,N1508_10_r_8;
wire N1371_0_r_14,N1508_0_r_14,N1507_6_r_14,N1508_6_r_14,G42_7_r_14,n_572_7_r_14,n_573_7_r_14,n_549_7_r_14,n_569_7_r_14,n_452_7_r_14,N6147_9_r_14,N6134_9_r_14,I_BUFF_1_9_r_14,N3_8_l_14,n47_14,n4_7_r_14,n26_14,n27_14,n28_14,n29_14,n30_14,n31_14,n32_14,n33_14,n34_14,n35_14,n36_14,n37_14,n38_14,n39_14,n40_14,n41_14,n42_14,n43_14,n44_14,n45_14,n46_14,N1508_0_r_8,N1372_1_r_8,I_BUFF_1_9_r_8,N1372_10_r_8,N3_8_l_8,n8_8,n53_8,n29_8,N3_8_r_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8,n38_8,n39_8,n40_8,n41_8,n42_8,n43_8,n44_8,n45_8,n46_8,n47_8,n48_8,n49_8,n50_8,n51_8,n52_8;
nor I_0(N1371_0_r_14,n47_14,n30_14);
nor I_1(N1508_0_r_14,n30_14,n41_14);
nor I_2(N1507_6_r_14,n37_14,n44_14);
nor I_3(N1508_6_r_14,n30_14,n39_14);
DFFARX1 I_4(n4_7_r_14,blif_clk_net_8_r_8,n8_8,G42_7_r_14,);
nor I_5(n_572_7_r_14,n28_14,n29_14);
nand I_6(n_573_7_r_14,n26_14,n27_14);
nor I_7(n_549_7_r_14,n31_14,n32_14);
nand I_8(n_569_7_r_14,n26_14,n30_14);
nor I_9(n_452_7_r_14,n47_14,n28_14);
nor I_10(N6147_9_r_14,n36_14,n37_14);
nor I_11(N6134_9_r_14,n28_14,n36_14);
not I_12(I_BUFF_1_9_r_14,n26_14);
and I_13(N3_8_l_14,IN_6_8_l_14,n38_14);
DFFARX1 I_14(N3_8_l_14,blif_clk_net_8_r_8,n8_8,n47_14,);
nor I_15(n4_7_r_14,n47_14,n35_14);
nand I_16(n26_14,IN_1_10_l_14,IN_2_10_l_14);
not I_17(n27_14,n28_14);
nor I_18(n28_14,IN_2_0_l_14,n43_14);
not I_19(n29_14,n33_14);
not I_20(n30_14,n31_14);
nor I_21(n31_14,IN_1_3_l_14,n46_14);
and I_22(n32_14,n33_14,n34_14);
nand I_23(n33_14,I_BUFF_1_9_r_14,n45_14);
nor I_24(n34_14,n42_14,n43_14);
nor I_25(n35_14,IN_1_8_l_14,IN_3_8_l_14);
nor I_26(n36_14,n47_14,n34_14);
not I_27(n37_14,n35_14);
nand I_28(n38_14,IN_2_8_l_14,IN_3_8_l_14);
nand I_29(n39_14,n29_14,n40_14);
nand I_30(n40_14,n27_14,n37_14);
nor I_31(n41_14,I_BUFF_1_9_r_14,n34_14);
nor I_32(n42_14,IN_3_0_l_14,IN_4_0_l_14);
not I_33(n43_14,IN_1_0_l_14);
nor I_34(n44_14,n27_14,n33_14);
or I_35(n45_14,IN_3_10_l_14,IN_4_10_l_14);
or I_36(n46_14,IN_2_3_l_14,IN_3_3_l_14);
nor I_37(N1371_0_r_8,n46_8,n51_8);
not I_38(N1508_0_r_8,n46_8);
nor I_39(N1372_1_r_8,n37_8,n49_8);
and I_40(N1508_1_r_8,N1372_1_r_8,n29_8);
nor I_41(N1507_6_r_8,n47_8,n48_8);
nor I_42(N1508_6_r_8,n37_8,n38_8);
nor I_43(n_42_8_r_8,I_BUFF_1_9_r_8,n53_8);
DFFARX1 I_44(N3_8_r_8,blif_clk_net_8_r_8,n8_8,G199_8_r_8,);
nor I_45(N6147_9_r_8,n29_8,n30_8);
nor I_46(N6134_9_r_8,n30_8,n31_8);
not I_47(I_BUFF_1_9_r_8,n35_8);
nor I_48(N1372_10_r_8,n46_8,n49_8);
nor I_49(N1508_10_r_8,n40_8,n41_8);
and I_50(N3_8_l_8,n36_8,N1508_0_r_14);
not I_51(n8_8,blif_reset_net_8_r_8);
DFFARX1 I_52(N3_8_l_8,blif_clk_net_8_r_8,n8_8,n53_8,);
not I_53(n29_8,n53_8);
nor I_54(N3_8_r_8,n33_8,n34_8);
and I_55(n30_8,n32_8,n33_8);
nor I_56(n31_8,N1371_0_r_14,N1507_6_r_14);
nand I_57(n32_8,n42_8,n_569_7_r_14);
or I_58(n33_8,n46_8,N1371_0_r_14);
nor I_59(n34_8,n32_8,n35_8);
nand I_60(n35_8,n44_8,n_549_7_r_14);
nand I_61(n36_8,N1371_0_r_14,N1508_6_r_14);
not I_62(n37_8,n31_8);
nand I_63(n38_8,N1508_0_r_8,n39_8);
nand I_64(n39_8,n33_8,n50_8);
and I_65(n40_8,n32_8,n35_8);
not I_66(n41_8,N1372_10_r_8);
and I_67(n42_8,n43_8,N6147_9_r_14);
nand I_68(n43_8,n44_8,n45_8);
nand I_69(n44_8,G42_7_r_14,N1507_6_r_14);
not I_70(n45_8,n_549_7_r_14);
nand I_71(n46_8,n_573_7_r_14,n_452_7_r_14);
not I_72(n47_8,n39_8);
nor I_73(n48_8,n35_8,n49_8);
not I_74(n49_8,n51_8);
nand I_75(n50_8,I_BUFF_1_9_r_8,n51_8);
nor I_76(n51_8,n52_8,n_572_7_r_14);
or I_77(n52_8,N1508_0_r_14,N6134_9_r_14);
endmodule


