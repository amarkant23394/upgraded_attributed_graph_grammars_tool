module test_I13177(I11296,I1477,I11768,I11847,I13409,I1470,I11327,I13177);
input I11296,I1477,I11768,I11847,I13409,I1470,I11327;
output I13177;
wire I11302,I11278,I8827,I13460,I11624,I13197,I13542,I13296,I13426,I11272,I13508,I13491,I11310,I11864;
nand I_0(I13177,I13296,I13542);
DFFARX1 I_1(I11864,I1470,I11310,,,I11302,);
DFFARX1 I_2(I11624,I1470,I11310,,,I11278,);
DFFARX1 I_3(I1470,,,I8827,);
not I_4(I13460,I13426);
nand I_5(I11624,I11327,I8827);
not I_6(I13197,I1477);
nor I_7(I13542,I13508,I13460);
nor I_8(I13296,I11278,I11302);
DFFARX1 I_9(I13409,I1470,I13197,,,I13426,);
DFFARX1 I_10(I11768,I1470,I11310,,,I11272,);
and I_11(I13508,I13491,I11272);
DFFARX1 I_12(I11296,I1470,I13197,,,I13491,);
not I_13(I11310,I1477);
and I_14(I11864,I11624,I11847);
endmodule


