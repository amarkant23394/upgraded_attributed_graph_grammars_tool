module test_final(G1_0_l_4,G2_0_l_4,IN_2_0_l_4,IN_4_0_l_4,IN_5_0_l_4,IN_7_0_l_4,IN_8_0_l_4,IN_10_0_l_4,IN_11_0_l_4,IN_1_5_l_4,IN_2_5_l_4,blif_clk_net_1_r_0,blif_reset_net_1_r_0,G42_1_r_0,n_572_1_r_0,n_573_1_r_0,n_549_1_r_0,n_42_2_r_0,G199_2_r_0,G199_4_r_0,G214_4_r_0);
input G1_0_l_4,G2_0_l_4,IN_2_0_l_4,IN_4_0_l_4,IN_5_0_l_4,IN_7_0_l_4,IN_8_0_l_4,IN_10_0_l_4,IN_11_0_l_4,IN_1_5_l_4,IN_2_5_l_4,blif_clk_net_1_r_0,blif_reset_net_1_r_0;
output G42_1_r_0,n_572_1_r_0,n_573_1_r_0,n_549_1_r_0,n_42_2_r_0,G199_2_r_0,G199_4_r_0,G214_4_r_0;
wire G42_1_r_4,n_572_1_r_4,n_573_1_r_4,n_549_1_r_4,n_569_1_r_4,ACVQN2_3_r_4,n_266_and_0_3_r_4,ACVQN1_5_r_4,P6_5_r_4,n_431_0_l_4,G78_0_l_4,ACVQN1_5_l_4,n16_4,n17_internal_4,n17_4,n4_1_r_4,n19_4,n15_internal_4,n15_4,P6_5_r_internal_4,n20_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n_569_1_r_0,n4_1_l_0,n6_0,n37_0,n38_0,n20_0,ACVQN1_3_l_0,n4_1_r_0,N3_2_r_0,N1_4_r_0,n2_0,n21_0,n22_0,n23_0,n24_0,n25_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0;
DFFARX1 I_0(n4_1_r_4,blif_clk_net_1_r_0,n6_0,G42_1_r_4,);
nor I_1(n_572_1_r_4,G78_0_l_4,n17_4);
nand I_2(n_573_1_r_4,G2_0_l_4,n16_4);
nor I_3(n_549_1_r_4,n22_4,n23_4);
nand I_4(n_569_1_r_4,n20_4,n21_4);
DFFARX1 I_5(n19_4,blif_clk_net_1_r_0,n6_0,ACVQN2_3_r_4,);
nor I_6(n_266_and_0_3_r_4,n15_4,n29_4);
DFFARX1 I_7(n19_4,blif_clk_net_1_r_0,n6_0,ACVQN1_5_r_4,);
not I_8(P6_5_r_4,P6_5_r_internal_4);
or I_9(n_431_0_l_4,IN_8_0_l_4,n26_4);
DFFARX1 I_10(n_431_0_l_4,blif_clk_net_1_r_0,n6_0,G78_0_l_4,);
DFFARX1 I_11(IN_2_5_l_4,blif_clk_net_1_r_0,n6_0,ACVQN1_5_l_4,);
not I_12(n16_4,ACVQN1_5_l_4);
DFFARX1 I_13(IN_1_5_l_4,blif_clk_net_1_r_0,n6_0,n17_internal_4,);
not I_14(n17_4,n17_internal_4);
nor I_15(n4_1_r_4,n30_4,n31_4);
nand I_16(n19_4,G1_0_l_4,n33_4);
DFFARX1 I_17(G78_0_l_4,blif_clk_net_1_r_0,n6_0,n15_internal_4,);
not I_18(n15_4,n15_internal_4);
DFFARX1 I_19(ACVQN1_5_l_4,blif_clk_net_1_r_0,n6_0,P6_5_r_internal_4,);
and I_20(n20_4,IN_11_0_l_4,n16_4);
nor I_21(n21_4,G2_0_l_4,IN_10_0_l_4);
nand I_22(n22_4,G78_0_l_4,n25_4);
nand I_23(n23_4,IN_11_0_l_4,n24_4);
not I_24(n24_4,G2_0_l_4);
not I_25(n25_4,IN_10_0_l_4);
and I_26(n26_4,IN_2_0_l_4,n27_4);
nor I_27(n27_4,IN_4_0_l_4,n28_4);
not I_28(n28_4,G1_0_l_4);
not I_29(n29_4,n30_4);
nand I_30(n30_4,IN_7_0_l_4,n32_4);
nand I_31(n31_4,IN_11_0_l_4,n25_4);
nor I_32(n32_4,G2_0_l_4,n33_4);
not I_33(n33_4,IN_5_0_l_4);
DFFARX1 I_34(n4_1_r_0,blif_clk_net_1_r_0,n6_0,G42_1_r_0,);
nor I_35(n_572_1_r_0,n23_0,ACVQN2_3_r_4);
nand I_36(n_573_1_r_0,n21_0,n22_0);
nand I_37(n_549_1_r_0,n_569_1_r_0,n24_0);
nand I_38(n_569_1_r_0,n21_0,n26_0);
nor I_39(n_42_2_r_0,n27_0,n28_0);
DFFARX1 I_40(N3_2_r_0,blif_clk_net_1_r_0,n6_0,G199_2_r_0,);
DFFARX1 I_41(N1_4_r_0,blif_clk_net_1_r_0,n6_0,G199_4_r_0,);
DFFARX1 I_42(n2_0,blif_clk_net_1_r_0,n6_0,G214_4_r_0,);
nor I_43(n4_1_l_0,G42_1_r_4,n_573_1_r_4);
not I_44(n6_0,blif_reset_net_1_r_0);
DFFARX1 I_45(n4_1_l_0,blif_clk_net_1_r_0,n6_0,n37_0,);
DFFARX1 I_46(n_549_1_r_4,blif_clk_net_1_r_0,n6_0,n38_0,);
not I_47(n20_0,n38_0);
DFFARX1 I_48(n_572_1_r_4,blif_clk_net_1_r_0,n6_0,ACVQN1_3_l_0,);
nor I_49(n4_1_r_0,n23_0,n_266_and_0_3_r_4);
nor I_50(N3_2_r_0,n31_0,n32_0);
nor I_51(N1_4_r_0,n29_0,n32_0);
not I_52(n2_0,n31_0);
nor I_53(n21_0,n37_0,n_569_1_r_4);
not I_54(n22_0,ACVQN2_3_r_4);
nand I_55(n23_0,n20_0,n30_0);
nand I_56(n24_0,n38_0,n25_0);
nor I_57(n25_0,n_569_1_r_4,n_266_and_0_3_r_4);
not I_58(n26_0,n_266_and_0_3_r_4);
not I_59(n27_0,n29_0);
nor I_60(n28_0,ACVQN1_5_r_4,P6_5_r_4);
nand I_61(n29_0,n26_0,n33_0);
not I_62(n30_0,n_569_1_r_4);
nand I_63(n31_0,ACVQN1_3_l_0,n_572_1_r_4);
and I_64(n32_0,n35_0,n36_0);
nand I_65(n33_0,n34_0,G42_1_r_4);
not I_66(n34_0,P6_5_r_4);
nor I_67(n35_0,n_573_1_r_4,P6_5_r_4);
nor I_68(n36_0,ACVQN2_3_r_4,ACVQN1_5_r_4);
endmodule


