module test_I13525(I1477,I11689,I11429,I1470,I11284,I11751,I13525);
input I1477,I11689,I11429,I1470,I11284,I11751;
output I13525;
wire I11296,I11768,I11559,I11287,I11281,I11593,I13197,I13409,I13392,I13426,I11272,I13508,I13491,I11310;
nand I_0(I11296,I11559,I11689);
and I_1(I11768,I11429,I11751);
DFFARX1 I_2(I1470,I11310,,,I11559,);
nor I_3(I13525,I13508,I13426);
DFFARX1 I_4(I1470,I11310,,,I11287,);
not I_5(I11281,I11593);
DFFARX1 I_6(I11559,I1470,I11310,,,I11593,);
not I_7(I13197,I1477);
and I_8(I13409,I13392,I11281);
nand I_9(I13392,I11287,I11284);
DFFARX1 I_10(I13409,I1470,I13197,,,I13426,);
DFFARX1 I_11(I11768,I1470,I11310,,,I11272,);
and I_12(I13508,I13491,I11272);
DFFARX1 I_13(I11296,I1470,I13197,,,I13491,);
not I_14(I11310,I1477);
endmodule


