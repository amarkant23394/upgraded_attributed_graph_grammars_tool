module test_I2827(I1351,I1407,I2827);
input I1351,I1407;
output I2827;
wire I2776;
nor I_0(I2827,I2776,I1351);
not I_1(I2776,I1407);
endmodule


