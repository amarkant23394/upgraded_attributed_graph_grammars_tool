module test_I3732(I1294,I1301,I3732);
input I1294,I1301;
output I3732;
wire I3396,I2554,I2866,I3379,I2548,I2583,I3246,I2945,I3715,I3698;
not I_0(I3396,I3379);
not I_1(I2554,I2866);
DFFARX1 I_2(I1294,I2583,,,I2866,);
not I_3(I3379,I2548);
DFFARX1 I_4(I2945,I1294,I2583,,,I2548,);
not I_5(I2583,I1301);
not I_6(I3246,I1301);
DFFARX1 I_7(I1294,I2583,,,I2945,);
not I_8(I3715,I3698);
nor I_9(I3732,I3715,I3396);
DFFARX1 I_10(I2554,I1294,I3246,,,I3698,);
endmodule


