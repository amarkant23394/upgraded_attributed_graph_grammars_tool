module test_final(G18_1_l_13,G15_1_l_13,IN_1_1_l_13,IN_4_1_l_13,IN_5_1_l_13,IN_7_1_l_13,IN_9_1_l_13,IN_10_1_l_13,IN_1_3_l_13,IN_2_3_l_13,IN_4_3_l_13,blif_clk_net_1_r_14,blif_reset_net_1_r_14,G42_1_r_14,n_572_1_r_14,n_573_1_r_14,n_549_1_r_14,n_569_1_r_14,n_42_2_r_14,G199_2_r_14,ACVQN1_5_r_14,P6_5_r_14);
input G18_1_l_13,G15_1_l_13,IN_1_1_l_13,IN_4_1_l_13,IN_5_1_l_13,IN_7_1_l_13,IN_9_1_l_13,IN_10_1_l_13,IN_1_3_l_13,IN_2_3_l_13,IN_4_3_l_13,blif_clk_net_1_r_14,blif_reset_net_1_r_14;
output G42_1_r_14,n_572_1_r_14,n_573_1_r_14,n_549_1_r_14,n_569_1_r_14,n_42_2_r_14,G199_2_r_14,ACVQN1_5_r_14,P6_5_r_14;
wire G42_1_r_13,n_572_1_r_13,n_573_1_r_13,n_549_1_r_13,n_569_1_r_13,n_452_1_r_13,ACVQN2_3_r_13,n_266_and_0_3_r_13,ACVQN1_5_r_13,P6_5_r_13,n4_1_l_13,n17_internal_13,n17_13,n28_13,ACVQN1_3_l_13,n4_1_r_13,n_266_and_0_3_l_13,n_573_1_l_13,n14_internal_13,n14_13,n_549_1_l_13,n_569_1_l_13,P6_5_r_internal_13,n18_13,n19_13,n20_13,n21_13,n22_13,n23_13,n24_13,n25_13,n26_13,n27_13,n_452_1_r_14,n4_1_l_14,n3_14,n15_internal_14,n15_14,ACVQN2_3_l_14,ACVQN1_3_l_14,N3_2_r_14,n_572_1_l_14,P6_5_r_internal_14,n16_14,n17_14,n18_14,n19_14,n20_14,n21_14,n22_14,n23_14,n24_14,n25_14,n26_14,n27_14,n28_14;
DFFARX1 I_0(n4_1_r_13,blif_clk_net_1_r_14,n3_14,G42_1_r_13,);
nor I_1(n_572_1_r_13,n28_13,n_569_1_l_13);
nand I_2(n_573_1_r_13,n18_13,n19_13);
nand I_3(n_549_1_r_13,n_569_1_r_13,n22_13);
nand I_4(n_569_1_r_13,n17_13,n18_13);
nor I_5(n_452_1_r_13,n_573_1_l_13,n25_13);
DFFARX1 I_6(n_266_and_0_3_l_13,blif_clk_net_1_r_14,n3_14,ACVQN2_3_r_13,);
nor I_7(n_266_and_0_3_r_13,n17_13,n14_13);
DFFARX1 I_8(n_549_1_l_13,blif_clk_net_1_r_14,n3_14,ACVQN1_5_r_13,);
not I_9(P6_5_r_13,P6_5_r_internal_13);
nor I_10(n4_1_l_13,G18_1_l_13,IN_1_1_l_13);
DFFARX1 I_11(n4_1_l_13,blif_clk_net_1_r_14,n3_14,n17_internal_13,);
not I_12(n17_13,n17_internal_13);
DFFARX1 I_13(IN_1_3_l_13,blif_clk_net_1_r_14,n3_14,n28_13,);
DFFARX1 I_14(IN_2_3_l_13,blif_clk_net_1_r_14,n3_14,ACVQN1_3_l_13,);
nor I_15(n4_1_r_13,n_573_1_l_13,n_549_1_l_13);
and I_16(n_266_and_0_3_l_13,IN_4_3_l_13,ACVQN1_3_l_13);
nand I_17(n_573_1_l_13,n20_13,n24_13);
DFFARX1 I_18(n_573_1_l_13,blif_clk_net_1_r_14,n3_14,n14_internal_13,);
not I_19(n14_13,n14_internal_13);
and I_20(n_549_1_l_13,n21_13,n26_13);
nand I_21(n_569_1_l_13,n20_13,n21_13);
DFFARX1 I_22(n_569_1_l_13,blif_clk_net_1_r_14,n3_14,P6_5_r_internal_13,);
nand I_23(n18_13,n23_13,n24_13);
or I_24(n19_13,G15_1_l_13,IN_7_1_l_13);
not I_25(n20_13,IN_9_1_l_13);
not I_26(n21_13,IN_10_1_l_13);
nand I_27(n22_13,n17_13,n28_13);
not I_28(n23_13,G18_1_l_13);
not I_29(n24_13,IN_5_1_l_13);
nor I_30(n25_13,G15_1_l_13,IN_7_1_l_13);
nand I_31(n26_13,IN_4_1_l_13,n27_13);
not I_32(n27_13,G15_1_l_13);
DFFARX1 I_33(n_452_1_r_14,blif_clk_net_1_r_14,n3_14,G42_1_r_14,);
and I_34(n_572_1_r_14,n18_14,n19_14);
nand I_35(n_573_1_r_14,n16_14,n17_14);
nor I_36(n_549_1_r_14,n20_14,n21_14);
or I_37(n_569_1_r_14,n_572_1_l_14,n20_14);
nor I_38(n_452_1_r_14,n23_14,ACVQN1_5_r_13);
nor I_39(n_42_2_r_14,n20_14,n22_14);
DFFARX1 I_40(N3_2_r_14,blif_clk_net_1_r_14,n3_14,G199_2_r_14,);
DFFARX1 I_41(n_572_1_l_14,blif_clk_net_1_r_14,n3_14,ACVQN1_5_r_14,);
not I_42(P6_5_r_14,P6_5_r_internal_14);
nor I_43(n4_1_l_14,n_572_1_r_13,n_573_1_r_13);
not I_44(n3_14,blif_reset_net_1_r_14);
DFFARX1 I_45(n4_1_l_14,blif_clk_net_1_r_14,n3_14,n15_internal_14,);
not I_46(n15_14,n15_internal_14);
DFFARX1 I_47(G42_1_r_13,blif_clk_net_1_r_14,n3_14,ACVQN2_3_l_14,);
DFFARX1 I_48(P6_5_r_13,blif_clk_net_1_r_14,n3_14,ACVQN1_3_l_14,);
and I_49(N3_2_r_14,n26_14,n27_14);
nor I_50(n_572_1_l_14,n_266_and_0_3_r_13,G42_1_r_13);
DFFARX1 I_51(ACVQN2_3_l_14,blif_clk_net_1_r_14,n3_14,P6_5_r_internal_14,);
nor I_52(n16_14,n_452_1_r_13,ACVQN1_5_r_13);
not I_53(n17_14,n_572_1_l_14);
nor I_54(n18_14,n_549_1_r_13,n_452_1_r_13);
nand I_55(n19_14,ACVQN1_3_l_14,n_572_1_r_13);
nor I_56(n20_14,n_572_1_r_13,n_549_1_r_13);
nor I_57(n21_14,n15_14,n22_14);
nand I_58(n22_14,n24_14,n25_14);
nand I_59(n23_14,n15_14,n24_14);
not I_60(n24_14,n_452_1_r_13);
not I_61(n25_14,n_549_1_r_13);
nor I_62(n26_14,n20_14,ACVQN1_5_r_13);
nand I_63(n27_14,n28_14,ACVQN2_3_r_13);
not I_64(n28_14,n_266_and_0_3_r_13);
endmodule


