module test_I17515(I15628,I15579,I13749,I1470,I15611,I16162,I15798,I17515);
input I15628,I15579,I13749,I1470,I15611,I16162,I15798;
output I17515;
wire I17430,I15597,I15600,I15832,I15815,I17481,I17498;
not I_0(I17430,I15579);
nor I_1(I15597,I15832,I16162);
not I_2(I17515,I17498);
or I_3(I15600,I15832,I15815);
nand I_4(I15832,I15628,I13749);
DFFARX1 I_5(I15798,I1470,I15611,,,I15815,);
nor I_6(I17481,I17430,I15597);
nand I_7(I17498,I17481,I15600);
endmodule


