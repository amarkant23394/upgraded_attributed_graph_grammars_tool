module test_final(IN_1_1_l,IN_2_1_l,IN_3_1_l,G18_7_l,G15_7_l,IN_1_7_l,IN_4_7_l,IN_5_7_l,IN_7_7_l,IN_9_7_l,IN_10_7_l,IN_1_8_l,IN_2_8_l,IN_3_8_l,IN_6_8_l,blif_clk_net_7_r,blif_reset_net_7_r,N1371_0_r,N1508_0_r,N1372_1_r,N1508_1_r,N6147_2_r,N1507_6_r,N1508_6_r,G42_7_r,n_572_7_r,n_573_7_r,n_549_7_r,n_569_7_r,n_452_7_r);
input IN_1_1_l,IN_2_1_l,IN_3_1_l,G18_7_l,G15_7_l,IN_1_7_l,IN_4_7_l,IN_5_7_l,IN_7_7_l,IN_9_7_l,IN_10_7_l,IN_1_8_l,IN_2_8_l,IN_3_8_l,IN_6_8_l,blif_clk_net_7_r,blif_reset_net_7_r;
output N1371_0_r,N1508_0_r,N1372_1_r,N1508_1_r,N6147_2_r,N1507_6_r,N1508_6_r,G42_7_r,n_572_7_r,n_573_7_r,n_549_7_r,n_569_7_r,n_452_7_r;
wire N1372_1_l,N1508_1_l,n4_1_l,G42_7_l,n_87_7_l,n_572_7_l,n_573_7_l,n_549_7_l,n_569_7_l,n_452_7_l,n4_7_l,n7_7_l,n_42_8_l,G199_8_l,N3_8_l,n3_8_l,n3_0_r,n4_0_r,n4_1_r,n5_2_r,n6_2_r,N6138_2_r,n7_2_r,n6_6_r,n7_6_r,n8_6_r,n9_6_r,n_87_7_r,n4_7_r,n2_7_r,n7_7_r;
not I_0(N1372_1_l,n4_1_l);
nor I_1(N1508_1_l,IN_3_1_l,n4_1_l);
nand I_2(n4_1_l,IN_1_1_l,IN_2_1_l);
DFFARX1 I_3(n4_7_l,blif_clk_net_7_r,n2_7_r,G42_7_l,);
not I_4(n_87_7_l,G15_7_l);
nor I_5(n_572_7_l,G15_7_l,IN_7_7_l);
or I_6(n_573_7_l,IN_5_7_l,IN_9_7_l);
nor I_7(n_549_7_l,IN_10_7_l,n7_7_l);
or I_8(n_569_7_l,IN_9_7_l,IN_10_7_l);
nor I_9(n_452_7_l,G18_7_l,IN_5_7_l);
nor I_10(n4_7_l,G18_7_l,IN_1_7_l);
and I_11(n7_7_l,IN_4_7_l,n_87_7_l);
nor I_12(n_42_8_l,IN_1_8_l,IN_3_8_l);
DFFARX1 I_13(N3_8_l,blif_clk_net_7_r,n2_7_r,G199_8_l,);
and I_14(N3_8_l,IN_6_8_l,n3_8_l);
nand I_15(n3_8_l,IN_2_8_l,IN_3_8_l);
nor I_16(N1371_0_r,n4_0_r,n_42_8_l);
nor I_17(N1508_0_r,n3_0_r,n4_0_r);
nor I_18(n3_0_r,n_572_7_l,n_549_7_l);
not I_19(n4_0_r,G199_8_l);
not I_20(N1372_1_r,n4_1_r);
nor I_21(N1508_1_r,n4_1_r,G42_7_l);
nand I_22(n4_1_r,n_572_7_l,n_573_7_l);
nor I_23(N6147_2_r,n5_2_r,n6_2_r);
nor I_24(n5_2_r,n7_2_r,N1508_1_l);
not I_25(n6_2_r,N6138_2_r);
nor I_26(N6138_2_r,n_573_7_l,n_569_7_l);
nor I_27(n7_2_r,N1372_1_l,n_572_7_l);
nor I_28(N1507_6_r,n8_6_r,n9_6_r);
and I_29(N1508_6_r,n6_6_r,G42_7_l);
nor I_30(n6_6_r,n7_6_r,n8_6_r);
not I_31(n7_6_r,N1372_1_l);
nor I_32(n8_6_r,n9_6_r,n_573_7_l);
and I_33(n9_6_r,N1508_1_l,N1372_1_l);
DFFARX1 I_34(n4_7_r,blif_clk_net_7_r,n2_7_r,G42_7_r,);
not I_35(n_87_7_r,n_452_7_l);
nor I_36(n_572_7_r,n_569_7_l,n_452_7_l);
or I_37(n_573_7_r,n_549_7_l,n_42_8_l);
nor I_38(n_549_7_r,n7_7_r,N1508_1_l);
or I_39(n_569_7_r,n_549_7_l,N1508_1_l);
nor I_40(n_452_7_r,G42_7_l,n_42_8_l);
nor I_41(n4_7_r,n_452_7_l,G42_7_l);
not I_42(n2_7_r,blif_reset_net_7_r);
and I_43(n7_7_r,n_87_7_r,G199_8_l);
endmodule


