module test_I15611(I1477,I15611);
input I1477;
output I15611;
wire ;
not I_0(I15611,I1477);
endmodule


