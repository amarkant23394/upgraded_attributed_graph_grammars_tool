module test_final(IN_1_0_l_0,IN_2_0_l_0,IN_4_0_l_0,IN_1_1_l_0,IN_2_1_l_0,IN_3_1_l_0,IN_6_1_l_0,IN_1_5_l_0,IN_2_5_l_0,IN_3_5_l_0,IN_6_5_l_0,blif_clk_net_3_r_10,blif_reset_net_3_r_10,n_429_or_0_3_r_10,G78_3_r_10,n_576_3_r_10,n_102_3_r_10,n_547_3_r_10,G42_4_r_10,n_572_4_r_10,n_573_4_r_10,n_549_4_r_10,n_569_4_r_10,n_452_4_r_10);
input IN_1_0_l_0,IN_2_0_l_0,IN_4_0_l_0,IN_1_1_l_0,IN_2_1_l_0,IN_3_1_l_0,IN_6_1_l_0,IN_1_5_l_0,IN_2_5_l_0,IN_3_5_l_0,IN_6_5_l_0,blif_clk_net_3_r_10,blif_reset_net_3_r_10;
output n_429_or_0_3_r_10,G78_3_r_10,n_576_3_r_10,n_102_3_r_10,n_547_3_r_10,G42_4_r_10,n_572_4_r_10,n_573_4_r_10,n_549_4_r_10,n_569_4_r_10,n_452_4_r_10;
wire n_429_or_0_3_r_0,G78_3_r_0,n_576_3_r_0,n_102_3_r_0,n_547_3_r_0,G42_4_r_0,n_572_4_r_0,n_573_4_r_0,n_549_4_r_0,n_569_4_r_0,n_452_4_r_0,ACVQN2_0_l_0,n_266_and_0_0_l_0,ACVQN1_0_l_0,N1_1_l_0,G199_1_l_0,G214_1_l_0,n3_1_l_0,n_42_5_l_0,N3_5_l_0,G199_5_l_0,n3_5_l_0,n12_3_r_0,n_431_3_r_0,n11_3_r_0,n13_3_r_0,n14_3_r_0,n15_3_r_0,n16_3_r_0,n4_4_r_0,n_87_4_r_0,n7_4_r_0,n2_3_r_10,ACVQN2_0_l_10,n_266_and_0_0_l_10,ACVQN1_0_l_10,n4_4_l_10,G42_4_l_10,n_87_4_l_10,n_572_4_l_10,n_573_4_l_10,n_549_4_l_10,n7_4_l_10,n_569_4_l_10,n_452_4_l_10,n12_3_r_10,n_431_3_r_10,n11_3_r_10,n13_3_r_10,n14_3_r_10,n15_3_r_10,n16_3_r_10,n4_4_r_10,n_87_4_r_10,n7_4_r_10;
nand I_0(n_429_or_0_3_r_0,ACVQN2_0_l_0,n12_3_r_0);
DFFARX1 I_1(n_431_3_r_0,blif_clk_net_3_r_10,n2_3_r_10,G78_3_r_0,);
nand I_2(n_576_3_r_0,n_266_and_0_0_l_0,n11_3_r_0);
not I_3(n_102_3_r_0,n_42_5_l_0);
nand I_4(n_547_3_r_0,ACVQN2_0_l_0,n13_3_r_0);
DFFARX1 I_5(n4_4_r_0,blif_clk_net_3_r_10,n2_3_r_10,G42_4_r_0,);
nor I_6(n_572_4_r_0,G199_1_l_0,G199_5_l_0);
or I_7(n_573_4_r_0,n_42_5_l_0,G199_5_l_0);
nor I_8(n_549_4_r_0,n_266_and_0_0_l_0,n7_4_r_0);
or I_9(n_569_4_r_0,n_266_and_0_0_l_0,n_42_5_l_0);
nor I_10(n_452_4_r_0,ACVQN2_0_l_0,G199_5_l_0);
DFFARX1 I_11(IN_1_0_l_0,blif_clk_net_3_r_10,n2_3_r_10,ACVQN2_0_l_0,);
and I_12(n_266_and_0_0_l_0,IN_4_0_l_0,ACVQN1_0_l_0);
DFFARX1 I_13(IN_2_0_l_0,blif_clk_net_3_r_10,n2_3_r_10,ACVQN1_0_l_0,);
and I_14(N1_1_l_0,IN_6_1_l_0,n3_1_l_0);
DFFARX1 I_15(N1_1_l_0,blif_clk_net_3_r_10,n2_3_r_10,G199_1_l_0,);
DFFARX1 I_16(IN_3_1_l_0,blif_clk_net_3_r_10,n2_3_r_10,G214_1_l_0,);
nand I_17(n3_1_l_0,IN_1_1_l_0,IN_2_1_l_0);
nor I_18(n_42_5_l_0,IN_1_5_l_0,IN_3_5_l_0);
and I_19(N3_5_l_0,IN_6_5_l_0,n3_5_l_0);
DFFARX1 I_20(N3_5_l_0,blif_clk_net_3_r_10,n2_3_r_10,G199_5_l_0,);
nand I_21(n3_5_l_0,IN_2_5_l_0,IN_3_5_l_0);
not I_22(n12_3_r_0,G199_1_l_0);
or I_23(n_431_3_r_0,n_266_and_0_0_l_0,n14_3_r_0);
nor I_24(n11_3_r_0,G214_1_l_0,n12_3_r_0);
nor I_25(n13_3_r_0,G214_1_l_0,n_42_5_l_0);
and I_26(n14_3_r_0,n_42_5_l_0,n15_3_r_0);
nor I_27(n15_3_r_0,G199_1_l_0,n16_3_r_0);
not I_28(n16_3_r_0,ACVQN2_0_l_0);
nor I_29(n4_4_r_0,ACVQN2_0_l_0,G214_1_l_0);
not I_30(n_87_4_r_0,G199_5_l_0);
and I_31(n7_4_r_0,ACVQN2_0_l_0,n_87_4_r_0);
nand I_32(n_429_or_0_3_r_10,n_266_and_0_0_l_10,n12_3_r_10);
DFFARX1 I_33(n_431_3_r_10,blif_clk_net_3_r_10,n2_3_r_10,G78_3_r_10,);
nand I_34(n_576_3_r_10,ACVQN2_0_l_10,n11_3_r_10);
not I_35(n_102_3_r_10,G42_4_l_10);
nand I_36(n_547_3_r_10,n_569_4_l_10,n13_3_r_10);
DFFARX1 I_37(n4_4_r_10,blif_clk_net_3_r_10,n2_3_r_10,G42_4_r_10,);
nor I_38(n_572_4_r_10,ACVQN2_0_l_10,n_573_4_l_10);
or I_39(n_573_4_r_10,n_569_4_l_10,n_452_4_l_10);
nor I_40(n_549_4_r_10,n_572_4_l_10,n7_4_r_10);
or I_41(n_569_4_r_10,n_572_4_l_10,n_569_4_l_10);
nor I_42(n_452_4_r_10,n_266_and_0_0_l_10,n_452_4_l_10);
not I_43(n2_3_r_10,blif_reset_net_3_r_10);
DFFARX1 I_44(n_547_3_r_0,blif_clk_net_3_r_10,n2_3_r_10,ACVQN2_0_l_10,);
and I_45(n_266_and_0_0_l_10,ACVQN1_0_l_10,n_572_4_r_0);
DFFARX1 I_46(n_102_3_r_0,blif_clk_net_3_r_10,n2_3_r_10,ACVQN1_0_l_10,);
nor I_47(n4_4_l_10,n_429_or_0_3_r_0,n_569_4_r_0);
DFFARX1 I_48(n4_4_l_10,blif_clk_net_3_r_10,n2_3_r_10,G42_4_l_10,);
not I_49(n_87_4_l_10,n_452_4_r_0);
nor I_50(n_572_4_l_10,n_549_4_r_0,n_452_4_r_0);
or I_51(n_573_4_l_10,G78_3_r_0,n_573_4_r_0);
nor I_52(n_549_4_l_10,n7_4_l_10,G42_4_r_0);
and I_53(n7_4_l_10,n_87_4_l_10,n_576_3_r_0);
or I_54(n_569_4_l_10,G42_4_r_0,n_573_4_r_0);
nor I_55(n_452_4_l_10,n_429_or_0_3_r_0,G78_3_r_0);
not I_56(n12_3_r_10,n_549_4_l_10);
or I_57(n_431_3_r_10,n_572_4_l_10,n14_3_r_10);
nor I_58(n11_3_r_10,G42_4_l_10,n12_3_r_10);
nor I_59(n13_3_r_10,G42_4_l_10,n_549_4_l_10);
and I_60(n14_3_r_10,ACVQN2_0_l_10,n15_3_r_10);
nor I_61(n15_3_r_10,n_573_4_l_10,n16_3_r_10);
not I_62(n16_3_r_10,n_266_and_0_0_l_10);
nor I_63(n4_4_r_10,n_266_and_0_0_l_10,G42_4_l_10);
not I_64(n_87_4_r_10,ACVQN2_0_l_10);
and I_65(n7_4_r_10,n_452_4_l_10,n_87_4_r_10);
endmodule


