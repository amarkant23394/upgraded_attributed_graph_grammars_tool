module test_I9483(I8202,I1477,I8561,I1470,I9483);
input I8202,I1477,I8561,I1470;
output I9483;
wire I9508,I9542,I8216,I8199,I8623,I9816,I8705,I8184,I9525,I8193,I9491;
nand I_0(I9508,I8199,I8202);
DFFARX1 I_1(I9525,I1470,I9491,,,I9542,);
not I_2(I8216,I1477);
DFFARX1 I_3(I1470,I8216,,,I8199,);
DFFARX1 I_4(I1470,I8216,,,I8623,);
DFFARX1 I_5(I8193,I1470,I9491,,,I9816,);
DFFARX1 I_6(I8623,I1470,I8216,,,I8705,);
nor I_7(I9483,I9816,I9542);
DFFARX1 I_8(I8561,I1470,I8216,,,I8184,);
and I_9(I9525,I9508,I8184);
not I_10(I8193,I8705);
not I_11(I9491,I1477);
endmodule


