module test_I2730(I1447,I1477,I1470,I2730);
input I1447,I1477,I1470;
output I2730;
wire I2759,I3076;
not I_0(I2730,I3076);
not I_1(I2759,I1477);
DFFARX1 I_2(I1447,I1470,I2759,,,I3076,);
endmodule


