module test_I7799(I6640,I1477,I6363,I1470,I6705,I7799);
input I6640,I1477,I6363,I1470,I6705;
output I7799;
wire I6781,I7765,I6722,I6329,I6380,I7782,I6312,I6411,I6291,I6303,I7748,I6306;
DFFARX1 I_0(I1470,I6329,,,I6781,);
or I_1(I7799,I7782,I6306);
nor I_2(I7765,I7748,I6303);
or I_3(I6722,I6705,I6640);
not I_4(I6329,I1477);
DFFARX1 I_5(I6363,I1470,I6329,,,I6380,);
and I_6(I7782,I7765,I6312);
DFFARX1 I_7(I6722,I1470,I6329,,,I6312,);
DFFARX1 I_8(I6380,I1470,I6329,,,I6411,);
DFFARX1 I_9(I6705,I1470,I6329,,,I6291,);
DFFARX1 I_10(I6781,I1470,I6329,,,I6303,);
not I_11(I7748,I6291);
not I_12(I6306,I6411);
endmodule


