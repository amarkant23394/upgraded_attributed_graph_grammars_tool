module test_I11491(I9131,I1477,I1470,I8964,I6896,I11491);
input I9131,I1477,I1470,I8964,I6896;
output I11491;
wire I9148,I8827,I8862,I9179,I9258;
and I_0(I9148,I8964,I9131);
not I_1(I11491,I8827);
DFFARX1 I_2(I9258,I1470,I8862,,,I8827,);
not I_3(I8862,I1477);
DFFARX1 I_4(I6896,I1470,I8862,,,I9179,);
or I_5(I9258,I9179,I9148);
endmodule


