module test_I17092(I14982,I1477,I1470,I17092);
input I14982,I1477,I1470;
output I17092;
wire I12619,I12670,I12584,I15047,I15064,I14954,I16818,I12587;
not I_0(I12619,I1477);
DFFARX1 I_1(I1470,I12619,,,I12670,);
and I_2(I12584,I12670);
nor I_3(I15047,I14982,I12584);
nand I_4(I15064,I15047,I12587);
not I_5(I14954,I15064);
DFFARX1 I_6(I14954,I1470,I16818,,,I17092,);
not I_7(I16818,I1477);
DFFARX1 I_8(I12670,I1470,I12619,,,I12587,);
endmodule


