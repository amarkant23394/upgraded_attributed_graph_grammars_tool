module test_I1475(I1271,I1247,I1475);
input I1271,I1247;
output I1475;
wire ;
nand I_0(I1475,I1247,I1271);
endmodule


