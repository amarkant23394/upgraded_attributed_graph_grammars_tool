module test_final(IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_4_l_4,IN_2_4_l_4,IN_3_4_l_4,IN_4_4_l_4,IN_5_4_l_4,IN_1_9_l_4,IN_2_9_l_4,IN_3_9_l_4,IN_4_9_l_4,IN_5_9_l_4,blif_clk_net_5_r_9,blif_reset_net_5_r_9,N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,G78_5_r_9,n_576_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9);
input IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_4_l_4,IN_2_4_l_4,IN_3_4_l_4,IN_4_4_l_4,IN_5_4_l_4,IN_1_9_l_4,IN_2_9_l_4,IN_3_9_l_4,IN_4_9_l_4,IN_5_9_l_4,blif_clk_net_5_r_9,blif_reset_net_5_r_9;
output N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,G78_5_r_9,n_576_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9;
wire N1371_0_r_4,N1508_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_573_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6147_9_r_4,N6134_9_r_4,I_BUFF_1_9_r_4,n4_7_r_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4,n38_4,n39_4,n40_4,n41_4,n_429_or_0_5_r_9,n_102_5_r_9,I_BUFF_1_9_r_9,n4_7_l_9,n10_9,n62_9,N3_8_l_9,n63_9,n38_9,n_431_5_r_9,N3_8_r_9,n39_9,n40_9,n41_9,n42_9,n43_9,n44_9,n45_9,n46_9,n47_9,n48_9,n49_9,n50_9,n51_9,n52_9,n53_9,n54_9,n55_9,n56_9,n57_9,n58_9,n59_9,n60_9,n61_9;
nor I_0(N1371_0_r_4,IN_1_9_l_4,n25_4);
not I_1(N1508_0_r_4,n25_4);
nor I_2(N1507_6_r_4,n32_4,n33_4);
nor I_3(N1508_6_r_4,n22_4,n29_4);
DFFARX1 I_4(n4_7_r_4,blif_clk_net_5_r_9,n10_9,G42_7_r_4,);
not I_5(n_572_7_r_4,n_573_7_r_4);
nand I_6(n_573_7_r_4,n21_4,n22_4);
nor I_7(n_549_7_r_4,IN_1_9_l_4,n24_4);
nand I_8(n_569_7_r_4,n22_4,n23_4);
nor I_9(n_452_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4);
not I_10(N6147_9_r_4,n28_4);
nor I_11(N6134_9_r_4,N1508_0_r_4,n28_4);
not I_12(I_BUFF_1_9_r_4,n21_4);
nor I_13(n4_7_r_4,IN_1_9_l_4,N6147_9_r_4);
nand I_14(n21_4,n39_4,n40_4);
or I_15(n22_4,IN_5_9_l_4,n31_4);
not I_16(n23_4,IN_1_9_l_4);
nor I_17(n24_4,n25_4,n26_4);
nand I_18(n25_4,IN_1_4_l_4,IN_2_4_l_4);
nand I_19(n26_4,n21_4,n27_4);
nand I_20(n27_4,n36_4,n37_4);
nand I_21(n28_4,IN_2_9_l_4,n38_4);
nand I_22(n29_4,N1508_0_r_4,n30_4);
nand I_23(n30_4,n34_4,n35_4);
nor I_24(n31_4,IN_3_9_l_4,IN_4_9_l_4);
not I_25(n32_4,n30_4);
nor I_26(n33_4,n21_4,n28_4);
nand I_27(n34_4,N6147_9_r_4,I_BUFF_1_9_r_4);
nand I_28(n35_4,N1508_0_r_4,n27_4);
not I_29(n36_4,IN_5_4_l_4);
nand I_30(n37_4,IN_3_4_l_4,IN_4_4_l_4);
or I_31(n38_4,IN_3_9_l_4,IN_4_9_l_4);
nor I_32(n39_4,IN_1_2_l_4,IN_2_2_l_4);
or I_33(n40_4,IN_5_2_l_4,n41_4);
nor I_34(n41_4,IN_3_2_l_4,IN_4_2_l_4);
nor I_35(N6147_2_r_9,n62_9,n46_9);
not I_36(N1372_4_r_9,n59_9);
nor I_37(N1508_4_r_9,n58_9,n59_9);
nand I_38(n_429_or_0_5_r_9,n_431_5_r_9,n42_9);
DFFARX1 I_39(n_431_5_r_9,blif_clk_net_5_r_9,n10_9,G78_5_r_9,);
nand I_40(n_576_5_r_9,n39_9,n40_9);
not I_41(n_102_5_r_9,I_BUFF_1_9_r_9);
nand I_42(n_547_5_r_9,n43_9,N1507_6_r_4);
and I_43(n_42_8_r_9,n44_9,n_549_7_r_4);
DFFARX1 I_44(N3_8_r_9,blif_clk_net_5_r_9,n10_9,G199_8_r_9,);
nor I_45(N6147_9_r_9,n41_9,n45_9);
nor I_46(N6134_9_r_9,n45_9,n51_9);
nor I_47(I_BUFF_1_9_r_9,n41_9,N1507_6_r_4);
nor I_48(n4_7_l_9,n_549_7_r_4,n_572_7_r_4);
not I_49(n10_9,blif_reset_net_5_r_9);
DFFARX1 I_50(n4_7_l_9,blif_clk_net_5_r_9,n10_9,n62_9,);
and I_51(N3_8_l_9,n57_9,G42_7_r_4);
DFFARX1 I_52(N3_8_l_9,blif_clk_net_5_r_9,n10_9,n63_9,);
not I_53(n38_9,n63_9);
nor I_54(n_431_5_r_9,N6134_9_r_4,N1508_6_r_4);
nor I_55(N3_8_r_9,n_102_5_r_9,n53_9);
nor I_56(n39_9,I_BUFF_1_9_r_9,n42_9);
not I_57(n40_9,n41_9);
nand I_58(n41_9,N1371_0_r_4,n_549_7_r_4);
nor I_59(n42_9,n_452_7_r_4,N1507_6_r_4);
nor I_60(n43_9,n63_9,n41_9);
nor I_61(n44_9,n_452_7_r_4,G42_7_r_4);
and I_62(n45_9,n52_9,n_569_7_r_4);
nor I_63(n46_9,n47_9,n48_9);
nor I_64(n47_9,n49_9,n50_9);
not I_65(n48_9,n_429_or_0_5_r_9);
not I_66(n49_9,n42_9);
or I_67(n50_9,n63_9,n51_9);
nor I_68(n51_9,N1371_0_r_4,N1508_6_r_4);
nor I_69(n52_9,n49_9,N1508_6_r_4);
nor I_70(n53_9,n54_9,n55_9);
nor I_71(n54_9,n56_9,N1508_6_r_4);
or I_72(n55_9,n44_9,N1507_6_r_4);
not I_73(n56_9,n_569_7_r_4);
nand I_74(n57_9,N1508_6_r_4,n_572_7_r_4);
nor I_75(n58_9,n62_9,n60_9);
nand I_76(n59_9,n51_9,n61_9);
nor I_77(n60_9,n38_9,n44_9);
nor I_78(n61_9,n_549_7_r_4,G42_7_r_4);
endmodule


