module test_final(IN_1_0_l_1,IN_2_0_l_1,IN_3_0_l_1,IN_4_0_l_1,IN_1_1_l_1,IN_2_1_l_1,IN_3_1_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_3_3_l_1,IN_1_6_l_1,IN_2_6_l_1,IN_3_6_l_1,IN_4_6_l_1,IN_5_6_l_1,blif_clk_net_7_r_12,blif_reset_net_7_r_12,N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_549_7_r_12,n_569_7_r_12,N6147_9_r_12);
input IN_1_0_l_1,IN_2_0_l_1,IN_3_0_l_1,IN_4_0_l_1,IN_1_1_l_1,IN_2_1_l_1,IN_3_1_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_3_3_l_1,IN_1_6_l_1,IN_2_6_l_1,IN_3_6_l_1,IN_4_6_l_1,IN_5_6_l_1,blif_clk_net_7_r_12,blif_reset_net_7_r_12;
output N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_549_7_r_12,n_569_7_r_12,N6147_9_r_12;
wire N1371_0_r_1,N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,n_452_7_r_1,N6147_9_r_1,N6134_9_r_1,I_BUFF_1_9_r_1,n4_7_r_1,n29_1,n30_1,n31_1,n32_1,n33_1,n34_1,n35_1,n36_1,n37_1,n38_1,n39_1,n40_1,n41_1,n42_1,n43_1,n44_1,n45_1,n46_1,n47_1,n48_1,n49_1,n50_1,n51_1,n52_1,n53_1,n54_1,n55_1,n_573_7_r_12,n_452_7_r_12,N6134_9_r_12,I_BUFF_1_9_r_12,n1_12,n8_12,n23_12,n24_12,n25_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12,n41_12,n42_12;
and I_0(N1371_0_r_1,I_BUFF_1_9_r_1,n55_1);
nor I_1(N1508_0_r_1,n40_1,n44_1);
nor I_2(N1507_6_r_1,n43_1,n49_1);
nor I_3(N1508_6_r_1,n41_1,n42_1);
DFFARX1 I_4(n4_7_r_1,blif_clk_net_7_r_12,n8_12,G42_7_r_1,);
nor I_5(n_572_7_r_1,n29_1,n30_1);
not I_6(n_573_7_r_1,n_452_7_r_1);
nor I_7(n_549_7_r_1,N1371_0_r_1,n31_1);
or I_8(n_569_7_r_1,n30_1,n31_1);
nor I_9(n_452_7_r_1,n30_1,n32_1);
nor I_10(N6147_9_r_1,n35_1,n36_1);
nand I_11(N6134_9_r_1,n38_1,n39_1);
not I_12(I_BUFF_1_9_r_1,n40_1);
nor I_13(n4_7_r_1,I_BUFF_1_9_r_1,n30_1);
nor I_14(n29_1,IN_2_0_l_1,n34_1);
nor I_15(n30_1,n33_1,n34_1);
nor I_16(n31_1,IN_1_3_l_1,n54_1);
not I_17(n32_1,n48_1);
nor I_18(n33_1,IN_3_0_l_1,IN_4_0_l_1);
not I_19(n34_1,IN_1_0_l_1);
nor I_20(n35_1,I_BUFF_1_9_r_1,n37_1);
not I_21(n36_1,n29_1);
not I_22(n37_1,n41_1);
nand I_23(n38_1,IN_3_1_l_1,I_BUFF_1_9_r_1);
nand I_24(n39_1,n37_1,n40_1);
nand I_25(n40_1,IN_1_1_l_1,IN_2_1_l_1);
nand I_26(n41_1,IN_5_6_l_1,n52_1);
or I_27(n42_1,n36_1,n43_1);
nor I_28(n43_1,n32_1,n49_1);
nand I_29(n44_1,n45_1,n46_1);
nand I_30(n45_1,n47_1,n48_1);
not I_31(n46_1,IN_3_1_l_1);
not I_32(n47_1,n31_1);
nand I_33(n48_1,IN_2_6_l_1,n50_1);
nor I_34(n49_1,n41_1,n47_1);
and I_35(n50_1,IN_1_6_l_1,n51_1);
nand I_36(n51_1,n52_1,n53_1);
nand I_37(n52_1,IN_3_6_l_1,IN_4_6_l_1);
not I_38(n53_1,IN_5_6_l_1);
or I_39(n54_1,IN_2_3_l_1,IN_3_3_l_1);
nor I_40(n55_1,IN_3_1_l_1,n29_1);
nor I_41(N1371_0_r_12,I_BUFF_1_9_r_12,n36_12);
nand I_42(N1508_0_r_12,n30_12,n37_12);
nor I_43(N1507_6_r_12,n25_12,n39_12);
nor I_44(N1508_6_r_12,n25_12,n29_12);
DFFARX1 I_45(n1_12,blif_clk_net_7_r_12,n8_12,G42_7_r_12,);
nor I_46(n_572_7_r_12,n23_12,n24_12);
nand I_47(n_573_7_r_12,n_452_7_r_12,n25_12);
nand I_48(n_549_7_r_12,n27_12,n28_12);
nand I_49(n_569_7_r_12,n25_12,n26_12);
nand I_50(n_452_7_r_12,N1507_6_r_1,N1508_6_r_1);
nand I_51(N6147_9_r_12,n30_12,n31_12);
nor I_52(N6134_9_r_12,n35_12,n36_12);
not I_53(I_BUFF_1_9_r_12,n_452_7_r_12);
not I_54(n1_12,n_573_7_r_12);
not I_55(n8_12,blif_reset_net_7_r_12);
not I_56(n23_12,n36_12);
nor I_57(n24_12,n_452_7_r_12,n_573_7_r_1);
nand I_58(n25_12,n23_12,n40_12);
not I_59(n26_12,n35_12);
not I_60(n27_12,N6134_9_r_12);
nand I_61(n28_12,n26_12,n29_12);
not I_62(n29_12,n24_12);
nand I_63(n30_12,n33_12,n41_12);
nand I_64(n31_12,n32_12,n33_12);
nor I_65(n32_12,n26_12,n34_12);
nor I_66(n33_12,n_572_7_r_1,n_573_7_r_1);
nor I_67(n34_12,n42_12,N6134_9_r_1);
nor I_68(n35_12,n38_12,G42_7_r_1);
nand I_69(n36_12,G42_7_r_1,n_549_7_r_1);
nand I_70(n37_12,n23_12,n35_12);
or I_71(n38_12,N1508_0_r_1,N1508_6_r_1);
not I_72(n39_12,n30_12);
or I_73(n40_12,n_569_7_r_1,N1507_6_r_1);
nor I_74(n41_12,n34_12,n36_12);
nor I_75(n42_12,N1508_0_r_1,N6147_9_r_1);
endmodule


