module test_final(IN_1_2_l_3,IN_2_2_l_3,IN_3_2_l_3,IN_4_2_l_3,IN_5_2_l_3,IN_1_6_l_3,IN_2_6_l_3,IN_3_6_l_3,IN_4_6_l_3,IN_5_6_l_3,IN_1_9_l_3,IN_2_9_l_3,IN_3_9_l_3,IN_4_9_l_3,IN_5_9_l_3,blif_clk_net_5_r_7,blif_reset_net_5_r_7,N1371_0_r_7,N1508_0_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_547_5_r_7,G42_7_r_7,n_572_7_r_7,n_573_7_r_7,n_549_7_r_7,n_569_7_r_7);
input IN_1_2_l_3,IN_2_2_l_3,IN_3_2_l_3,IN_4_2_l_3,IN_5_2_l_3,IN_1_6_l_3,IN_2_6_l_3,IN_3_6_l_3,IN_4_6_l_3,IN_5_6_l_3,IN_1_9_l_3,IN_2_9_l_3,IN_3_9_l_3,IN_4_9_l_3,IN_5_9_l_3,blif_clk_net_5_r_7,blif_reset_net_5_r_7;
output N1371_0_r_7,N1508_0_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_547_5_r_7,G42_7_r_7,n_572_7_r_7,n_573_7_r_7,n_549_7_r_7,n_569_7_r_7;
wire N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_572_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6147_9_r_3,N6134_9_r_3,I_BUFF_1_9_r_3,n4_7_r_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3,n40_3,n41_3,n42_3,n43_3,n44_3,n45_3,n46_3,n47_3,n48_3,n49_3,n50_3,n51_3,n_102_5_r_7,n_452_7_r_7,n4_7_l_7,n6_7,n53_7,n30_7,N3_8_l_7,n54_7,n_431_5_r_7,n4_7_r_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7,n43_7,n44_7,n45_7,n46_7,n47_7,n48_7,n49_7,n50_7,n51_7,n52_7;
not I_0(N1372_1_r_3,n40_3);
nor I_1(N1508_1_r_3,N6147_9_r_3,n40_3);
nor I_2(N1507_6_r_3,n31_3,n42_3);
nor I_3(N1508_6_r_3,n30_3,n38_3);
DFFARX1 I_4(n4_7_r_3,blif_clk_net_5_r_7,n6_7,G42_7_r_3,);
nor I_5(n_572_7_r_3,I_BUFF_1_9_r_3,n35_3);
nand I_6(n_573_7_r_3,n30_3,n31_3);
nor I_7(n_549_7_r_3,N6147_9_r_3,n33_3);
nand I_8(n_569_7_r_3,n30_3,n32_3);
nor I_9(n_452_7_r_3,IN_1_9_l_3,n35_3);
not I_10(N6147_9_r_3,n32_3);
nor I_11(N6134_9_r_3,n36_3,n37_3);
not I_12(I_BUFF_1_9_r_3,n45_3);
nor I_13(n4_7_r_3,IN_1_9_l_3,I_BUFF_1_9_r_3);
not I_14(n30_3,n39_3);
not I_15(n31_3,n35_3);
nand I_16(n32_3,IN_5_6_l_3,n41_3);
nor I_17(n33_3,I_BUFF_1_9_r_3,n34_3);
nand I_18(n34_3,IN_2_6_l_3,n46_3);
nor I_19(n35_3,n43_3,n44_3);
not I_20(n36_3,n34_3);
nor I_21(n37_3,IN_1_9_l_3,N6147_9_r_3);
or I_22(n38_3,n_572_7_r_3,n34_3);
nor I_23(n39_3,IN_5_9_l_3,n44_3);
nand I_24(n40_3,IN_1_9_l_3,n39_3);
nand I_25(n41_3,IN_3_6_l_3,IN_4_6_l_3);
nor I_26(n42_3,n34_3,n45_3);
not I_27(n43_3,IN_2_9_l_3);
nor I_28(n44_3,IN_3_9_l_3,IN_4_9_l_3);
nand I_29(n45_3,n49_3,n50_3);
and I_30(n46_3,IN_1_6_l_3,n47_3);
nand I_31(n47_3,n41_3,n48_3);
not I_32(n48_3,IN_5_6_l_3);
nor I_33(n49_3,IN_1_2_l_3,IN_2_2_l_3);
or I_34(n50_3,IN_5_2_l_3,n51_3);
nor I_35(n51_3,IN_3_2_l_3,IN_4_2_l_3);
nor I_36(N1371_0_r_7,n53_7,n52_7);
nor I_37(N1508_0_r_7,n51_7,n52_7);
nand I_38(n_429_or_0_5_r_7,n43_7,n48_7);
DFFARX1 I_39(n_431_5_r_7,blif_clk_net_5_r_7,n6_7,G78_5_r_7,);
nand I_40(n_576_5_r_7,n31_7,n32_7);
nor I_41(n_102_5_r_7,n_549_7_r_3,N1508_6_r_3);
nand I_42(n_547_5_r_7,n31_7,n38_7);
DFFARX1 I_43(n4_7_r_7,blif_clk_net_5_r_7,n6_7,G42_7_r_7,);
nor I_44(n_572_7_r_7,n54_7,n33_7);
nand I_45(n_573_7_r_7,n_102_5_r_7,n_452_7_r_7);
nor I_46(n_549_7_r_7,n53_7,n36_7);
nand I_47(n_569_7_r_7,n_102_5_r_7,n30_7);
nand I_48(n_452_7_r_7,G42_7_r_3,n_452_7_r_3);
nor I_49(n4_7_l_7,N1508_1_r_3,N1508_6_r_3);
not I_50(n6_7,blif_reset_net_5_r_7);
DFFARX1 I_51(n4_7_l_7,blif_clk_net_5_r_7,n6_7,n53_7,);
not I_52(n30_7,n53_7);
and I_53(N3_8_l_7,n50_7,G42_7_r_3);
DFFARX1 I_54(N3_8_l_7,blif_clk_net_5_r_7,n6_7,n54_7,);
nand I_55(n_431_5_r_7,n40_7,n41_7);
nor I_56(n4_7_r_7,n54_7,n49_7);
and I_57(n31_7,n_102_5_r_7,n39_7);
not I_58(n32_7,N1508_6_r_3);
nor I_59(n33_7,n34_7,N1372_1_r_3);
and I_60(n34_7,n35_7,n_569_7_r_3);
not I_61(n35_7,N1507_6_r_3);
nor I_62(n36_7,n37_7,N1508_6_r_3);
or I_63(n37_7,n54_7,N1508_6_r_3);
or I_64(n38_7,N1372_1_r_3,n_573_7_r_3);
nor I_65(n39_7,n_452_7_r_7,N1507_6_r_3);
nand I_66(n40_7,n46_7,n47_7);
nand I_67(n41_7,n42_7,n43_7);
nor I_68(n42_7,n44_7,n45_7);
nor I_69(n43_7,N1372_1_r_3,n_573_7_r_3);
nor I_70(n44_7,N1507_6_r_3,N6134_9_r_3);
nor I_71(n45_7,n_549_7_r_3,N1372_1_r_3);
nand I_72(n46_7,n35_7,n_569_7_r_3);
not I_73(n47_7,N1372_1_r_3);
or I_74(n48_7,n_452_7_r_7,N1507_6_r_3);
not I_75(n49_7,n_452_7_r_7);
nand I_76(n50_7,n_573_7_r_3,N1508_1_r_3);
and I_77(n51_7,n_452_7_r_7,n45_7);
not I_78(n52_7,n44_7);
endmodule


