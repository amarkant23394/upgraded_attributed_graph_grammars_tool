module test_I17157(I15064,I1477,I15276,I15109,I14942,I1470,I17157);
input I15064,I1477,I15276,I15109,I14942,I1470;
output I17157;
wire I14954,I15310,I14965,I17047,I17013,I17030,I14933,I14939,I17092,I16818,I17109,I14930,I15293,I15341;
not I_0(I14954,I15064);
and I_1(I15310,I15276,I15293);
not I_2(I14965,I1477);
nand I_3(I17157,I17109,I17047);
DFFARX1 I_4(I17030,I1470,I16818,,,I17047,);
nand I_5(I17013,I14942,I14939);
and I_6(I17030,I17013,I14930);
DFFARX1 I_7(I15310,I1470,I14965,,,I14933,);
DFFARX1 I_8(I1470,I14965,,,I14939,);
DFFARX1 I_9(I14954,I1470,I16818,,,I17092,);
not I_10(I16818,I1477);
and I_11(I17109,I17092,I14933);
and I_12(I14930,I15109,I15341);
nand I_13(I15293,I15276);
DFFARX1 I_14(I15276,I1470,I14965,,,I15341,);
endmodule


