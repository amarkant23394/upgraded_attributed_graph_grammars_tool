module test_final(IN_1_1_l_2,IN_2_1_l_2,IN_3_1_l_2,G18_7_l_2,G15_7_l_2,IN_1_7_l_2,IN_4_7_l_2,IN_5_7_l_2,IN_7_7_l_2,IN_9_7_l_2,IN_10_7_l_2,IN_1_8_l_2,IN_2_8_l_2,IN_3_8_l_2,IN_6_8_l_2,blif_clk_net_7_r_5,blif_reset_net_7_r_5,N1371_0_r_5,N1508_0_r_5,N1372_1_r_5,N1508_1_r_5,N6147_2_r_5,N1507_6_r_5,N1508_6_r_5,G42_7_r_5,n_572_7_r_5,n_573_7_r_5,n_569_7_r_5,n_452_7_r_5);
input IN_1_1_l_2,IN_2_1_l_2,IN_3_1_l_2,G18_7_l_2,G15_7_l_2,IN_1_7_l_2,IN_4_7_l_2,IN_5_7_l_2,IN_7_7_l_2,IN_9_7_l_2,IN_10_7_l_2,IN_1_8_l_2,IN_2_8_l_2,IN_3_8_l_2,IN_6_8_l_2,blif_clk_net_7_r_5,blif_reset_net_7_r_5;
output N1371_0_r_5,N1508_0_r_5,N1372_1_r_5,N1508_1_r_5,N6147_2_r_5,N1507_6_r_5,N1508_6_r_5,G42_7_r_5,n_572_7_r_5,n_573_7_r_5,n_569_7_r_5,n_452_7_r_5;
wire N1371_0_r_2,N1508_0_r_2,N1372_1_r_2,N1508_1_r_2,N6147_2_r_2,N1507_6_r_2,N1508_6_r_2,G42_7_r_2,n_572_7_r_2,n_573_7_r_2,n_549_7_r_2,n_569_7_r_2,n_452_7_r_2,n4_7_l_2,n59_2,n33_2,N3_8_l_2,n32_internal_2,n32_2,n4_7_r_2,n34_2,n35_2,n36_2,n37_2,n38_2,n39_2,n40_2,n41_2,n42_2,n43_2,n44_2,n45_2,n46_2,n47_2,n48_2,n49_2,n50_2,n51_2,n52_2,n53_2,n54_2,n55_2,n56_2,n57_2,n58_2,n_549_7_r_5,n4_7_r_5,n7_5,n26_5,n27_5,n28_5,n29_5,n30_5,n31_5,n32_5,n33_5,n34_5,n35_5,n36_5,n37_5,n38_5,n39_5,n40_5,n41_5,n42_5,n43_5,n44_5,n45_5,n46_5,n47_5;
nor I_0(N1371_0_r_2,n32_2,n35_2);
nor I_1(N1508_0_r_2,n32_2,n55_2);
not I_2(N1372_1_r_2,n54_2);
nor I_3(N1508_1_r_2,n59_2,n54_2);
nor I_4(N6147_2_r_2,n42_2,n43_2);
nor I_5(N1507_6_r_2,n40_2,n53_2);
nor I_6(N1508_6_r_2,n33_2,n50_2);
DFFARX1 I_7(n4_7_r_2,blif_clk_net_7_r_5,n7_5,G42_7_r_2,);
nor I_8(n_572_7_r_2,n36_2,n37_2);
or I_9(n_573_7_r_2,n34_2,n35_2);
nor I_10(n_549_7_r_2,n40_2,n41_2);
nand I_11(n_569_7_r_2,n38_2,n39_2);
nor I_12(n_452_7_r_2,n59_2,n35_2);
nor I_13(n4_7_l_2,G18_7_l_2,IN_1_7_l_2);
DFFARX1 I_14(n4_7_l_2,blif_clk_net_7_r_5,n7_5,n59_2,);
not I_15(n33_2,n59_2);
and I_16(N3_8_l_2,IN_6_8_l_2,n49_2);
DFFARX1 I_17(N3_8_l_2,blif_clk_net_7_r_5,n7_5,n32_internal_2,);
not I_18(n32_2,n32_internal_2);
nor I_19(n4_7_r_2,n59_2,n36_2);
not I_20(n34_2,n39_2);
nor I_21(n35_2,IN_1_8_l_2,IN_3_8_l_2);
nor I_22(n36_2,G18_7_l_2,IN_5_7_l_2);
or I_23(n37_2,IN_9_7_l_2,IN_10_7_l_2);
not I_24(n38_2,n40_2);
nand I_25(n39_2,n45_2,n57_2);
nor I_26(n40_2,IN_3_1_l_2,n47_2);
nor I_27(n41_2,n32_2,n36_2);
not I_28(n42_2,n53_2);
nand I_29(n43_2,n44_2,n45_2);
nand I_30(n44_2,n38_2,n46_2);
not I_31(n45_2,IN_10_7_l_2);
nand I_32(n46_2,n47_2,n48_2);
nand I_33(n47_2,IN_1_1_l_2,IN_2_1_l_2);
or I_34(n48_2,G15_7_l_2,IN_7_7_l_2);
nand I_35(n49_2,IN_2_8_l_2,IN_3_8_l_2);
nand I_36(n50_2,n51_2,n52_2);
not I_37(n51_2,n47_2);
nand I_38(n52_2,n38_2,n53_2);
nor I_39(n53_2,IN_5_7_l_2,IN_9_7_l_2);
nand I_40(n54_2,n42_2,n56_2);
nor I_41(n55_2,n34_2,n56_2);
nor I_42(n56_2,G15_7_l_2,IN_7_7_l_2);
nand I_43(n57_2,IN_4_7_l_2,n58_2);
not I_44(n58_2,G15_7_l_2);
nor I_45(N1371_0_r_5,n28_5,n46_5);
nand I_46(N1508_0_r_5,n26_5,n43_5);
not I_47(N1372_1_r_5,n43_5);
nor I_48(N1508_1_r_5,n30_5,n43_5);
nor I_49(N6147_2_r_5,n29_5,n32_5);
nor I_50(N1507_6_r_5,n26_5,n44_5);
nor I_51(N1508_6_r_5,n27_5,n37_5);
DFFARX1 I_52(n4_7_r_5,blif_clk_net_7_r_5,n7_5,G42_7_r_5,);
and I_53(n_572_7_r_5,n27_5,n28_5);
nand I_54(n_573_7_r_5,n26_5,n27_5);
nand I_55(n_549_7_r_5,N1508_0_r_2,n_549_7_r_2);
nand I_56(n_569_7_r_5,n_549_7_r_5,n26_5);
not I_57(n_452_7_r_5,n29_5);
nor I_58(n4_7_r_5,n30_5,n31_5);
not I_59(n7_5,blif_reset_net_7_r_5);
not I_60(n26_5,n35_5);
nand I_61(n27_5,n40_5,n41_5);
nand I_62(n28_5,N1371_0_r_2,n_452_7_r_2);
nand I_63(n29_5,n27_5,n33_5);
nor I_64(n30_5,n45_5,N1508_6_r_2);
not I_65(n31_5,n_549_7_r_5);
nor I_66(n32_5,n34_5,n35_5);
not I_67(n33_5,n30_5);
nor I_68(n34_5,n31_5,n36_5);
nor I_69(n35_5,n28_5,N1508_0_r_2);
not I_70(n36_5,n28_5);
nand I_71(n37_5,n36_5,n38_5);
nand I_72(n38_5,n26_5,n39_5);
nand I_73(n39_5,n30_5,n31_5);
nor I_74(n40_5,N1372_1_r_2,n_569_7_r_2);
or I_75(n41_5,n42_5,N1371_0_r_2);
nor I_76(n42_5,N1508_1_r_2,n_572_7_r_2);
nand I_77(n43_5,n36_5,n46_5);
nor I_78(n44_5,n_549_7_r_5,n33_5);
or I_79(n45_5,N6147_2_r_2,n_573_7_r_2);
and I_80(n46_5,n31_5,n47_5);
or I_81(n47_5,N1507_6_r_2,G42_7_r_2);
endmodule


