module test_I4979(I1477,I1470,I2695,I2146,I4979);
input I1477,I1470,I2695,I2146;
output I4979;
wire I2181,I4544,I4869,I2149,I4962,I4708,I4742,I4725,I2164,I2263,I2158;
nor I_0(I4979,I4742,I4962);
not I_1(I2181,I1477);
not I_2(I4544,I1477);
DFFARX1 I_3(I2149,I1470,I4544,,,I4869,);
DFFARX1 I_4(I2695,I1470,I2181,,,I2149,);
not I_5(I4962,I4869);
nand I_6(I4708,I2146,I2164);
DFFARX1 I_7(I4725,I1470,I4544,,,I4742,);
and I_8(I4725,I4708,I2158);
DFFARX1 I_9(I1470,I2181,,,I2164,);
DFFARX1 I_10(I1470,I2181,,,I2263,);
not I_11(I2158,I2263);
endmodule


