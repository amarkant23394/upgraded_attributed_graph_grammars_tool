module test_I14438(I11296,I11429,I1477,I1470,I11395,I14438);
input I11296,I11429,I1477,I1470,I11395;
output I14438;
wire I13601,I13197,I11299,I11768,I11272,I13186,I13508,I13491,I11310,I13159;
DFFARX1 I_0(I11299,I1470,I13197,,,I13601,);
not I_1(I13197,I1477);
nor I_2(I11299,I11395,I11429);
and I_3(I11768,I11429);
DFFARX1 I_4(I11768,I1470,I11310,,,I11272,);
nor I_5(I13186,I13601,I13508);
and I_6(I13508,I13491,I11272);
DFFARX1 I_7(I11296,I1470,I13197,,,I13491,);
not I_8(I11310,I1477);
DFFARX1 I_9(I13508,I1470,I13197,,,I13159,);
nor I_10(I14438,I13159,I13186);
endmodule


