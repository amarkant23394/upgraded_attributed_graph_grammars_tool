module test_I10459(I8107,I1477,I6321,I7714,I10086,I1470,I7915,I10459);
input I8107,I1477,I6321,I7714,I10086,I1470,I7915;
output I10459;
wire I10253,I10120,I7538,I10219,I7532,I7731,I10052,I7977,I10349,I7946,I10236,I7535,I10332,I10270,I7550,I7570,I10103;
nor I_0(I10253,I10103,I10236);
nor I_1(I10120,I7538,I7535);
DFFARX1 I_2(I7915,I1470,I7570,,,I7538,);
DFFARX1 I_3(I1470,I10052,,,I10219,);
DFFARX1 I_4(I8107,I1470,I7570,,,I7532,);
not I_5(I7731,I7714);
not I_6(I10052,I1477);
DFFARX1 I_7(I6321,I1470,I7570,,,I7977,);
and I_8(I10349,I10332,I7550);
DFFARX1 I_9(I1470,I7570,,,I7946,);
not I_10(I10236,I10219);
and I_11(I7535,I7714,I7946);
DFFARX1 I_12(I7532,I1470,I10052,,,I10332,);
or I_13(I10459,I10349,I10270);
and I_14(I10270,I10120,I10253);
nand I_15(I7550,I7977,I7731);
not I_16(I7570,I1477);
DFFARX1 I_17(I10086,I1470,I10052,,,I10103,);
endmodule


