module test_I9049(I1477,I7461,I5070,I1470,I6881,I6958,I9049);
input I1477,I7461,I5070,I1470,I6881,I6958;
output I9049;
wire I8998,I9032,I7365,I7026,I5067,I9015,I6907,I7348,I7269,I6890,I6899,I6869;
not I_0(I8998,I6881);
and I_1(I9032,I9015,I6890);
or I_2(I9049,I9032,I6869);
and I_3(I7365,I7026,I7348);
not I_4(I7026,I5070);
DFFARX1 I_5(I1470,,,I5067,);
nor I_6(I9015,I8998,I6899);
not I_7(I6907,I1477);
nand I_8(I7348,I7269,I6958);
DFFARX1 I_9(I5067,I1470,I6907,,,I7269,);
not I_10(I6890,I7269);
DFFARX1 I_11(I7461,I1470,I6907,,,I6899,);
DFFARX1 I_12(I7365,I1470,I6907,,,I6869,);
endmodule


