module test_I1319(I1223,I1255,I1526,I1294,I1239,I1207,I1301,I1319);
input I1223,I1255,I1526,I1294,I1239,I1207,I1301;
output I1319;
wire I1410,I1560,I1622,I1749,I1543,I1342,I1393,I1639;
nor I_0(I1410,I1223,I1239);
DFFARX1 I_1(I1749,I1294,I1342,,,I1319,);
and I_2(I1560,I1410,I1543);
DFFARX1 I_3(I1255,I1294,I1342,,,I1622,);
or I_4(I1749,I1639,I1560);
nor I_5(I1543,I1393,I1526);
not I_6(I1342,I1301);
DFFARX1 I_7(I1294,I1342,,,I1393,);
and I_8(I1639,I1622,I1207);
endmodule


