module test_final(IN_1_1_l_9,IN_2_1_l_9,IN_3_1_l_9,G18_7_l_9,G15_7_l_9,IN_1_7_l_9,IN_4_7_l_9,IN_5_7_l_9,IN_7_7_l_9,IN_9_7_l_9,IN_10_7_l_9,IN_1_8_l_9,IN_2_8_l_9,IN_3_8_l_9,IN_6_8_l_9,blif_clk_net_8_r_10,blif_reset_net_8_r_10,N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10);
input IN_1_1_l_9,IN_2_1_l_9,IN_3_1_l_9,G18_7_l_9,G15_7_l_9,IN_1_7_l_9,IN_4_7_l_9,IN_5_7_l_9,IN_7_7_l_9,IN_9_7_l_9,IN_10_7_l_9,IN_1_8_l_9,IN_2_8_l_9,IN_3_8_l_9,IN_6_8_l_9,blif_clk_net_8_r_10,blif_reset_net_8_r_10;
output N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10;
wire N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,n_429_or_0_5_r_9,G78_5_r_9,n_576_5_r_9,n_102_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9,I_BUFF_1_9_r_9,n4_7_l_9,n62_9,N3_8_l_9,n63_9,n38_9,n_431_5_r_9,N3_8_r_9,n39_9,n40_9,n41_9,n42_9,n43_9,n44_9,n45_9,n46_9,n47_9,n48_9,n49_9,n50_9,n51_9,n52_9,n53_9,n54_9,n55_9,n56_9,n57_9,n58_9,n59_9,n60_9,n61_9,N1372_4_r_10,I_BUFF_1_9_r_10,N3_8_r_10,n11_10,n35_10,n36_10,n37_10,n38_10,n39_10,n40_10,n41_10,n42_10,n43_10,n44_10,n45_10,n46_10,n47_10,n48_10,n49_10,n50_10,n51_10,n52_10,n53_10,n54_10,n55_10,n56_10,n57_10,n58_10,n59_10,n60_10,n61_10,n62_10,n63_10,n64_10;
nor I_0(N6147_2_r_9,n62_9,n46_9);
not I_1(N1372_4_r_9,n59_9);
nor I_2(N1508_4_r_9,n58_9,n59_9);
nand I_3(n_429_or_0_5_r_9,n_431_5_r_9,n42_9);
DFFARX1 I_4(n_431_5_r_9,blif_clk_net_8_r_10,n11_10,G78_5_r_9,);
nand I_5(n_576_5_r_9,n39_9,n40_9);
not I_6(n_102_5_r_9,I_BUFF_1_9_r_9);
nand I_7(n_547_5_r_9,IN_3_1_l_9,n43_9);
and I_8(n_42_8_r_9,G18_7_l_9,n44_9);
DFFARX1 I_9(N3_8_r_9,blif_clk_net_8_r_10,n11_10,G199_8_r_9,);
nor I_10(N6147_9_r_9,n41_9,n45_9);
nor I_11(N6134_9_r_9,n45_9,n51_9);
nor I_12(I_BUFF_1_9_r_9,IN_3_1_l_9,n41_9);
nor I_13(n4_7_l_9,G18_7_l_9,IN_1_7_l_9);
DFFARX1 I_14(n4_7_l_9,blif_clk_net_8_r_10,n11_10,n62_9,);
and I_15(N3_8_l_9,IN_6_8_l_9,n57_9);
DFFARX1 I_16(N3_8_l_9,blif_clk_net_8_r_10,n11_10,n63_9,);
not I_17(n38_9,n63_9);
nor I_18(n_431_5_r_9,G15_7_l_9,IN_7_7_l_9);
nor I_19(N3_8_r_9,n_102_5_r_9,n53_9);
nor I_20(n39_9,I_BUFF_1_9_r_9,n42_9);
not I_21(n40_9,n41_9);
nand I_22(n41_9,IN_1_1_l_9,IN_2_1_l_9);
nor I_23(n42_9,IN_9_7_l_9,IN_10_7_l_9);
nor I_24(n43_9,n63_9,n41_9);
nor I_25(n44_9,IN_5_7_l_9,IN_9_7_l_9);
and I_26(n45_9,IN_4_7_l_9,n52_9);
nor I_27(n46_9,n47_9,n48_9);
nor I_28(n47_9,n49_9,n50_9);
not I_29(n48_9,n_429_or_0_5_r_9);
not I_30(n49_9,n42_9);
or I_31(n50_9,n63_9,n51_9);
nor I_32(n51_9,IN_1_8_l_9,IN_3_8_l_9);
nor I_33(n52_9,G15_7_l_9,n49_9);
nor I_34(n53_9,n54_9,n55_9);
nor I_35(n54_9,G15_7_l_9,n56_9);
or I_36(n55_9,IN_10_7_l_9,n44_9);
not I_37(n56_9,IN_4_7_l_9);
nand I_38(n57_9,IN_2_8_l_9,IN_3_8_l_9);
nor I_39(n58_9,n62_9,n60_9);
nand I_40(n59_9,n51_9,n61_9);
nor I_41(n60_9,n38_9,n44_9);
nor I_42(n61_9,G18_7_l_9,IN_5_7_l_9);
nor I_43(N1371_0_r_10,n37_10,n38_10);
nor I_44(N1508_0_r_10,n37_10,n58_10);
nand I_45(N6147_2_r_10,n39_10,n40_10);
not I_46(N6147_3_r_10,n39_10);
nor I_47(N1372_4_r_10,n46_10,n49_10);
nor I_48(N1508_4_r_10,n51_10,n52_10);
nor I_49(N1507_6_r_10,n49_10,n60_10);
nor I_50(N1508_6_r_10,n49_10,n50_10);
nor I_51(n_42_8_r_10,I_BUFF_1_9_r_10,n35_10);
DFFARX1 I_52(N3_8_r_10,blif_clk_net_8_r_10,n11_10,G199_8_r_10,);
nor I_53(N6147_9_r_10,n36_10,n37_10);
nor I_54(N6134_9_r_10,I_BUFF_1_9_r_10,n46_10);
not I_55(I_BUFF_1_9_r_10,n48_10);
nor I_56(N3_8_r_10,n44_10,n47_10);
not I_57(n11_10,blif_reset_net_8_r_10);
not I_58(n35_10,n49_10);
nor I_59(n36_10,I_BUFF_1_9_r_10,n38_10);
not I_60(n37_10,N1508_4_r_9);
not I_61(n38_10,n46_10);
nand I_62(n39_10,n43_10,n44_10);
nand I_63(n40_10,I_BUFF_1_9_r_10,n41_10);
nor I_64(n41_10,n42_10,N1508_4_r_9);
not I_65(n42_10,n44_10);
nor I_66(n43_10,n45_10,N1508_4_r_9);
nand I_67(n44_10,n54_10,N1372_4_r_9);
nor I_68(n45_10,n59_10,G199_8_r_9);
nand I_69(n46_10,n61_10,N6147_9_r_9);
nor I_70(n47_10,n46_10,n48_10);
nand I_71(n48_10,n62_10,n63_10);
nand I_72(n49_10,n56_10,G78_5_r_9);
not I_73(n50_10,n45_10);
nor I_74(n51_10,n42_10,n53_10);
not I_75(n52_10,N1372_4_r_10);
nor I_76(n53_10,n48_10,n50_10);
and I_77(n54_10,n55_10,n_576_5_r_9);
nand I_78(n55_10,n56_10,n57_10);
nand I_79(n56_10,N6134_9_r_9,N6147_2_r_9);
not I_80(n57_10,G78_5_r_9);
nor I_81(n58_10,n35_10,n45_10);
nor I_82(n59_10,N1508_4_r_9,n_576_5_r_9);
nor I_83(n60_10,n37_10,n46_10);
or I_84(n61_10,N1508_4_r_9,n_576_5_r_9);
nor I_85(n62_10,n_547_5_r_9,n_42_8_r_9);
or I_86(n63_10,n64_10,N6147_2_r_9);
nor I_87(n64_10,N1372_4_r_9,G78_5_r_9);
endmodule


