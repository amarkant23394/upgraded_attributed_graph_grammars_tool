module test_I12442(I7550,I1477,I1470,I12442);
input I7550,I1477,I1470;
output I12442;
wire I10349,I10038,I12425,I10538,I10490,I11973,I10103,I10332;
and I_0(I10349,I10332,I7550);
nand I_1(I10038,I10349,I10538);
DFFARX1 I_2(I10038,I1470,I11973,,,I12425,);
nor I_3(I10538,I10490,I10103);
DFFARX1 I_4(I1470,,,I10490,);
not I_5(I11973,I1477);
not I_6(I12442,I12425);
DFFARX1 I_7(I1470,,,I10103,);
DFFARX1 I_8(I1470,,,I10332,);
endmodule


