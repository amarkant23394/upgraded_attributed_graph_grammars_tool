module test_final(G1_0_l_11,G2_0_l_11,IN_2_0_l_11,IN_4_0_l_11,IN_5_0_l_11,IN_7_0_l_11,IN_8_0_l_11,IN_10_0_l_11,IN_11_0_l_11,IN_1_5_l_11,IN_2_5_l_11,blif_clk_net_1_r_12,blif_reset_net_1_r_12,G42_1_r_12,n_572_1_r_12,n_573_1_r_12,n_549_1_r_12,n_42_2_r_12,G199_2_r_12,ACVQN1_5_r_12,P6_5_r_12);
input G1_0_l_11,G2_0_l_11,IN_2_0_l_11,IN_4_0_l_11,IN_5_0_l_11,IN_7_0_l_11,IN_8_0_l_11,IN_10_0_l_11,IN_11_0_l_11,IN_1_5_l_11,IN_2_5_l_11,blif_clk_net_1_r_12,blif_reset_net_1_r_12;
output G42_1_r_12,n_572_1_r_12,n_573_1_r_12,n_549_1_r_12,n_42_2_r_12,G199_2_r_12,ACVQN1_5_r_12,P6_5_r_12;
wire G42_1_r_11,n_572_1_r_11,n_573_1_r_11,n_549_1_r_11,n_569_1_r_11,n_452_1_r_11,n_42_2_r_11,G199_2_r_11,ACVQN2_3_r_11,n_266_and_0_3_r_11,n_431_0_l_11,n43_11,n26_11,n44_11,n45_11,n27_11,n4_1_r_11,N3_2_r_11,n24_11,n25_11,n20_internal_11,n20_11,n28_11,n29_11,n30_11,n31_11,n32_11,n33_11,n34_11,n35_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11,n_431_0_l_12,n8_12,n41_12,ACVQN1_5_l_12,n22_12,n42_12,n4_1_r_12,N3_2_r_12,n3_12,P6_5_r_internal_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12;
DFFARX1 I_0(n4_1_r_11,blif_clk_net_1_r_12,n8_12,G42_1_r_11,);
nor I_1(n_572_1_r_11,n29_11,n30_11);
nand I_2(n_573_1_r_11,n26_11,n28_11);
nor I_3(n_549_1_r_11,n27_11,n32_11);
nand I_4(n_569_1_r_11,n45_11,n28_11);
nor I_5(n_452_1_r_11,n43_11,n44_11);
nor I_6(n_42_2_r_11,n35_11,n36_11);
DFFARX1 I_7(N3_2_r_11,blif_clk_net_1_r_12,n8_12,G199_2_r_11,);
DFFARX1 I_8(n24_11,blif_clk_net_1_r_12,n8_12,ACVQN2_3_r_11,);
nor I_9(n_266_and_0_3_r_11,n20_11,n37_11);
or I_10(n_431_0_l_11,IN_8_0_l_11,n33_11);
DFFARX1 I_11(n_431_0_l_11,blif_clk_net_1_r_12,n8_12,n43_11,);
not I_12(n26_11,n43_11);
DFFARX1 I_13(IN_2_5_l_11,blif_clk_net_1_r_12,n8_12,n44_11,);
DFFARX1 I_14(IN_1_5_l_11,blif_clk_net_1_r_12,n8_12,n45_11,);
not I_15(n27_11,n45_11);
nor I_16(n4_1_r_11,n44_11,n25_11);
nor I_17(N3_2_r_11,n45_11,n40_11);
nand I_18(n24_11,IN_11_0_l_11,n39_11);
nand I_19(n25_11,IN_7_0_l_11,n38_11);
DFFARX1 I_20(n25_11,blif_clk_net_1_r_12,n8_12,n20_internal_11,);
not I_21(n20_11,n20_internal_11);
not I_22(n28_11,n25_11);
not I_23(n29_11,G1_0_l_11);
nand I_24(n30_11,n26_11,n31_11);
not I_25(n31_11,IN_5_0_l_11);
and I_26(n32_11,n26_11,n44_11);
and I_27(n33_11,IN_2_0_l_11,n34_11);
nor I_28(n34_11,IN_4_0_l_11,n29_11);
not I_29(n35_11,G2_0_l_11);
nand I_30(n36_11,G1_0_l_11,n31_11);
nor I_31(n37_11,IN_5_0_l_11,n29_11);
nor I_32(n38_11,G2_0_l_11,n31_11);
nor I_33(n39_11,G2_0_l_11,IN_10_0_l_11);
nor I_34(n40_11,G2_0_l_11,n41_11);
nor I_35(n41_11,IN_10_0_l_11,n42_11);
not I_36(n42_11,IN_11_0_l_11);
DFFARX1 I_37(n4_1_r_12,blif_clk_net_1_r_12,n8_12,G42_1_r_12,);
nor I_38(n_572_1_r_12,n29_12,n30_12);
nand I_39(n_573_1_r_12,n26_12,n27_12);
nor I_40(n_549_1_r_12,n33_12,n34_12);
and I_41(n_42_2_r_12,n42_12,n39_12);
DFFARX1 I_42(N3_2_r_12,blif_clk_net_1_r_12,n8_12,G199_2_r_12,);
DFFARX1 I_43(n3_12,blif_clk_net_1_r_12,n8_12,ACVQN1_5_r_12,);
not I_44(P6_5_r_12,P6_5_r_internal_12);
or I_45(n_431_0_l_12,n36_12,ACVQN2_3_r_11);
not I_46(n8_12,blif_reset_net_1_r_12);
DFFARX1 I_47(n_431_0_l_12,blif_clk_net_1_r_12,n8_12,n41_12,);
DFFARX1 I_48(n_452_1_r_11,blif_clk_net_1_r_12,n8_12,ACVQN1_5_l_12,);
not I_49(n22_12,ACVQN1_5_l_12);
DFFARX1 I_50(G42_1_r_11,blif_clk_net_1_r_12,n8_12,n42_12,);
nor I_51(n4_1_r_12,n41_12,n31_12);
nor I_52(N3_2_r_12,n22_12,n40_12);
not I_53(n3_12,n39_12);
DFFARX1 I_54(ACVQN1_5_l_12,blif_clk_net_1_r_12,n8_12,P6_5_r_internal_12,);
and I_55(n26_12,n_573_1_r_11,G199_2_r_11);
nor I_56(n27_12,n28_12,n29_12);
not I_57(n28_12,G42_1_r_11);
nand I_58(n29_12,n31_12,n32_12);
nand I_59(n30_12,n42_12,G42_1_r_11);
not I_60(n31_12,n_569_1_r_11);
not I_61(n32_12,n_549_1_r_11);
nand I_62(n33_12,n31_12,n35_12);
nand I_63(n34_12,n_573_1_r_11,G199_2_r_11);
nand I_64(n35_12,n41_12,n42_12);
and I_65(n36_12,n37_12,n_266_and_0_3_r_11);
nor I_66(n37_12,n38_12,n_572_1_r_11);
not I_67(n38_12,n_42_2_r_11);
nor I_68(n39_12,n38_12,G199_2_r_11);
nor I_69(n40_12,n39_12,n_569_1_r_11);
endmodule


