module test_I2759(I1477,I2759);
input I1477;
output I2759;
wire ;
not I_0(I2759,I1477);
endmodule


