module test_final(IN_1_2_l_13,IN_2_2_l_13,G1_3_l_13,G2_3_l_13,IN_2_3_l_13,IN_4_3_l_13,IN_5_3_l_13,IN_7_3_l_13,IN_8_3_l_13,IN_10_3_l_13,IN_11_3_l_13,blif_clk_net_3_r_0,blif_reset_net_3_r_0,n_429_or_0_3_r_0,G78_3_r_0,n_576_3_r_0,n_102_3_r_0,n_547_3_r_0,G42_4_r_0,n_572_4_r_0,n_573_4_r_0,n_549_4_r_0,n_569_4_r_0,n_452_4_r_0);
input IN_1_2_l_13,IN_2_2_l_13,G1_3_l_13,G2_3_l_13,IN_2_3_l_13,IN_4_3_l_13,IN_5_3_l_13,IN_7_3_l_13,IN_8_3_l_13,IN_10_3_l_13,IN_11_3_l_13,blif_clk_net_3_r_0,blif_reset_net_3_r_0;
output n_429_or_0_3_r_0,G78_3_r_0,n_576_3_r_0,n_102_3_r_0,n_547_3_r_0,G42_4_r_0,n_572_4_r_0,n_573_4_r_0,n_549_4_r_0,n_569_4_r_0,n_452_4_r_0;
wire n_429_or_0_3_r_13,G78_3_r_13,n_576_3_r_13,n_102_3_r_13,n_547_3_r_13,G42_4_r_13,n_572_4_r_13,n_573_4_r_13,n_549_4_r_13,n_569_4_r_13,n_452_4_r_13,ACVQN1_2_l_13,P6_2_l_13,P6_internal_2_l_13,n_429_or_0_3_l_13,n12_3_l_13,n_431_3_l_13,G78_3_l_13,n_576_3_l_13,n11_3_l_13,n_102_3_l_13,n_547_3_l_13,n13_3_l_13,n14_3_l_13,n15_3_l_13,n16_3_l_13,n12_3_r_13,n_431_3_r_13,n11_3_r_13,n13_3_r_13,n14_3_r_13,n15_3_r_13,n16_3_r_13,n4_4_r_13,n_87_4_r_13,n7_4_r_13,n2_3_r_0,ACVQN2_0_l_0,n_266_and_0_0_l_0,ACVQN1_0_l_0,N1_1_l_0,G199_1_l_0,G214_1_l_0,n3_1_l_0,n_42_5_l_0,N3_5_l_0,G199_5_l_0,n3_5_l_0,n12_3_r_0,n_431_3_r_0,n11_3_r_0,n13_3_r_0,n14_3_r_0,n15_3_r_0,n16_3_r_0,n4_4_r_0,n_87_4_r_0,n7_4_r_0;
nand I_0(n_429_or_0_3_r_13,n_429_or_0_3_l_13,n12_3_r_13);
DFFARX1 I_1(n_431_3_r_13,blif_clk_net_3_r_0,n2_3_r_0,G78_3_r_13,);
nand I_2(n_576_3_r_13,n_547_3_l_13,n11_3_r_13);
not I_3(n_102_3_r_13,ACVQN1_2_l_13);
nand I_4(n_547_3_r_13,P6_2_l_13,n13_3_r_13);
DFFARX1 I_5(n4_4_r_13,blif_clk_net_3_r_0,n2_3_r_0,G42_4_r_13,);
nor I_6(n_572_4_r_13,P6_2_l_13,n_429_or_0_3_l_13);
or I_7(n_573_4_r_13,ACVQN1_2_l_13,G78_3_l_13);
nor I_8(n_549_4_r_13,n_429_or_0_3_l_13,n7_4_r_13);
or I_9(n_569_4_r_13,n_429_or_0_3_l_13,G78_3_l_13);
nor I_10(n_452_4_r_13,ACVQN1_2_l_13,P6_2_l_13);
DFFARX1 I_11(IN_2_2_l_13,blif_clk_net_3_r_0,n2_3_r_0,ACVQN1_2_l_13,);
not I_12(P6_2_l_13,P6_internal_2_l_13);
DFFARX1 I_13(IN_1_2_l_13,blif_clk_net_3_r_0,n2_3_r_0,P6_internal_2_l_13,);
nand I_14(n_429_or_0_3_l_13,G1_3_l_13,n12_3_l_13);
not I_15(n12_3_l_13,IN_5_3_l_13);
or I_16(n_431_3_l_13,IN_8_3_l_13,n14_3_l_13);
DFFARX1 I_17(n_431_3_l_13,blif_clk_net_3_r_0,n2_3_r_0,G78_3_l_13,);
nand I_18(n_576_3_l_13,IN_7_3_l_13,n11_3_l_13);
nor I_19(n11_3_l_13,G2_3_l_13,n12_3_l_13);
not I_20(n_102_3_l_13,G2_3_l_13);
nand I_21(n_547_3_l_13,IN_11_3_l_13,n13_3_l_13);
nor I_22(n13_3_l_13,G2_3_l_13,IN_10_3_l_13);
and I_23(n14_3_l_13,IN_2_3_l_13,n15_3_l_13);
nor I_24(n15_3_l_13,IN_4_3_l_13,n16_3_l_13);
not I_25(n16_3_l_13,G1_3_l_13);
not I_26(n12_3_r_13,n_102_3_l_13);
or I_27(n_431_3_r_13,ACVQN1_2_l_13,n14_3_r_13);
nor I_28(n11_3_r_13,ACVQN1_2_l_13,n12_3_r_13);
nor I_29(n13_3_r_13,ACVQN1_2_l_13,n_576_3_l_13);
and I_30(n14_3_r_13,n_102_3_l_13,n15_3_r_13);
nor I_31(n15_3_r_13,G78_3_l_13,n16_3_r_13);
not I_32(n16_3_r_13,n_429_or_0_3_l_13);
nor I_33(n4_4_r_13,P6_2_l_13,n_547_3_l_13);
not I_34(n_87_4_r_13,P6_2_l_13);
and I_35(n7_4_r_13,n_576_3_l_13,n_87_4_r_13);
nand I_36(n_429_or_0_3_r_0,ACVQN2_0_l_0,n12_3_r_0);
DFFARX1 I_37(n_431_3_r_0,blif_clk_net_3_r_0,n2_3_r_0,G78_3_r_0,);
nand I_38(n_576_3_r_0,n_266_and_0_0_l_0,n11_3_r_0);
not I_39(n_102_3_r_0,n_42_5_l_0);
nand I_40(n_547_3_r_0,ACVQN2_0_l_0,n13_3_r_0);
DFFARX1 I_41(n4_4_r_0,blif_clk_net_3_r_0,n2_3_r_0,G42_4_r_0,);
nor I_42(n_572_4_r_0,G199_1_l_0,G199_5_l_0);
or I_43(n_573_4_r_0,n_42_5_l_0,G199_5_l_0);
nor I_44(n_549_4_r_0,n_266_and_0_0_l_0,n7_4_r_0);
or I_45(n_569_4_r_0,n_266_and_0_0_l_0,n_42_5_l_0);
nor I_46(n_452_4_r_0,ACVQN2_0_l_0,G199_5_l_0);
not I_47(n2_3_r_0,blif_reset_net_3_r_0);
DFFARX1 I_48(n_576_3_r_13,blif_clk_net_3_r_0,n2_3_r_0,ACVQN2_0_l_0,);
and I_49(n_266_and_0_0_l_0,ACVQN1_0_l_0,n_547_3_r_13);
DFFARX1 I_50(n_549_4_r_13,blif_clk_net_3_r_0,n2_3_r_0,ACVQN1_0_l_0,);
and I_51(N1_1_l_0,n3_1_l_0,n_569_4_r_13);
DFFARX1 I_52(N1_1_l_0,blif_clk_net_3_r_0,n2_3_r_0,G199_1_l_0,);
DFFARX1 I_53(n_452_4_r_13,blif_clk_net_3_r_0,n2_3_r_0,G214_1_l_0,);
nand I_54(n3_1_l_0,G42_4_r_13,n_572_4_r_13);
nor I_55(n_42_5_l_0,G78_3_r_13,n_573_4_r_13);
and I_56(N3_5_l_0,n3_5_l_0,n_102_3_r_13);
DFFARX1 I_57(N3_5_l_0,blif_clk_net_3_r_0,n2_3_r_0,G199_5_l_0,);
nand I_58(n3_5_l_0,n_429_or_0_3_r_13,G78_3_r_13);
not I_59(n12_3_r_0,G199_1_l_0);
or I_60(n_431_3_r_0,n_266_and_0_0_l_0,n14_3_r_0);
nor I_61(n11_3_r_0,G214_1_l_0,n12_3_r_0);
nor I_62(n13_3_r_0,G214_1_l_0,n_42_5_l_0);
and I_63(n14_3_r_0,n_42_5_l_0,n15_3_r_0);
nor I_64(n15_3_r_0,G199_1_l_0,n16_3_r_0);
not I_65(n16_3_r_0,ACVQN2_0_l_0);
nor I_66(n4_4_r_0,ACVQN2_0_l_0,G214_1_l_0);
not I_67(n_87_4_r_0,G199_5_l_0);
and I_68(n7_4_r_0,ACVQN2_0_l_0,n_87_4_r_0);
endmodule


