module test_I5751_rst(I1477_rst,I5751_rst);
,I5751_rst);
input I1477_rst;
output I5751_rst;
wire ;
not I_0(I5751_rst,I1477_rst);
endmodule


