module test_I3975(I2878,I1477,I1470,I2793,I1335,I3975);
input I2878,I1477,I1470,I2793,I1335;
output I3975;
wire I2730,I2721,I2810,I4017,I3124,I2727,I4000,I3076,I4308,I4034,I2724,I3983;
not I_0(I2730,I3076);
nand I_1(I2721,I2878);
nor I_2(I3975,I4308,I4034);
nand I_3(I2810,I2793,I1335);
and I_4(I4017,I4000,I2730);
nor I_5(I3124,I3076,I2878);
nand I_6(I2727,I2810,I3124);
nand I_7(I4000,I2721,I2724);
DFFARX1 I_8(I1470,,,I3076,);
DFFARX1 I_9(I2727,I1470,I3983,,,I4308,);
DFFARX1 I_10(I4017,I1470,I3983,,,I4034,);
DFFARX1 I_11(I1470,,,I2724,);
not I_12(I3983,I1477);
endmodule


