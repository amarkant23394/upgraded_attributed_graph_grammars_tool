module Benchmark_testing10000(I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1804,I1812,I1820,I1828,I1836,I1844,I1852,I1860,I1868,I1876,I1884,I1892,I1900,I1908,I1916,I1924,I1932,I1940,I1948,I1956,I1964,I1972,I1980,I1988,I1996,I2004,I2012,I2020,I2028,I2036,I2044,I2052,I2060,I2067,I2074,I3291,I3282,I3279,I3285,I3273,I3267,I3288,I3276,I3270,I74895,I74892,I74877,I74889,I74883,I74871,I74880,I74886,I74874,I90577,I90580,I90562,I90571,I90583,I90574,I90565,I90568,I90586,I128799,I128802,I128778,I128790,I128805,I128793,I128787,I128781,I128784,I128796,I135701,I135683,I135686,I135695,I135698,I135692,I135680,I135689,I140863,I140851,I140872,I140848,I140869,I140860,I140866,I140857,I140854,I146065,I146053,I146074,I146050,I146071,I146062,I146068,I146059,I146056,I164094,I164073,I164079,I164088,I164091,I164070,I164085,I164082,I164076);
input I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1804,I1812,I1820,I1828,I1836,I1844,I1852,I1860,I1868,I1876,I1884,I1892,I1900,I1908,I1916,I1924,I1932,I1940,I1948,I1956,I1964,I1972,I1980,I1988,I1996,I2004,I2012,I2020,I2028,I2036,I2044,I2052,I2060,I2067,I2074;
output I3291,I3282,I3279,I3285,I3273,I3267,I3288,I3276,I3270,I74895,I74892,I74877,I74889,I74883,I74871,I74880,I74886,I74874,I90577,I90580,I90562,I90571,I90583,I90574,I90565,I90568,I90586,I128799,I128802,I128778,I128790,I128805,I128793,I128787,I128781,I128784,I128796,I135701,I135683,I135686,I135695,I135698,I135692,I135680,I135689,I140863,I140851,I140872,I140848,I140869,I140860,I140866,I140857,I140854,I146065,I146053,I146074,I146050,I146071,I146062,I146068,I146059,I146056,I164094,I164073,I164079,I164088,I164091,I164070,I164085,I164082,I164076;
wire I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1804,I1812,I1820,I1828,I1836,I1844,I1852,I1860,I1868,I1876,I1884,I1892,I1900,I1908,I1916,I1924,I1932,I1940,I1948,I1956,I1964,I1972,I1980,I1988,I1996,I2004,I2012,I2020,I2028,I2036,I2044,I2052,I2060,I2067,I2074,I2106,I33411,I2132,I2140,I2157,I2098,I33417,I2197,I2205,I2222,I33426,I2239,I33420,I2256,I2273,I2077,I2304,I2321,I2338,I33423,I33429,I2080,I2369,I2386,I33432,I2403,I33408,I2420,I2437,I2454,I2089,I2485,I33414,I2502,I2519,I2095,I2550,I2092,I2581,I2607,I2615,I2632,I2086,I2083,I2701,I14346,I2727,I2735,I14337,I2752,I2693,I14358,I2792,I2800,I2817,I14334,I2834,I2851,I2868,I2672,I2899,I2916,I2933,I14343,I2675,I2964,I2981,I14355,I2998,I14352,I3015,I3032,I3049,I2684,I3080,I14349,I3097,I3114,I2690,I3145,I2687,I3176,I14340,I3202,I3210,I3227,I2681,I2678,I3299,I161195,I3325,I3342,I3350,I3367,I161198,I161192,I3384,I161201,I3410,I161189,I3455,I3463,I161204,I3480,I161180,I3520,I3528,I3573,I161183,I3590,I3616,I3624,I3655,I3672,I161186,I3689,I3706,I3723,I3754,I3826,I32819,I3852,I3869,I3877,I3894,I32837,I32822,I3911,I32825,I3937,I3818,I3809,I32813,I3982,I3990,I32816,I4007,I3806,I32828,I4047,I4055,I3812,I3800,I4100,I32834,I32831,I4117,I4143,I4151,I3794,I4182,I4199,I4216,I4233,I4250,I3815,I4281,I3803,I3797,I4353,I61305,I4379,I4396,I4404,I4421,I61308,I4438,I61329,I4464,I4345,I4336,I61317,I4509,I4517,I61320,I4534,I4333,I61326,I4574,I4582,I4339,I4327,I4627,I61323,I61311,I4644,I61314,I4670,I4678,I4321,I4709,I4726,I61332,I4743,I4760,I4777,I4342,I4808,I4330,I4324,I4880,I92302,I4906,I4923,I4931,I4948,I92317,I92320,I4965,I92299,I4991,I4872,I4863,I92305,I5036,I5044,I92311,I5061,I4860,I5101,I5109,I4866,I4854,I5154,I92314,I92296,I5171,I92308,I5197,I5205,I4848,I5236,I5253,I5270,I5287,I5304,I4869,I5335,I4857,I4851,I5407,I57575,I5433,I5450,I5458,I5475,I57572,I57566,I5492,I57560,I5518,I5399,I5390,I57548,I5563,I5571,I57557,I5588,I5387,I57554,I5628,I5636,I5393,I5381,I5681,I57551,I57569,I5698,I5724,I5732,I5375,I5763,I5780,I57563,I5797,I5814,I5831,I5396,I5862,I5384,I5378,I5934,I50197,I5960,I5977,I5985,I6002,I50194,I50188,I6019,I50182,I6045,I5926,I5917,I50170,I6090,I6098,I50179,I6115,I5914,I50176,I6155,I6163,I5920,I5908,I6208,I50173,I50191,I6225,I6251,I6259,I5902,I6290,I6307,I50185,I6324,I6341,I6358,I5923,I6389,I5911,I5905,I6461,I106024,I6487,I6504,I6512,I6529,I106015,I106036,I6546,I106018,I6572,I6453,I6444,I6617,I6625,I106033,I6642,I6441,I106027,I6682,I6690,I6447,I6435,I6735,I106021,I106030,I6752,I6778,I6786,I6429,I6817,I6834,I6851,I6868,I6885,I6450,I6916,I6438,I6432,I6988,I50724,I7014,I7031,I7039,I7056,I50721,I50715,I7073,I50709,I7099,I6980,I6971,I50697,I7144,I7152,I50706,I7169,I6968,I50703,I7209,I7217,I6974,I6962,I7262,I50700,I50718,I7279,I7305,I7313,I6956,I7344,I7361,I50712,I7378,I7395,I7412,I6977,I7443,I6965,I6959,I7515,I70715,I7541,I7558,I7566,I7583,I70721,I70709,I7600,I70706,I7626,I7507,I7498,I70718,I7671,I7679,I70712,I7696,I7495,I70730,I7736,I7744,I7501,I7489,I7789,I70724,I70727,I7806,I7832,I7840,I7483,I7871,I7888,I7905,I7922,I7939,I7504,I7970,I7492,I7486,I8042,I87678,I8068,I8085,I8093,I8110,I87693,I87696,I8127,I87675,I8153,I8034,I8025,I87681,I8198,I8206,I87687,I8223,I8022,I8263,I8271,I8028,I8016,I8316,I87690,I87672,I8333,I87684,I8359,I8367,I8010,I8398,I8415,I8432,I8449,I8466,I8031,I8497,I8019,I8013,I8569,I100394,I8595,I8612,I8620,I8637,I100409,I100412,I8654,I100391,I8680,I8561,I8552,I100397,I8725,I8733,I100403,I8750,I8549,I8790,I8798,I8555,I8543,I8843,I100406,I100388,I8860,I100400,I8886,I8894,I8537,I8925,I8942,I8959,I8976,I8993,I8558,I9024,I8546,I8540,I9096,I160617,I9122,I9139,I9147,I9164,I160620,I160614,I9181,I160623,I9207,I9088,I9079,I160611,I9252,I9260,I160626,I9277,I9076,I160602,I9317,I9325,I9082,I9070,I9370,I160605,I9387,I9413,I9421,I9064,I9452,I9469,I160608,I9486,I9503,I9520,I9085,I9551,I9073,I9067,I9623,I53359,I9649,I9657,I9674,I53341,I53356,I9691,I53332,I9717,I53335,I9734,I9742,I53350,I9759,I9591,I9790,I9807,I9603,I53353,I9847,I9612,I9869,I53344,I9886,I53338,I9912,I9929,I9615,I9951,I9600,I9982,I53347,I9999,I10016,I10033,I9609,I10064,I9597,I9606,I9594,I10150,I98088,I10176,I10184,I10201,I98079,I98097,I10218,I98076,I10244,I10261,I10269,I98082,I10286,I10118,I10317,I10334,I10130,I10374,I10139,I10396,I98094,I98085,I10413,I98100,I10439,I10456,I10142,I10478,I10127,I10509,I98091,I10526,I10543,I10560,I10136,I10591,I10124,I10133,I10121,I10677,I85369,I10703,I10711,I10728,I85381,I85366,I10745,I85360,I10771,I85375,I10788,I10796,I85363,I10813,I10645,I10844,I10861,I10657,I85372,I10901,I10666,I10923,I85378,I85384,I10940,I10966,I10983,I10669,I11005,I10654,I11036,I11053,I11070,I11087,I10663,I11118,I10651,I10660,I10648,I11204,I11230,I11238,I11255,I11272,I11298,I11315,I11323,I11340,I11172,I11371,I11388,I11184,I11428,I11193,I11450,I11467,I11493,I11510,I11196,I11532,I11181,I11563,I11580,I11597,I11614,I11190,I11645,I11178,I11187,I11175,I11731,I112875,I11757,I11765,I11782,I112872,I112887,I11799,I112869,I11825,I112866,I11842,I11850,I11867,I11699,I11898,I11915,I11711,I11955,I11720,I11977,I112881,I11994,I112884,I12020,I12037,I11723,I12059,I11708,I12090,I112878,I12107,I12124,I12141,I11717,I12172,I11705,I11714,I11702,I12258,I168111,I12284,I12292,I12309,I168105,I168126,I12326,I168102,I12352,I168123,I12369,I12377,I168120,I12394,I12226,I12425,I12442,I12238,I168108,I12482,I12247,I12504,I168117,I168114,I12521,I168099,I12547,I12564,I12250,I12586,I12235,I12617,I12634,I12651,I12668,I12244,I12699,I12232,I12241,I12229,I12785,I67307,I12811,I12819,I12836,I67301,I67292,I12853,I67313,I12879,I67295,I12896,I12904,I67289,I12921,I12753,I12952,I12969,I12765,I13009,I12774,I13031,I67316,I67298,I13048,I67304,I13074,I13091,I12777,I13113,I12762,I13144,I67310,I13161,I13178,I13195,I12771,I13226,I12759,I12768,I12756,I13312,I69519,I13338,I13346,I13363,I69540,I69534,I13380,I69516,I13406,I13423,I13431,I69528,I13448,I13280,I13479,I13496,I13292,I69525,I13536,I13301,I13558,I69531,I69522,I13575,I13601,I13618,I13304,I13640,I13289,I13671,I69537,I13688,I13705,I13722,I13298,I13753,I13286,I13295,I13283,I13839,I162357,I13865,I13873,I13890,I162360,I162354,I13907,I162351,I13933,I162336,I13950,I13958,I162345,I13975,I13807,I14006,I14023,I13819,I14063,I13828,I14085,I162339,I162342,I14102,I162348,I14128,I14145,I13831,I14167,I13816,I14198,I14215,I14232,I14249,I13825,I14280,I13813,I13822,I13810,I14366,I14392,I14400,I14417,I14434,I14460,I14477,I14485,I14502,I14533,I14550,I14590,I14612,I14629,I14655,I14672,I14694,I14725,I14742,I14759,I14776,I14807,I14893,I83635,I14919,I14927,I14944,I83647,I83632,I14961,I83626,I14987,I83641,I15004,I15012,I83629,I15029,I14861,I15060,I15077,I14873,I83638,I15117,I14882,I15139,I83644,I83650,I15156,I15182,I15199,I14885,I15221,I14870,I15252,I15269,I15286,I15303,I14879,I15334,I14867,I14876,I14864,I15420,I15446,I15454,I15471,I15488,I15514,I15531,I15539,I15556,I15388,I15587,I15604,I15400,I15644,I15409,I15666,I15683,I15709,I15726,I15412,I15748,I15397,I15779,I15796,I15813,I15830,I15406,I15861,I15394,I15403,I15391,I15947,I79589,I15973,I15981,I15998,I79601,I79586,I16015,I79580,I16041,I79595,I16058,I16066,I79583,I16083,I15915,I16114,I16131,I15927,I79592,I16171,I15936,I16193,I79598,I79604,I16210,I16236,I16253,I15939,I16275,I15924,I16306,I16323,I16340,I16357,I15933,I16388,I15921,I15930,I15918,I16474,I136244,I16500,I16508,I16525,I136241,I136247,I16542,I16568,I16585,I16593,I16610,I16442,I16641,I16658,I16454,I136250,I16698,I16463,I16720,I136253,I136262,I16737,I136256,I16763,I16780,I16466,I16802,I16451,I16833,I136259,I16850,I16867,I16884,I16460,I16915,I16448,I16457,I16445,I17001,I53886,I17027,I17035,I17052,I53868,I53883,I17069,I53859,I17095,I53862,I17112,I17120,I53877,I17137,I16969,I17168,I17185,I16981,I53880,I17225,I16990,I17247,I53871,I17264,I53865,I17290,I17307,I16993,I17329,I16978,I17360,I53874,I17377,I17394,I17411,I16987,I17442,I16975,I16984,I16972,I17528,I151836,I17554,I17562,I17579,I151851,I151830,I17596,I151833,I17622,I151854,I17639,I17647,I17664,I17496,I17695,I17712,I17508,I17752,I17517,I17774,I151842,I151839,I17791,I151845,I17817,I17834,I17520,I17856,I17505,I17887,I151848,I17904,I17921,I17938,I17514,I17969,I17502,I17511,I17499,I18055,I74279,I18081,I18089,I18106,I74300,I74294,I18123,I74276,I18149,I18166,I18174,I74288,I18191,I18023,I18222,I18239,I18035,I74285,I18279,I18044,I18301,I74291,I74282,I18318,I18344,I18361,I18047,I18383,I18032,I18414,I74297,I18431,I18448,I18465,I18041,I18496,I18029,I18038,I18026,I18582,I18608,I18616,I18633,I18650,I18676,I18693,I18701,I18718,I18550,I18749,I18766,I18562,I18806,I18571,I18828,I18845,I18871,I18888,I18574,I18910,I18559,I18941,I18958,I18975,I18992,I18568,I19023,I18556,I18565,I18553,I19109,I26875,I19135,I19143,I19160,I26869,I26863,I19177,I26884,I19203,I26881,I19220,I19228,I26878,I19245,I19077,I19276,I19293,I19089,I19333,I19098,I19355,I26866,I19372,I26887,I19398,I19415,I19101,I19437,I19086,I19468,I26872,I19485,I19502,I19519,I19095,I19550,I19083,I19092,I19080,I19636,I84791,I19662,I19670,I19687,I84803,I84788,I19704,I84782,I19730,I84797,I19747,I19755,I84785,I19772,I19604,I19803,I19820,I19616,I84794,I19860,I19625,I19882,I84800,I84806,I19899,I19925,I19942,I19628,I19964,I19613,I19995,I20012,I20029,I20046,I19622,I20077,I19610,I19619,I19607,I20163,I34610,I20189,I20197,I20214,I34604,I34598,I20231,I34619,I20257,I34616,I20274,I20282,I34613,I20299,I20131,I20330,I20347,I20143,I20387,I20152,I20409,I34601,I20426,I34622,I20452,I20469,I20155,I20491,I20140,I20522,I34607,I20539,I20556,I20573,I20149,I20604,I20137,I20146,I20134,I20690,I75469,I20716,I20724,I20741,I75490,I75484,I20758,I75466,I20784,I20801,I20809,I75478,I20826,I20658,I20857,I20874,I20670,I75475,I20914,I20679,I20936,I75481,I75472,I20953,I20979,I20996,I20682,I21018,I20667,I21049,I75487,I21066,I21083,I21100,I20676,I21131,I20664,I20673,I20661,I21217,I25090,I21243,I21251,I21268,I25084,I25078,I21285,I25099,I21311,I25096,I21328,I21336,I25093,I21353,I21185,I21384,I21401,I21197,I21441,I21206,I21463,I25081,I21480,I25102,I21506,I21523,I21209,I21545,I21194,I21576,I25087,I21593,I21610,I21627,I21203,I21658,I21191,I21200,I21188,I21744,I178821,I21770,I21778,I21795,I178815,I178836,I21812,I178812,I21838,I178833,I21855,I21863,I178830,I21880,I21712,I21911,I21928,I21724,I178818,I21968,I21733,I21990,I178827,I178824,I22007,I178809,I22033,I22050,I21736,I22072,I21721,I22103,I22120,I22137,I22154,I21730,I22185,I21718,I21727,I21715,I22271,I102712,I22297,I22305,I22322,I102703,I102721,I22339,I102700,I22365,I22382,I22390,I102706,I22407,I22239,I22438,I22455,I22251,I22495,I22260,I22517,I102718,I102709,I22534,I102724,I22560,I22577,I22263,I22599,I22248,I22630,I102715,I22647,I22664,I22681,I22257,I22712,I22245,I22254,I22242,I22798,I43873,I22824,I22832,I22849,I43855,I43870,I22866,I43846,I22892,I43849,I22909,I22917,I43864,I22934,I22766,I22965,I22982,I22778,I43867,I23022,I22787,I23044,I43858,I23061,I43852,I23087,I23104,I22790,I23126,I22775,I23157,I43861,I23174,I23191,I23208,I22784,I23239,I22772,I22781,I22769,I23328,I23354,I23362,I23388,I23396,I23413,I23430,I23305,I23461,I23299,I23492,I23509,I23526,I23543,I23560,I23577,I23314,I23311,I23317,I23636,I23653,I23670,I23696,I23296,I23727,I23735,I23320,I23766,I23783,I23800,I23302,I23831,I23848,I23293,I23308,I23920,I89418,I23946,I23963,I23912,I23985,I89415,I24011,I24019,I24036,I89421,I24053,I89406,I24070,I24087,I89409,I24104,I89430,I24121,I89427,I24138,I23888,I24169,I24186,I24203,I24220,I23900,I23894,I24265,I23909,I23903,I24310,I24327,I89412,I24344,I89424,I24361,I24387,I24395,I23897,I23891,I24449,I24457,I23906,I24515,I52278,I24541,I24558,I24507,I24580,I52293,I24606,I24614,I24631,I52290,I24648,I24665,I24682,I52287,I24699,I52302,I24716,I52299,I24733,I24483,I24764,I24781,I24798,I24815,I24495,I24489,I24860,I52296,I24504,I24498,I24905,I24922,I52284,I24939,I52305,I24956,I52281,I24982,I24990,I24492,I24486,I25044,I25052,I24501,I25110,I124271,I25136,I25153,I25175,I124280,I25201,I25209,I25226,I124268,I25243,I124259,I25260,I25277,I124265,I25294,I124283,I25311,I124256,I25328,I25359,I25376,I25393,I25410,I25455,I124262,I25500,I25517,I124274,I25534,I25551,I124277,I25577,I25585,I25639,I25647,I25705,I44373,I25731,I25748,I25697,I25770,I44388,I25796,I25804,I25821,I44385,I25838,I25855,I25872,I44382,I25889,I44397,I25906,I44394,I25923,I25673,I25954,I25971,I25988,I26005,I25685,I25679,I26050,I44391,I25694,I25688,I26095,I26112,I44379,I26129,I44400,I26146,I44376,I26172,I26180,I25682,I25676,I26234,I26242,I25691,I26300,I67857,I26326,I26343,I26292,I26365,I67845,I26391,I26399,I26416,I67854,I26433,I67851,I26450,I26467,I67842,I26484,I67848,I26501,I67833,I26518,I26268,I26549,I26566,I26583,I26600,I26280,I26274,I26645,I26289,I26283,I26690,I26707,I67839,I26724,I67836,I26741,I67860,I26767,I26775,I26277,I26271,I26829,I26837,I26286,I26895,I163495,I26921,I26938,I26960,I163507,I26986,I26994,I27011,I163501,I27028,I163513,I27045,I27062,I163498,I27079,I163510,I27096,I163492,I27113,I27144,I27161,I27178,I27195,I27240,I163504,I27285,I27302,I27319,I27336,I163516,I27362,I27370,I27424,I27432,I27490,I104967,I27516,I27533,I27482,I27555,I104961,I27581,I27589,I27606,I104979,I27623,I27640,I27657,I27674,I104973,I27691,I104964,I27708,I27458,I27739,I27756,I27773,I27790,I27470,I27464,I27835,I104976,I27479,I27473,I27880,I27897,I104982,I27914,I27931,I104970,I27957,I27965,I27467,I27461,I28019,I28027,I27476,I28085,I49116,I28111,I28128,I28077,I28150,I49131,I28176,I28184,I28201,I49128,I28218,I28235,I28252,I49125,I28269,I49140,I28286,I49137,I28303,I28053,I28334,I28351,I28368,I28385,I28065,I28059,I28430,I49134,I28074,I28068,I28475,I28492,I49122,I28509,I49143,I28526,I49119,I28552,I28560,I28062,I28056,I28614,I28622,I28071,I28680,I28706,I28723,I28672,I28745,I28771,I28779,I28796,I28813,I28830,I28847,I28864,I28881,I28898,I28648,I28929,I28946,I28963,I28980,I28660,I28654,I29025,I28669,I28663,I29070,I29087,I29104,I29121,I29147,I29155,I28657,I28651,I29209,I29217,I28666,I29275,I29301,I29318,I29267,I29340,I29366,I29374,I29391,I29408,I29425,I29442,I29459,I29476,I29493,I29243,I29524,I29541,I29558,I29575,I29255,I29249,I29620,I29264,I29258,I29665,I29682,I29699,I29716,I29742,I29750,I29252,I29246,I29804,I29812,I29261,I29870,I89996,I29896,I29913,I29862,I29935,I89993,I29961,I29969,I29986,I89999,I30003,I89984,I30020,I30037,I89987,I30054,I90008,I30071,I90005,I30088,I29838,I30119,I30136,I30153,I30170,I29850,I29844,I30215,I29859,I29853,I30260,I30277,I89990,I30294,I90002,I30311,I30337,I30345,I29847,I29841,I30399,I30407,I29856,I30465,I174665,I30491,I30508,I30457,I30530,I174656,I30556,I30564,I30581,I174650,I30598,I174644,I30615,I30632,I174671,I30649,I30666,I174668,I30683,I30433,I30714,I30731,I30748,I30765,I30445,I30439,I30810,I174653,I30454,I30448,I30855,I30872,I174659,I30889,I174662,I30906,I174647,I30932,I30940,I30442,I30436,I30994,I31002,I30451,I31060,I68401,I31086,I31103,I31052,I31125,I68389,I31151,I31159,I31176,I68398,I31193,I68395,I31210,I31227,I68386,I31244,I68392,I31261,I68377,I31278,I31028,I31309,I31326,I31343,I31360,I31040,I31034,I31405,I31049,I31043,I31450,I31467,I68383,I31484,I68380,I31501,I68404,I31527,I31535,I31037,I31031,I31589,I31597,I31046,I31655,I31681,I31698,I31647,I31720,I31746,I31754,I31771,I31788,I31805,I31822,I31839,I31856,I31873,I31623,I31904,I31921,I31938,I31955,I31635,I31629,I32000,I31644,I31638,I32045,I32062,I32079,I32096,I32122,I32130,I31632,I31626,I32184,I32192,I31641,I32250,I91730,I32276,I32293,I32242,I32315,I91727,I32341,I32349,I32366,I91733,I32383,I91718,I32400,I32417,I91721,I32434,I91742,I32451,I91739,I32468,I32218,I32499,I32516,I32533,I32550,I32230,I32224,I32595,I32239,I32233,I32640,I32657,I91724,I32674,I91736,I32691,I32717,I32725,I32227,I32221,I32779,I32787,I32236,I32845,I32871,I32888,I32910,I32936,I32944,I32961,I32978,I32995,I33012,I33029,I33046,I33063,I33094,I33111,I33128,I33145,I33190,I33235,I33252,I33269,I33286,I33312,I33320,I33374,I33382,I33440,I104440,I33466,I33483,I33505,I104434,I33531,I33539,I33556,I104452,I33573,I33590,I33607,I33624,I104446,I33641,I104437,I33658,I33689,I33706,I33723,I33740,I33785,I104449,I33830,I33847,I104455,I33864,I33881,I104443,I33907,I33915,I33969,I33977,I34035,I132317,I34061,I34078,I34027,I34100,I132326,I34126,I34134,I34151,I132320,I34168,I132314,I34185,I34202,I132329,I34219,I34236,I132323,I34253,I34003,I34284,I34301,I34318,I34335,I34015,I34009,I34380,I34024,I34018,I34425,I34442,I132335,I34459,I132332,I34476,I34502,I34510,I34012,I34006,I34564,I34572,I34021,I34630,I103290,I34656,I34673,I34695,I103287,I34721,I34729,I34746,I103293,I34763,I103278,I34780,I34797,I103281,I34814,I103302,I34831,I103299,I34848,I34879,I34896,I34913,I34930,I34975,I35020,I35037,I103284,I35054,I103296,I35071,I35097,I35105,I35159,I35167,I35225,I101556,I35251,I35268,I35217,I35290,I101553,I35316,I35324,I35341,I101559,I35358,I101544,I35375,I35392,I101547,I35409,I101568,I35426,I101565,I35443,I35193,I35474,I35491,I35508,I35525,I35205,I35199,I35570,I35214,I35208,I35615,I35632,I101550,I35649,I101562,I35666,I35692,I35700,I35202,I35196,I35754,I35762,I35211,I35820,I125563,I35846,I35863,I35812,I35885,I125572,I35911,I35919,I35936,I125560,I35953,I125551,I35970,I35987,I125557,I36004,I125575,I36021,I125548,I36038,I35788,I36069,I36086,I36103,I36120,I35800,I35794,I36165,I125554,I35809,I35803,I36210,I36227,I125566,I36244,I36261,I125569,I36287,I36295,I35797,I35791,I36349,I36357,I35806,I36415,I47535,I36441,I36458,I36407,I36480,I47550,I36506,I36514,I36531,I47547,I36548,I36565,I36582,I47544,I36599,I47559,I36616,I47556,I36633,I36383,I36664,I36681,I36698,I36715,I36395,I36389,I36760,I47553,I36404,I36398,I36805,I36822,I47541,I36839,I47562,I36856,I47538,I36882,I36890,I36392,I36386,I36944,I36952,I36401,I37010,I37036,I37053,I37002,I37075,I37101,I37109,I37126,I37143,I37160,I37177,I37194,I37211,I37228,I36978,I37259,I37276,I37293,I37310,I36990,I36984,I37355,I36999,I36993,I37400,I37417,I37434,I37451,I37477,I37485,I36987,I36981,I37539,I37547,I36996,I37605,I173475,I37631,I37648,I37597,I37670,I173466,I37696,I37704,I37721,I173460,I37738,I173454,I37755,I37772,I173481,I37789,I37806,I173478,I37823,I37573,I37854,I37871,I37888,I37905,I37585,I37579,I37950,I173463,I37594,I37588,I37995,I38012,I173469,I38029,I173472,I38046,I173457,I38072,I38080,I37582,I37576,I38134,I38142,I37591,I38200,I175855,I38226,I38243,I38192,I38265,I175846,I38291,I38299,I38316,I175840,I38333,I175834,I38350,I38367,I175861,I38384,I38401,I175858,I38418,I38168,I38449,I38466,I38483,I38500,I38180,I38174,I38545,I175843,I38189,I38183,I38590,I38607,I175849,I38624,I175852,I38641,I175837,I38667,I38675,I38177,I38171,I38729,I38737,I38186,I38795,I38821,I38838,I38787,I38860,I38886,I38894,I38911,I38928,I38945,I38962,I38979,I38996,I39013,I38763,I39044,I39061,I39078,I39095,I38775,I38769,I39140,I38784,I38778,I39185,I39202,I39219,I39236,I39262,I39270,I38772,I38766,I39324,I39332,I38781,I39390,I39416,I39433,I39382,I39455,I39481,I39489,I39506,I39523,I39540,I39557,I39574,I39591,I39608,I39358,I39639,I39656,I39673,I39690,I39370,I39364,I39735,I39379,I39373,I39780,I39797,I39814,I39831,I39857,I39865,I39367,I39361,I39919,I39927,I39376,I39985,I40011,I40028,I39977,I40050,I40076,I40084,I40101,I40118,I40135,I40152,I40169,I40186,I40203,I39953,I40234,I40251,I40268,I40285,I39965,I39959,I40330,I39974,I39968,I40375,I40392,I40409,I40426,I40452,I40460,I39962,I39956,I40514,I40522,I39971,I40580,I42792,I40606,I40623,I40572,I40645,I42807,I40671,I40679,I40696,I42804,I40713,I40730,I40747,I42801,I40764,I42816,I40781,I42813,I40798,I40548,I40829,I40846,I40863,I40880,I40560,I40554,I40925,I42810,I40569,I40563,I40970,I40987,I42798,I41004,I42819,I41021,I42795,I41047,I41055,I40557,I40551,I41109,I41117,I40566,I41175,I152408,I41201,I41218,I41167,I41240,I41266,I41274,I41291,I152411,I41308,I152423,I41325,I41342,I152429,I41359,I152420,I41376,I152426,I41393,I41143,I41424,I41441,I41458,I41475,I41155,I41149,I41520,I152417,I41164,I41158,I41565,I41582,I152414,I41599,I152432,I41616,I41642,I41650,I41152,I41146,I41704,I41712,I41161,I41773,I41799,I41807,I41824,I41850,I41741,I41872,I41898,I41906,I41923,I41949,I41765,I41971,I41747,I42011,I42028,I42036,I42053,I41750,I42084,I42101,I42127,I42135,I41738,I41756,I42180,I42197,I41759,I41744,I41753,I41762,I42300,I147784,I42326,I42334,I147799,I42351,I147802,I42377,I42268,I42399,I147808,I42425,I42433,I147790,I42450,I42476,I42292,I42498,I42274,I147787,I42538,I42555,I42563,I42580,I42277,I42611,I147793,I42628,I147805,I42654,I42662,I42265,I42283,I42707,I147796,I42724,I42286,I42271,I42280,I42289,I42827,I42853,I42861,I42878,I42904,I42926,I42952,I42960,I42977,I43003,I43025,I43065,I43082,I43090,I43107,I43138,I43155,I43181,I43189,I43234,I43251,I43354,I97510,I43380,I43388,I97501,I97516,I43405,I97522,I43431,I43322,I43453,I97507,I43479,I43487,I43504,I43530,I43346,I43552,I43328,I97504,I43592,I43609,I43617,I43634,I43331,I43665,I97498,I97513,I43682,I43708,I43716,I43319,I43337,I43761,I97519,I43778,I43340,I43325,I43334,I43343,I43881,I140270,I43907,I43915,I140285,I43932,I140288,I43958,I43980,I140294,I44006,I44014,I140276,I44031,I44057,I44079,I140273,I44119,I44136,I44144,I44161,I44192,I140279,I44209,I140291,I44235,I44243,I44288,I140282,I44305,I44408,I115215,I44434,I44442,I115212,I115230,I44459,I115221,I44485,I44507,I115236,I44533,I44541,I115218,I44558,I44584,I44606,I115224,I44646,I44663,I44671,I44688,I44719,I115239,I44736,I115227,I44762,I44770,I44815,I115233,I44832,I44935,I145472,I44961,I44969,I145487,I44986,I145490,I45012,I44903,I45034,I145496,I45060,I45068,I145478,I45085,I45111,I44927,I45133,I44909,I145475,I45173,I45190,I45198,I45215,I44912,I45246,I145481,I45263,I145493,I45289,I45297,I44900,I44918,I45342,I145484,I45359,I44921,I44906,I44915,I44924,I45462,I45488,I45496,I45513,I45539,I45430,I45561,I45587,I45595,I45612,I45638,I45454,I45660,I45436,I45700,I45717,I45725,I45742,I45439,I45773,I45790,I45816,I45824,I45427,I45445,I45869,I45886,I45448,I45433,I45442,I45451,I45989,I164663,I46015,I46023,I164660,I164651,I46040,I164648,I46066,I45957,I46088,I164657,I46114,I46122,I164666,I46139,I46165,I45981,I46187,I45963,I164669,I46227,I46244,I46252,I46269,I45966,I46300,I164654,I46317,I164672,I46343,I46351,I45954,I45972,I46396,I46413,I45975,I45960,I45969,I45978,I46516,I144316,I46542,I46550,I144331,I46567,I144334,I46593,I46484,I46615,I144340,I46641,I46649,I144322,I46666,I46692,I46508,I46714,I46490,I144319,I46754,I46771,I46779,I46796,I46493,I46827,I144325,I46844,I144337,I46870,I46878,I46481,I46499,I46923,I144328,I46940,I46502,I46487,I46496,I46505,I47043,I156812,I47069,I47077,I156794,I156818,I47094,I156809,I47120,I47011,I47142,I156815,I47168,I47176,I156803,I47193,I47219,I47035,I47241,I47017,I47281,I47298,I47306,I47323,I47020,I47354,I156800,I156797,I47371,I156806,I47397,I47405,I47008,I47026,I47450,I47467,I47029,I47014,I47023,I47032,I47570,I47596,I47604,I47621,I47647,I47669,I47695,I47703,I47720,I47746,I47768,I47808,I47825,I47833,I47850,I47881,I47898,I47924,I47932,I47977,I47994,I48097,I162929,I48123,I48131,I162926,I162917,I48148,I162914,I48174,I48065,I48196,I162923,I48222,I48230,I162932,I48247,I48273,I48089,I48295,I48071,I162935,I48335,I48352,I48360,I48377,I48074,I48408,I162920,I48425,I162938,I48451,I48459,I48062,I48080,I48504,I48521,I48083,I48068,I48077,I48086,I48624,I149518,I48650,I48658,I149533,I48675,I149536,I48701,I48592,I48723,I149542,I48749,I48757,I149524,I48774,I48800,I48616,I48822,I48598,I149521,I48862,I48879,I48887,I48904,I48601,I48935,I149527,I48952,I149539,I48978,I48986,I48589,I48607,I49031,I149530,I49048,I48610,I48595,I48604,I48613,I49151,I130634,I49177,I49185,I130631,I49202,I130643,I49228,I49250,I49276,I49284,I130649,I49301,I49327,I49349,I130637,I49389,I49406,I49414,I49431,I49462,I130646,I130652,I49479,I49505,I49513,I49558,I130640,I49575,I49678,I108653,I49704,I49712,I108656,I108650,I49729,I108662,I49755,I49646,I49777,I108665,I49803,I49811,I49828,I49854,I49670,I49876,I49652,I108668,I49916,I49933,I49941,I49958,I49655,I49989,I108659,I50006,I50032,I50040,I49643,I49661,I50085,I108671,I50102,I49664,I49649,I49658,I49667,I50205,I171690,I50231,I50239,I171669,I50256,I171696,I50282,I50304,I171684,I50330,I50338,I171687,I50355,I50381,I50403,I171678,I50443,I50460,I50468,I50485,I50516,I171675,I171672,I50533,I171693,I50559,I50567,I50612,I171681,I50629,I50732,I109707,I50758,I50766,I109710,I109704,I50783,I109716,I50809,I50831,I109719,I50857,I50865,I50882,I50908,I50930,I109722,I50970,I50987,I50995,I51012,I51043,I109713,I51060,I51086,I51094,I51139,I109725,I51156,I51259,I51285,I51293,I51310,I51336,I51227,I51358,I51384,I51392,I51409,I51435,I51251,I51457,I51233,I51497,I51514,I51522,I51539,I51236,I51570,I51587,I51613,I51621,I51224,I51242,I51666,I51683,I51245,I51230,I51239,I51248,I51786,I84219,I51812,I51820,I84204,I84207,I51837,I84222,I51863,I51754,I51885,I84216,I51911,I51919,I51936,I51962,I51778,I51984,I51760,I84213,I52024,I52041,I52049,I52066,I51763,I52097,I84228,I52114,I84225,I52140,I52148,I51751,I51769,I52193,I84210,I52210,I51772,I51757,I51766,I51775,I52313,I113923,I52339,I52347,I113920,I113938,I52364,I113929,I52390,I52412,I113944,I52438,I52446,I113926,I52463,I52489,I52511,I113932,I52551,I52568,I52576,I52593,I52624,I113947,I52641,I113935,I52667,I52675,I52720,I113941,I52737,I52840,I106545,I52866,I52874,I106548,I106542,I52891,I106554,I52917,I52808,I52939,I106557,I52965,I52973,I52990,I53016,I52832,I53038,I52814,I106560,I53078,I53095,I53103,I53120,I52817,I53151,I106551,I53168,I53194,I53202,I52805,I52823,I53247,I106563,I53264,I52826,I52811,I52820,I52829,I53367,I165819,I53393,I53401,I165816,I165807,I53418,I165804,I53444,I53466,I165813,I53492,I53500,I165822,I53517,I53543,I53565,I165825,I53605,I53622,I53630,I53647,I53678,I165810,I53695,I165828,I53721,I53729,I53774,I53791,I53894,I53920,I53928,I53945,I53971,I53993,I54019,I54027,I54044,I54070,I54092,I54132,I54149,I54157,I54174,I54205,I54222,I54248,I54256,I54301,I54318,I54421,I54447,I54455,I54472,I54498,I54389,I54520,I54546,I54554,I54571,I54597,I54413,I54619,I54395,I54659,I54676,I54684,I54701,I54398,I54732,I54749,I54775,I54783,I54386,I54404,I54828,I54845,I54407,I54392,I54401,I54410,I54948,I177045,I54974,I54982,I177024,I54999,I177051,I55025,I54916,I55047,I177039,I55073,I55081,I177042,I55098,I55124,I54940,I55146,I54922,I177033,I55186,I55203,I55211,I55228,I54925,I55259,I177030,I177027,I55276,I177048,I55302,I55310,I54913,I54931,I55355,I177036,I55372,I54934,I54919,I54928,I54937,I55475,I78439,I55501,I55509,I78424,I78427,I55526,I78442,I55552,I55443,I55574,I78436,I55600,I55608,I55625,I55651,I55467,I55673,I55449,I78433,I55713,I55730,I55738,I55755,I55452,I55786,I78448,I55803,I78445,I55829,I55837,I55440,I55458,I55882,I78430,I55899,I55461,I55446,I55455,I55464,I56002,I68924,I56028,I56036,I68936,I56053,I68921,I56079,I55970,I56101,I68945,I56127,I56135,I68942,I56152,I56178,I55994,I56200,I55976,I68933,I56240,I56257,I56265,I56282,I55979,I56313,I68930,I56330,I68939,I56356,I56364,I55967,I55985,I56409,I68927,I56426,I55988,I55973,I55982,I55991,I56529,I56555,I56563,I56580,I56606,I56497,I56628,I56654,I56662,I56679,I56705,I56521,I56727,I56503,I56767,I56784,I56792,I56809,I56506,I56840,I56857,I56883,I56891,I56494,I56512,I56936,I56953,I56515,I56500,I56509,I56518,I57056,I118445,I57082,I57090,I118442,I118460,I57107,I118451,I57133,I57024,I57155,I118466,I57181,I57189,I118448,I57206,I57232,I57048,I57254,I57030,I118454,I57294,I57311,I57319,I57336,I57033,I57367,I118469,I57384,I118457,I57410,I57418,I57021,I57039,I57463,I118463,I57480,I57042,I57027,I57036,I57045,I57583,I57609,I57617,I57634,I57660,I57682,I57708,I57716,I57733,I57759,I57781,I57821,I57838,I57846,I57863,I57894,I57911,I57937,I57945,I57990,I58007,I58110,I117153,I58136,I58144,I117150,I117168,I58161,I117159,I58187,I58078,I58209,I117174,I58235,I58243,I117156,I58260,I58286,I58102,I58308,I58084,I117162,I58348,I58365,I58373,I58390,I58087,I58421,I117177,I58438,I117165,I58464,I58472,I58075,I58093,I58517,I117171,I58534,I58096,I58081,I58090,I58099,I58637,I62949,I58663,I58671,I62961,I62940,I58688,I62964,I58714,I58605,I58736,I62955,I58762,I58770,I62937,I58787,I58813,I58629,I58835,I58611,I62952,I58875,I58892,I58900,I58917,I58614,I58948,I62943,I58965,I62946,I58991,I58999,I58602,I58620,I59044,I62958,I59061,I58623,I58608,I58617,I58626,I59164,I138539,I59190,I59207,I59156,I59229,I59246,I138551,I59263,I138542,I59289,I59297,I138560,I59323,I59331,I138536,I59348,I59135,I138554,I59388,I59396,I59129,I59144,I59441,I138548,I138545,I59458,I138557,I59484,I59132,I59506,I59523,I59540,I59147,I59571,I59588,I59138,I59619,I59141,I59153,I59150,I59708,I59734,I59751,I59700,I59773,I59790,I59807,I59833,I59841,I59867,I59875,I59892,I59679,I59932,I59940,I59673,I59688,I59985,I60002,I60028,I59676,I60050,I60067,I60084,I59691,I60115,I60132,I59682,I60163,I59685,I59697,I59694,I60252,I100969,I60278,I60295,I60244,I60317,I60334,I100990,I100981,I60351,I60377,I60385,I100975,I60411,I60419,I100972,I60436,I60223,I100966,I60476,I60484,I60217,I60232,I60529,I100978,I60546,I100987,I60572,I60220,I60594,I60611,I60628,I60235,I60659,I60676,I100984,I60226,I60707,I60229,I60241,I60238,I60796,I155709,I60822,I60839,I60788,I60861,I60878,I155721,I155724,I60895,I155727,I60921,I60929,I155712,I60955,I60963,I155718,I60980,I60767,I155706,I61020,I61028,I60761,I60776,I61073,I155730,I61090,I155715,I61116,I60764,I61138,I61155,I61172,I60779,I61203,I61220,I60770,I61251,I60773,I60785,I60782,I61340,I143163,I61366,I61383,I61405,I61422,I143175,I61439,I143166,I61465,I61473,I143184,I61499,I61507,I143160,I61524,I143178,I61564,I61572,I61617,I143172,I143169,I61634,I143181,I61660,I61682,I61699,I61716,I61747,I61764,I61795,I61884,I142585,I61910,I61927,I61876,I61949,I61966,I142597,I61983,I142588,I62009,I62017,I142606,I62043,I62051,I142582,I62068,I61855,I142600,I62108,I62116,I61849,I61864,I62161,I142594,I142591,I62178,I142603,I62204,I61852,I62226,I62243,I62260,I61867,I62291,I62308,I61858,I62339,I61861,I61873,I61870,I62428,I62454,I62471,I62420,I62493,I62510,I62527,I62553,I62561,I62587,I62595,I62612,I62399,I62652,I62660,I62393,I62408,I62705,I62722,I62748,I62396,I62770,I62787,I62804,I62411,I62835,I62852,I62402,I62883,I62405,I62417,I62414,I62972,I107081,I62998,I63015,I63037,I63054,I107075,I107072,I63071,I107087,I63097,I63105,I63131,I63139,I107069,I63156,I63196,I63204,I63249,I107084,I107078,I63266,I63292,I63314,I63331,I63348,I63379,I63396,I107090,I63427,I63516,I63542,I63559,I63508,I63581,I63598,I63615,I63641,I63649,I63675,I63683,I63700,I63487,I63740,I63748,I63481,I63496,I63793,I63810,I63836,I63484,I63858,I63875,I63892,I63499,I63923,I63940,I63490,I63971,I63493,I63505,I63502,I64060,I64086,I64103,I64052,I64125,I64142,I64159,I64185,I64193,I64219,I64227,I64244,I64031,I64284,I64292,I64025,I64040,I64337,I64354,I64380,I64028,I64402,I64419,I64436,I64043,I64467,I64484,I64034,I64515,I64037,I64049,I64046,I64604,I64630,I64647,I64596,I64669,I64686,I64703,I64729,I64737,I64763,I64771,I64788,I64575,I64828,I64836,I64569,I64584,I64881,I64898,I64924,I64572,I64946,I64963,I64980,I64587,I65011,I65028,I64578,I65059,I64581,I64593,I64590,I65148,I65174,I65191,I65140,I65213,I65230,I65247,I65273,I65281,I65307,I65315,I65332,I65119,I65372,I65380,I65113,I65128,I65425,I65442,I65468,I65116,I65490,I65507,I65524,I65131,I65555,I65572,I65122,I65603,I65125,I65137,I65134,I65692,I65718,I65735,I65684,I65757,I65774,I65791,I65817,I65825,I65851,I65859,I65876,I65663,I65916,I65924,I65657,I65672,I65969,I65986,I66012,I65660,I66034,I66051,I66068,I65675,I66099,I66116,I65666,I66147,I65669,I65681,I65678,I66236,I127492,I66262,I66279,I66228,I66301,I66318,I127507,I127495,I66335,I127486,I66361,I66369,I127498,I66395,I66403,I127489,I66420,I66207,I127504,I66460,I66468,I66201,I66216,I66513,I127513,I127501,I66530,I127510,I66556,I66204,I66578,I66595,I66612,I66219,I66643,I66660,I66210,I66691,I66213,I66225,I66222,I66780,I147209,I66806,I66823,I66772,I66845,I66862,I147221,I66879,I147212,I66905,I66913,I147230,I66939,I66947,I147206,I66964,I66751,I147224,I67004,I67012,I66745,I66760,I67057,I147218,I147215,I67074,I147227,I67100,I66748,I67122,I67139,I67156,I66763,I67187,I67204,I66754,I67235,I66757,I66769,I66766,I67324,I115864,I67350,I67367,I67389,I67406,I115879,I115867,I67423,I115858,I67449,I67457,I115870,I67483,I67491,I115861,I67508,I115876,I67548,I67556,I67601,I115885,I115873,I67618,I115882,I67644,I67666,I67683,I67700,I67731,I67748,I67779,I67868,I67894,I67911,I67933,I67950,I67967,I67993,I68001,I68027,I68035,I68052,I68092,I68100,I68145,I68162,I68188,I68210,I68227,I68244,I68275,I68292,I68323,I68412,I68438,I68455,I68477,I68494,I68511,I68537,I68545,I68571,I68579,I68596,I68636,I68644,I68689,I68706,I68732,I68754,I68771,I68788,I68819,I68836,I68867,I68953,I110240,I68979,I68996,I110237,I69027,I69035,I69052,I69069,I110234,I69086,I110249,I69103,I69120,I69137,I69168,I110243,I69185,I110231,I69202,I69247,I69264,I69295,I110252,I69312,I69343,I69360,I110246,I69377,I69403,I69411,I69442,I69459,I69490,I69548,I69574,I69591,I69622,I69630,I69647,I69664,I69681,I69698,I69715,I69732,I69763,I69780,I69797,I69842,I69859,I69890,I69907,I69938,I69955,I69972,I69998,I70006,I70037,I70054,I70085,I70143,I70169,I70186,I70135,I70217,I70225,I70242,I70259,I70276,I70293,I70310,I70327,I70132,I70358,I70375,I70392,I70117,I70129,I70437,I70454,I70123,I70485,I70502,I70111,I70533,I70550,I70567,I70593,I70601,I70120,I70632,I70649,I70126,I70680,I70114,I70738,I70764,I70781,I70812,I70820,I70837,I70854,I70871,I70888,I70905,I70922,I70953,I70970,I70987,I71032,I71049,I71080,I71097,I71128,I71145,I71162,I71188,I71196,I71227,I71244,I71275,I71333,I80739,I71359,I71376,I71325,I80751,I71407,I71415,I80736,I71432,I71449,I80754,I71466,I80745,I71483,I71500,I71517,I71322,I71548,I80757,I71565,I80760,I71582,I71307,I71319,I71627,I71644,I71313,I71675,I71692,I71301,I71723,I80748,I71740,I80742,I71757,I71783,I71791,I71310,I71822,I71839,I71316,I71870,I71304,I71928,I71954,I71971,I71920,I72002,I72010,I72027,I72044,I72061,I72078,I72095,I72112,I71917,I72143,I72160,I72177,I71902,I71914,I72222,I72239,I71908,I72270,I72287,I71896,I72318,I72335,I72352,I72378,I72386,I71905,I72417,I72434,I71911,I72465,I71899,I72523,I135119,I72549,I72566,I72515,I135122,I72597,I72605,I135125,I72622,I72639,I135137,I72656,I135128,I72673,I72690,I72707,I72512,I72738,I135134,I72755,I72772,I72497,I72509,I72817,I72834,I72503,I72865,I72882,I72491,I72913,I135131,I72930,I72947,I135140,I72973,I72981,I72500,I73012,I73029,I72506,I73060,I72494,I73118,I73144,I73161,I73110,I73192,I73200,I73217,I73234,I73251,I73268,I73285,I73302,I73107,I73333,I73350,I73367,I73092,I73104,I73412,I73429,I73098,I73460,I73477,I73086,I73508,I73525,I73542,I73568,I73576,I73095,I73607,I73624,I73101,I73655,I73089,I73713,I119749,I73739,I73756,I73705,I119737,I73787,I73795,I119734,I73812,I73829,I119746,I73846,I119743,I73863,I73880,I73897,I73702,I73928,I119752,I73945,I119755,I73962,I73687,I73699,I74007,I74024,I73693,I74055,I119758,I74072,I73681,I74103,I119761,I74120,I119740,I74137,I74163,I74171,I73690,I74202,I74219,I73696,I74250,I73684,I74308,I87103,I74334,I74351,I87097,I74382,I74390,I87094,I74407,I74424,I87106,I74441,I87109,I74458,I74475,I74492,I74523,I87118,I74540,I87112,I74557,I74602,I74619,I74650,I87100,I74667,I74698,I87115,I74715,I74732,I74758,I74766,I74797,I74814,I74845,I74903,I92883,I74929,I74946,I92877,I74977,I74985,I92874,I75002,I75019,I92886,I75036,I92889,I75053,I75070,I75087,I75118,I92898,I75135,I92892,I75152,I75197,I75214,I75245,I92880,I75262,I75293,I92895,I75310,I75327,I75353,I75361,I75392,I75409,I75440,I75498,I75524,I75541,I75572,I75580,I75597,I75614,I75631,I75648,I75665,I75682,I75713,I75730,I75747,I75792,I75809,I75840,I75857,I75888,I75905,I75922,I75948,I75956,I75987,I76004,I76035,I76093,I76119,I76136,I76085,I76167,I76175,I76192,I76209,I76226,I76243,I76260,I76277,I76082,I76308,I76325,I76342,I76067,I76079,I76387,I76404,I76073,I76435,I76452,I76061,I76483,I76500,I76517,I76543,I76551,I76070,I76582,I76599,I76076,I76630,I76064,I76688,I154074,I76714,I76731,I76680,I154089,I76762,I76770,I154098,I76787,I76804,I154077,I76821,I154083,I76838,I76855,I76872,I76677,I76903,I154095,I76920,I154092,I76937,I76662,I76674,I76982,I76999,I76668,I77030,I77047,I76656,I77078,I154086,I77095,I154080,I77112,I77138,I77146,I76665,I77177,I77194,I76671,I77225,I76659,I77283,I105497,I77309,I77326,I77275,I105494,I77357,I77365,I77382,I77399,I105491,I77416,I105506,I77433,I77450,I77467,I77272,I77498,I105500,I77515,I105488,I77532,I77257,I77269,I77577,I77594,I77263,I77625,I105509,I77642,I77251,I77673,I77690,I105503,I77707,I77733,I77741,I77260,I77772,I77789,I77266,I77820,I77254,I77878,I124908,I77904,I77912,I124905,I77938,I77946,I124902,I77963,I124929,I77980,I77997,I124917,I78014,I77864,I78045,I78062,I78079,I124923,I78096,I124914,I77861,I77852,I78141,I77855,I77849,I78186,I124911,I78203,I78220,I77858,I78251,I124926,I78268,I124920,I78285,I78311,I78319,I77846,I77870,I78364,I78381,I78398,I77867,I78456,I78482,I78490,I78516,I78524,I78541,I78558,I78575,I78592,I78623,I78640,I78657,I78674,I78719,I78764,I78781,I78798,I78829,I78846,I78863,I78889,I78897,I78942,I78959,I78976,I79034,I79060,I79068,I79094,I79102,I79119,I79136,I79153,I79170,I79020,I79201,I79218,I79235,I79252,I79017,I79008,I79297,I79011,I79005,I79342,I79359,I79376,I79014,I79407,I79424,I79441,I79467,I79475,I79002,I79026,I79520,I79537,I79554,I79023,I79612,I131774,I79638,I79646,I131765,I79672,I79680,I131759,I79697,I131771,I79714,I79731,I131762,I79748,I79779,I79796,I79813,I131768,I79830,I131753,I79875,I79920,I79937,I79954,I79985,I131756,I80002,I80019,I80045,I80053,I80098,I80115,I80132,I80190,I80216,I80224,I80250,I80258,I80275,I80292,I80309,I80326,I80176,I80357,I80374,I80391,I80408,I80173,I80164,I80453,I80167,I80161,I80498,I80515,I80532,I80170,I80563,I80580,I80597,I80623,I80631,I80158,I80182,I80676,I80693,I80710,I80179,I80768,I128138,I80794,I80802,I128135,I80828,I80836,I128132,I80853,I128159,I80870,I80887,I128147,I80904,I80935,I80952,I80969,I128153,I80986,I128144,I81031,I81076,I128141,I81093,I81110,I81141,I128156,I81158,I128150,I81175,I81201,I81209,I81254,I81271,I81288,I81346,I81372,I81380,I81406,I81414,I81431,I81448,I81465,I81482,I81332,I81513,I81530,I81547,I81564,I81329,I81320,I81609,I81323,I81317,I81654,I81671,I81688,I81326,I81719,I81736,I81753,I81779,I81787,I81314,I81338,I81832,I81849,I81866,I81335,I81924,I81950,I81958,I81984,I81992,I82009,I82026,I82043,I82060,I81910,I82091,I82108,I82125,I82142,I81907,I81898,I82187,I81901,I81895,I82232,I82249,I82266,I81904,I82297,I82314,I82331,I82357,I82365,I81892,I81916,I82410,I82427,I82444,I81913,I82502,I122970,I82528,I82536,I122967,I82562,I82570,I122964,I82587,I122991,I82604,I82621,I122979,I82638,I82488,I82669,I82686,I82703,I122985,I82720,I122976,I82485,I82476,I82765,I82479,I82473,I82810,I122973,I82827,I82844,I82482,I82875,I122988,I82892,I122982,I82909,I82935,I82943,I82470,I82494,I82988,I83005,I83022,I82491,I83080,I175239,I83106,I83114,I83140,I83148,I175263,I83165,I175245,I83182,I83199,I175260,I83216,I83066,I83247,I83264,I83281,I175242,I83298,I175251,I83063,I83054,I83343,I83057,I83051,I83388,I175248,I83405,I83422,I83060,I83453,I175257,I83470,I175266,I83487,I175254,I83513,I83521,I83048,I83072,I83566,I83583,I83600,I83069,I83658,I144894,I83684,I83692,I144900,I83718,I83726,I83743,I144897,I83760,I83777,I144915,I83794,I83825,I83842,I83859,I144918,I83876,I83921,I83966,I144903,I83983,I84000,I84031,I144909,I84048,I144906,I84065,I144912,I84091,I84099,I84144,I84161,I84178,I84236,I159532,I84262,I84270,I159526,I84296,I84304,I159535,I84321,I159514,I84338,I84355,I159523,I84372,I84403,I84420,I84437,I159538,I84454,I159517,I84499,I84544,I159520,I84561,I84578,I84609,I159529,I84626,I84643,I84669,I84677,I84722,I84739,I84756,I84814,I161770,I84840,I84848,I161782,I84874,I84882,I161773,I84899,I161761,I84916,I84933,I161758,I84950,I84981,I84998,I85015,I161764,I85032,I85077,I85122,I161779,I85139,I85156,I85187,I161767,I85204,I85221,I161776,I85247,I85255,I85300,I85317,I85334,I85392,I94608,I85418,I85426,I94620,I85452,I85460,I94611,I85477,I94614,I85494,I85511,I94617,I85528,I85559,I85576,I85593,I85610,I94623,I85655,I85700,I94629,I85717,I85734,I85765,I85782,I94626,I85799,I94632,I85825,I85833,I85878,I85895,I85912,I85970,I85996,I86004,I86030,I86038,I86055,I86072,I86089,I86106,I85956,I86137,I86154,I86171,I86188,I85953,I85944,I86233,I85947,I85941,I86278,I86295,I86312,I85950,I86343,I86360,I86377,I86403,I86411,I85938,I85962,I86456,I86473,I86490,I85959,I86548,I86574,I86582,I86599,I86616,I86642,I86650,I86676,I86684,I86701,I86718,I86735,I86531,I86775,I86783,I86800,I86817,I86834,I86534,I86865,I86882,I86908,I86916,I86516,I86947,I86525,I86978,I86995,I86537,I87026,I86528,I86519,I86522,I86540,I87126,I119112,I87152,I87160,I87177,I119088,I119103,I87194,I119115,I87220,I87228,I119100,I119091,I87254,I87262,I87279,I87296,I87313,I87353,I87361,I87378,I87395,I87412,I87443,I119106,I119097,I87460,I119109,I87486,I87494,I87525,I87556,I87573,I87604,I119094,I87704,I166397,I87730,I87738,I87755,I166385,I166403,I87772,I166394,I87798,I87806,I166409,I166406,I87832,I87840,I87857,I87874,I87891,I166388,I87931,I87939,I87956,I87973,I87990,I88021,I166382,I88038,I166391,I88064,I88072,I88103,I88134,I88151,I88182,I166400,I88282,I121696,I88308,I88316,I88333,I121672,I121687,I88350,I121699,I88376,I88384,I121684,I121675,I88410,I88418,I88435,I88452,I88469,I88265,I88509,I88517,I88534,I88551,I88568,I88268,I88599,I121690,I121681,I88616,I121693,I88642,I88650,I88250,I88681,I88259,I88712,I88729,I88271,I88760,I121678,I88262,I88253,I88256,I88274,I88860,I122342,I88886,I88894,I88911,I122318,I122333,I88928,I122345,I88954,I88962,I122330,I122321,I88988,I88996,I89013,I89030,I89047,I88843,I89087,I89095,I89112,I89129,I89146,I88846,I89177,I122336,I122327,I89194,I122339,I89220,I89228,I88828,I89259,I88837,I89290,I89307,I88849,I89338,I122324,I88840,I88831,I88834,I88852,I89438,I89464,I89472,I89489,I89506,I89532,I89540,I89566,I89574,I89591,I89608,I89625,I89665,I89673,I89690,I89707,I89724,I89755,I89772,I89798,I89806,I89837,I89868,I89885,I89916,I90016,I90042,I90050,I90067,I90084,I90110,I90118,I90144,I90152,I90169,I90186,I90203,I90243,I90251,I90268,I90285,I90302,I90333,I90350,I90376,I90384,I90415,I90446,I90463,I90494,I90594,I90620,I90628,I90645,I90662,I90688,I90696,I90722,I90730,I90747,I90764,I90781,I90821,I90829,I90846,I90863,I90880,I90911,I90928,I90954,I90962,I90993,I91024,I91041,I91072,I91172,I91198,I91206,I91223,I91240,I91266,I91274,I91300,I91308,I91325,I91342,I91359,I91155,I91399,I91407,I91424,I91441,I91458,I91158,I91489,I91506,I91532,I91540,I91140,I91571,I91149,I91602,I91619,I91161,I91650,I91152,I91143,I91146,I91164,I91750,I132881,I91776,I91784,I91801,I132878,I132896,I91818,I132893,I91844,I91852,I132875,I91878,I91886,I91903,I91920,I91937,I132887,I91977,I91985,I92002,I92019,I92036,I92067,I132890,I92084,I92110,I92118,I92149,I92180,I92197,I92228,I132884,I92328,I92354,I92362,I92379,I92396,I92422,I92430,I92456,I92464,I92481,I92498,I92515,I92555,I92563,I92580,I92597,I92614,I92645,I92662,I92688,I92696,I92727,I92758,I92775,I92806,I92906,I116528,I92932,I92940,I92957,I116504,I116519,I92974,I116531,I93000,I93008,I116516,I116507,I93034,I93042,I93059,I93076,I93093,I93133,I93141,I93158,I93175,I93192,I93223,I116522,I116513,I93240,I116525,I93266,I93274,I93305,I93336,I93353,I93384,I116510,I93484,I129448,I93510,I93518,I93535,I129424,I129439,I93552,I129451,I93578,I93586,I129436,I129427,I93612,I93620,I93637,I93654,I93671,I93467,I93711,I93719,I93736,I93753,I93770,I93470,I93801,I129442,I129433,I93818,I129445,I93844,I93852,I93452,I93883,I93461,I93914,I93931,I93473,I93962,I129430,I93464,I93455,I93458,I93476,I94062,I94088,I94096,I94113,I94130,I94156,I94164,I94190,I94198,I94215,I94232,I94249,I94045,I94289,I94297,I94314,I94331,I94348,I94048,I94379,I94396,I94422,I94430,I94030,I94461,I94039,I94492,I94509,I94051,I94540,I94042,I94033,I94036,I94054,I94640,I148958,I94666,I94674,I94691,I148940,I148952,I94708,I148955,I94734,I94742,I148949,I148946,I94768,I94776,I94793,I94810,I94827,I148964,I94867,I94875,I94892,I94909,I94926,I94957,I148943,I94974,I95000,I95008,I95039,I95070,I95087,I95118,I148961,I95218,I95244,I95252,I95269,I95286,I95312,I95320,I95346,I95354,I95371,I95388,I95405,I95201,I95445,I95453,I95470,I95487,I95504,I95204,I95535,I95552,I95578,I95586,I95186,I95617,I95195,I95648,I95665,I95207,I95696,I95198,I95189,I95192,I95210,I95796,I177646,I95822,I95830,I95847,I177631,I177619,I95864,I177634,I95890,I95898,I177637,I95924,I95932,I95949,I95966,I95983,I95779,I177625,I96023,I96031,I96048,I96065,I96082,I95782,I96113,I177622,I177628,I96130,I177643,I96156,I96164,I95764,I96195,I95773,I96226,I96243,I95785,I96274,I177640,I95776,I95767,I95770,I95788,I96374,I96400,I96408,I96425,I96442,I96468,I96476,I96502,I96510,I96527,I96544,I96561,I96357,I96601,I96609,I96626,I96643,I96660,I96360,I96691,I96708,I96734,I96742,I96342,I96773,I96351,I96804,I96821,I96363,I96852,I96354,I96345,I96348,I96366,I96952,I96978,I96986,I97003,I97020,I97046,I97054,I97080,I97088,I97105,I97122,I97139,I96935,I97179,I97187,I97204,I97221,I97238,I96938,I97269,I97286,I97312,I97320,I96920,I97351,I96929,I97382,I97399,I96941,I97430,I96932,I96923,I96926,I96944,I97530,I133442,I97556,I97564,I97581,I133439,I133457,I97598,I133454,I97624,I97632,I133436,I97658,I97666,I97683,I97700,I97717,I133448,I97757,I97765,I97782,I97799,I97816,I97847,I133451,I97864,I97890,I97898,I97929,I97960,I97977,I98008,I133445,I98108,I126218,I98134,I98142,I98159,I126194,I126209,I98176,I126221,I98202,I98210,I126206,I126197,I98236,I98244,I98261,I98278,I98295,I98335,I98343,I98360,I98377,I98394,I98425,I126212,I126203,I98442,I126215,I98468,I98476,I98507,I98538,I98555,I98586,I126200,I98686,I98712,I98720,I98737,I98754,I98780,I98788,I98814,I98822,I98839,I98856,I98873,I98669,I98913,I98921,I98938,I98955,I98972,I98672,I99003,I99020,I99046,I99054,I98654,I99085,I98663,I99116,I99133,I98675,I99164,I98666,I98657,I98660,I98678,I99264,I137976,I99290,I99298,I99315,I137958,I137970,I99332,I137973,I99358,I99366,I137967,I137964,I99392,I99400,I99417,I99434,I99451,I99247,I137982,I99491,I99499,I99516,I99533,I99550,I99250,I99581,I137961,I99598,I99624,I99632,I99232,I99663,I99241,I99694,I99711,I99253,I99742,I137979,I99244,I99235,I99238,I99256,I99842,I158970,I99868,I99876,I99893,I158973,I158982,I99910,I158985,I99936,I99944,I158994,I158976,I99970,I99978,I99995,I100012,I100029,I99825,I100069,I100077,I100094,I100111,I100128,I99828,I100159,I158991,I100176,I158988,I100202,I100210,I99810,I100241,I99819,I100272,I100289,I99831,I100320,I158979,I99822,I99813,I99816,I99834,I100420,I111300,I100446,I100454,I100471,I111288,I111306,I100488,I111303,I100514,I100522,I111294,I111291,I100548,I100556,I100573,I100590,I100607,I111285,I100647,I100655,I100672,I100689,I100706,I100737,I100754,I100780,I100788,I100819,I100850,I100867,I100898,I111297,I100998,I167531,I101024,I101032,I101049,I167516,I167504,I101066,I167519,I101092,I101100,I167522,I101126,I101134,I101151,I101168,I101185,I167510,I101225,I101233,I101250,I101267,I101284,I101315,I167507,I167513,I101332,I167528,I101358,I101366,I101397,I101428,I101445,I101476,I167525,I101576,I150114,I101602,I101610,I101627,I150096,I150108,I101644,I150111,I101670,I101678,I150105,I150102,I101704,I101712,I101729,I101746,I101763,I150120,I101803,I101811,I101828,I101845,I101862,I101893,I150099,I101910,I101936,I101944,I101975,I102006,I102023,I102054,I150117,I102154,I150692,I102180,I102188,I102205,I150674,I150686,I102222,I150689,I102248,I102256,I150683,I150680,I102282,I102290,I102307,I102324,I102341,I102137,I150698,I102381,I102389,I102406,I102423,I102440,I102140,I102471,I150677,I102488,I102514,I102522,I102122,I102553,I102131,I102584,I102601,I102143,I102632,I150695,I102134,I102125,I102128,I102146,I102732,I102758,I102766,I102783,I102800,I102826,I102834,I102860,I102868,I102885,I102902,I102919,I102959,I102967,I102984,I103001,I103018,I103049,I103066,I103092,I103100,I103131,I103162,I103179,I103210,I103310,I103336,I103344,I103361,I103378,I103404,I103412,I103438,I103446,I103463,I103480,I103497,I103537,I103545,I103562,I103579,I103596,I103627,I103644,I103670,I103678,I103709,I103740,I103757,I103788,I103888,I172291,I103914,I103922,I103939,I172276,I172264,I103956,I172279,I103982,I103990,I172282,I104016,I104024,I104041,I104058,I104075,I103871,I172270,I104115,I104123,I104140,I104157,I104174,I103874,I104205,I172267,I172273,I104222,I172288,I104248,I104256,I103856,I104287,I103865,I104318,I104335,I103877,I104366,I172285,I103868,I103859,I103862,I103880,I104463,I104489,I104497,I104514,I104531,I104557,I104588,I104596,I104613,I104639,I104647,I104687,I104723,I104740,I104766,I104774,I104791,I104822,I104839,I104856,I104887,I104918,I104935,I104990,I171089,I105016,I105024,I105041,I171086,I171095,I105058,I171074,I105084,I171077,I105115,I105123,I171092,I105140,I105166,I105174,I171098,I105214,I105250,I171080,I171101,I105267,I171083,I105293,I105301,I105318,I105349,I105366,I105383,I105414,I105445,I105462,I105517,I105543,I105551,I105568,I105585,I105611,I105642,I105650,I105667,I105693,I105701,I105741,I105777,I105794,I105820,I105828,I105845,I105876,I105893,I105910,I105941,I105972,I105989,I106044,I169304,I106070,I106078,I106095,I169301,I169310,I106112,I169289,I106138,I169292,I106169,I106177,I169307,I106194,I106220,I106228,I169313,I106268,I106304,I169295,I169316,I106321,I169298,I106347,I106355,I106372,I106403,I106420,I106437,I106468,I106499,I106516,I106571,I168709,I106597,I106605,I106622,I168706,I168715,I106639,I168694,I106665,I168697,I106696,I106704,I168712,I106721,I106747,I106755,I168718,I106795,I106831,I168700,I168721,I106848,I168703,I106874,I106882,I106899,I106930,I106947,I106964,I106995,I107026,I107043,I107098,I143756,I107124,I107132,I107149,I143738,I107166,I143744,I107192,I143741,I107223,I107231,I143750,I107248,I107274,I107282,I143762,I107322,I107358,I143753,I143747,I107375,I107401,I107409,I107426,I107457,I143759,I107474,I107491,I107522,I107553,I107570,I107625,I107651,I107659,I107676,I107693,I107719,I107614,I107750,I107758,I107775,I107801,I107809,I107617,I107849,I107608,I107599,I107885,I107902,I107928,I107936,I107953,I107602,I107984,I108001,I108018,I107611,I108049,I107596,I108080,I108097,I107605,I108152,I108178,I108186,I108203,I108220,I108246,I108141,I108277,I108285,I108302,I108328,I108336,I108144,I108376,I108135,I108126,I108412,I108429,I108455,I108463,I108480,I108129,I108511,I108528,I108545,I108138,I108576,I108123,I108607,I108624,I108132,I108679,I108705,I108713,I108730,I108747,I108773,I108804,I108812,I108829,I108855,I108863,I108903,I108939,I108956,I108982,I108990,I109007,I109038,I109055,I109072,I109103,I109134,I109151,I109206,I109232,I109240,I109257,I109274,I109300,I109195,I109331,I109339,I109356,I109382,I109390,I109198,I109430,I109189,I109180,I109466,I109483,I109509,I109517,I109534,I109183,I109565,I109582,I109599,I109192,I109630,I109177,I109661,I109678,I109186,I109733,I109759,I109767,I109784,I109801,I109827,I109858,I109866,I109883,I109909,I109917,I109957,I109993,I110010,I110036,I110044,I110061,I110092,I110109,I110126,I110157,I110188,I110205,I110260,I172874,I110286,I110294,I110311,I172871,I172880,I110328,I172859,I110354,I172862,I110385,I110393,I172877,I110410,I110436,I110444,I172883,I110484,I110520,I172865,I172886,I110537,I172868,I110563,I110571,I110588,I110619,I110636,I110653,I110684,I110715,I110732,I110787,I169899,I110813,I110821,I110838,I169896,I169905,I110855,I169884,I110881,I110776,I169887,I110912,I110920,I169902,I110937,I110963,I110971,I110779,I169908,I111011,I110770,I110761,I111047,I169890,I169911,I111064,I169893,I111090,I111098,I111115,I110764,I111146,I111163,I111180,I110773,I111211,I110758,I111242,I111259,I110767,I111314,I111340,I111348,I111365,I111382,I111408,I111439,I111447,I111464,I111490,I111498,I111538,I111574,I111591,I111617,I111625,I111642,I111673,I111690,I111707,I111738,I111769,I111786,I111841,I111867,I111875,I111892,I111909,I111935,I111830,I111966,I111974,I111991,I112017,I112025,I111833,I112065,I111824,I111815,I112101,I112118,I112144,I112152,I112169,I111818,I112200,I112217,I112234,I111827,I112265,I111812,I112296,I112313,I111821,I112368,I137398,I112394,I112402,I112419,I137380,I112436,I137386,I112462,I112357,I137383,I112493,I112501,I137392,I112518,I112544,I112552,I112360,I137404,I112592,I112351,I112342,I112628,I137395,I137389,I112645,I112671,I112679,I112696,I112345,I112727,I137401,I112744,I112761,I112354,I112792,I112339,I112823,I112840,I112348,I112895,I146646,I112921,I112929,I112946,I146628,I112963,I146634,I112989,I146631,I113020,I113028,I146640,I113045,I113071,I113079,I146652,I113119,I113155,I146643,I146637,I113172,I113198,I113206,I113223,I113254,I146649,I113271,I113288,I113319,I113350,I113367,I113422,I160070,I113448,I113456,I113473,I160076,I160058,I113490,I160067,I113516,I113411,I160073,I113547,I113555,I160061,I113572,I113598,I113606,I113414,I160079,I113646,I113405,I113396,I113682,I160064,I113699,I160082,I113725,I113733,I113750,I113399,I113781,I113798,I113815,I113408,I113846,I113393,I113877,I113894,I113402,I113955,I113981,I113998,I114006,I114023,I114040,I114057,I114074,I114091,I114122,I114139,I114170,I114187,I114204,I114235,I114275,I114283,I114300,I114317,I114334,I114365,I114382,I114399,I114425,I114447,I114464,I114495,I114540,I114601,I114627,I114644,I114652,I114669,I114686,I114703,I114720,I114737,I114587,I114768,I114785,I114590,I114816,I114833,I114850,I114566,I114881,I114578,I114921,I114929,I114946,I114963,I114980,I114593,I115011,I115028,I115045,I115071,I114581,I115093,I115110,I114575,I115141,I114569,I114572,I115186,I114584,I115247,I115273,I115290,I115298,I115315,I115332,I115349,I115366,I115383,I115414,I115431,I115462,I115479,I115496,I115527,I115567,I115575,I115592,I115609,I115626,I115657,I115674,I115691,I115717,I115739,I115756,I115787,I115832,I115893,I115919,I115936,I115944,I115961,I115978,I115995,I116012,I116029,I116060,I116077,I116108,I116125,I116142,I116173,I116213,I116221,I116238,I116255,I116272,I116303,I116320,I116337,I116363,I116385,I116402,I116433,I116478,I116539,I116565,I116582,I116590,I116607,I116624,I116641,I116658,I116675,I116706,I116723,I116754,I116771,I116788,I116819,I116859,I116867,I116884,I116901,I116918,I116949,I116966,I116983,I117009,I117031,I117048,I117079,I117124,I117185,I117211,I117228,I117236,I117253,I117270,I117287,I117304,I117321,I117352,I117369,I117400,I117417,I117434,I117465,I117505,I117513,I117530,I117547,I117564,I117595,I117612,I117629,I117655,I117677,I117694,I117725,I117770,I117831,I157356,I117857,I157362,I117874,I117882,I117899,I157359,I117916,I157338,I117933,I157341,I117950,I157347,I117967,I117817,I117998,I118015,I117820,I118046,I118063,I118080,I117796,I118111,I117808,I118151,I118159,I118176,I118193,I157350,I118210,I117823,I118241,I118258,I157344,I118275,I157353,I118301,I117811,I118323,I118340,I117805,I118371,I117799,I117802,I118416,I117814,I118477,I118503,I118520,I118528,I118545,I118562,I118579,I118596,I118613,I118644,I118661,I118692,I118709,I118726,I118757,I118797,I118805,I118822,I118839,I118856,I118887,I118904,I118921,I118947,I118969,I118986,I119017,I119062,I119123,I119149,I119166,I119174,I119191,I119208,I119225,I119242,I119259,I119290,I119307,I119338,I119355,I119372,I119403,I119443,I119451,I119468,I119485,I119502,I119533,I119550,I119567,I119593,I119615,I119632,I119663,I119708,I119769,I119795,I119812,I119820,I119837,I119854,I119871,I119888,I119905,I119936,I119953,I119984,I120001,I120018,I120049,I120089,I120097,I120114,I120131,I120148,I120179,I120196,I120213,I120239,I120261,I120278,I120309,I120354,I120415,I176429,I120441,I176453,I120458,I120466,I120483,I176435,I120500,I176444,I120517,I120534,I176450,I120551,I120401,I120582,I120599,I120404,I120630,I120647,I176447,I120664,I120380,I120695,I120392,I120735,I120743,I120760,I120777,I176441,I120794,I120407,I120825,I176432,I120842,I176456,I120859,I176438,I120885,I120395,I120907,I120924,I120389,I120955,I120383,I120386,I121000,I120398,I121061,I121087,I121104,I121112,I121129,I121146,I121163,I121180,I121197,I121047,I121228,I121245,I121050,I121276,I121293,I121310,I121026,I121341,I121038,I121381,I121389,I121406,I121423,I121440,I121053,I121471,I121488,I121505,I121531,I121041,I121553,I121570,I121035,I121601,I121029,I121032,I121646,I121044,I121707,I121733,I121750,I121758,I121775,I121792,I121809,I121826,I121843,I121874,I121891,I121922,I121939,I121956,I121987,I122027,I122035,I122052,I122069,I122086,I122117,I122134,I122151,I122177,I122199,I122216,I122247,I122292,I122353,I122379,I122396,I122404,I122421,I122438,I122455,I122472,I122489,I122520,I122537,I122568,I122585,I122602,I122633,I122673,I122681,I122698,I122715,I122732,I122763,I122780,I122797,I122823,I122845,I122862,I122893,I122938,I122999,I123025,I123042,I123050,I123067,I123084,I123101,I123118,I123135,I123166,I123183,I123214,I123231,I123248,I123279,I123319,I123327,I123344,I123361,I123378,I123409,I123426,I123443,I123469,I123491,I123508,I123539,I123584,I123645,I123671,I123688,I123696,I123713,I123730,I123747,I123764,I123781,I123631,I123812,I123829,I123634,I123860,I123877,I123894,I123610,I123925,I123622,I123965,I123973,I123990,I124007,I124024,I123637,I124055,I124072,I124089,I124115,I123625,I124137,I124154,I123619,I124185,I123613,I123616,I124230,I123628,I124291,I141444,I124317,I141426,I124334,I124342,I124359,I141435,I124376,I141447,I124393,I141429,I124410,I141438,I124427,I124458,I124475,I124506,I124523,I141450,I124540,I124571,I124611,I124619,I124636,I124653,I124670,I124701,I141432,I124718,I141441,I124735,I124761,I124783,I124800,I124831,I124876,I124937,I124963,I124980,I124988,I125005,I125022,I125039,I125056,I125073,I125104,I125121,I125152,I125169,I125186,I125217,I125257,I125265,I125282,I125299,I125316,I125347,I125364,I125381,I125407,I125429,I125446,I125477,I125522,I125583,I125609,I125626,I125634,I125651,I125668,I125685,I125702,I125719,I125750,I125767,I125798,I125815,I125832,I125863,I125903,I125911,I125928,I125945,I125962,I125993,I126010,I126027,I126053,I126075,I126092,I126123,I126168,I126229,I126255,I126272,I126280,I126297,I126314,I126331,I126348,I126365,I126396,I126413,I126444,I126461,I126478,I126509,I126549,I126557,I126574,I126591,I126608,I126639,I126656,I126673,I126699,I126721,I126738,I126769,I126814,I126875,I126901,I126918,I126926,I126943,I126960,I126977,I126994,I127011,I126861,I127042,I127059,I126864,I127090,I127107,I127124,I126840,I127155,I126852,I127195,I127203,I127220,I127237,I127254,I126867,I127285,I127302,I127319,I127345,I126855,I127367,I127384,I126849,I127415,I126843,I126846,I127460,I126858,I127521,I134558,I127547,I134561,I127564,I127572,I127589,I127606,I134570,I127623,I134579,I127640,I134567,I127657,I127688,I127705,I127736,I127753,I134573,I127770,I127801,I127841,I127849,I127866,I127883,I134564,I127900,I127931,I134576,I127948,I127965,I127991,I128013,I128030,I128061,I128106,I128167,I128193,I128210,I128218,I128235,I128252,I128269,I128286,I128303,I128334,I128351,I128382,I128399,I128416,I128447,I128487,I128495,I128512,I128529,I128546,I128577,I128594,I128611,I128637,I128659,I128676,I128707,I128752,I128813,I128839,I128856,I128864,I128881,I128898,I128915,I128932,I128949,I128980,I128997,I129028,I129045,I129062,I129093,I129133,I129141,I129158,I129175,I129192,I129223,I129240,I129257,I129283,I129305,I129322,I129353,I129398,I129459,I136820,I129485,I136802,I129502,I129510,I129527,I136811,I129544,I136823,I129561,I136805,I129578,I136814,I129595,I129626,I129643,I129674,I129691,I136826,I129708,I129739,I129779,I129787,I129804,I129821,I129838,I129869,I136808,I129886,I136817,I129903,I129929,I129951,I129968,I129999,I130044,I130099,I130125,I130142,I130091,I130164,I130190,I130198,I130215,I130232,I130249,I130266,I130283,I130300,I130073,I130331,I130076,I130362,I130379,I130396,I130413,I130085,I130444,I130088,I130082,I130489,I130506,I130523,I130549,I130557,I130070,I130588,I130605,I130079,I130660,I152992,I130686,I130703,I130725,I152998,I130751,I130759,I153007,I130776,I130793,I152986,I130810,I152989,I130827,I130844,I153001,I130861,I130892,I130923,I152995,I130940,I130957,I130974,I131005,I131050,I153010,I131067,I131084,I153004,I131110,I131118,I131149,I131166,I131221,I153536,I131247,I131264,I131213,I131286,I153542,I131312,I131320,I153551,I131337,I131354,I153530,I131371,I153533,I131388,I131405,I153545,I131422,I131195,I131453,I131198,I131484,I153539,I131501,I131518,I131535,I131207,I131566,I131210,I131204,I131611,I153554,I131628,I131645,I153548,I131671,I131679,I131192,I131710,I131727,I131201,I131782,I131808,I131825,I131847,I131873,I131881,I131898,I131915,I131932,I131949,I131966,I131983,I132014,I132045,I132062,I132079,I132096,I132127,I132172,I132189,I132206,I132232,I132240,I132271,I132288,I132343,I132369,I132386,I132408,I132434,I132442,I132459,I132476,I132493,I132510,I132527,I132544,I132575,I132606,I132623,I132640,I132657,I132688,I132733,I132750,I132767,I132793,I132801,I132832,I132849,I132904,I132930,I132947,I132969,I132995,I133003,I133020,I133037,I133054,I133071,I133088,I133105,I133136,I133167,I133184,I133201,I133218,I133249,I133294,I133311,I133328,I133354,I133362,I133393,I133410,I133465,I133491,I133508,I133530,I133556,I133564,I133581,I133598,I133615,I133632,I133649,I133666,I133697,I133728,I133745,I133762,I133779,I133810,I133855,I133872,I133889,I133915,I133923,I133954,I133971,I134026,I142019,I134052,I134069,I134018,I134091,I142010,I134117,I134125,I142007,I134142,I134159,I142016,I134176,I142025,I134193,I134210,I142004,I134227,I134000,I134258,I134003,I134289,I142013,I134306,I134323,I134340,I134012,I134371,I134015,I134009,I134416,I142028,I134433,I134450,I142022,I134476,I134484,I133997,I134515,I134532,I134006,I134587,I165229,I134613,I134630,I134652,I165226,I134678,I134686,I165232,I134703,I134720,I165241,I134737,I165235,I134754,I134771,I165247,I134788,I134819,I134850,I165244,I134867,I134884,I134901,I134932,I134977,I165238,I134994,I165250,I135011,I135037,I135045,I135076,I135093,I135148,I135174,I135191,I135213,I135239,I135247,I135264,I135281,I135298,I135315,I135332,I135349,I135380,I135411,I135428,I135445,I135462,I135493,I135538,I135555,I135572,I135598,I135606,I135637,I135654,I135709,I166964,I135735,I135752,I135774,I166949,I135800,I135808,I166958,I135825,I135842,I166952,I135859,I166970,I166967,I135876,I135893,I166943,I135910,I135941,I135972,I166946,I135989,I136006,I136023,I136054,I136099,I136116,I166961,I136133,I166955,I136159,I136167,I136198,I136215,I136270,I136296,I136313,I136335,I136361,I136369,I136386,I136403,I136420,I136437,I136454,I136471,I136502,I136533,I136550,I136567,I136584,I136615,I136660,I136677,I136694,I136720,I136728,I136759,I136776,I136834,I136860,I136868,I136908,I136916,I136933,I136950,I136990,I137012,I137029,I137055,I137063,I137080,I137097,I137114,I137131,I137176,I137207,I137224,I137250,I137258,I137289,I137306,I137323,I137340,I137412,I137438,I137446,I137486,I137494,I137511,I137528,I137568,I137590,I137607,I137633,I137641,I137658,I137675,I137692,I137709,I137754,I137785,I137802,I137828,I137836,I137867,I137884,I137901,I137918,I137990,I138016,I138024,I138064,I138072,I138089,I138106,I138146,I138168,I138185,I138211,I138219,I138236,I138253,I138270,I138287,I138332,I138363,I138380,I138406,I138414,I138445,I138462,I138479,I138496,I138568,I138594,I138602,I138642,I138650,I138667,I138684,I138724,I138746,I138763,I138789,I138797,I138814,I138831,I138848,I138865,I138910,I138941,I138958,I138984,I138992,I139023,I139040,I139057,I139074,I139146,I139172,I139180,I139129,I139220,I139228,I139245,I139262,I139117,I139302,I139138,I139324,I139341,I139367,I139375,I139392,I139409,I139426,I139443,I139114,I139135,I139488,I139126,I139519,I139536,I139562,I139570,I139132,I139601,I139618,I139635,I139652,I139123,I139120,I139724,I139750,I139758,I139707,I139798,I139806,I139823,I139840,I139695,I139880,I139716,I139902,I139919,I139945,I139953,I139970,I139987,I140004,I140021,I139692,I139713,I140066,I139704,I140097,I140114,I140140,I140148,I139710,I140179,I140196,I140213,I140230,I139701,I139698,I140302,I140328,I140336,I140376,I140384,I140401,I140418,I140458,I140480,I140497,I140523,I140531,I140548,I140565,I140582,I140599,I140644,I140675,I140692,I140718,I140726,I140757,I140774,I140791,I140808,I140880,I140906,I140914,I140954,I140962,I140979,I140996,I141036,I141058,I141075,I141101,I141109,I141126,I141143,I141160,I141177,I141222,I141253,I141270,I141296,I141304,I141335,I141352,I141369,I141386,I141458,I141484,I141492,I141532,I141540,I141557,I141574,I141614,I141636,I141653,I141679,I141687,I141704,I141721,I141738,I141755,I141800,I141831,I141848,I141874,I141882,I141913,I141930,I141947,I141964,I142036,I142062,I142070,I142110,I142118,I142135,I142152,I142192,I142214,I142231,I142257,I142265,I142282,I142299,I142316,I142333,I142378,I142409,I142426,I142452,I142460,I142491,I142508,I142525,I142542,I142614,I142640,I142648,I142688,I142696,I142713,I142730,I142770,I142792,I142809,I142835,I142843,I142860,I142877,I142894,I142911,I142956,I142987,I143004,I143030,I143038,I143069,I143086,I143103,I143120,I143192,I143218,I143226,I143266,I143274,I143291,I143308,I143348,I143370,I143387,I143413,I143421,I143438,I143455,I143472,I143489,I143534,I143565,I143582,I143608,I143616,I143647,I143664,I143681,I143698,I143770,I143796,I143804,I143844,I143852,I143869,I143886,I143926,I143948,I143965,I143991,I143999,I144016,I144033,I144050,I144067,I144112,I144143,I144160,I144186,I144194,I144225,I144242,I144259,I144276,I144348,I144374,I144382,I144422,I144430,I144447,I144464,I144504,I144526,I144543,I144569,I144577,I144594,I144611,I144628,I144645,I144690,I144721,I144738,I144764,I144772,I144803,I144820,I144837,I144854,I144926,I144952,I144960,I145000,I145008,I145025,I145042,I145082,I145104,I145121,I145147,I145155,I145172,I145189,I145206,I145223,I145268,I145299,I145316,I145342,I145350,I145381,I145398,I145415,I145432,I145504,I145530,I145538,I145578,I145586,I145603,I145620,I145660,I145682,I145699,I145725,I145733,I145750,I145767,I145784,I145801,I145846,I145877,I145894,I145920,I145928,I145959,I145976,I145993,I146010,I146082,I146108,I146116,I146156,I146164,I146181,I146198,I146238,I146260,I146277,I146303,I146311,I146328,I146345,I146362,I146379,I146424,I146455,I146472,I146498,I146506,I146537,I146554,I146571,I146588,I146660,I146686,I146694,I146734,I146742,I146759,I146776,I146816,I146838,I146855,I146881,I146889,I146906,I146923,I146940,I146957,I147002,I147033,I147050,I147076,I147084,I147115,I147132,I147149,I147166,I147238,I147264,I147272,I147312,I147320,I147337,I147354,I147394,I147416,I147433,I147459,I147467,I147484,I147501,I147518,I147535,I147580,I147611,I147628,I147654,I147662,I147693,I147710,I147727,I147744,I147816,I147842,I147850,I147890,I147898,I147915,I147932,I147972,I147994,I148011,I148037,I148045,I148062,I148079,I148096,I148113,I148158,I148189,I148206,I148232,I148240,I148271,I148288,I148305,I148322,I148394,I148420,I148428,I148377,I148468,I148476,I148493,I148510,I148365,I148550,I148386,I148572,I148589,I148615,I148623,I148640,I148657,I148674,I148691,I148362,I148383,I148736,I148374,I148767,I148784,I148810,I148818,I148380,I148849,I148866,I148883,I148900,I148371,I148368,I148972,I148998,I149006,I149046,I149054,I149071,I149088,I149128,I149150,I149167,I149193,I149201,I149218,I149235,I149252,I149269,I149314,I149345,I149362,I149388,I149396,I149427,I149444,I149461,I149478,I149550,I149576,I149584,I149624,I149632,I149649,I149666,I149706,I149728,I149745,I149771,I149779,I149796,I149813,I149830,I149847,I149892,I149923,I149940,I149966,I149974,I150005,I150022,I150039,I150056,I150128,I150154,I150162,I150202,I150210,I150227,I150244,I150284,I150306,I150323,I150349,I150357,I150374,I150391,I150408,I150425,I150470,I150501,I150518,I150544,I150552,I150583,I150600,I150617,I150634,I150706,I170506,I150732,I150740,I170488,I170479,I150780,I150788,I170494,I150805,I170482,I150822,I150862,I150884,I170491,I150901,I150927,I150935,I150952,I170500,I150969,I150986,I151003,I151048,I170503,I151079,I151096,I170497,I170485,I151122,I151130,I151161,I151178,I151195,I151212,I151284,I151310,I151318,I151267,I151358,I151366,I151383,I151400,I151255,I151440,I151276,I151462,I151479,I151505,I151513,I151530,I151547,I151564,I151581,I151252,I151273,I151626,I151264,I151657,I151674,I151700,I151708,I151270,I151739,I151756,I151773,I151790,I151261,I151258,I151862,I151888,I151896,I151936,I151944,I151961,I151978,I152018,I152040,I152057,I152083,I152091,I152108,I152125,I152142,I152159,I152204,I152235,I152252,I152278,I152286,I152317,I152334,I152351,I152368,I152440,I158447,I152466,I152474,I158441,I158426,I152514,I152522,I158432,I152539,I158444,I152556,I152596,I152618,I152635,I152661,I152669,I152686,I158450,I152703,I158438,I152720,I152737,I152782,I158429,I152813,I152830,I158435,I152856,I152864,I152895,I152912,I152929,I152946,I153018,I153044,I153052,I153078,I153095,I153117,I153134,I153151,I153168,I153185,I153216,I153233,I153250,I153267,I153312,I153329,I153346,I153405,I153431,I153439,I153456,I153473,I153504,I153562,I153588,I153596,I153622,I153639,I153661,I153678,I153695,I153712,I153729,I153760,I153777,I153794,I153811,I153856,I153873,I153890,I153949,I153975,I153983,I154000,I154017,I154048,I154106,I154132,I154140,I154166,I154183,I154205,I154222,I154239,I154256,I154273,I154304,I154321,I154338,I154355,I154400,I154417,I154434,I154493,I154519,I154527,I154544,I154561,I154592,I154650,I154676,I154684,I154710,I154727,I154642,I154749,I154766,I154783,I154800,I154817,I154621,I154848,I154865,I154882,I154899,I154624,I154639,I154944,I154961,I154978,I154636,I154633,I154630,I155037,I155063,I155071,I155088,I155105,I154618,I155136,I154627,I155194,I178241,I155220,I155228,I178226,I178220,I155254,I155271,I155186,I155293,I178214,I155310,I178235,I155327,I178223,I155344,I155361,I155165,I155392,I178232,I155409,I178238,I155426,I178229,I155443,I155168,I155183,I155488,I178217,I155505,I155522,I155180,I155177,I155174,I155581,I155607,I155615,I155632,I155649,I155162,I155680,I155171,I155738,I155764,I155772,I155798,I155815,I155837,I155854,I155871,I155888,I155905,I155936,I155953,I155970,I155987,I156032,I156049,I156066,I156125,I156151,I156159,I156176,I156193,I156224,I156282,I156308,I156316,I156342,I156359,I156274,I156381,I156398,I156415,I156432,I156449,I156253,I156480,I156497,I156514,I156531,I156256,I156271,I156576,I156593,I156610,I156268,I156265,I156262,I156669,I156695,I156703,I156720,I156737,I156250,I156768,I156259,I156826,I156852,I156860,I156886,I156903,I156925,I156942,I156959,I156976,I156993,I157024,I157041,I157058,I157075,I157120,I157137,I157154,I157213,I157239,I157247,I157264,I157281,I157312,I157370,I157396,I157404,I157430,I157447,I157469,I157486,I157503,I157520,I157537,I157568,I157585,I157602,I157619,I157664,I157681,I157698,I157757,I157783,I157791,I157808,I157825,I157856,I157914,I157940,I157948,I157974,I157991,I157906,I158013,I158030,I158047,I158064,I158081,I157885,I158112,I158129,I158146,I158163,I157888,I157903,I158208,I158225,I158242,I157900,I157897,I157894,I158301,I158327,I158335,I158352,I158369,I157882,I158400,I157891,I158458,I158484,I158492,I158518,I158535,I158557,I158574,I158591,I158608,I158625,I158656,I158673,I158690,I158707,I158752,I158769,I158786,I158845,I158871,I158879,I158896,I158913,I158944,I159002,I159028,I159036,I159062,I159079,I159101,I159118,I159135,I159152,I159169,I159200,I159217,I159234,I159251,I159296,I159313,I159330,I159389,I159415,I159423,I159440,I159457,I159488,I159546,I159572,I159580,I159606,I159623,I159645,I159662,I159679,I159696,I159713,I159744,I159761,I159778,I159795,I159840,I159857,I159874,I159933,I159959,I159967,I159984,I160001,I160032,I160090,I174076,I160116,I160124,I174061,I174055,I160150,I160167,I160189,I174049,I160206,I174070,I160223,I174058,I160240,I160257,I160288,I174067,I160305,I174073,I160322,I174064,I160339,I160384,I174052,I160401,I160418,I160477,I160503,I160511,I160528,I160545,I160576,I160634,I160660,I160668,I160685,I160711,I160719,I160736,I160753,I160770,I160787,I160818,I160835,I160852,I160883,I160900,I160940,I160948,I160979,I160996,I161013,I161030,I161061,I161092,I161118,I161140,I161212,I161238,I161246,I161263,I161289,I161297,I161314,I161331,I161348,I161365,I161396,I161413,I161430,I161461,I161478,I161518,I161526,I161557,I161574,I161591,I161608,I161639,I161670,I161696,I161718,I161790,I161816,I161824,I161841,I161867,I161875,I161892,I161909,I161926,I161943,I161974,I161991,I162008,I162039,I162056,I162096,I162104,I162135,I162152,I162169,I162186,I162217,I162248,I162274,I162296,I162368,I162394,I162402,I162419,I162445,I162453,I162470,I162487,I162504,I162521,I162552,I162569,I162586,I162617,I162634,I162674,I162682,I162713,I162730,I162747,I162764,I162795,I162826,I162852,I162874,I162946,I162972,I162980,I162997,I163023,I163031,I163048,I163065,I163082,I163099,I163130,I163147,I163164,I163195,I163212,I163252,I163260,I163291,I163308,I163325,I163342,I163373,I163404,I163430,I163452,I163524,I163550,I163558,I163575,I163601,I163609,I163626,I163643,I163660,I163677,I163708,I163725,I163742,I163773,I163790,I163830,I163838,I163869,I163886,I163903,I163920,I163951,I163982,I164008,I164030,I164102,I164128,I164136,I164153,I164179,I164187,I164204,I164221,I164238,I164255,I164286,I164303,I164320,I164351,I164368,I164408,I164416,I164447,I164464,I164481,I164498,I164529,I164560,I164586,I164608,I164680,I164706,I164714,I164731,I164757,I164765,I164782,I164799,I164816,I164833,I164864,I164881,I164898,I164929,I164946,I164986,I164994,I165025,I165042,I165059,I165076,I165107,I165138,I165164,I165186,I165258,I165284,I165292,I165309,I165335,I165343,I165360,I165377,I165394,I165411,I165442,I165459,I165476,I165507,I165524,I165564,I165572,I165603,I165620,I165637,I165654,I165685,I165716,I165742,I165764,I165836,I165862,I165870,I165887,I165913,I165921,I165938,I165955,I165972,I165989,I166020,I166037,I166054,I166085,I166102,I166142,I166150,I166181,I166198,I166215,I166232,I166263,I166294,I166320,I166342,I166417,I166443,I166451,I166468,I166494,I166502,I166519,I166536,I166567,I166598,I166615,I166632,I166649,I166666,I166697,I166756,I166773,I166799,I166821,I166847,I166855,I166872,I166903,I166978,I167004,I167012,I167029,I167055,I167063,I167080,I167097,I167128,I167159,I167176,I167193,I167210,I167227,I167258,I167317,I167334,I167360,I167382,I167408,I167416,I167433,I167464,I167539,I167565,I167582,I167590,I167635,I167652,I167669,I167686,I167703,I167720,I167737,I167768,I167785,I167830,I167847,I167864,I167895,I167921,I167929,I167960,I167977,I167994,I168020,I168028,I168045,I168134,I168160,I168177,I168185,I168230,I168247,I168264,I168281,I168298,I168315,I168332,I168363,I168380,I168425,I168442,I168459,I168490,I168516,I168524,I168555,I168572,I168589,I168615,I168623,I168640,I168729,I168755,I168772,I168780,I168825,I168842,I168859,I168876,I168893,I168910,I168927,I168958,I168975,I169020,I169037,I169054,I169085,I169111,I169119,I169150,I169167,I169184,I169210,I169218,I169235,I169324,I169350,I169367,I169375,I169420,I169437,I169454,I169471,I169488,I169505,I169522,I169553,I169570,I169615,I169632,I169649,I169680,I169706,I169714,I169745,I169762,I169779,I169805,I169813,I169830,I169919,I169945,I169962,I169970,I170015,I170032,I170049,I170066,I170083,I170100,I170117,I170148,I170165,I170210,I170227,I170244,I170275,I170301,I170309,I170340,I170357,I170374,I170400,I170408,I170425,I170514,I170540,I170557,I170565,I170610,I170627,I170644,I170661,I170678,I170695,I170712,I170743,I170760,I170805,I170822,I170839,I170870,I170896,I170904,I170935,I170952,I170969,I170995,I171003,I171020,I171109,I171135,I171152,I171160,I171205,I171222,I171239,I171256,I171273,I171290,I171307,I171338,I171355,I171400,I171417,I171434,I171465,I171491,I171499,I171530,I171547,I171564,I171590,I171598,I171615,I171704,I171730,I171747,I171755,I171800,I171817,I171834,I171851,I171868,I171885,I171902,I171933,I171950,I171995,I172012,I172029,I172060,I172086,I172094,I172125,I172142,I172159,I172185,I172193,I172210,I172299,I172325,I172342,I172350,I172395,I172412,I172429,I172446,I172463,I172480,I172497,I172528,I172545,I172590,I172607,I172624,I172655,I172681,I172689,I172720,I172737,I172754,I172780,I172788,I172805,I172894,I172920,I172937,I172945,I172990,I173007,I173024,I173041,I173058,I173075,I173092,I173123,I173140,I173185,I173202,I173219,I173250,I173276,I173284,I173315,I173332,I173349,I173375,I173383,I173400,I173489,I173515,I173532,I173540,I173585,I173602,I173619,I173636,I173653,I173670,I173687,I173718,I173735,I173780,I173797,I173814,I173845,I173871,I173879,I173910,I173927,I173944,I173970,I173978,I173995,I174084,I174110,I174127,I174135,I174180,I174197,I174214,I174231,I174248,I174265,I174282,I174313,I174330,I174375,I174392,I174409,I174440,I174466,I174474,I174505,I174522,I174539,I174565,I174573,I174590,I174679,I174705,I174722,I174730,I174775,I174792,I174809,I174826,I174843,I174860,I174877,I174908,I174925,I174970,I174987,I175004,I175035,I175061,I175069,I175100,I175117,I175134,I175160,I175168,I175185,I175274,I175300,I175317,I175325,I175370,I175387,I175404,I175421,I175438,I175455,I175472,I175503,I175520,I175565,I175582,I175599,I175630,I175656,I175664,I175695,I175712,I175729,I175755,I175763,I175780,I175869,I175895,I175912,I175920,I175965,I175982,I175999,I176016,I176033,I176050,I176067,I176098,I176115,I176160,I176177,I176194,I176225,I176251,I176259,I176290,I176307,I176324,I176350,I176358,I176375,I176464,I176490,I176507,I176515,I176560,I176577,I176594,I176611,I176628,I176645,I176662,I176693,I176710,I176755,I176772,I176789,I176820,I176846,I176854,I176885,I176902,I176919,I176945,I176953,I176970,I177059,I177085,I177102,I177110,I177155,I177172,I177189,I177206,I177223,I177240,I177257,I177288,I177305,I177350,I177367,I177384,I177415,I177441,I177449,I177480,I177497,I177514,I177540,I177548,I177565,I177654,I177680,I177697,I177705,I177750,I177767,I177784,I177801,I177818,I177835,I177852,I177883,I177900,I177945,I177962,I177979,I178010,I178036,I178044,I178075,I178092,I178109,I178135,I178143,I178160,I178249,I178275,I178292,I178300,I178345,I178362,I178379,I178396,I178413,I178430,I178447,I178478,I178495,I178540,I178557,I178574,I178605,I178631,I178639,I178670,I178687,I178704,I178730,I178738,I178755,I178844,I178870,I178887,I178895,I178940,I178957,I178974,I178991,I179008,I179025,I179042,I179073,I179090,I179135,I179152,I179169,I179200,I179226,I179234,I179265,I179282,I179299,I179325,I179333,I179350;
not I_0 (I2106,I2074);
DFFARX1 I_1 (I33411,I2067,I2106,I2132,);
nand I_2 (I2140,I2132,I33411);
not I_3 (I2157,I2140);
DFFARX1 I_4 (I2157,I2067,I2106,I2098,);
DFFARX1 I_5 (I33417,I2067,I2106,I2197,);
not I_6 (I2205,I2197);
not I_7 (I2222,I33426);
not I_8 (I2239,I33420);
nand I_9 (I2256,I2205,I2239);
nor I_10 (I2273,I2256,I33426);
DFFARX1 I_11 (I2273,I2067,I2106,I2077,);
nor I_12 (I2304,I33420,I33426);
nand I_13 (I2321,I2197,I2304);
nor I_14 (I2338,I33423,I33429);
nor I_15 (I2080,I2256,I33423);
not I_16 (I2369,I33423);
not I_17 (I2386,I33432);
nand I_18 (I2403,I2386,I33408);
nand I_19 (I2420,I2222,I2403);
not I_20 (I2437,I2420);
nor I_21 (I2454,I33432,I33429);
nor I_22 (I2089,I2437,I2454);
nor I_23 (I2485,I33414,I33432);
and I_24 (I2502,I2485,I2338);
nor I_25 (I2519,I2420,I2502);
DFFARX1 I_26 (I2519,I2067,I2106,I2095,);
nor I_27 (I2550,I2140,I2502);
DFFARX1 I_28 (I2550,I2067,I2106,I2092,);
nor I_29 (I2581,I33414,I33408);
DFFARX1 I_30 (I2581,I2067,I2106,I2607,);
nor I_31 (I2615,I2607,I33420);
nand I_32 (I2632,I2615,I2222);
nand I_33 (I2086,I2632,I2321);
nand I_34 (I2083,I2615,I2369);
not I_35 (I2701,I2074);
DFFARX1 I_36 (I14346,I2067,I2701,I2727,);
nand I_37 (I2735,I2727,I14337);
not I_38 (I2752,I2735);
DFFARX1 I_39 (I2752,I2067,I2701,I2693,);
DFFARX1 I_40 (I14358,I2067,I2701,I2792,);
not I_41 (I2800,I2792);
not I_42 (I2817,I14334);
not I_43 (I2834,I14334);
nand I_44 (I2851,I2800,I2834);
nor I_45 (I2868,I2851,I14334);
DFFARX1 I_46 (I2868,I2067,I2701,I2672,);
nor I_47 (I2899,I14334,I14334);
nand I_48 (I2916,I2792,I2899);
nor I_49 (I2933,I14343,I14337);
nor I_50 (I2675,I2851,I14343);
not I_51 (I2964,I14343);
not I_52 (I2981,I14355);
nand I_53 (I2998,I2981,I14352);
nand I_54 (I3015,I2817,I2998);
not I_55 (I3032,I3015);
nor I_56 (I3049,I14355,I14337);
nor I_57 (I2684,I3032,I3049);
nor I_58 (I3080,I14349,I14355);
and I_59 (I3097,I3080,I2933);
nor I_60 (I3114,I3015,I3097);
DFFARX1 I_61 (I3114,I2067,I2701,I2690,);
nor I_62 (I3145,I2735,I3097);
DFFARX1 I_63 (I3145,I2067,I2701,I2687,);
nor I_64 (I3176,I14349,I14340);
DFFARX1 I_65 (I3176,I2067,I2701,I3202,);
nor I_66 (I3210,I3202,I14334);
nand I_67 (I3227,I3210,I2817);
nand I_68 (I2681,I3227,I2916);
nand I_69 (I2678,I3210,I2964);
not I_70 (I3299,I2074);
DFFARX1 I_71 (I161195,I2067,I3299,I3325,);
DFFARX1 I_72 (I3325,I2067,I3299,I3342,);
not I_73 (I3350,I3342);
nand I_74 (I3367,I161198,I161192);
and I_75 (I3384,I3367,I161201);
DFFARX1 I_76 (I3384,I2067,I3299,I3410,);
DFFARX1 I_77 (I3410,I2067,I3299,I3291,);
DFFARX1 I_78 (I3410,I2067,I3299,I3282,);
DFFARX1 I_79 (I161189,I2067,I3299,I3455,);
nand I_80 (I3463,I3455,I161204);
not I_81 (I3480,I3463);
nor I_82 (I3279,I3325,I3480);
DFFARX1 I_83 (I161180,I2067,I3299,I3520,);
not I_84 (I3528,I3520);
nor I_85 (I3285,I3528,I3350);
nand I_86 (I3273,I3528,I3463);
nand I_87 (I3573,I161183,I161183);
and I_88 (I3590,I3573,I161180);
DFFARX1 I_89 (I3590,I2067,I3299,I3616,);
nor I_90 (I3624,I3616,I3325);
DFFARX1 I_91 (I3624,I2067,I3299,I3267,);
not I_92 (I3655,I3616);
nor I_93 (I3672,I161186,I161183);
not I_94 (I3689,I3672);
nor I_95 (I3706,I3463,I3689);
nor I_96 (I3723,I3655,I3706);
DFFARX1 I_97 (I3723,I2067,I3299,I3288,);
nor I_98 (I3754,I3616,I3689);
nor I_99 (I3276,I3480,I3754);
nor I_100 (I3270,I3616,I3672);
not I_101 (I3826,I2074);
DFFARX1 I_102 (I32819,I2067,I3826,I3852,);
DFFARX1 I_103 (I3852,I2067,I3826,I3869,);
not I_104 (I3877,I3869);
nand I_105 (I3894,I32837,I32822);
and I_106 (I3911,I3894,I32825);
DFFARX1 I_107 (I3911,I2067,I3826,I3937,);
DFFARX1 I_108 (I3937,I2067,I3826,I3818,);
DFFARX1 I_109 (I3937,I2067,I3826,I3809,);
DFFARX1 I_110 (I32813,I2067,I3826,I3982,);
nand I_111 (I3990,I3982,I32816);
not I_112 (I4007,I3990);
nor I_113 (I3806,I3852,I4007);
DFFARX1 I_114 (I32828,I2067,I3826,I4047,);
not I_115 (I4055,I4047);
nor I_116 (I3812,I4055,I3877);
nand I_117 (I3800,I4055,I3990);
nand I_118 (I4100,I32834,I32831);
and I_119 (I4117,I4100,I32816);
DFFARX1 I_120 (I4117,I2067,I3826,I4143,);
nor I_121 (I4151,I4143,I3852);
DFFARX1 I_122 (I4151,I2067,I3826,I3794,);
not I_123 (I4182,I4143);
nor I_124 (I4199,I32813,I32831);
not I_125 (I4216,I4199);
nor I_126 (I4233,I3990,I4216);
nor I_127 (I4250,I4182,I4233);
DFFARX1 I_128 (I4250,I2067,I3826,I3815,);
nor I_129 (I4281,I4143,I4216);
nor I_130 (I3803,I4007,I4281);
nor I_131 (I3797,I4143,I4199);
not I_132 (I4353,I2074);
DFFARX1 I_133 (I61305,I2067,I4353,I4379,);
DFFARX1 I_134 (I4379,I2067,I4353,I4396,);
not I_135 (I4404,I4396);
nand I_136 (I4421,I61305,I61308);
and I_137 (I4438,I4421,I61329);
DFFARX1 I_138 (I4438,I2067,I4353,I4464,);
DFFARX1 I_139 (I4464,I2067,I4353,I4345,);
DFFARX1 I_140 (I4464,I2067,I4353,I4336,);
DFFARX1 I_141 (I61317,I2067,I4353,I4509,);
nand I_142 (I4517,I4509,I61320);
not I_143 (I4534,I4517);
nor I_144 (I4333,I4379,I4534);
DFFARX1 I_145 (I61326,I2067,I4353,I4574,);
not I_146 (I4582,I4574);
nor I_147 (I4339,I4582,I4404);
nand I_148 (I4327,I4582,I4517);
nand I_149 (I4627,I61323,I61311);
and I_150 (I4644,I4627,I61314);
DFFARX1 I_151 (I4644,I2067,I4353,I4670,);
nor I_152 (I4678,I4670,I4379);
DFFARX1 I_153 (I4678,I2067,I4353,I4321,);
not I_154 (I4709,I4670);
nor I_155 (I4726,I61332,I61311);
not I_156 (I4743,I4726);
nor I_157 (I4760,I4517,I4743);
nor I_158 (I4777,I4709,I4760);
DFFARX1 I_159 (I4777,I2067,I4353,I4342,);
nor I_160 (I4808,I4670,I4743);
nor I_161 (I4330,I4534,I4808);
nor I_162 (I4324,I4670,I4726);
not I_163 (I4880,I2074);
DFFARX1 I_164 (I92302,I2067,I4880,I4906,);
DFFARX1 I_165 (I4906,I2067,I4880,I4923,);
not I_166 (I4931,I4923);
nand I_167 (I4948,I92317,I92320);
and I_168 (I4965,I4948,I92299);
DFFARX1 I_169 (I4965,I2067,I4880,I4991,);
DFFARX1 I_170 (I4991,I2067,I4880,I4872,);
DFFARX1 I_171 (I4991,I2067,I4880,I4863,);
DFFARX1 I_172 (I92305,I2067,I4880,I5036,);
nand I_173 (I5044,I5036,I92311);
not I_174 (I5061,I5044);
nor I_175 (I4860,I4906,I5061);
DFFARX1 I_176 (I92299,I2067,I4880,I5101,);
not I_177 (I5109,I5101);
nor I_178 (I4866,I5109,I4931);
nand I_179 (I4854,I5109,I5044);
nand I_180 (I5154,I92314,I92296);
and I_181 (I5171,I5154,I92308);
DFFARX1 I_182 (I5171,I2067,I4880,I5197,);
nor I_183 (I5205,I5197,I4906);
DFFARX1 I_184 (I5205,I2067,I4880,I4848,);
not I_185 (I5236,I5197);
nor I_186 (I5253,I92296,I92296);
not I_187 (I5270,I5253);
nor I_188 (I5287,I5044,I5270);
nor I_189 (I5304,I5236,I5287);
DFFARX1 I_190 (I5304,I2067,I4880,I4869,);
nor I_191 (I5335,I5197,I5270);
nor I_192 (I4857,I5061,I5335);
nor I_193 (I4851,I5197,I5253);
not I_194 (I5407,I2074);
DFFARX1 I_195 (I57575,I2067,I5407,I5433,);
DFFARX1 I_196 (I5433,I2067,I5407,I5450,);
not I_197 (I5458,I5450);
nand I_198 (I5475,I57572,I57566);
and I_199 (I5492,I5475,I57560);
DFFARX1 I_200 (I5492,I2067,I5407,I5518,);
DFFARX1 I_201 (I5518,I2067,I5407,I5399,);
DFFARX1 I_202 (I5518,I2067,I5407,I5390,);
DFFARX1 I_203 (I57548,I2067,I5407,I5563,);
nand I_204 (I5571,I5563,I57557);
not I_205 (I5588,I5571);
nor I_206 (I5387,I5433,I5588);
DFFARX1 I_207 (I57554,I2067,I5407,I5628,);
not I_208 (I5636,I5628);
nor I_209 (I5393,I5636,I5458);
nand I_210 (I5381,I5636,I5571);
nand I_211 (I5681,I57551,I57569);
and I_212 (I5698,I5681,I57548);
DFFARX1 I_213 (I5698,I2067,I5407,I5724,);
nor I_214 (I5732,I5724,I5433);
DFFARX1 I_215 (I5732,I2067,I5407,I5375,);
not I_216 (I5763,I5724);
nor I_217 (I5780,I57563,I57569);
not I_218 (I5797,I5780);
nor I_219 (I5814,I5571,I5797);
nor I_220 (I5831,I5763,I5814);
DFFARX1 I_221 (I5831,I2067,I5407,I5396,);
nor I_222 (I5862,I5724,I5797);
nor I_223 (I5384,I5588,I5862);
nor I_224 (I5378,I5724,I5780);
not I_225 (I5934,I2074);
DFFARX1 I_226 (I50197,I2067,I5934,I5960,);
DFFARX1 I_227 (I5960,I2067,I5934,I5977,);
not I_228 (I5985,I5977);
nand I_229 (I6002,I50194,I50188);
and I_230 (I6019,I6002,I50182);
DFFARX1 I_231 (I6019,I2067,I5934,I6045,);
DFFARX1 I_232 (I6045,I2067,I5934,I5926,);
DFFARX1 I_233 (I6045,I2067,I5934,I5917,);
DFFARX1 I_234 (I50170,I2067,I5934,I6090,);
nand I_235 (I6098,I6090,I50179);
not I_236 (I6115,I6098);
nor I_237 (I5914,I5960,I6115);
DFFARX1 I_238 (I50176,I2067,I5934,I6155,);
not I_239 (I6163,I6155);
nor I_240 (I5920,I6163,I5985);
nand I_241 (I5908,I6163,I6098);
nand I_242 (I6208,I50173,I50191);
and I_243 (I6225,I6208,I50170);
DFFARX1 I_244 (I6225,I2067,I5934,I6251,);
nor I_245 (I6259,I6251,I5960);
DFFARX1 I_246 (I6259,I2067,I5934,I5902,);
not I_247 (I6290,I6251);
nor I_248 (I6307,I50185,I50191);
not I_249 (I6324,I6307);
nor I_250 (I6341,I6098,I6324);
nor I_251 (I6358,I6290,I6341);
DFFARX1 I_252 (I6358,I2067,I5934,I5923,);
nor I_253 (I6389,I6251,I6324);
nor I_254 (I5911,I6115,I6389);
nor I_255 (I5905,I6251,I6307);
not I_256 (I6461,I2074);
DFFARX1 I_257 (I106024,I2067,I6461,I6487,);
DFFARX1 I_258 (I6487,I2067,I6461,I6504,);
not I_259 (I6512,I6504);
nand I_260 (I6529,I106015,I106036);
and I_261 (I6546,I6529,I106018);
DFFARX1 I_262 (I6546,I2067,I6461,I6572,);
DFFARX1 I_263 (I6572,I2067,I6461,I6453,);
DFFARX1 I_264 (I6572,I2067,I6461,I6444,);
DFFARX1 I_265 (I106018,I2067,I6461,I6617,);
nand I_266 (I6625,I6617,I106033);
not I_267 (I6642,I6625);
nor I_268 (I6441,I6487,I6642);
DFFARX1 I_269 (I106027,I2067,I6461,I6682,);
not I_270 (I6690,I6682);
nor I_271 (I6447,I6690,I6512);
nand I_272 (I6435,I6690,I6625);
nand I_273 (I6735,I106021,I106030);
and I_274 (I6752,I6735,I106015);
DFFARX1 I_275 (I6752,I2067,I6461,I6778,);
nor I_276 (I6786,I6778,I6487);
DFFARX1 I_277 (I6786,I2067,I6461,I6429,);
not I_278 (I6817,I6778);
nor I_279 (I6834,I106021,I106030);
not I_280 (I6851,I6834);
nor I_281 (I6868,I6625,I6851);
nor I_282 (I6885,I6817,I6868);
DFFARX1 I_283 (I6885,I2067,I6461,I6450,);
nor I_284 (I6916,I6778,I6851);
nor I_285 (I6438,I6642,I6916);
nor I_286 (I6432,I6778,I6834);
not I_287 (I6988,I2074);
DFFARX1 I_288 (I50724,I2067,I6988,I7014,);
DFFARX1 I_289 (I7014,I2067,I6988,I7031,);
not I_290 (I7039,I7031);
nand I_291 (I7056,I50721,I50715);
and I_292 (I7073,I7056,I50709);
DFFARX1 I_293 (I7073,I2067,I6988,I7099,);
DFFARX1 I_294 (I7099,I2067,I6988,I6980,);
DFFARX1 I_295 (I7099,I2067,I6988,I6971,);
DFFARX1 I_296 (I50697,I2067,I6988,I7144,);
nand I_297 (I7152,I7144,I50706);
not I_298 (I7169,I7152);
nor I_299 (I6968,I7014,I7169);
DFFARX1 I_300 (I50703,I2067,I6988,I7209,);
not I_301 (I7217,I7209);
nor I_302 (I6974,I7217,I7039);
nand I_303 (I6962,I7217,I7152);
nand I_304 (I7262,I50700,I50718);
and I_305 (I7279,I7262,I50697);
DFFARX1 I_306 (I7279,I2067,I6988,I7305,);
nor I_307 (I7313,I7305,I7014);
DFFARX1 I_308 (I7313,I2067,I6988,I6956,);
not I_309 (I7344,I7305);
nor I_310 (I7361,I50712,I50718);
not I_311 (I7378,I7361);
nor I_312 (I7395,I7152,I7378);
nor I_313 (I7412,I7344,I7395);
DFFARX1 I_314 (I7412,I2067,I6988,I6977,);
nor I_315 (I7443,I7305,I7378);
nor I_316 (I6965,I7169,I7443);
nor I_317 (I6959,I7305,I7361);
not I_318 (I7515,I2074);
DFFARX1 I_319 (I70715,I2067,I7515,I7541,);
DFFARX1 I_320 (I7541,I2067,I7515,I7558,);
not I_321 (I7566,I7558);
nand I_322 (I7583,I70721,I70709);
and I_323 (I7600,I7583,I70706);
DFFARX1 I_324 (I7600,I2067,I7515,I7626,);
DFFARX1 I_325 (I7626,I2067,I7515,I7507,);
DFFARX1 I_326 (I7626,I2067,I7515,I7498,);
DFFARX1 I_327 (I70718,I2067,I7515,I7671,);
nand I_328 (I7679,I7671,I70712);
not I_329 (I7696,I7679);
nor I_330 (I7495,I7541,I7696);
DFFARX1 I_331 (I70730,I2067,I7515,I7736,);
not I_332 (I7744,I7736);
nor I_333 (I7501,I7744,I7566);
nand I_334 (I7489,I7744,I7679);
nand I_335 (I7789,I70724,I70727);
and I_336 (I7806,I7789,I70709);
DFFARX1 I_337 (I7806,I2067,I7515,I7832,);
nor I_338 (I7840,I7832,I7541);
DFFARX1 I_339 (I7840,I2067,I7515,I7483,);
not I_340 (I7871,I7832);
nor I_341 (I7888,I70706,I70727);
not I_342 (I7905,I7888);
nor I_343 (I7922,I7679,I7905);
nor I_344 (I7939,I7871,I7922);
DFFARX1 I_345 (I7939,I2067,I7515,I7504,);
nor I_346 (I7970,I7832,I7905);
nor I_347 (I7492,I7696,I7970);
nor I_348 (I7486,I7832,I7888);
not I_349 (I8042,I2074);
DFFARX1 I_350 (I87678,I2067,I8042,I8068,);
DFFARX1 I_351 (I8068,I2067,I8042,I8085,);
not I_352 (I8093,I8085);
nand I_353 (I8110,I87693,I87696);
and I_354 (I8127,I8110,I87675);
DFFARX1 I_355 (I8127,I2067,I8042,I8153,);
DFFARX1 I_356 (I8153,I2067,I8042,I8034,);
DFFARX1 I_357 (I8153,I2067,I8042,I8025,);
DFFARX1 I_358 (I87681,I2067,I8042,I8198,);
nand I_359 (I8206,I8198,I87687);
not I_360 (I8223,I8206);
nor I_361 (I8022,I8068,I8223);
DFFARX1 I_362 (I87675,I2067,I8042,I8263,);
not I_363 (I8271,I8263);
nor I_364 (I8028,I8271,I8093);
nand I_365 (I8016,I8271,I8206);
nand I_366 (I8316,I87690,I87672);
and I_367 (I8333,I8316,I87684);
DFFARX1 I_368 (I8333,I2067,I8042,I8359,);
nor I_369 (I8367,I8359,I8068);
DFFARX1 I_370 (I8367,I2067,I8042,I8010,);
not I_371 (I8398,I8359);
nor I_372 (I8415,I87672,I87672);
not I_373 (I8432,I8415);
nor I_374 (I8449,I8206,I8432);
nor I_375 (I8466,I8398,I8449);
DFFARX1 I_376 (I8466,I2067,I8042,I8031,);
nor I_377 (I8497,I8359,I8432);
nor I_378 (I8019,I8223,I8497);
nor I_379 (I8013,I8359,I8415);
not I_380 (I8569,I2074);
DFFARX1 I_381 (I100394,I2067,I8569,I8595,);
DFFARX1 I_382 (I8595,I2067,I8569,I8612,);
not I_383 (I8620,I8612);
nand I_384 (I8637,I100409,I100412);
and I_385 (I8654,I8637,I100391);
DFFARX1 I_386 (I8654,I2067,I8569,I8680,);
DFFARX1 I_387 (I8680,I2067,I8569,I8561,);
DFFARX1 I_388 (I8680,I2067,I8569,I8552,);
DFFARX1 I_389 (I100397,I2067,I8569,I8725,);
nand I_390 (I8733,I8725,I100403);
not I_391 (I8750,I8733);
nor I_392 (I8549,I8595,I8750);
DFFARX1 I_393 (I100391,I2067,I8569,I8790,);
not I_394 (I8798,I8790);
nor I_395 (I8555,I8798,I8620);
nand I_396 (I8543,I8798,I8733);
nand I_397 (I8843,I100406,I100388);
and I_398 (I8860,I8843,I100400);
DFFARX1 I_399 (I8860,I2067,I8569,I8886,);
nor I_400 (I8894,I8886,I8595);
DFFARX1 I_401 (I8894,I2067,I8569,I8537,);
not I_402 (I8925,I8886);
nor I_403 (I8942,I100388,I100388);
not I_404 (I8959,I8942);
nor I_405 (I8976,I8733,I8959);
nor I_406 (I8993,I8925,I8976);
DFFARX1 I_407 (I8993,I2067,I8569,I8558,);
nor I_408 (I9024,I8886,I8959);
nor I_409 (I8546,I8750,I9024);
nor I_410 (I8540,I8886,I8942);
not I_411 (I9096,I2074);
DFFARX1 I_412 (I160617,I2067,I9096,I9122,);
DFFARX1 I_413 (I9122,I2067,I9096,I9139,);
not I_414 (I9147,I9139);
nand I_415 (I9164,I160620,I160614);
and I_416 (I9181,I9164,I160623);
DFFARX1 I_417 (I9181,I2067,I9096,I9207,);
DFFARX1 I_418 (I9207,I2067,I9096,I9088,);
DFFARX1 I_419 (I9207,I2067,I9096,I9079,);
DFFARX1 I_420 (I160611,I2067,I9096,I9252,);
nand I_421 (I9260,I9252,I160626);
not I_422 (I9277,I9260);
nor I_423 (I9076,I9122,I9277);
DFFARX1 I_424 (I160602,I2067,I9096,I9317,);
not I_425 (I9325,I9317);
nor I_426 (I9082,I9325,I9147);
nand I_427 (I9070,I9325,I9260);
nand I_428 (I9370,I160605,I160605);
and I_429 (I9387,I9370,I160602);
DFFARX1 I_430 (I9387,I2067,I9096,I9413,);
nor I_431 (I9421,I9413,I9122);
DFFARX1 I_432 (I9421,I2067,I9096,I9064,);
not I_433 (I9452,I9413);
nor I_434 (I9469,I160608,I160605);
not I_435 (I9486,I9469);
nor I_436 (I9503,I9260,I9486);
nor I_437 (I9520,I9452,I9503);
DFFARX1 I_438 (I9520,I2067,I9096,I9085,);
nor I_439 (I9551,I9413,I9486);
nor I_440 (I9073,I9277,I9551);
nor I_441 (I9067,I9413,I9469);
not I_442 (I9623,I2074);
DFFARX1 I_443 (I53359,I2067,I9623,I9649,);
not I_444 (I9657,I9649);
nand I_445 (I9674,I53341,I53356);
and I_446 (I9691,I9674,I53332);
DFFARX1 I_447 (I9691,I2067,I9623,I9717,);
DFFARX1 I_448 (I53335,I2067,I9623,I9734,);
and I_449 (I9742,I9734,I53350);
nor I_450 (I9759,I9717,I9742);
DFFARX1 I_451 (I9759,I2067,I9623,I9591,);
nand I_452 (I9790,I9734,I53350);
nand I_453 (I9807,I9657,I9790);
not I_454 (I9603,I9807);
DFFARX1 I_455 (I53353,I2067,I9623,I9847,);
DFFARX1 I_456 (I9847,I2067,I9623,I9612,);
nand I_457 (I9869,I53332,I53344);
and I_458 (I9886,I9869,I53338);
DFFARX1 I_459 (I9886,I2067,I9623,I9912,);
DFFARX1 I_460 (I9912,I2067,I9623,I9929,);
not I_461 (I9615,I9929);
not I_462 (I9951,I9912);
nand I_463 (I9600,I9951,I9790);
nor I_464 (I9982,I53347,I53344);
not I_465 (I9999,I9982);
nor I_466 (I10016,I9951,I9999);
nor I_467 (I10033,I9657,I10016);
DFFARX1 I_468 (I10033,I2067,I9623,I9609,);
nor I_469 (I10064,I9717,I9999);
nor I_470 (I9597,I9912,I10064);
nor I_471 (I9606,I9847,I9982);
nor I_472 (I9594,I9717,I9982);
not I_473 (I10150,I2074);
DFFARX1 I_474 (I98088,I2067,I10150,I10176,);
not I_475 (I10184,I10176);
nand I_476 (I10201,I98079,I98097);
and I_477 (I10218,I10201,I98076);
DFFARX1 I_478 (I10218,I2067,I10150,I10244,);
DFFARX1 I_479 (I98079,I2067,I10150,I10261,);
and I_480 (I10269,I10261,I98082);
nor I_481 (I10286,I10244,I10269);
DFFARX1 I_482 (I10286,I2067,I10150,I10118,);
nand I_483 (I10317,I10261,I98082);
nand I_484 (I10334,I10184,I10317);
not I_485 (I10130,I10334);
DFFARX1 I_486 (I98076,I2067,I10150,I10374,);
DFFARX1 I_487 (I10374,I2067,I10150,I10139,);
nand I_488 (I10396,I98094,I98085);
and I_489 (I10413,I10396,I98100);
DFFARX1 I_490 (I10413,I2067,I10150,I10439,);
DFFARX1 I_491 (I10439,I2067,I10150,I10456,);
not I_492 (I10142,I10456);
not I_493 (I10478,I10439);
nand I_494 (I10127,I10478,I10317);
nor I_495 (I10509,I98091,I98085);
not I_496 (I10526,I10509);
nor I_497 (I10543,I10478,I10526);
nor I_498 (I10560,I10184,I10543);
DFFARX1 I_499 (I10560,I2067,I10150,I10136,);
nor I_500 (I10591,I10244,I10526);
nor I_501 (I10124,I10439,I10591);
nor I_502 (I10133,I10374,I10509);
nor I_503 (I10121,I10244,I10509);
not I_504 (I10677,I2074);
DFFARX1 I_505 (I85369,I2067,I10677,I10703,);
not I_506 (I10711,I10703);
nand I_507 (I10728,I85381,I85366);
and I_508 (I10745,I10728,I85360);
DFFARX1 I_509 (I10745,I2067,I10677,I10771,);
DFFARX1 I_510 (I85375,I2067,I10677,I10788,);
and I_511 (I10796,I10788,I85363);
nor I_512 (I10813,I10771,I10796);
DFFARX1 I_513 (I10813,I2067,I10677,I10645,);
nand I_514 (I10844,I10788,I85363);
nand I_515 (I10861,I10711,I10844);
not I_516 (I10657,I10861);
DFFARX1 I_517 (I85372,I2067,I10677,I10901,);
DFFARX1 I_518 (I10901,I2067,I10677,I10666,);
nand I_519 (I10923,I85378,I85384);
and I_520 (I10940,I10923,I85360);
DFFARX1 I_521 (I10940,I2067,I10677,I10966,);
DFFARX1 I_522 (I10966,I2067,I10677,I10983,);
not I_523 (I10669,I10983);
not I_524 (I11005,I10966);
nand I_525 (I10654,I11005,I10844);
nor I_526 (I11036,I85363,I85384);
not I_527 (I11053,I11036);
nor I_528 (I11070,I11005,I11053);
nor I_529 (I11087,I10711,I11070);
DFFARX1 I_530 (I11087,I2067,I10677,I10663,);
nor I_531 (I11118,I10771,I11053);
nor I_532 (I10651,I10966,I11118);
nor I_533 (I10660,I10901,I11036);
nor I_534 (I10648,I10771,I11036);
not I_535 (I11204,I2074);
DFFARX1 I_536 (I2092,I2067,I11204,I11230,);
not I_537 (I11238,I11230);
nand I_538 (I11255,I2077,I2077);
and I_539 (I11272,I11255,I2098);
DFFARX1 I_540 (I11272,I2067,I11204,I11298,);
DFFARX1 I_541 (I2080,I2067,I11204,I11315,);
and I_542 (I11323,I11315,I2089);
nor I_543 (I11340,I11298,I11323);
DFFARX1 I_544 (I11340,I2067,I11204,I11172,);
nand I_545 (I11371,I11315,I2089);
nand I_546 (I11388,I11238,I11371);
not I_547 (I11184,I11388);
DFFARX1 I_548 (I2083,I2067,I11204,I11428,);
DFFARX1 I_549 (I11428,I2067,I11204,I11193,);
nand I_550 (I11450,I2086,I2095);
and I_551 (I11467,I11450,I2080);
DFFARX1 I_552 (I11467,I2067,I11204,I11493,);
DFFARX1 I_553 (I11493,I2067,I11204,I11510,);
not I_554 (I11196,I11510);
not I_555 (I11532,I11493);
nand I_556 (I11181,I11532,I11371);
nor I_557 (I11563,I2083,I2095);
not I_558 (I11580,I11563);
nor I_559 (I11597,I11532,I11580);
nor I_560 (I11614,I11238,I11597);
DFFARX1 I_561 (I11614,I2067,I11204,I11190,);
nor I_562 (I11645,I11298,I11580);
nor I_563 (I11178,I11493,I11645);
nor I_564 (I11187,I11428,I11563);
nor I_565 (I11175,I11298,I11563);
not I_566 (I11731,I2074);
DFFARX1 I_567 (I112875,I2067,I11731,I11757,);
not I_568 (I11765,I11757);
nand I_569 (I11782,I112872,I112887);
and I_570 (I11799,I11782,I112869);
DFFARX1 I_571 (I11799,I2067,I11731,I11825,);
DFFARX1 I_572 (I112866,I2067,I11731,I11842,);
and I_573 (I11850,I11842,I112866);
nor I_574 (I11867,I11825,I11850);
DFFARX1 I_575 (I11867,I2067,I11731,I11699,);
nand I_576 (I11898,I11842,I112866);
nand I_577 (I11915,I11765,I11898);
not I_578 (I11711,I11915);
DFFARX1 I_579 (I112869,I2067,I11731,I11955,);
DFFARX1 I_580 (I11955,I2067,I11731,I11720,);
nand I_581 (I11977,I112881,I112872);
and I_582 (I11994,I11977,I112884);
DFFARX1 I_583 (I11994,I2067,I11731,I12020,);
DFFARX1 I_584 (I12020,I2067,I11731,I12037,);
not I_585 (I11723,I12037);
not I_586 (I12059,I12020);
nand I_587 (I11708,I12059,I11898);
nor I_588 (I12090,I112878,I112872);
not I_589 (I12107,I12090);
nor I_590 (I12124,I12059,I12107);
nor I_591 (I12141,I11765,I12124);
DFFARX1 I_592 (I12141,I2067,I11731,I11717,);
nor I_593 (I12172,I11825,I12107);
nor I_594 (I11705,I12020,I12172);
nor I_595 (I11714,I11955,I12090);
nor I_596 (I11702,I11825,I12090);
not I_597 (I12258,I2074);
DFFARX1 I_598 (I168111,I2067,I12258,I12284,);
not I_599 (I12292,I12284);
nand I_600 (I12309,I168105,I168126);
and I_601 (I12326,I12309,I168102);
DFFARX1 I_602 (I12326,I2067,I12258,I12352,);
DFFARX1 I_603 (I168123,I2067,I12258,I12369,);
and I_604 (I12377,I12369,I168120);
nor I_605 (I12394,I12352,I12377);
DFFARX1 I_606 (I12394,I2067,I12258,I12226,);
nand I_607 (I12425,I12369,I168120);
nand I_608 (I12442,I12292,I12425);
not I_609 (I12238,I12442);
DFFARX1 I_610 (I168108,I2067,I12258,I12482,);
DFFARX1 I_611 (I12482,I2067,I12258,I12247,);
nand I_612 (I12504,I168117,I168114);
and I_613 (I12521,I12504,I168099);
DFFARX1 I_614 (I12521,I2067,I12258,I12547,);
DFFARX1 I_615 (I12547,I2067,I12258,I12564,);
not I_616 (I12250,I12564);
not I_617 (I12586,I12547);
nand I_618 (I12235,I12586,I12425);
nor I_619 (I12617,I168099,I168114);
not I_620 (I12634,I12617);
nor I_621 (I12651,I12586,I12634);
nor I_622 (I12668,I12292,I12651);
DFFARX1 I_623 (I12668,I2067,I12258,I12244,);
nor I_624 (I12699,I12352,I12634);
nor I_625 (I12232,I12547,I12699);
nor I_626 (I12241,I12482,I12617);
nor I_627 (I12229,I12352,I12617);
not I_628 (I12785,I2074);
DFFARX1 I_629 (I67307,I2067,I12785,I12811,);
not I_630 (I12819,I12811);
nand I_631 (I12836,I67301,I67292);
and I_632 (I12853,I12836,I67313);
DFFARX1 I_633 (I12853,I2067,I12785,I12879,);
DFFARX1 I_634 (I67295,I2067,I12785,I12896,);
and I_635 (I12904,I12896,I67289);
nor I_636 (I12921,I12879,I12904);
DFFARX1 I_637 (I12921,I2067,I12785,I12753,);
nand I_638 (I12952,I12896,I67289);
nand I_639 (I12969,I12819,I12952);
not I_640 (I12765,I12969);
DFFARX1 I_641 (I67289,I2067,I12785,I13009,);
DFFARX1 I_642 (I13009,I2067,I12785,I12774,);
nand I_643 (I13031,I67316,I67298);
and I_644 (I13048,I13031,I67304);
DFFARX1 I_645 (I13048,I2067,I12785,I13074,);
DFFARX1 I_646 (I13074,I2067,I12785,I13091,);
not I_647 (I12777,I13091);
not I_648 (I13113,I13074);
nand I_649 (I12762,I13113,I12952);
nor I_650 (I13144,I67310,I67298);
not I_651 (I13161,I13144);
nor I_652 (I13178,I13113,I13161);
nor I_653 (I13195,I12819,I13178);
DFFARX1 I_654 (I13195,I2067,I12785,I12771,);
nor I_655 (I13226,I12879,I13161);
nor I_656 (I12759,I13074,I13226);
nor I_657 (I12768,I13009,I13144);
nor I_658 (I12756,I12879,I13144);
not I_659 (I13312,I2074);
DFFARX1 I_660 (I69519,I2067,I13312,I13338,);
not I_661 (I13346,I13338);
nand I_662 (I13363,I69540,I69534);
and I_663 (I13380,I13363,I69516);
DFFARX1 I_664 (I13380,I2067,I13312,I13406,);
DFFARX1 I_665 (I69519,I2067,I13312,I13423,);
and I_666 (I13431,I13423,I69528);
nor I_667 (I13448,I13406,I13431);
DFFARX1 I_668 (I13448,I2067,I13312,I13280,);
nand I_669 (I13479,I13423,I69528);
nand I_670 (I13496,I13346,I13479);
not I_671 (I13292,I13496);
DFFARX1 I_672 (I69525,I2067,I13312,I13536,);
DFFARX1 I_673 (I13536,I2067,I13312,I13301,);
nand I_674 (I13558,I69531,I69522);
and I_675 (I13575,I13558,I69516);
DFFARX1 I_676 (I13575,I2067,I13312,I13601,);
DFFARX1 I_677 (I13601,I2067,I13312,I13618,);
not I_678 (I13304,I13618);
not I_679 (I13640,I13601);
nand I_680 (I13289,I13640,I13479);
nor I_681 (I13671,I69537,I69522);
not I_682 (I13688,I13671);
nor I_683 (I13705,I13640,I13688);
nor I_684 (I13722,I13346,I13705);
DFFARX1 I_685 (I13722,I2067,I13312,I13298,);
nor I_686 (I13753,I13406,I13688);
nor I_687 (I13286,I13601,I13753);
nor I_688 (I13295,I13536,I13671);
nor I_689 (I13283,I13406,I13671);
not I_690 (I13839,I2074);
DFFARX1 I_691 (I162357,I2067,I13839,I13865,);
not I_692 (I13873,I13865);
nand I_693 (I13890,I162360,I162354);
and I_694 (I13907,I13890,I162351);
DFFARX1 I_695 (I13907,I2067,I13839,I13933,);
DFFARX1 I_696 (I162336,I2067,I13839,I13950,);
and I_697 (I13958,I13950,I162345);
nor I_698 (I13975,I13933,I13958);
DFFARX1 I_699 (I13975,I2067,I13839,I13807,);
nand I_700 (I14006,I13950,I162345);
nand I_701 (I14023,I13873,I14006);
not I_702 (I13819,I14023);
DFFARX1 I_703 (I162336,I2067,I13839,I14063,);
DFFARX1 I_704 (I14063,I2067,I13839,I13828,);
nand I_705 (I14085,I162339,I162342);
and I_706 (I14102,I14085,I162348);
DFFARX1 I_707 (I14102,I2067,I13839,I14128,);
DFFARX1 I_708 (I14128,I2067,I13839,I14145,);
not I_709 (I13831,I14145);
not I_710 (I14167,I14128);
nand I_711 (I13816,I14167,I14006);
nor I_712 (I14198,I162339,I162342);
not I_713 (I14215,I14198);
nor I_714 (I14232,I14167,I14215);
nor I_715 (I14249,I13873,I14232);
DFFARX1 I_716 (I14249,I2067,I13839,I13825,);
nor I_717 (I14280,I13933,I14215);
nor I_718 (I13813,I14128,I14280);
nor I_719 (I13822,I14063,I14198);
nor I_720 (I13810,I13933,I14198);
not I_721 (I14366,I2074);
DFFARX1 I_722 (I7507,I2067,I14366,I14392,);
not I_723 (I14400,I14392);
nand I_724 (I14417,I7495,I7501);
and I_725 (I14434,I14417,I7504);
DFFARX1 I_726 (I14434,I2067,I14366,I14460,);
DFFARX1 I_727 (I7486,I2067,I14366,I14477,);
and I_728 (I14485,I14477,I7492);
nor I_729 (I14502,I14460,I14485);
DFFARX1 I_730 (I14502,I2067,I14366,I14334,);
nand I_731 (I14533,I14477,I7492);
nand I_732 (I14550,I14400,I14533);
not I_733 (I14346,I14550);
DFFARX1 I_734 (I7486,I2067,I14366,I14590,);
DFFARX1 I_735 (I14590,I2067,I14366,I14355,);
nand I_736 (I14612,I7489,I7483);
and I_737 (I14629,I14612,I7498);
DFFARX1 I_738 (I14629,I2067,I14366,I14655,);
DFFARX1 I_739 (I14655,I2067,I14366,I14672,);
not I_740 (I14358,I14672);
not I_741 (I14694,I14655);
nand I_742 (I14343,I14694,I14533);
nor I_743 (I14725,I7483,I7483);
not I_744 (I14742,I14725);
nor I_745 (I14759,I14694,I14742);
nor I_746 (I14776,I14400,I14759);
DFFARX1 I_747 (I14776,I2067,I14366,I14352,);
nor I_748 (I14807,I14460,I14742);
nor I_749 (I14340,I14655,I14807);
nor I_750 (I14349,I14590,I14725);
nor I_751 (I14337,I14460,I14725);
not I_752 (I14893,I2074);
DFFARX1 I_753 (I83635,I2067,I14893,I14919,);
not I_754 (I14927,I14919);
nand I_755 (I14944,I83647,I83632);
and I_756 (I14961,I14944,I83626);
DFFARX1 I_757 (I14961,I2067,I14893,I14987,);
DFFARX1 I_758 (I83641,I2067,I14893,I15004,);
and I_759 (I15012,I15004,I83629);
nor I_760 (I15029,I14987,I15012);
DFFARX1 I_761 (I15029,I2067,I14893,I14861,);
nand I_762 (I15060,I15004,I83629);
nand I_763 (I15077,I14927,I15060);
not I_764 (I14873,I15077);
DFFARX1 I_765 (I83638,I2067,I14893,I15117,);
DFFARX1 I_766 (I15117,I2067,I14893,I14882,);
nand I_767 (I15139,I83644,I83650);
and I_768 (I15156,I15139,I83626);
DFFARX1 I_769 (I15156,I2067,I14893,I15182,);
DFFARX1 I_770 (I15182,I2067,I14893,I15199,);
not I_771 (I14885,I15199);
not I_772 (I15221,I15182);
nand I_773 (I14870,I15221,I15060);
nor I_774 (I15252,I83629,I83650);
not I_775 (I15269,I15252);
nor I_776 (I15286,I15221,I15269);
nor I_777 (I15303,I14927,I15286);
DFFARX1 I_778 (I15303,I2067,I14893,I14879,);
nor I_779 (I15334,I14987,I15269);
nor I_780 (I14867,I15182,I15334);
nor I_781 (I14876,I15117,I15252);
nor I_782 (I14864,I14987,I15252);
not I_783 (I15420,I2074);
DFFARX1 I_784 (I1820,I2067,I15420,I15446,);
not I_785 (I15454,I15446);
nand I_786 (I15471,I1668,I1956);
and I_787 (I15488,I15471,I1828);
DFFARX1 I_788 (I15488,I2067,I15420,I15514,);
DFFARX1 I_789 (I1644,I2067,I15420,I15531,);
and I_790 (I15539,I15531,I1548);
nor I_791 (I15556,I15514,I15539);
DFFARX1 I_792 (I15556,I2067,I15420,I15388,);
nand I_793 (I15587,I15531,I1548);
nand I_794 (I15604,I15454,I15587);
not I_795 (I15400,I15604);
DFFARX1 I_796 (I1980,I2067,I15420,I15644,);
DFFARX1 I_797 (I15644,I2067,I15420,I15409,);
nand I_798 (I15666,I1732,I1756);
and I_799 (I15683,I15666,I1516);
DFFARX1 I_800 (I15683,I2067,I15420,I15709,);
DFFARX1 I_801 (I15709,I2067,I15420,I15726,);
not I_802 (I15412,I15726);
not I_803 (I15748,I15709);
nand I_804 (I15397,I15748,I15587);
nor I_805 (I15779,I1636,I1756);
not I_806 (I15796,I15779);
nor I_807 (I15813,I15748,I15796);
nor I_808 (I15830,I15454,I15813);
DFFARX1 I_809 (I15830,I2067,I15420,I15406,);
nor I_810 (I15861,I15514,I15796);
nor I_811 (I15394,I15709,I15861);
nor I_812 (I15403,I15644,I15779);
nor I_813 (I15391,I15514,I15779);
not I_814 (I15947,I2074);
DFFARX1 I_815 (I79589,I2067,I15947,I15973,);
not I_816 (I15981,I15973);
nand I_817 (I15998,I79601,I79586);
and I_818 (I16015,I15998,I79580);
DFFARX1 I_819 (I16015,I2067,I15947,I16041,);
DFFARX1 I_820 (I79595,I2067,I15947,I16058,);
and I_821 (I16066,I16058,I79583);
nor I_822 (I16083,I16041,I16066);
DFFARX1 I_823 (I16083,I2067,I15947,I15915,);
nand I_824 (I16114,I16058,I79583);
nand I_825 (I16131,I15981,I16114);
not I_826 (I15927,I16131);
DFFARX1 I_827 (I79592,I2067,I15947,I16171,);
DFFARX1 I_828 (I16171,I2067,I15947,I15936,);
nand I_829 (I16193,I79598,I79604);
and I_830 (I16210,I16193,I79580);
DFFARX1 I_831 (I16210,I2067,I15947,I16236,);
DFFARX1 I_832 (I16236,I2067,I15947,I16253,);
not I_833 (I15939,I16253);
not I_834 (I16275,I16236);
nand I_835 (I15924,I16275,I16114);
nor I_836 (I16306,I79583,I79604);
not I_837 (I16323,I16306);
nor I_838 (I16340,I16275,I16323);
nor I_839 (I16357,I15981,I16340);
DFFARX1 I_840 (I16357,I2067,I15947,I15933,);
nor I_841 (I16388,I16041,I16323);
nor I_842 (I15921,I16236,I16388);
nor I_843 (I15930,I16171,I16306);
nor I_844 (I15918,I16041,I16306);
not I_845 (I16474,I2074);
DFFARX1 I_846 (I136244,I2067,I16474,I16500,);
not I_847 (I16508,I16500);
nand I_848 (I16525,I136241,I136247);
and I_849 (I16542,I16525,I136244);
DFFARX1 I_850 (I16542,I2067,I16474,I16568,);
DFFARX1 I_851 (I136247,I2067,I16474,I16585,);
and I_852 (I16593,I16585,I136241);
nor I_853 (I16610,I16568,I16593);
DFFARX1 I_854 (I16610,I2067,I16474,I16442,);
nand I_855 (I16641,I16585,I136241);
nand I_856 (I16658,I16508,I16641);
not I_857 (I16454,I16658);
DFFARX1 I_858 (I136250,I2067,I16474,I16698,);
DFFARX1 I_859 (I16698,I2067,I16474,I16463,);
nand I_860 (I16720,I136253,I136262);
and I_861 (I16737,I16720,I136256);
DFFARX1 I_862 (I16737,I2067,I16474,I16763,);
DFFARX1 I_863 (I16763,I2067,I16474,I16780,);
not I_864 (I16466,I16780);
not I_865 (I16802,I16763);
nand I_866 (I16451,I16802,I16641);
nor I_867 (I16833,I136259,I136262);
not I_868 (I16850,I16833);
nor I_869 (I16867,I16802,I16850);
nor I_870 (I16884,I16508,I16867);
DFFARX1 I_871 (I16884,I2067,I16474,I16460,);
nor I_872 (I16915,I16568,I16850);
nor I_873 (I16448,I16763,I16915);
nor I_874 (I16457,I16698,I16833);
nor I_875 (I16445,I16568,I16833);
not I_876 (I17001,I2074);
DFFARX1 I_877 (I53886,I2067,I17001,I17027,);
not I_878 (I17035,I17027);
nand I_879 (I17052,I53868,I53883);
and I_880 (I17069,I17052,I53859);
DFFARX1 I_881 (I17069,I2067,I17001,I17095,);
DFFARX1 I_882 (I53862,I2067,I17001,I17112,);
and I_883 (I17120,I17112,I53877);
nor I_884 (I17137,I17095,I17120);
DFFARX1 I_885 (I17137,I2067,I17001,I16969,);
nand I_886 (I17168,I17112,I53877);
nand I_887 (I17185,I17035,I17168);
not I_888 (I16981,I17185);
DFFARX1 I_889 (I53880,I2067,I17001,I17225,);
DFFARX1 I_890 (I17225,I2067,I17001,I16990,);
nand I_891 (I17247,I53859,I53871);
and I_892 (I17264,I17247,I53865);
DFFARX1 I_893 (I17264,I2067,I17001,I17290,);
DFFARX1 I_894 (I17290,I2067,I17001,I17307,);
not I_895 (I16993,I17307);
not I_896 (I17329,I17290);
nand I_897 (I16978,I17329,I17168);
nor I_898 (I17360,I53874,I53871);
not I_899 (I17377,I17360);
nor I_900 (I17394,I17329,I17377);
nor I_901 (I17411,I17035,I17394);
DFFARX1 I_902 (I17411,I2067,I17001,I16987,);
nor I_903 (I17442,I17095,I17377);
nor I_904 (I16975,I17290,I17442);
nor I_905 (I16984,I17225,I17360);
nor I_906 (I16972,I17095,I17360);
not I_907 (I17528,I2074);
DFFARX1 I_908 (I151836,I2067,I17528,I17554,);
not I_909 (I17562,I17554);
nand I_910 (I17579,I151851,I151830);
and I_911 (I17596,I17579,I151833);
DFFARX1 I_912 (I17596,I2067,I17528,I17622,);
DFFARX1 I_913 (I151854,I2067,I17528,I17639,);
and I_914 (I17647,I17639,I151833);
nor I_915 (I17664,I17622,I17647);
DFFARX1 I_916 (I17664,I2067,I17528,I17496,);
nand I_917 (I17695,I17639,I151833);
nand I_918 (I17712,I17562,I17695);
not I_919 (I17508,I17712);
DFFARX1 I_920 (I151830,I2067,I17528,I17752,);
DFFARX1 I_921 (I17752,I2067,I17528,I17517,);
nand I_922 (I17774,I151842,I151839);
and I_923 (I17791,I17774,I151845);
DFFARX1 I_924 (I17791,I2067,I17528,I17817,);
DFFARX1 I_925 (I17817,I2067,I17528,I17834,);
not I_926 (I17520,I17834);
not I_927 (I17856,I17817);
nand I_928 (I17505,I17856,I17695);
nor I_929 (I17887,I151848,I151839);
not I_930 (I17904,I17887);
nor I_931 (I17921,I17856,I17904);
nor I_932 (I17938,I17562,I17921);
DFFARX1 I_933 (I17938,I2067,I17528,I17514,);
nor I_934 (I17969,I17622,I17904);
nor I_935 (I17502,I17817,I17969);
nor I_936 (I17511,I17752,I17887);
nor I_937 (I17499,I17622,I17887);
not I_938 (I18055,I2074);
DFFARX1 I_939 (I74279,I2067,I18055,I18081,);
not I_940 (I18089,I18081);
nand I_941 (I18106,I74300,I74294);
and I_942 (I18123,I18106,I74276);
DFFARX1 I_943 (I18123,I2067,I18055,I18149,);
DFFARX1 I_944 (I74279,I2067,I18055,I18166,);
and I_945 (I18174,I18166,I74288);
nor I_946 (I18191,I18149,I18174);
DFFARX1 I_947 (I18191,I2067,I18055,I18023,);
nand I_948 (I18222,I18166,I74288);
nand I_949 (I18239,I18089,I18222);
not I_950 (I18035,I18239);
DFFARX1 I_951 (I74285,I2067,I18055,I18279,);
DFFARX1 I_952 (I18279,I2067,I18055,I18044,);
nand I_953 (I18301,I74291,I74282);
and I_954 (I18318,I18301,I74276);
DFFARX1 I_955 (I18318,I2067,I18055,I18344,);
DFFARX1 I_956 (I18344,I2067,I18055,I18361,);
not I_957 (I18047,I18361);
not I_958 (I18383,I18344);
nand I_959 (I18032,I18383,I18222);
nor I_960 (I18414,I74297,I74282);
not I_961 (I18431,I18414);
nor I_962 (I18448,I18383,I18431);
nor I_963 (I18465,I18089,I18448);
DFFARX1 I_964 (I18465,I2067,I18055,I18041,);
nor I_965 (I18496,I18149,I18431);
nor I_966 (I18029,I18344,I18496);
nor I_967 (I18038,I18279,I18414);
nor I_968 (I18026,I18149,I18414);
not I_969 (I18582,I2074);
DFFARX1 I_970 (I1748,I2067,I18582,I18608,);
not I_971 (I18616,I18608);
nand I_972 (I18633,I1420,I1364);
and I_973 (I18650,I18633,I1404);
DFFARX1 I_974 (I18650,I2067,I18582,I18676,);
DFFARX1 I_975 (I1964,I2067,I18582,I18693,);
and I_976 (I18701,I18693,I1628);
nor I_977 (I18718,I18676,I18701);
DFFARX1 I_978 (I18718,I2067,I18582,I18550,);
nand I_979 (I18749,I18693,I1628);
nand I_980 (I18766,I18616,I18749);
not I_981 (I18562,I18766);
DFFARX1 I_982 (I1692,I2067,I18582,I18806,);
DFFARX1 I_983 (I18806,I2067,I18582,I18571,);
nand I_984 (I18828,I1540,I1932);
and I_985 (I18845,I18828,I1988);
DFFARX1 I_986 (I18845,I2067,I18582,I18871,);
DFFARX1 I_987 (I18871,I2067,I18582,I18888,);
not I_988 (I18574,I18888);
not I_989 (I18910,I18871);
nand I_990 (I18559,I18910,I18749);
nor I_991 (I18941,I1908,I1932);
not I_992 (I18958,I18941);
nor I_993 (I18975,I18910,I18958);
nor I_994 (I18992,I18616,I18975);
DFFARX1 I_995 (I18992,I2067,I18582,I18568,);
nor I_996 (I19023,I18676,I18958);
nor I_997 (I18556,I18871,I19023);
nor I_998 (I18565,I18806,I18941);
nor I_999 (I18553,I18676,I18941);
not I_1000 (I19109,I2074);
DFFARX1 I_1001 (I26875,I2067,I19109,I19135,);
not I_1002 (I19143,I19135);
nand I_1003 (I19160,I26869,I26863);
and I_1004 (I19177,I19160,I26884);
DFFARX1 I_1005 (I19177,I2067,I19109,I19203,);
DFFARX1 I_1006 (I26881,I2067,I19109,I19220,);
and I_1007 (I19228,I19220,I26878);
nor I_1008 (I19245,I19203,I19228);
DFFARX1 I_1009 (I19245,I2067,I19109,I19077,);
nand I_1010 (I19276,I19220,I26878);
nand I_1011 (I19293,I19143,I19276);
not I_1012 (I19089,I19293);
DFFARX1 I_1013 (I26863,I2067,I19109,I19333,);
DFFARX1 I_1014 (I19333,I2067,I19109,I19098,);
nand I_1015 (I19355,I26866,I26866);
and I_1016 (I19372,I19355,I26887);
DFFARX1 I_1017 (I19372,I2067,I19109,I19398,);
DFFARX1 I_1018 (I19398,I2067,I19109,I19415,);
not I_1019 (I19101,I19415);
not I_1020 (I19437,I19398);
nand I_1021 (I19086,I19437,I19276);
nor I_1022 (I19468,I26872,I26866);
not I_1023 (I19485,I19468);
nor I_1024 (I19502,I19437,I19485);
nor I_1025 (I19519,I19143,I19502);
DFFARX1 I_1026 (I19519,I2067,I19109,I19095,);
nor I_1027 (I19550,I19203,I19485);
nor I_1028 (I19083,I19398,I19550);
nor I_1029 (I19092,I19333,I19468);
nor I_1030 (I19080,I19203,I19468);
not I_1031 (I19636,I2074);
DFFARX1 I_1032 (I84791,I2067,I19636,I19662,);
not I_1033 (I19670,I19662);
nand I_1034 (I19687,I84803,I84788);
and I_1035 (I19704,I19687,I84782);
DFFARX1 I_1036 (I19704,I2067,I19636,I19730,);
DFFARX1 I_1037 (I84797,I2067,I19636,I19747,);
and I_1038 (I19755,I19747,I84785);
nor I_1039 (I19772,I19730,I19755);
DFFARX1 I_1040 (I19772,I2067,I19636,I19604,);
nand I_1041 (I19803,I19747,I84785);
nand I_1042 (I19820,I19670,I19803);
not I_1043 (I19616,I19820);
DFFARX1 I_1044 (I84794,I2067,I19636,I19860,);
DFFARX1 I_1045 (I19860,I2067,I19636,I19625,);
nand I_1046 (I19882,I84800,I84806);
and I_1047 (I19899,I19882,I84782);
DFFARX1 I_1048 (I19899,I2067,I19636,I19925,);
DFFARX1 I_1049 (I19925,I2067,I19636,I19942,);
not I_1050 (I19628,I19942);
not I_1051 (I19964,I19925);
nand I_1052 (I19613,I19964,I19803);
nor I_1053 (I19995,I84785,I84806);
not I_1054 (I20012,I19995);
nor I_1055 (I20029,I19964,I20012);
nor I_1056 (I20046,I19670,I20029);
DFFARX1 I_1057 (I20046,I2067,I19636,I19622,);
nor I_1058 (I20077,I19730,I20012);
nor I_1059 (I19610,I19925,I20077);
nor I_1060 (I19619,I19860,I19995);
nor I_1061 (I19607,I19730,I19995);
not I_1062 (I20163,I2074);
DFFARX1 I_1063 (I34610,I2067,I20163,I20189,);
not I_1064 (I20197,I20189);
nand I_1065 (I20214,I34604,I34598);
and I_1066 (I20231,I20214,I34619);
DFFARX1 I_1067 (I20231,I2067,I20163,I20257,);
DFFARX1 I_1068 (I34616,I2067,I20163,I20274,);
and I_1069 (I20282,I20274,I34613);
nor I_1070 (I20299,I20257,I20282);
DFFARX1 I_1071 (I20299,I2067,I20163,I20131,);
nand I_1072 (I20330,I20274,I34613);
nand I_1073 (I20347,I20197,I20330);
not I_1074 (I20143,I20347);
DFFARX1 I_1075 (I34598,I2067,I20163,I20387,);
DFFARX1 I_1076 (I20387,I2067,I20163,I20152,);
nand I_1077 (I20409,I34601,I34601);
and I_1078 (I20426,I20409,I34622);
DFFARX1 I_1079 (I20426,I2067,I20163,I20452,);
DFFARX1 I_1080 (I20452,I2067,I20163,I20469,);
not I_1081 (I20155,I20469);
not I_1082 (I20491,I20452);
nand I_1083 (I20140,I20491,I20330);
nor I_1084 (I20522,I34607,I34601);
not I_1085 (I20539,I20522);
nor I_1086 (I20556,I20491,I20539);
nor I_1087 (I20573,I20197,I20556);
DFFARX1 I_1088 (I20573,I2067,I20163,I20149,);
nor I_1089 (I20604,I20257,I20539);
nor I_1090 (I20137,I20452,I20604);
nor I_1091 (I20146,I20387,I20522);
nor I_1092 (I20134,I20257,I20522);
not I_1093 (I20690,I2074);
DFFARX1 I_1094 (I75469,I2067,I20690,I20716,);
not I_1095 (I20724,I20716);
nand I_1096 (I20741,I75490,I75484);
and I_1097 (I20758,I20741,I75466);
DFFARX1 I_1098 (I20758,I2067,I20690,I20784,);
DFFARX1 I_1099 (I75469,I2067,I20690,I20801,);
and I_1100 (I20809,I20801,I75478);
nor I_1101 (I20826,I20784,I20809);
DFFARX1 I_1102 (I20826,I2067,I20690,I20658,);
nand I_1103 (I20857,I20801,I75478);
nand I_1104 (I20874,I20724,I20857);
not I_1105 (I20670,I20874);
DFFARX1 I_1106 (I75475,I2067,I20690,I20914,);
DFFARX1 I_1107 (I20914,I2067,I20690,I20679,);
nand I_1108 (I20936,I75481,I75472);
and I_1109 (I20953,I20936,I75466);
DFFARX1 I_1110 (I20953,I2067,I20690,I20979,);
DFFARX1 I_1111 (I20979,I2067,I20690,I20996,);
not I_1112 (I20682,I20996);
not I_1113 (I21018,I20979);
nand I_1114 (I20667,I21018,I20857);
nor I_1115 (I21049,I75487,I75472);
not I_1116 (I21066,I21049);
nor I_1117 (I21083,I21018,I21066);
nor I_1118 (I21100,I20724,I21083);
DFFARX1 I_1119 (I21100,I2067,I20690,I20676,);
nor I_1120 (I21131,I20784,I21066);
nor I_1121 (I20664,I20979,I21131);
nor I_1122 (I20673,I20914,I21049);
nor I_1123 (I20661,I20784,I21049);
not I_1124 (I21217,I2074);
DFFARX1 I_1125 (I25090,I2067,I21217,I21243,);
not I_1126 (I21251,I21243);
nand I_1127 (I21268,I25084,I25078);
and I_1128 (I21285,I21268,I25099);
DFFARX1 I_1129 (I21285,I2067,I21217,I21311,);
DFFARX1 I_1130 (I25096,I2067,I21217,I21328,);
and I_1131 (I21336,I21328,I25093);
nor I_1132 (I21353,I21311,I21336);
DFFARX1 I_1133 (I21353,I2067,I21217,I21185,);
nand I_1134 (I21384,I21328,I25093);
nand I_1135 (I21401,I21251,I21384);
not I_1136 (I21197,I21401);
DFFARX1 I_1137 (I25078,I2067,I21217,I21441,);
DFFARX1 I_1138 (I21441,I2067,I21217,I21206,);
nand I_1139 (I21463,I25081,I25081);
and I_1140 (I21480,I21463,I25102);
DFFARX1 I_1141 (I21480,I2067,I21217,I21506,);
DFFARX1 I_1142 (I21506,I2067,I21217,I21523,);
not I_1143 (I21209,I21523);
not I_1144 (I21545,I21506);
nand I_1145 (I21194,I21545,I21384);
nor I_1146 (I21576,I25087,I25081);
not I_1147 (I21593,I21576);
nor I_1148 (I21610,I21545,I21593);
nor I_1149 (I21627,I21251,I21610);
DFFARX1 I_1150 (I21627,I2067,I21217,I21203,);
nor I_1151 (I21658,I21311,I21593);
nor I_1152 (I21191,I21506,I21658);
nor I_1153 (I21200,I21441,I21576);
nor I_1154 (I21188,I21311,I21576);
not I_1155 (I21744,I2074);
DFFARX1 I_1156 (I178821,I2067,I21744,I21770,);
not I_1157 (I21778,I21770);
nand I_1158 (I21795,I178815,I178836);
and I_1159 (I21812,I21795,I178812);
DFFARX1 I_1160 (I21812,I2067,I21744,I21838,);
DFFARX1 I_1161 (I178833,I2067,I21744,I21855,);
and I_1162 (I21863,I21855,I178830);
nor I_1163 (I21880,I21838,I21863);
DFFARX1 I_1164 (I21880,I2067,I21744,I21712,);
nand I_1165 (I21911,I21855,I178830);
nand I_1166 (I21928,I21778,I21911);
not I_1167 (I21724,I21928);
DFFARX1 I_1168 (I178818,I2067,I21744,I21968,);
DFFARX1 I_1169 (I21968,I2067,I21744,I21733,);
nand I_1170 (I21990,I178827,I178824);
and I_1171 (I22007,I21990,I178809);
DFFARX1 I_1172 (I22007,I2067,I21744,I22033,);
DFFARX1 I_1173 (I22033,I2067,I21744,I22050,);
not I_1174 (I21736,I22050);
not I_1175 (I22072,I22033);
nand I_1176 (I21721,I22072,I21911);
nor I_1177 (I22103,I178809,I178824);
not I_1178 (I22120,I22103);
nor I_1179 (I22137,I22072,I22120);
nor I_1180 (I22154,I21778,I22137);
DFFARX1 I_1181 (I22154,I2067,I21744,I21730,);
nor I_1182 (I22185,I21838,I22120);
nor I_1183 (I21718,I22033,I22185);
nor I_1184 (I21727,I21968,I22103);
nor I_1185 (I21715,I21838,I22103);
not I_1186 (I22271,I2074);
DFFARX1 I_1187 (I102712,I2067,I22271,I22297,);
not I_1188 (I22305,I22297);
nand I_1189 (I22322,I102703,I102721);
and I_1190 (I22339,I22322,I102700);
DFFARX1 I_1191 (I22339,I2067,I22271,I22365,);
DFFARX1 I_1192 (I102703,I2067,I22271,I22382,);
and I_1193 (I22390,I22382,I102706);
nor I_1194 (I22407,I22365,I22390);
DFFARX1 I_1195 (I22407,I2067,I22271,I22239,);
nand I_1196 (I22438,I22382,I102706);
nand I_1197 (I22455,I22305,I22438);
not I_1198 (I22251,I22455);
DFFARX1 I_1199 (I102700,I2067,I22271,I22495,);
DFFARX1 I_1200 (I22495,I2067,I22271,I22260,);
nand I_1201 (I22517,I102718,I102709);
and I_1202 (I22534,I22517,I102724);
DFFARX1 I_1203 (I22534,I2067,I22271,I22560,);
DFFARX1 I_1204 (I22560,I2067,I22271,I22577,);
not I_1205 (I22263,I22577);
not I_1206 (I22599,I22560);
nand I_1207 (I22248,I22599,I22438);
nor I_1208 (I22630,I102715,I102709);
not I_1209 (I22647,I22630);
nor I_1210 (I22664,I22599,I22647);
nor I_1211 (I22681,I22305,I22664);
DFFARX1 I_1212 (I22681,I2067,I22271,I22257,);
nor I_1213 (I22712,I22365,I22647);
nor I_1214 (I22245,I22560,I22712);
nor I_1215 (I22254,I22495,I22630);
nor I_1216 (I22242,I22365,I22630);
not I_1217 (I22798,I2074);
DFFARX1 I_1218 (I43873,I2067,I22798,I22824,);
not I_1219 (I22832,I22824);
nand I_1220 (I22849,I43855,I43870);
and I_1221 (I22866,I22849,I43846);
DFFARX1 I_1222 (I22866,I2067,I22798,I22892,);
DFFARX1 I_1223 (I43849,I2067,I22798,I22909,);
and I_1224 (I22917,I22909,I43864);
nor I_1225 (I22934,I22892,I22917);
DFFARX1 I_1226 (I22934,I2067,I22798,I22766,);
nand I_1227 (I22965,I22909,I43864);
nand I_1228 (I22982,I22832,I22965);
not I_1229 (I22778,I22982);
DFFARX1 I_1230 (I43867,I2067,I22798,I23022,);
DFFARX1 I_1231 (I23022,I2067,I22798,I22787,);
nand I_1232 (I23044,I43846,I43858);
and I_1233 (I23061,I23044,I43852);
DFFARX1 I_1234 (I23061,I2067,I22798,I23087,);
DFFARX1 I_1235 (I23087,I2067,I22798,I23104,);
not I_1236 (I22790,I23104);
not I_1237 (I23126,I23087);
nand I_1238 (I22775,I23126,I22965);
nor I_1239 (I23157,I43861,I43858);
not I_1240 (I23174,I23157);
nor I_1241 (I23191,I23126,I23174);
nor I_1242 (I23208,I22832,I23191);
DFFARX1 I_1243 (I23208,I2067,I22798,I22784,);
nor I_1244 (I23239,I22892,I23174);
nor I_1245 (I22772,I23087,I23239);
nor I_1246 (I22781,I23022,I23157);
nor I_1247 (I22769,I22892,I23157);
not I_1248 (I23328,I2074);
DFFARX1 I_1249 (I1588,I2067,I23328,I23354,);
not I_1250 (I23362,I23354);
DFFARX1 I_1251 (I2044,I2067,I23328,I23388,);
not I_1252 (I23396,I1868);
or I_1253 (I23413,I1532,I1868);
nor I_1254 (I23430,I23388,I1532);
nand I_1255 (I23305,I23396,I23430);
nor I_1256 (I23461,I1660,I1532);
nand I_1257 (I23299,I23461,I23396);
not I_1258 (I23492,I1804);
nand I_1259 (I23509,I23396,I23492);
nor I_1260 (I23526,I1700,I1740);
not I_1261 (I23543,I23526);
nor I_1262 (I23560,I23543,I23509);
nor I_1263 (I23577,I23461,I23560);
DFFARX1 I_1264 (I23577,I2067,I23328,I23314,);
nor I_1265 (I23311,I23526,I23413);
DFFARX1 I_1266 (I23526,I2067,I23328,I23317,);
nor I_1267 (I23636,I23492,I1700);
nor I_1268 (I23653,I23636,I1868);
nor I_1269 (I23670,I1764,I1780);
DFFARX1 I_1270 (I23670,I2067,I23328,I23696,);
nor I_1271 (I23296,I23696,I23653);
DFFARX1 I_1272 (I23696,I2067,I23328,I23727,);
nand I_1273 (I23735,I23727,I1436);
nor I_1274 (I23320,I23362,I23735);
not I_1275 (I23766,I23696);
nand I_1276 (I23783,I23766,I1436);
nor I_1277 (I23800,I23362,I23783);
nor I_1278 (I23302,I23388,I23800);
nor I_1279 (I23831,I1764,I1660);
nor I_1280 (I23848,I23388,I23831);
DFFARX1 I_1281 (I23848,I2067,I23328,I23293,);
and I_1282 (I23308,I23461,I1764);
not I_1283 (I23920,I2074);
DFFARX1 I_1284 (I89418,I2067,I23920,I23946,);
DFFARX1 I_1285 (I23946,I2067,I23920,I23963,);
not I_1286 (I23912,I23963);
not I_1287 (I23985,I23946);
DFFARX1 I_1288 (I89415,I2067,I23920,I24011,);
not I_1289 (I24019,I24011);
and I_1290 (I24036,I23985,I89421);
not I_1291 (I24053,I89406);
nand I_1292 (I24070,I24053,I89421);
not I_1293 (I24087,I89409);
nor I_1294 (I24104,I24087,I89430);
nand I_1295 (I24121,I24104,I89427);
nor I_1296 (I24138,I24121,I24070);
DFFARX1 I_1297 (I24138,I2067,I23920,I23888,);
not I_1298 (I24169,I24121);
not I_1299 (I24186,I89430);
nand I_1300 (I24203,I24186,I89421);
nor I_1301 (I24220,I89430,I89406);
nand I_1302 (I23900,I24036,I24220);
nand I_1303 (I23894,I23985,I89430);
nand I_1304 (I24265,I24087,I89406);
DFFARX1 I_1305 (I24265,I2067,I23920,I23909,);
DFFARX1 I_1306 (I24265,I2067,I23920,I23903,);
not I_1307 (I24310,I89406);
nor I_1308 (I24327,I24310,I89412);
and I_1309 (I24344,I24327,I89424);
or I_1310 (I24361,I24344,I89409);
DFFARX1 I_1311 (I24361,I2067,I23920,I24387,);
nand I_1312 (I24395,I24387,I24053);
nor I_1313 (I23897,I24395,I24203);
nor I_1314 (I23891,I24387,I24019);
DFFARX1 I_1315 (I24387,I2067,I23920,I24449,);
not I_1316 (I24457,I24449);
nor I_1317 (I23906,I24457,I24169);
not I_1318 (I24515,I2074);
DFFARX1 I_1319 (I52278,I2067,I24515,I24541,);
DFFARX1 I_1320 (I24541,I2067,I24515,I24558,);
not I_1321 (I24507,I24558);
not I_1322 (I24580,I24541);
DFFARX1 I_1323 (I52293,I2067,I24515,I24606,);
not I_1324 (I24614,I24606);
and I_1325 (I24631,I24580,I52290);
not I_1326 (I24648,I52278);
nand I_1327 (I24665,I24648,I52290);
not I_1328 (I24682,I52287);
nor I_1329 (I24699,I24682,I52302);
nand I_1330 (I24716,I24699,I52299);
nor I_1331 (I24733,I24716,I24665);
DFFARX1 I_1332 (I24733,I2067,I24515,I24483,);
not I_1333 (I24764,I24716);
not I_1334 (I24781,I52302);
nand I_1335 (I24798,I24781,I52290);
nor I_1336 (I24815,I52302,I52278);
nand I_1337 (I24495,I24631,I24815);
nand I_1338 (I24489,I24580,I52302);
nand I_1339 (I24860,I24682,I52296);
DFFARX1 I_1340 (I24860,I2067,I24515,I24504,);
DFFARX1 I_1341 (I24860,I2067,I24515,I24498,);
not I_1342 (I24905,I52296);
nor I_1343 (I24922,I24905,I52284);
and I_1344 (I24939,I24922,I52305);
or I_1345 (I24956,I24939,I52281);
DFFARX1 I_1346 (I24956,I2067,I24515,I24982,);
nand I_1347 (I24990,I24982,I24648);
nor I_1348 (I24492,I24990,I24798);
nor I_1349 (I24486,I24982,I24614);
DFFARX1 I_1350 (I24982,I2067,I24515,I25044,);
not I_1351 (I25052,I25044);
nor I_1352 (I24501,I25052,I24764);
not I_1353 (I25110,I2074);
DFFARX1 I_1354 (I124271,I2067,I25110,I25136,);
DFFARX1 I_1355 (I25136,I2067,I25110,I25153,);
not I_1356 (I25102,I25153);
not I_1357 (I25175,I25136);
DFFARX1 I_1358 (I124280,I2067,I25110,I25201,);
not I_1359 (I25209,I25201);
and I_1360 (I25226,I25175,I124268);
not I_1361 (I25243,I124259);
nand I_1362 (I25260,I25243,I124268);
not I_1363 (I25277,I124265);
nor I_1364 (I25294,I25277,I124283);
nand I_1365 (I25311,I25294,I124256);
nor I_1366 (I25328,I25311,I25260);
DFFARX1 I_1367 (I25328,I2067,I25110,I25078,);
not I_1368 (I25359,I25311);
not I_1369 (I25376,I124283);
nand I_1370 (I25393,I25376,I124268);
nor I_1371 (I25410,I124283,I124259);
nand I_1372 (I25090,I25226,I25410);
nand I_1373 (I25084,I25175,I124283);
nand I_1374 (I25455,I25277,I124262);
DFFARX1 I_1375 (I25455,I2067,I25110,I25099,);
DFFARX1 I_1376 (I25455,I2067,I25110,I25093,);
not I_1377 (I25500,I124262);
nor I_1378 (I25517,I25500,I124274);
and I_1379 (I25534,I25517,I124256);
or I_1380 (I25551,I25534,I124277);
DFFARX1 I_1381 (I25551,I2067,I25110,I25577,);
nand I_1382 (I25585,I25577,I25243);
nor I_1383 (I25087,I25585,I25393);
nor I_1384 (I25081,I25577,I25209);
DFFARX1 I_1385 (I25577,I2067,I25110,I25639,);
not I_1386 (I25647,I25639);
nor I_1387 (I25096,I25647,I25359);
not I_1388 (I25705,I2074);
DFFARX1 I_1389 (I44373,I2067,I25705,I25731,);
DFFARX1 I_1390 (I25731,I2067,I25705,I25748,);
not I_1391 (I25697,I25748);
not I_1392 (I25770,I25731);
DFFARX1 I_1393 (I44388,I2067,I25705,I25796,);
not I_1394 (I25804,I25796);
and I_1395 (I25821,I25770,I44385);
not I_1396 (I25838,I44373);
nand I_1397 (I25855,I25838,I44385);
not I_1398 (I25872,I44382);
nor I_1399 (I25889,I25872,I44397);
nand I_1400 (I25906,I25889,I44394);
nor I_1401 (I25923,I25906,I25855);
DFFARX1 I_1402 (I25923,I2067,I25705,I25673,);
not I_1403 (I25954,I25906);
not I_1404 (I25971,I44397);
nand I_1405 (I25988,I25971,I44385);
nor I_1406 (I26005,I44397,I44373);
nand I_1407 (I25685,I25821,I26005);
nand I_1408 (I25679,I25770,I44397);
nand I_1409 (I26050,I25872,I44391);
DFFARX1 I_1410 (I26050,I2067,I25705,I25694,);
DFFARX1 I_1411 (I26050,I2067,I25705,I25688,);
not I_1412 (I26095,I44391);
nor I_1413 (I26112,I26095,I44379);
and I_1414 (I26129,I26112,I44400);
or I_1415 (I26146,I26129,I44376);
DFFARX1 I_1416 (I26146,I2067,I25705,I26172,);
nand I_1417 (I26180,I26172,I25838);
nor I_1418 (I25682,I26180,I25988);
nor I_1419 (I25676,I26172,I25804);
DFFARX1 I_1420 (I26172,I2067,I25705,I26234,);
not I_1421 (I26242,I26234);
nor I_1422 (I25691,I26242,I25954);
not I_1423 (I26300,I2074);
DFFARX1 I_1424 (I67857,I2067,I26300,I26326,);
DFFARX1 I_1425 (I26326,I2067,I26300,I26343,);
not I_1426 (I26292,I26343);
not I_1427 (I26365,I26326);
DFFARX1 I_1428 (I67845,I2067,I26300,I26391,);
not I_1429 (I26399,I26391);
and I_1430 (I26416,I26365,I67854);
not I_1431 (I26433,I67851);
nand I_1432 (I26450,I26433,I67854);
not I_1433 (I26467,I67842);
nor I_1434 (I26484,I26467,I67848);
nand I_1435 (I26501,I26484,I67833);
nor I_1436 (I26518,I26501,I26450);
DFFARX1 I_1437 (I26518,I2067,I26300,I26268,);
not I_1438 (I26549,I26501);
not I_1439 (I26566,I67848);
nand I_1440 (I26583,I26566,I67854);
nor I_1441 (I26600,I67848,I67851);
nand I_1442 (I26280,I26416,I26600);
nand I_1443 (I26274,I26365,I67848);
nand I_1444 (I26645,I26467,I67833);
DFFARX1 I_1445 (I26645,I2067,I26300,I26289,);
DFFARX1 I_1446 (I26645,I2067,I26300,I26283,);
not I_1447 (I26690,I67833);
nor I_1448 (I26707,I26690,I67839);
and I_1449 (I26724,I26707,I67836);
or I_1450 (I26741,I26724,I67860);
DFFARX1 I_1451 (I26741,I2067,I26300,I26767,);
nand I_1452 (I26775,I26767,I26433);
nor I_1453 (I26277,I26775,I26583);
nor I_1454 (I26271,I26767,I26399);
DFFARX1 I_1455 (I26767,I2067,I26300,I26829,);
not I_1456 (I26837,I26829);
nor I_1457 (I26286,I26837,I26549);
not I_1458 (I26895,I2074);
DFFARX1 I_1459 (I163495,I2067,I26895,I26921,);
DFFARX1 I_1460 (I26921,I2067,I26895,I26938,);
not I_1461 (I26887,I26938);
not I_1462 (I26960,I26921);
DFFARX1 I_1463 (I163507,I2067,I26895,I26986,);
not I_1464 (I26994,I26986);
and I_1465 (I27011,I26960,I163501);
not I_1466 (I27028,I163513);
nand I_1467 (I27045,I27028,I163501);
not I_1468 (I27062,I163498);
nor I_1469 (I27079,I27062,I163510);
nand I_1470 (I27096,I27079,I163492);
nor I_1471 (I27113,I27096,I27045);
DFFARX1 I_1472 (I27113,I2067,I26895,I26863,);
not I_1473 (I27144,I27096);
not I_1474 (I27161,I163510);
nand I_1475 (I27178,I27161,I163501);
nor I_1476 (I27195,I163510,I163513);
nand I_1477 (I26875,I27011,I27195);
nand I_1478 (I26869,I26960,I163510);
nand I_1479 (I27240,I27062,I163504);
DFFARX1 I_1480 (I27240,I2067,I26895,I26884,);
DFFARX1 I_1481 (I27240,I2067,I26895,I26878,);
not I_1482 (I27285,I163504);
nor I_1483 (I27302,I27285,I163495);
and I_1484 (I27319,I27302,I163492);
or I_1485 (I27336,I27319,I163516);
DFFARX1 I_1486 (I27336,I2067,I26895,I27362,);
nand I_1487 (I27370,I27362,I27028);
nor I_1488 (I26872,I27370,I27178);
nor I_1489 (I26866,I27362,I26994);
DFFARX1 I_1490 (I27362,I2067,I26895,I27424,);
not I_1491 (I27432,I27424);
nor I_1492 (I26881,I27432,I27144);
not I_1493 (I27490,I2074);
DFFARX1 I_1494 (I104967,I2067,I27490,I27516,);
DFFARX1 I_1495 (I27516,I2067,I27490,I27533,);
not I_1496 (I27482,I27533);
not I_1497 (I27555,I27516);
DFFARX1 I_1498 (I104961,I2067,I27490,I27581,);
not I_1499 (I27589,I27581);
and I_1500 (I27606,I27555,I104979);
not I_1501 (I27623,I104967);
nand I_1502 (I27640,I27623,I104979);
not I_1503 (I27657,I104961);
nor I_1504 (I27674,I27657,I104973);
nand I_1505 (I27691,I27674,I104964);
nor I_1506 (I27708,I27691,I27640);
DFFARX1 I_1507 (I27708,I2067,I27490,I27458,);
not I_1508 (I27739,I27691);
not I_1509 (I27756,I104973);
nand I_1510 (I27773,I27756,I104979);
nor I_1511 (I27790,I104973,I104967);
nand I_1512 (I27470,I27606,I27790);
nand I_1513 (I27464,I27555,I104973);
nand I_1514 (I27835,I27657,I104976);
DFFARX1 I_1515 (I27835,I2067,I27490,I27479,);
DFFARX1 I_1516 (I27835,I2067,I27490,I27473,);
not I_1517 (I27880,I104976);
nor I_1518 (I27897,I27880,I104982);
and I_1519 (I27914,I27897,I104964);
or I_1520 (I27931,I27914,I104970);
DFFARX1 I_1521 (I27931,I2067,I27490,I27957,);
nand I_1522 (I27965,I27957,I27623);
nor I_1523 (I27467,I27965,I27773);
nor I_1524 (I27461,I27957,I27589);
DFFARX1 I_1525 (I27957,I2067,I27490,I28019,);
not I_1526 (I28027,I28019);
nor I_1527 (I27476,I28027,I27739);
not I_1528 (I28085,I2074);
DFFARX1 I_1529 (I49116,I2067,I28085,I28111,);
DFFARX1 I_1530 (I28111,I2067,I28085,I28128,);
not I_1531 (I28077,I28128);
not I_1532 (I28150,I28111);
DFFARX1 I_1533 (I49131,I2067,I28085,I28176,);
not I_1534 (I28184,I28176);
and I_1535 (I28201,I28150,I49128);
not I_1536 (I28218,I49116);
nand I_1537 (I28235,I28218,I49128);
not I_1538 (I28252,I49125);
nor I_1539 (I28269,I28252,I49140);
nand I_1540 (I28286,I28269,I49137);
nor I_1541 (I28303,I28286,I28235);
DFFARX1 I_1542 (I28303,I2067,I28085,I28053,);
not I_1543 (I28334,I28286);
not I_1544 (I28351,I49140);
nand I_1545 (I28368,I28351,I49128);
nor I_1546 (I28385,I49140,I49116);
nand I_1547 (I28065,I28201,I28385);
nand I_1548 (I28059,I28150,I49140);
nand I_1549 (I28430,I28252,I49134);
DFFARX1 I_1550 (I28430,I2067,I28085,I28074,);
DFFARX1 I_1551 (I28430,I2067,I28085,I28068,);
not I_1552 (I28475,I49134);
nor I_1553 (I28492,I28475,I49122);
and I_1554 (I28509,I28492,I49143);
or I_1555 (I28526,I28509,I49119);
DFFARX1 I_1556 (I28526,I2067,I28085,I28552,);
nand I_1557 (I28560,I28552,I28218);
nor I_1558 (I28062,I28560,I28368);
nor I_1559 (I28056,I28552,I28184);
DFFARX1 I_1560 (I28552,I2067,I28085,I28614,);
not I_1561 (I28622,I28614);
nor I_1562 (I28071,I28622,I28334);
not I_1563 (I28680,I2074);
DFFARX1 I_1564 (I6980,I2067,I28680,I28706,);
DFFARX1 I_1565 (I28706,I2067,I28680,I28723,);
not I_1566 (I28672,I28723);
not I_1567 (I28745,I28706);
DFFARX1 I_1568 (I6956,I2067,I28680,I28771,);
not I_1569 (I28779,I28771);
and I_1570 (I28796,I28745,I6971);
not I_1571 (I28813,I6959);
nand I_1572 (I28830,I28813,I6971);
not I_1573 (I28847,I6962);
nor I_1574 (I28864,I28847,I6974);
nand I_1575 (I28881,I28864,I6965);
nor I_1576 (I28898,I28881,I28830);
DFFARX1 I_1577 (I28898,I2067,I28680,I28648,);
not I_1578 (I28929,I28881);
not I_1579 (I28946,I6974);
nand I_1580 (I28963,I28946,I6971);
nor I_1581 (I28980,I6974,I6959);
nand I_1582 (I28660,I28796,I28980);
nand I_1583 (I28654,I28745,I6974);
nand I_1584 (I29025,I28847,I6968);
DFFARX1 I_1585 (I29025,I2067,I28680,I28669,);
DFFARX1 I_1586 (I29025,I2067,I28680,I28663,);
not I_1587 (I29070,I6968);
nor I_1588 (I29087,I29070,I6959);
and I_1589 (I29104,I29087,I6956);
or I_1590 (I29121,I29104,I6977);
DFFARX1 I_1591 (I29121,I2067,I28680,I29147,);
nand I_1592 (I29155,I29147,I28813);
nor I_1593 (I28657,I29155,I28963);
nor I_1594 (I28651,I29147,I28779);
DFFARX1 I_1595 (I29147,I2067,I28680,I29209,);
not I_1596 (I29217,I29209);
nor I_1597 (I28666,I29217,I28929);
not I_1598 (I29275,I2074);
DFFARX1 I_1599 (I1396,I2067,I29275,I29301,);
DFFARX1 I_1600 (I29301,I2067,I29275,I29318,);
not I_1601 (I29267,I29318);
not I_1602 (I29340,I29301);
DFFARX1 I_1603 (I1940,I2067,I29275,I29366,);
not I_1604 (I29374,I29366);
and I_1605 (I29391,I29340,I2052);
not I_1606 (I29408,I2060);
nand I_1607 (I29425,I29408,I2052);
not I_1608 (I29442,I2028);
nor I_1609 (I29459,I29442,I1916);
nand I_1610 (I29476,I29459,I1788);
nor I_1611 (I29493,I29476,I29425);
DFFARX1 I_1612 (I29493,I2067,I29275,I29243,);
not I_1613 (I29524,I29476);
not I_1614 (I29541,I1916);
nand I_1615 (I29558,I29541,I2052);
nor I_1616 (I29575,I1916,I2060);
nand I_1617 (I29255,I29391,I29575);
nand I_1618 (I29249,I29340,I1916);
nand I_1619 (I29620,I29442,I1476);
DFFARX1 I_1620 (I29620,I2067,I29275,I29264,);
DFFARX1 I_1621 (I29620,I2067,I29275,I29258,);
not I_1622 (I29665,I1476);
nor I_1623 (I29682,I29665,I1380);
and I_1624 (I29699,I29682,I1580);
or I_1625 (I29716,I29699,I1524);
DFFARX1 I_1626 (I29716,I2067,I29275,I29742,);
nand I_1627 (I29750,I29742,I29408);
nor I_1628 (I29252,I29750,I29558);
nor I_1629 (I29246,I29742,I29374);
DFFARX1 I_1630 (I29742,I2067,I29275,I29804,);
not I_1631 (I29812,I29804);
nor I_1632 (I29261,I29812,I29524);
not I_1633 (I29870,I2074);
DFFARX1 I_1634 (I89996,I2067,I29870,I29896,);
DFFARX1 I_1635 (I29896,I2067,I29870,I29913,);
not I_1636 (I29862,I29913);
not I_1637 (I29935,I29896);
DFFARX1 I_1638 (I89993,I2067,I29870,I29961,);
not I_1639 (I29969,I29961);
and I_1640 (I29986,I29935,I89999);
not I_1641 (I30003,I89984);
nand I_1642 (I30020,I30003,I89999);
not I_1643 (I30037,I89987);
nor I_1644 (I30054,I30037,I90008);
nand I_1645 (I30071,I30054,I90005);
nor I_1646 (I30088,I30071,I30020);
DFFARX1 I_1647 (I30088,I2067,I29870,I29838,);
not I_1648 (I30119,I30071);
not I_1649 (I30136,I90008);
nand I_1650 (I30153,I30136,I89999);
nor I_1651 (I30170,I90008,I89984);
nand I_1652 (I29850,I29986,I30170);
nand I_1653 (I29844,I29935,I90008);
nand I_1654 (I30215,I30037,I89984);
DFFARX1 I_1655 (I30215,I2067,I29870,I29859,);
DFFARX1 I_1656 (I30215,I2067,I29870,I29853,);
not I_1657 (I30260,I89984);
nor I_1658 (I30277,I30260,I89990);
and I_1659 (I30294,I30277,I90002);
or I_1660 (I30311,I30294,I89987);
DFFARX1 I_1661 (I30311,I2067,I29870,I30337,);
nand I_1662 (I30345,I30337,I30003);
nor I_1663 (I29847,I30345,I30153);
nor I_1664 (I29841,I30337,I29969);
DFFARX1 I_1665 (I30337,I2067,I29870,I30399,);
not I_1666 (I30407,I30399);
nor I_1667 (I29856,I30407,I30119);
not I_1668 (I30465,I2074);
DFFARX1 I_1669 (I174665,I2067,I30465,I30491,);
DFFARX1 I_1670 (I30491,I2067,I30465,I30508,);
not I_1671 (I30457,I30508);
not I_1672 (I30530,I30491);
DFFARX1 I_1673 (I174656,I2067,I30465,I30556,);
not I_1674 (I30564,I30556);
and I_1675 (I30581,I30530,I174650);
not I_1676 (I30598,I174644);
nand I_1677 (I30615,I30598,I174650);
not I_1678 (I30632,I174671);
nor I_1679 (I30649,I30632,I174644);
nand I_1680 (I30666,I30649,I174668);
nor I_1681 (I30683,I30666,I30615);
DFFARX1 I_1682 (I30683,I2067,I30465,I30433,);
not I_1683 (I30714,I30666);
not I_1684 (I30731,I174644);
nand I_1685 (I30748,I30731,I174650);
nor I_1686 (I30765,I174644,I174644);
nand I_1687 (I30445,I30581,I30765);
nand I_1688 (I30439,I30530,I174644);
nand I_1689 (I30810,I30632,I174653);
DFFARX1 I_1690 (I30810,I2067,I30465,I30454,);
DFFARX1 I_1691 (I30810,I2067,I30465,I30448,);
not I_1692 (I30855,I174653);
nor I_1693 (I30872,I30855,I174659);
and I_1694 (I30889,I30872,I174662);
or I_1695 (I30906,I30889,I174647);
DFFARX1 I_1696 (I30906,I2067,I30465,I30932,);
nand I_1697 (I30940,I30932,I30598);
nor I_1698 (I30442,I30940,I30748);
nor I_1699 (I30436,I30932,I30564);
DFFARX1 I_1700 (I30932,I2067,I30465,I30994,);
not I_1701 (I31002,I30994);
nor I_1702 (I30451,I31002,I30714);
not I_1703 (I31060,I2074);
DFFARX1 I_1704 (I68401,I2067,I31060,I31086,);
DFFARX1 I_1705 (I31086,I2067,I31060,I31103,);
not I_1706 (I31052,I31103);
not I_1707 (I31125,I31086);
DFFARX1 I_1708 (I68389,I2067,I31060,I31151,);
not I_1709 (I31159,I31151);
and I_1710 (I31176,I31125,I68398);
not I_1711 (I31193,I68395);
nand I_1712 (I31210,I31193,I68398);
not I_1713 (I31227,I68386);
nor I_1714 (I31244,I31227,I68392);
nand I_1715 (I31261,I31244,I68377);
nor I_1716 (I31278,I31261,I31210);
DFFARX1 I_1717 (I31278,I2067,I31060,I31028,);
not I_1718 (I31309,I31261);
not I_1719 (I31326,I68392);
nand I_1720 (I31343,I31326,I68398);
nor I_1721 (I31360,I68392,I68395);
nand I_1722 (I31040,I31176,I31360);
nand I_1723 (I31034,I31125,I68392);
nand I_1724 (I31405,I31227,I68377);
DFFARX1 I_1725 (I31405,I2067,I31060,I31049,);
DFFARX1 I_1726 (I31405,I2067,I31060,I31043,);
not I_1727 (I31450,I68377);
nor I_1728 (I31467,I31450,I68383);
and I_1729 (I31484,I31467,I68380);
or I_1730 (I31501,I31484,I68404);
DFFARX1 I_1731 (I31501,I2067,I31060,I31527,);
nand I_1732 (I31535,I31527,I31193);
nor I_1733 (I31037,I31535,I31343);
nor I_1734 (I31031,I31527,I31159);
DFFARX1 I_1735 (I31527,I2067,I31060,I31589,);
not I_1736 (I31597,I31589);
nor I_1737 (I31046,I31597,I31309);
not I_1738 (I31655,I2074);
DFFARX1 I_1739 (I22775,I2067,I31655,I31681,);
DFFARX1 I_1740 (I31681,I2067,I31655,I31698,);
not I_1741 (I31647,I31698);
not I_1742 (I31720,I31681);
DFFARX1 I_1743 (I22769,I2067,I31655,I31746,);
not I_1744 (I31754,I31746);
and I_1745 (I31771,I31720,I22766);
not I_1746 (I31788,I22787);
nand I_1747 (I31805,I31788,I22766);
not I_1748 (I31822,I22781);
nor I_1749 (I31839,I31822,I22772);
nand I_1750 (I31856,I31839,I22778);
nor I_1751 (I31873,I31856,I31805);
DFFARX1 I_1752 (I31873,I2067,I31655,I31623,);
not I_1753 (I31904,I31856);
not I_1754 (I31921,I22772);
nand I_1755 (I31938,I31921,I22766);
nor I_1756 (I31955,I22772,I22787);
nand I_1757 (I31635,I31771,I31955);
nand I_1758 (I31629,I31720,I22772);
nand I_1759 (I32000,I31822,I22766);
DFFARX1 I_1760 (I32000,I2067,I31655,I31644,);
DFFARX1 I_1761 (I32000,I2067,I31655,I31638,);
not I_1762 (I32045,I22766);
nor I_1763 (I32062,I32045,I22784);
and I_1764 (I32079,I32062,I22790);
or I_1765 (I32096,I32079,I22769);
DFFARX1 I_1766 (I32096,I2067,I31655,I32122,);
nand I_1767 (I32130,I32122,I31788);
nor I_1768 (I31632,I32130,I31938);
nor I_1769 (I31626,I32122,I31754);
DFFARX1 I_1770 (I32122,I2067,I31655,I32184,);
not I_1771 (I32192,I32184);
nor I_1772 (I31641,I32192,I31904);
not I_1773 (I32250,I2074);
DFFARX1 I_1774 (I91730,I2067,I32250,I32276,);
DFFARX1 I_1775 (I32276,I2067,I32250,I32293,);
not I_1776 (I32242,I32293);
not I_1777 (I32315,I32276);
DFFARX1 I_1778 (I91727,I2067,I32250,I32341,);
not I_1779 (I32349,I32341);
and I_1780 (I32366,I32315,I91733);
not I_1781 (I32383,I91718);
nand I_1782 (I32400,I32383,I91733);
not I_1783 (I32417,I91721);
nor I_1784 (I32434,I32417,I91742);
nand I_1785 (I32451,I32434,I91739);
nor I_1786 (I32468,I32451,I32400);
DFFARX1 I_1787 (I32468,I2067,I32250,I32218,);
not I_1788 (I32499,I32451);
not I_1789 (I32516,I91742);
nand I_1790 (I32533,I32516,I91733);
nor I_1791 (I32550,I91742,I91718);
nand I_1792 (I32230,I32366,I32550);
nand I_1793 (I32224,I32315,I91742);
nand I_1794 (I32595,I32417,I91718);
DFFARX1 I_1795 (I32595,I2067,I32250,I32239,);
DFFARX1 I_1796 (I32595,I2067,I32250,I32233,);
not I_1797 (I32640,I91718);
nor I_1798 (I32657,I32640,I91724);
and I_1799 (I32674,I32657,I91736);
or I_1800 (I32691,I32674,I91721);
DFFARX1 I_1801 (I32691,I2067,I32250,I32717,);
nand I_1802 (I32725,I32717,I32383);
nor I_1803 (I32227,I32725,I32533);
nor I_1804 (I32221,I32717,I32349);
DFFARX1 I_1805 (I32717,I2067,I32250,I32779,);
not I_1806 (I32787,I32779);
nor I_1807 (I32236,I32787,I32499);
not I_1808 (I32845,I2074);
DFFARX1 I_1809 (I6453,I2067,I32845,I32871,);
DFFARX1 I_1810 (I32871,I2067,I32845,I32888,);
not I_1811 (I32837,I32888);
not I_1812 (I32910,I32871);
DFFARX1 I_1813 (I6429,I2067,I32845,I32936,);
not I_1814 (I32944,I32936);
and I_1815 (I32961,I32910,I6444);
not I_1816 (I32978,I6432);
nand I_1817 (I32995,I32978,I6444);
not I_1818 (I33012,I6435);
nor I_1819 (I33029,I33012,I6447);
nand I_1820 (I33046,I33029,I6438);
nor I_1821 (I33063,I33046,I32995);
DFFARX1 I_1822 (I33063,I2067,I32845,I32813,);
not I_1823 (I33094,I33046);
not I_1824 (I33111,I6447);
nand I_1825 (I33128,I33111,I6444);
nor I_1826 (I33145,I6447,I6432);
nand I_1827 (I32825,I32961,I33145);
nand I_1828 (I32819,I32910,I6447);
nand I_1829 (I33190,I33012,I6441);
DFFARX1 I_1830 (I33190,I2067,I32845,I32834,);
DFFARX1 I_1831 (I33190,I2067,I32845,I32828,);
not I_1832 (I33235,I6441);
nor I_1833 (I33252,I33235,I6432);
and I_1834 (I33269,I33252,I6429);
or I_1835 (I33286,I33269,I6450);
DFFARX1 I_1836 (I33286,I2067,I32845,I33312,);
nand I_1837 (I33320,I33312,I32978);
nor I_1838 (I32822,I33320,I33128);
nor I_1839 (I32816,I33312,I32944);
DFFARX1 I_1840 (I33312,I2067,I32845,I33374,);
not I_1841 (I33382,I33374);
nor I_1842 (I32831,I33382,I33094);
not I_1843 (I33440,I2074);
DFFARX1 I_1844 (I104440,I2067,I33440,I33466,);
DFFARX1 I_1845 (I33466,I2067,I33440,I33483,);
not I_1846 (I33432,I33483);
not I_1847 (I33505,I33466);
DFFARX1 I_1848 (I104434,I2067,I33440,I33531,);
not I_1849 (I33539,I33531);
and I_1850 (I33556,I33505,I104452);
not I_1851 (I33573,I104440);
nand I_1852 (I33590,I33573,I104452);
not I_1853 (I33607,I104434);
nor I_1854 (I33624,I33607,I104446);
nand I_1855 (I33641,I33624,I104437);
nor I_1856 (I33658,I33641,I33590);
DFFARX1 I_1857 (I33658,I2067,I33440,I33408,);
not I_1858 (I33689,I33641);
not I_1859 (I33706,I104446);
nand I_1860 (I33723,I33706,I104452);
nor I_1861 (I33740,I104446,I104440);
nand I_1862 (I33420,I33556,I33740);
nand I_1863 (I33414,I33505,I104446);
nand I_1864 (I33785,I33607,I104449);
DFFARX1 I_1865 (I33785,I2067,I33440,I33429,);
DFFARX1 I_1866 (I33785,I2067,I33440,I33423,);
not I_1867 (I33830,I104449);
nor I_1868 (I33847,I33830,I104455);
and I_1869 (I33864,I33847,I104437);
or I_1870 (I33881,I33864,I104443);
DFFARX1 I_1871 (I33881,I2067,I33440,I33907,);
nand I_1872 (I33915,I33907,I33573);
nor I_1873 (I33417,I33915,I33723);
nor I_1874 (I33411,I33907,I33539);
DFFARX1 I_1875 (I33907,I2067,I33440,I33969,);
not I_1876 (I33977,I33969);
nor I_1877 (I33426,I33977,I33689);
not I_1878 (I34035,I2074);
DFFARX1 I_1879 (I132317,I2067,I34035,I34061,);
DFFARX1 I_1880 (I34061,I2067,I34035,I34078,);
not I_1881 (I34027,I34078);
not I_1882 (I34100,I34061);
DFFARX1 I_1883 (I132326,I2067,I34035,I34126,);
not I_1884 (I34134,I34126);
and I_1885 (I34151,I34100,I132320);
not I_1886 (I34168,I132314);
nand I_1887 (I34185,I34168,I132320);
not I_1888 (I34202,I132329);
nor I_1889 (I34219,I34202,I132317);
nand I_1890 (I34236,I34219,I132323);
nor I_1891 (I34253,I34236,I34185);
DFFARX1 I_1892 (I34253,I2067,I34035,I34003,);
not I_1893 (I34284,I34236);
not I_1894 (I34301,I132317);
nand I_1895 (I34318,I34301,I132320);
nor I_1896 (I34335,I132317,I132314);
nand I_1897 (I34015,I34151,I34335);
nand I_1898 (I34009,I34100,I132317);
nand I_1899 (I34380,I34202,I132320);
DFFARX1 I_1900 (I34380,I2067,I34035,I34024,);
DFFARX1 I_1901 (I34380,I2067,I34035,I34018,);
not I_1902 (I34425,I132320);
nor I_1903 (I34442,I34425,I132335);
and I_1904 (I34459,I34442,I132332);
or I_1905 (I34476,I34459,I132314);
DFFARX1 I_1906 (I34476,I2067,I34035,I34502,);
nand I_1907 (I34510,I34502,I34168);
nor I_1908 (I34012,I34510,I34318);
nor I_1909 (I34006,I34502,I34134);
DFFARX1 I_1910 (I34502,I2067,I34035,I34564,);
not I_1911 (I34572,I34564);
nor I_1912 (I34021,I34572,I34284);
not I_1913 (I34630,I2074);
DFFARX1 I_1914 (I103290,I2067,I34630,I34656,);
DFFARX1 I_1915 (I34656,I2067,I34630,I34673,);
not I_1916 (I34622,I34673);
not I_1917 (I34695,I34656);
DFFARX1 I_1918 (I103287,I2067,I34630,I34721,);
not I_1919 (I34729,I34721);
and I_1920 (I34746,I34695,I103293);
not I_1921 (I34763,I103278);
nand I_1922 (I34780,I34763,I103293);
not I_1923 (I34797,I103281);
nor I_1924 (I34814,I34797,I103302);
nand I_1925 (I34831,I34814,I103299);
nor I_1926 (I34848,I34831,I34780);
DFFARX1 I_1927 (I34848,I2067,I34630,I34598,);
not I_1928 (I34879,I34831);
not I_1929 (I34896,I103302);
nand I_1930 (I34913,I34896,I103293);
nor I_1931 (I34930,I103302,I103278);
nand I_1932 (I34610,I34746,I34930);
nand I_1933 (I34604,I34695,I103302);
nand I_1934 (I34975,I34797,I103278);
DFFARX1 I_1935 (I34975,I2067,I34630,I34619,);
DFFARX1 I_1936 (I34975,I2067,I34630,I34613,);
not I_1937 (I35020,I103278);
nor I_1938 (I35037,I35020,I103284);
and I_1939 (I35054,I35037,I103296);
or I_1940 (I35071,I35054,I103281);
DFFARX1 I_1941 (I35071,I2067,I34630,I35097,);
nand I_1942 (I35105,I35097,I34763);
nor I_1943 (I34607,I35105,I34913);
nor I_1944 (I34601,I35097,I34729);
DFFARX1 I_1945 (I35097,I2067,I34630,I35159,);
not I_1946 (I35167,I35159);
nor I_1947 (I34616,I35167,I34879);
not I_1948 (I35225,I2074);
DFFARX1 I_1949 (I101556,I2067,I35225,I35251,);
DFFARX1 I_1950 (I35251,I2067,I35225,I35268,);
not I_1951 (I35217,I35268);
not I_1952 (I35290,I35251);
DFFARX1 I_1953 (I101553,I2067,I35225,I35316,);
not I_1954 (I35324,I35316);
and I_1955 (I35341,I35290,I101559);
not I_1956 (I35358,I101544);
nand I_1957 (I35375,I35358,I101559);
not I_1958 (I35392,I101547);
nor I_1959 (I35409,I35392,I101568);
nand I_1960 (I35426,I35409,I101565);
nor I_1961 (I35443,I35426,I35375);
DFFARX1 I_1962 (I35443,I2067,I35225,I35193,);
not I_1963 (I35474,I35426);
not I_1964 (I35491,I101568);
nand I_1965 (I35508,I35491,I101559);
nor I_1966 (I35525,I101568,I101544);
nand I_1967 (I35205,I35341,I35525);
nand I_1968 (I35199,I35290,I101568);
nand I_1969 (I35570,I35392,I101544);
DFFARX1 I_1970 (I35570,I2067,I35225,I35214,);
DFFARX1 I_1971 (I35570,I2067,I35225,I35208,);
not I_1972 (I35615,I101544);
nor I_1973 (I35632,I35615,I101550);
and I_1974 (I35649,I35632,I101562);
or I_1975 (I35666,I35649,I101547);
DFFARX1 I_1976 (I35666,I2067,I35225,I35692,);
nand I_1977 (I35700,I35692,I35358);
nor I_1978 (I35202,I35700,I35508);
nor I_1979 (I35196,I35692,I35324);
DFFARX1 I_1980 (I35692,I2067,I35225,I35754,);
not I_1981 (I35762,I35754);
nor I_1982 (I35211,I35762,I35474);
not I_1983 (I35820,I2074);
DFFARX1 I_1984 (I125563,I2067,I35820,I35846,);
DFFARX1 I_1985 (I35846,I2067,I35820,I35863,);
not I_1986 (I35812,I35863);
not I_1987 (I35885,I35846);
DFFARX1 I_1988 (I125572,I2067,I35820,I35911,);
not I_1989 (I35919,I35911);
and I_1990 (I35936,I35885,I125560);
not I_1991 (I35953,I125551);
nand I_1992 (I35970,I35953,I125560);
not I_1993 (I35987,I125557);
nor I_1994 (I36004,I35987,I125575);
nand I_1995 (I36021,I36004,I125548);
nor I_1996 (I36038,I36021,I35970);
DFFARX1 I_1997 (I36038,I2067,I35820,I35788,);
not I_1998 (I36069,I36021);
not I_1999 (I36086,I125575);
nand I_2000 (I36103,I36086,I125560);
nor I_2001 (I36120,I125575,I125551);
nand I_2002 (I35800,I35936,I36120);
nand I_2003 (I35794,I35885,I125575);
nand I_2004 (I36165,I35987,I125554);
DFFARX1 I_2005 (I36165,I2067,I35820,I35809,);
DFFARX1 I_2006 (I36165,I2067,I35820,I35803,);
not I_2007 (I36210,I125554);
nor I_2008 (I36227,I36210,I125566);
and I_2009 (I36244,I36227,I125548);
or I_2010 (I36261,I36244,I125569);
DFFARX1 I_2011 (I36261,I2067,I35820,I36287,);
nand I_2012 (I36295,I36287,I35953);
nor I_2013 (I35797,I36295,I36103);
nor I_2014 (I35791,I36287,I35919);
DFFARX1 I_2015 (I36287,I2067,I35820,I36349,);
not I_2016 (I36357,I36349);
nor I_2017 (I35806,I36357,I36069);
not I_2018 (I36415,I2074);
DFFARX1 I_2019 (I47535,I2067,I36415,I36441,);
DFFARX1 I_2020 (I36441,I2067,I36415,I36458,);
not I_2021 (I36407,I36458);
not I_2022 (I36480,I36441);
DFFARX1 I_2023 (I47550,I2067,I36415,I36506,);
not I_2024 (I36514,I36506);
and I_2025 (I36531,I36480,I47547);
not I_2026 (I36548,I47535);
nand I_2027 (I36565,I36548,I47547);
not I_2028 (I36582,I47544);
nor I_2029 (I36599,I36582,I47559);
nand I_2030 (I36616,I36599,I47556);
nor I_2031 (I36633,I36616,I36565);
DFFARX1 I_2032 (I36633,I2067,I36415,I36383,);
not I_2033 (I36664,I36616);
not I_2034 (I36681,I47559);
nand I_2035 (I36698,I36681,I47547);
nor I_2036 (I36715,I47559,I47535);
nand I_2037 (I36395,I36531,I36715);
nand I_2038 (I36389,I36480,I47559);
nand I_2039 (I36760,I36582,I47553);
DFFARX1 I_2040 (I36760,I2067,I36415,I36404,);
DFFARX1 I_2041 (I36760,I2067,I36415,I36398,);
not I_2042 (I36805,I47553);
nor I_2043 (I36822,I36805,I47541);
and I_2044 (I36839,I36822,I47562);
or I_2045 (I36856,I36839,I47538);
DFFARX1 I_2046 (I36856,I2067,I36415,I36882,);
nand I_2047 (I36890,I36882,I36548);
nor I_2048 (I36392,I36890,I36698);
nor I_2049 (I36386,I36882,I36514);
DFFARX1 I_2050 (I36882,I2067,I36415,I36944,);
not I_2051 (I36952,I36944);
nor I_2052 (I36401,I36952,I36664);
not I_2053 (I37010,I2074);
DFFARX1 I_2054 (I22248,I2067,I37010,I37036,);
DFFARX1 I_2055 (I37036,I2067,I37010,I37053,);
not I_2056 (I37002,I37053);
not I_2057 (I37075,I37036);
DFFARX1 I_2058 (I22242,I2067,I37010,I37101,);
not I_2059 (I37109,I37101);
and I_2060 (I37126,I37075,I22239);
not I_2061 (I37143,I22260);
nand I_2062 (I37160,I37143,I22239);
not I_2063 (I37177,I22254);
nor I_2064 (I37194,I37177,I22245);
nand I_2065 (I37211,I37194,I22251);
nor I_2066 (I37228,I37211,I37160);
DFFARX1 I_2067 (I37228,I2067,I37010,I36978,);
not I_2068 (I37259,I37211);
not I_2069 (I37276,I22245);
nand I_2070 (I37293,I37276,I22239);
nor I_2071 (I37310,I22245,I22260);
nand I_2072 (I36990,I37126,I37310);
nand I_2073 (I36984,I37075,I22245);
nand I_2074 (I37355,I37177,I22239);
DFFARX1 I_2075 (I37355,I2067,I37010,I36999,);
DFFARX1 I_2076 (I37355,I2067,I37010,I36993,);
not I_2077 (I37400,I22239);
nor I_2078 (I37417,I37400,I22257);
and I_2079 (I37434,I37417,I22263);
or I_2080 (I37451,I37434,I22242);
DFFARX1 I_2081 (I37451,I2067,I37010,I37477,);
nand I_2082 (I37485,I37477,I37143);
nor I_2083 (I36987,I37485,I37293);
nor I_2084 (I36981,I37477,I37109);
DFFARX1 I_2085 (I37477,I2067,I37010,I37539,);
not I_2086 (I37547,I37539);
nor I_2087 (I36996,I37547,I37259);
not I_2088 (I37605,I2074);
DFFARX1 I_2089 (I173475,I2067,I37605,I37631,);
DFFARX1 I_2090 (I37631,I2067,I37605,I37648,);
not I_2091 (I37597,I37648);
not I_2092 (I37670,I37631);
DFFARX1 I_2093 (I173466,I2067,I37605,I37696,);
not I_2094 (I37704,I37696);
and I_2095 (I37721,I37670,I173460);
not I_2096 (I37738,I173454);
nand I_2097 (I37755,I37738,I173460);
not I_2098 (I37772,I173481);
nor I_2099 (I37789,I37772,I173454);
nand I_2100 (I37806,I37789,I173478);
nor I_2101 (I37823,I37806,I37755);
DFFARX1 I_2102 (I37823,I2067,I37605,I37573,);
not I_2103 (I37854,I37806);
not I_2104 (I37871,I173454);
nand I_2105 (I37888,I37871,I173460);
nor I_2106 (I37905,I173454,I173454);
nand I_2107 (I37585,I37721,I37905);
nand I_2108 (I37579,I37670,I173454);
nand I_2109 (I37950,I37772,I173463);
DFFARX1 I_2110 (I37950,I2067,I37605,I37594,);
DFFARX1 I_2111 (I37950,I2067,I37605,I37588,);
not I_2112 (I37995,I173463);
nor I_2113 (I38012,I37995,I173469);
and I_2114 (I38029,I38012,I173472);
or I_2115 (I38046,I38029,I173457);
DFFARX1 I_2116 (I38046,I2067,I37605,I38072,);
nand I_2117 (I38080,I38072,I37738);
nor I_2118 (I37582,I38080,I37888);
nor I_2119 (I37576,I38072,I37704);
DFFARX1 I_2120 (I38072,I2067,I37605,I38134,);
not I_2121 (I38142,I38134);
nor I_2122 (I37591,I38142,I37854);
not I_2123 (I38200,I2074);
DFFARX1 I_2124 (I175855,I2067,I38200,I38226,);
DFFARX1 I_2125 (I38226,I2067,I38200,I38243,);
not I_2126 (I38192,I38243);
not I_2127 (I38265,I38226);
DFFARX1 I_2128 (I175846,I2067,I38200,I38291,);
not I_2129 (I38299,I38291);
and I_2130 (I38316,I38265,I175840);
not I_2131 (I38333,I175834);
nand I_2132 (I38350,I38333,I175840);
not I_2133 (I38367,I175861);
nor I_2134 (I38384,I38367,I175834);
nand I_2135 (I38401,I38384,I175858);
nor I_2136 (I38418,I38401,I38350);
DFFARX1 I_2137 (I38418,I2067,I38200,I38168,);
not I_2138 (I38449,I38401);
not I_2139 (I38466,I175834);
nand I_2140 (I38483,I38466,I175840);
nor I_2141 (I38500,I175834,I175834);
nand I_2142 (I38180,I38316,I38500);
nand I_2143 (I38174,I38265,I175834);
nand I_2144 (I38545,I38367,I175843);
DFFARX1 I_2145 (I38545,I2067,I38200,I38189,);
DFFARX1 I_2146 (I38545,I2067,I38200,I38183,);
not I_2147 (I38590,I175843);
nor I_2148 (I38607,I38590,I175849);
and I_2149 (I38624,I38607,I175852);
or I_2150 (I38641,I38624,I175837);
DFFARX1 I_2151 (I38641,I2067,I38200,I38667,);
nand I_2152 (I38675,I38667,I38333);
nor I_2153 (I38177,I38675,I38483);
nor I_2154 (I38171,I38667,I38299);
DFFARX1 I_2155 (I38667,I2067,I38200,I38729,);
not I_2156 (I38737,I38729);
nor I_2157 (I38186,I38737,I38449);
not I_2158 (I38795,I2074);
DFFARX1 I_2159 (I19613,I2067,I38795,I38821,);
DFFARX1 I_2160 (I38821,I2067,I38795,I38838,);
not I_2161 (I38787,I38838);
not I_2162 (I38860,I38821);
DFFARX1 I_2163 (I19607,I2067,I38795,I38886,);
not I_2164 (I38894,I38886);
and I_2165 (I38911,I38860,I19604);
not I_2166 (I38928,I19625);
nand I_2167 (I38945,I38928,I19604);
not I_2168 (I38962,I19619);
nor I_2169 (I38979,I38962,I19610);
nand I_2170 (I38996,I38979,I19616);
nor I_2171 (I39013,I38996,I38945);
DFFARX1 I_2172 (I39013,I2067,I38795,I38763,);
not I_2173 (I39044,I38996);
not I_2174 (I39061,I19610);
nand I_2175 (I39078,I39061,I19604);
nor I_2176 (I39095,I19610,I19625);
nand I_2177 (I38775,I38911,I39095);
nand I_2178 (I38769,I38860,I19610);
nand I_2179 (I39140,I38962,I19604);
DFFARX1 I_2180 (I39140,I2067,I38795,I38784,);
DFFARX1 I_2181 (I39140,I2067,I38795,I38778,);
not I_2182 (I39185,I19604);
nor I_2183 (I39202,I39185,I19622);
and I_2184 (I39219,I39202,I19628);
or I_2185 (I39236,I39219,I19607);
DFFARX1 I_2186 (I39236,I2067,I38795,I39262,);
nand I_2187 (I39270,I39262,I38928);
nor I_2188 (I38772,I39270,I39078);
nor I_2189 (I38766,I39262,I38894);
DFFARX1 I_2190 (I39262,I2067,I38795,I39324,);
not I_2191 (I39332,I39324);
nor I_2192 (I38781,I39332,I39044);
not I_2193 (I39390,I2074);
DFFARX1 I_2194 (I17505,I2067,I39390,I39416,);
DFFARX1 I_2195 (I39416,I2067,I39390,I39433,);
not I_2196 (I39382,I39433);
not I_2197 (I39455,I39416);
DFFARX1 I_2198 (I17499,I2067,I39390,I39481,);
not I_2199 (I39489,I39481);
and I_2200 (I39506,I39455,I17496);
not I_2201 (I39523,I17517);
nand I_2202 (I39540,I39523,I17496);
not I_2203 (I39557,I17511);
nor I_2204 (I39574,I39557,I17502);
nand I_2205 (I39591,I39574,I17508);
nor I_2206 (I39608,I39591,I39540);
DFFARX1 I_2207 (I39608,I2067,I39390,I39358,);
not I_2208 (I39639,I39591);
not I_2209 (I39656,I17502);
nand I_2210 (I39673,I39656,I17496);
nor I_2211 (I39690,I17502,I17517);
nand I_2212 (I39370,I39506,I39690);
nand I_2213 (I39364,I39455,I17502);
nand I_2214 (I39735,I39557,I17496);
DFFARX1 I_2215 (I39735,I2067,I39390,I39379,);
DFFARX1 I_2216 (I39735,I2067,I39390,I39373,);
not I_2217 (I39780,I17496);
nor I_2218 (I39797,I39780,I17514);
and I_2219 (I39814,I39797,I17520);
or I_2220 (I39831,I39814,I17499);
DFFARX1 I_2221 (I39831,I2067,I39390,I39857,);
nand I_2222 (I39865,I39857,I39523);
nor I_2223 (I39367,I39865,I39673);
nor I_2224 (I39361,I39857,I39489);
DFFARX1 I_2225 (I39857,I2067,I39390,I39919,);
not I_2226 (I39927,I39919);
nor I_2227 (I39376,I39927,I39639);
not I_2228 (I39985,I2074);
DFFARX1 I_2229 (I15924,I2067,I39985,I40011,);
DFFARX1 I_2230 (I40011,I2067,I39985,I40028,);
not I_2231 (I39977,I40028);
not I_2232 (I40050,I40011);
DFFARX1 I_2233 (I15918,I2067,I39985,I40076,);
not I_2234 (I40084,I40076);
and I_2235 (I40101,I40050,I15915);
not I_2236 (I40118,I15936);
nand I_2237 (I40135,I40118,I15915);
not I_2238 (I40152,I15930);
nor I_2239 (I40169,I40152,I15921);
nand I_2240 (I40186,I40169,I15927);
nor I_2241 (I40203,I40186,I40135);
DFFARX1 I_2242 (I40203,I2067,I39985,I39953,);
not I_2243 (I40234,I40186);
not I_2244 (I40251,I15921);
nand I_2245 (I40268,I40251,I15915);
nor I_2246 (I40285,I15921,I15936);
nand I_2247 (I39965,I40101,I40285);
nand I_2248 (I39959,I40050,I15921);
nand I_2249 (I40330,I40152,I15915);
DFFARX1 I_2250 (I40330,I2067,I39985,I39974,);
DFFARX1 I_2251 (I40330,I2067,I39985,I39968,);
not I_2252 (I40375,I15915);
nor I_2253 (I40392,I40375,I15933);
and I_2254 (I40409,I40392,I15939);
or I_2255 (I40426,I40409,I15918);
DFFARX1 I_2256 (I40426,I2067,I39985,I40452,);
nand I_2257 (I40460,I40452,I40118);
nor I_2258 (I39962,I40460,I40268);
nor I_2259 (I39956,I40452,I40084);
DFFARX1 I_2260 (I40452,I2067,I39985,I40514,);
not I_2261 (I40522,I40514);
nor I_2262 (I39971,I40522,I40234);
not I_2263 (I40580,I2074);
DFFARX1 I_2264 (I42792,I2067,I40580,I40606,);
DFFARX1 I_2265 (I40606,I2067,I40580,I40623,);
not I_2266 (I40572,I40623);
not I_2267 (I40645,I40606);
DFFARX1 I_2268 (I42807,I2067,I40580,I40671,);
not I_2269 (I40679,I40671);
and I_2270 (I40696,I40645,I42804);
not I_2271 (I40713,I42792);
nand I_2272 (I40730,I40713,I42804);
not I_2273 (I40747,I42801);
nor I_2274 (I40764,I40747,I42816);
nand I_2275 (I40781,I40764,I42813);
nor I_2276 (I40798,I40781,I40730);
DFFARX1 I_2277 (I40798,I2067,I40580,I40548,);
not I_2278 (I40829,I40781);
not I_2279 (I40846,I42816);
nand I_2280 (I40863,I40846,I42804);
nor I_2281 (I40880,I42816,I42792);
nand I_2282 (I40560,I40696,I40880);
nand I_2283 (I40554,I40645,I42816);
nand I_2284 (I40925,I40747,I42810);
DFFARX1 I_2285 (I40925,I2067,I40580,I40569,);
DFFARX1 I_2286 (I40925,I2067,I40580,I40563,);
not I_2287 (I40970,I42810);
nor I_2288 (I40987,I40970,I42798);
and I_2289 (I41004,I40987,I42819);
or I_2290 (I41021,I41004,I42795);
DFFARX1 I_2291 (I41021,I2067,I40580,I41047,);
nand I_2292 (I41055,I41047,I40713);
nor I_2293 (I40557,I41055,I40863);
nor I_2294 (I40551,I41047,I40679);
DFFARX1 I_2295 (I41047,I2067,I40580,I41109,);
not I_2296 (I41117,I41109);
nor I_2297 (I40566,I41117,I40829);
not I_2298 (I41175,I2074);
DFFARX1 I_2299 (I152408,I2067,I41175,I41201,);
DFFARX1 I_2300 (I41201,I2067,I41175,I41218,);
not I_2301 (I41167,I41218);
not I_2302 (I41240,I41201);
DFFARX1 I_2303 (I152408,I2067,I41175,I41266,);
not I_2304 (I41274,I41266);
and I_2305 (I41291,I41240,I152411);
not I_2306 (I41308,I152423);
nand I_2307 (I41325,I41308,I152411);
not I_2308 (I41342,I152429);
nor I_2309 (I41359,I41342,I152420);
nand I_2310 (I41376,I41359,I152426);
nor I_2311 (I41393,I41376,I41325);
DFFARX1 I_2312 (I41393,I2067,I41175,I41143,);
not I_2313 (I41424,I41376);
not I_2314 (I41441,I152420);
nand I_2315 (I41458,I41441,I152411);
nor I_2316 (I41475,I152420,I152423);
nand I_2317 (I41155,I41291,I41475);
nand I_2318 (I41149,I41240,I152420);
nand I_2319 (I41520,I41342,I152417);
DFFARX1 I_2320 (I41520,I2067,I41175,I41164,);
DFFARX1 I_2321 (I41520,I2067,I41175,I41158,);
not I_2322 (I41565,I152417);
nor I_2323 (I41582,I41565,I152414);
and I_2324 (I41599,I41582,I152432);
or I_2325 (I41616,I41599,I152411);
DFFARX1 I_2326 (I41616,I2067,I41175,I41642,);
nand I_2327 (I41650,I41642,I41308);
nor I_2328 (I41152,I41650,I41458);
nor I_2329 (I41146,I41642,I41274);
DFFARX1 I_2330 (I41642,I2067,I41175,I41704,);
not I_2331 (I41712,I41704);
nor I_2332 (I41161,I41712,I41424);
not I_2333 (I41773,I2074);
DFFARX1 I_2334 (I25673,I2067,I41773,I41799,);
nand I_2335 (I41807,I25673,I25679);
and I_2336 (I41824,I41807,I25697);
DFFARX1 I_2337 (I41824,I2067,I41773,I41850,);
nor I_2338 (I41741,I41850,I41799);
not I_2339 (I41872,I41850);
DFFARX1 I_2340 (I25685,I2067,I41773,I41898,);
nand I_2341 (I41906,I41898,I25682);
not I_2342 (I41923,I41906);
DFFARX1 I_2343 (I41923,I2067,I41773,I41949,);
not I_2344 (I41765,I41949);
nor I_2345 (I41971,I41799,I41906);
nor I_2346 (I41747,I41850,I41971);
DFFARX1 I_2347 (I25691,I2067,I41773,I42011,);
DFFARX1 I_2348 (I42011,I2067,I41773,I42028,);
not I_2349 (I42036,I42028);
not I_2350 (I42053,I42011);
nand I_2351 (I41750,I42053,I41872);
nand I_2352 (I42084,I25676,I25676);
and I_2353 (I42101,I42084,I25688);
DFFARX1 I_2354 (I42101,I2067,I41773,I42127,);
nor I_2355 (I42135,I42127,I41799);
DFFARX1 I_2356 (I42135,I2067,I41773,I41738,);
DFFARX1 I_2357 (I42127,I2067,I41773,I41756,);
nor I_2358 (I42180,I25694,I25676);
not I_2359 (I42197,I42180);
nor I_2360 (I41759,I42036,I42197);
nand I_2361 (I41744,I42053,I42197);
nor I_2362 (I41753,I41799,I42180);
DFFARX1 I_2363 (I42180,I2067,I41773,I41762,);
not I_2364 (I42300,I2074);
DFFARX1 I_2365 (I147784,I2067,I42300,I42326,);
nand I_2366 (I42334,I147799,I147784);
and I_2367 (I42351,I42334,I147802);
DFFARX1 I_2368 (I42351,I2067,I42300,I42377,);
nor I_2369 (I42268,I42377,I42326);
not I_2370 (I42399,I42377);
DFFARX1 I_2371 (I147808,I2067,I42300,I42425,);
nand I_2372 (I42433,I42425,I147790);
not I_2373 (I42450,I42433);
DFFARX1 I_2374 (I42450,I2067,I42300,I42476,);
not I_2375 (I42292,I42476);
nor I_2376 (I42498,I42326,I42433);
nor I_2377 (I42274,I42377,I42498);
DFFARX1 I_2378 (I147787,I2067,I42300,I42538,);
DFFARX1 I_2379 (I42538,I2067,I42300,I42555,);
not I_2380 (I42563,I42555);
not I_2381 (I42580,I42538);
nand I_2382 (I42277,I42580,I42399);
nand I_2383 (I42611,I147787,I147793);
and I_2384 (I42628,I42611,I147805);
DFFARX1 I_2385 (I42628,I2067,I42300,I42654,);
nor I_2386 (I42662,I42654,I42326);
DFFARX1 I_2387 (I42662,I2067,I42300,I42265,);
DFFARX1 I_2388 (I42654,I2067,I42300,I42283,);
nor I_2389 (I42707,I147796,I147793);
not I_2390 (I42724,I42707);
nor I_2391 (I42286,I42563,I42724);
nand I_2392 (I42271,I42580,I42724);
nor I_2393 (I42280,I42326,I42707);
DFFARX1 I_2394 (I42707,I2067,I42300,I42289,);
not I_2395 (I42827,I2074);
DFFARX1 I_2396 (I39953,I2067,I42827,I42853,);
nand I_2397 (I42861,I39953,I39959);
and I_2398 (I42878,I42861,I39977);
DFFARX1 I_2399 (I42878,I2067,I42827,I42904,);
nor I_2400 (I42795,I42904,I42853);
not I_2401 (I42926,I42904);
DFFARX1 I_2402 (I39965,I2067,I42827,I42952,);
nand I_2403 (I42960,I42952,I39962);
not I_2404 (I42977,I42960);
DFFARX1 I_2405 (I42977,I2067,I42827,I43003,);
not I_2406 (I42819,I43003);
nor I_2407 (I43025,I42853,I42960);
nor I_2408 (I42801,I42904,I43025);
DFFARX1 I_2409 (I39971,I2067,I42827,I43065,);
DFFARX1 I_2410 (I43065,I2067,I42827,I43082,);
not I_2411 (I43090,I43082);
not I_2412 (I43107,I43065);
nand I_2413 (I42804,I43107,I42926);
nand I_2414 (I43138,I39956,I39956);
and I_2415 (I43155,I43138,I39968);
DFFARX1 I_2416 (I43155,I2067,I42827,I43181,);
nor I_2417 (I43189,I43181,I42853);
DFFARX1 I_2418 (I43189,I2067,I42827,I42792,);
DFFARX1 I_2419 (I43181,I2067,I42827,I42810,);
nor I_2420 (I43234,I39974,I39956);
not I_2421 (I43251,I43234);
nor I_2422 (I42813,I43090,I43251);
nand I_2423 (I42798,I43107,I43251);
nor I_2424 (I42807,I42853,I43234);
DFFARX1 I_2425 (I43234,I2067,I42827,I42816,);
not I_2426 (I43354,I2074);
DFFARX1 I_2427 (I97510,I2067,I43354,I43380,);
nand I_2428 (I43388,I97501,I97516);
and I_2429 (I43405,I43388,I97522);
DFFARX1 I_2430 (I43405,I2067,I43354,I43431,);
nor I_2431 (I43322,I43431,I43380);
not I_2432 (I43453,I43431);
DFFARX1 I_2433 (I97507,I2067,I43354,I43479,);
nand I_2434 (I43487,I43479,I97501);
not I_2435 (I43504,I43487);
DFFARX1 I_2436 (I43504,I2067,I43354,I43530,);
not I_2437 (I43346,I43530);
nor I_2438 (I43552,I43380,I43487);
nor I_2439 (I43328,I43431,I43552);
DFFARX1 I_2440 (I97504,I2067,I43354,I43592,);
DFFARX1 I_2441 (I43592,I2067,I43354,I43609,);
not I_2442 (I43617,I43609);
not I_2443 (I43634,I43592);
nand I_2444 (I43331,I43634,I43453);
nand I_2445 (I43665,I97498,I97513);
and I_2446 (I43682,I43665,I97498);
DFFARX1 I_2447 (I43682,I2067,I43354,I43708,);
nor I_2448 (I43716,I43708,I43380);
DFFARX1 I_2449 (I43716,I2067,I43354,I43319,);
DFFARX1 I_2450 (I43708,I2067,I43354,I43337,);
nor I_2451 (I43761,I97519,I97513);
not I_2452 (I43778,I43761);
nor I_2453 (I43340,I43617,I43778);
nand I_2454 (I43325,I43634,I43778);
nor I_2455 (I43334,I43380,I43761);
DFFARX1 I_2456 (I43761,I2067,I43354,I43343,);
not I_2457 (I43881,I2074);
DFFARX1 I_2458 (I140270,I2067,I43881,I43907,);
nand I_2459 (I43915,I140285,I140270);
and I_2460 (I43932,I43915,I140288);
DFFARX1 I_2461 (I43932,I2067,I43881,I43958,);
nor I_2462 (I43849,I43958,I43907);
not I_2463 (I43980,I43958);
DFFARX1 I_2464 (I140294,I2067,I43881,I44006,);
nand I_2465 (I44014,I44006,I140276);
not I_2466 (I44031,I44014);
DFFARX1 I_2467 (I44031,I2067,I43881,I44057,);
not I_2468 (I43873,I44057);
nor I_2469 (I44079,I43907,I44014);
nor I_2470 (I43855,I43958,I44079);
DFFARX1 I_2471 (I140273,I2067,I43881,I44119,);
DFFARX1 I_2472 (I44119,I2067,I43881,I44136,);
not I_2473 (I44144,I44136);
not I_2474 (I44161,I44119);
nand I_2475 (I43858,I44161,I43980);
nand I_2476 (I44192,I140273,I140279);
and I_2477 (I44209,I44192,I140291);
DFFARX1 I_2478 (I44209,I2067,I43881,I44235,);
nor I_2479 (I44243,I44235,I43907);
DFFARX1 I_2480 (I44243,I2067,I43881,I43846,);
DFFARX1 I_2481 (I44235,I2067,I43881,I43864,);
nor I_2482 (I44288,I140282,I140279);
not I_2483 (I44305,I44288);
nor I_2484 (I43867,I44144,I44305);
nand I_2485 (I43852,I44161,I44305);
nor I_2486 (I43861,I43907,I44288);
DFFARX1 I_2487 (I44288,I2067,I43881,I43870,);
not I_2488 (I44408,I2074);
DFFARX1 I_2489 (I115215,I2067,I44408,I44434,);
nand I_2490 (I44442,I115212,I115230);
and I_2491 (I44459,I44442,I115221);
DFFARX1 I_2492 (I44459,I2067,I44408,I44485,);
nor I_2493 (I44376,I44485,I44434);
not I_2494 (I44507,I44485);
DFFARX1 I_2495 (I115236,I2067,I44408,I44533,);
nand I_2496 (I44541,I44533,I115218);
not I_2497 (I44558,I44541);
DFFARX1 I_2498 (I44558,I2067,I44408,I44584,);
not I_2499 (I44400,I44584);
nor I_2500 (I44606,I44434,I44541);
nor I_2501 (I44382,I44485,I44606);
DFFARX1 I_2502 (I115224,I2067,I44408,I44646,);
DFFARX1 I_2503 (I44646,I2067,I44408,I44663,);
not I_2504 (I44671,I44663);
not I_2505 (I44688,I44646);
nand I_2506 (I44385,I44688,I44507);
nand I_2507 (I44719,I115212,I115239);
and I_2508 (I44736,I44719,I115227);
DFFARX1 I_2509 (I44736,I2067,I44408,I44762,);
nor I_2510 (I44770,I44762,I44434);
DFFARX1 I_2511 (I44770,I2067,I44408,I44373,);
DFFARX1 I_2512 (I44762,I2067,I44408,I44391,);
nor I_2513 (I44815,I115233,I115239);
not I_2514 (I44832,I44815);
nor I_2515 (I44394,I44671,I44832);
nand I_2516 (I44379,I44688,I44832);
nor I_2517 (I44388,I44434,I44815);
DFFARX1 I_2518 (I44815,I2067,I44408,I44397,);
not I_2519 (I44935,I2074);
DFFARX1 I_2520 (I145472,I2067,I44935,I44961,);
nand I_2521 (I44969,I145487,I145472);
and I_2522 (I44986,I44969,I145490);
DFFARX1 I_2523 (I44986,I2067,I44935,I45012,);
nor I_2524 (I44903,I45012,I44961);
not I_2525 (I45034,I45012);
DFFARX1 I_2526 (I145496,I2067,I44935,I45060,);
nand I_2527 (I45068,I45060,I145478);
not I_2528 (I45085,I45068);
DFFARX1 I_2529 (I45085,I2067,I44935,I45111,);
not I_2530 (I44927,I45111);
nor I_2531 (I45133,I44961,I45068);
nor I_2532 (I44909,I45012,I45133);
DFFARX1 I_2533 (I145475,I2067,I44935,I45173,);
DFFARX1 I_2534 (I45173,I2067,I44935,I45190,);
not I_2535 (I45198,I45190);
not I_2536 (I45215,I45173);
nand I_2537 (I44912,I45215,I45034);
nand I_2538 (I45246,I145475,I145481);
and I_2539 (I45263,I45246,I145493);
DFFARX1 I_2540 (I45263,I2067,I44935,I45289,);
nor I_2541 (I45297,I45289,I44961);
DFFARX1 I_2542 (I45297,I2067,I44935,I44900,);
DFFARX1 I_2543 (I45289,I2067,I44935,I44918,);
nor I_2544 (I45342,I145484,I145481);
not I_2545 (I45359,I45342);
nor I_2546 (I44921,I45198,I45359);
nand I_2547 (I44906,I45215,I45359);
nor I_2548 (I44915,I44961,I45342);
DFFARX1 I_2549 (I45342,I2067,I44935,I44924,);
not I_2550 (I45462,I2074);
DFFARX1 I_2551 (I10121,I2067,I45462,I45488,);
nand I_2552 (I45496,I10133,I10142);
and I_2553 (I45513,I45496,I10121);
DFFARX1 I_2554 (I45513,I2067,I45462,I45539,);
nor I_2555 (I45430,I45539,I45488);
not I_2556 (I45561,I45539);
DFFARX1 I_2557 (I10136,I2067,I45462,I45587,);
nand I_2558 (I45595,I45587,I10124);
not I_2559 (I45612,I45595);
DFFARX1 I_2560 (I45612,I2067,I45462,I45638,);
not I_2561 (I45454,I45638);
nor I_2562 (I45660,I45488,I45595);
nor I_2563 (I45436,I45539,I45660);
DFFARX1 I_2564 (I10127,I2067,I45462,I45700,);
DFFARX1 I_2565 (I45700,I2067,I45462,I45717,);
not I_2566 (I45725,I45717);
not I_2567 (I45742,I45700);
nand I_2568 (I45439,I45742,I45561);
nand I_2569 (I45773,I10118,I10118);
and I_2570 (I45790,I45773,I10130);
DFFARX1 I_2571 (I45790,I2067,I45462,I45816,);
nor I_2572 (I45824,I45816,I45488);
DFFARX1 I_2573 (I45824,I2067,I45462,I45427,);
DFFARX1 I_2574 (I45816,I2067,I45462,I45445,);
nor I_2575 (I45869,I10139,I10118);
not I_2576 (I45886,I45869);
nor I_2577 (I45448,I45725,I45886);
nand I_2578 (I45433,I45742,I45886);
nor I_2579 (I45442,I45488,I45869);
DFFARX1 I_2580 (I45869,I2067,I45462,I45451,);
not I_2581 (I45989,I2074);
DFFARX1 I_2582 (I164663,I2067,I45989,I46015,);
nand I_2583 (I46023,I164660,I164651);
and I_2584 (I46040,I46023,I164648);
DFFARX1 I_2585 (I46040,I2067,I45989,I46066,);
nor I_2586 (I45957,I46066,I46015);
not I_2587 (I46088,I46066);
DFFARX1 I_2588 (I164657,I2067,I45989,I46114,);
nand I_2589 (I46122,I46114,I164666);
not I_2590 (I46139,I46122);
DFFARX1 I_2591 (I46139,I2067,I45989,I46165,);
not I_2592 (I45981,I46165);
nor I_2593 (I46187,I46015,I46122);
nor I_2594 (I45963,I46066,I46187);
DFFARX1 I_2595 (I164669,I2067,I45989,I46227,);
DFFARX1 I_2596 (I46227,I2067,I45989,I46244,);
not I_2597 (I46252,I46244);
not I_2598 (I46269,I46227);
nand I_2599 (I45966,I46269,I46088);
nand I_2600 (I46300,I164648,I164654);
and I_2601 (I46317,I46300,I164672);
DFFARX1 I_2602 (I46317,I2067,I45989,I46343,);
nor I_2603 (I46351,I46343,I46015);
DFFARX1 I_2604 (I46351,I2067,I45989,I45954,);
DFFARX1 I_2605 (I46343,I2067,I45989,I45972,);
nor I_2606 (I46396,I164651,I164654);
not I_2607 (I46413,I46396);
nor I_2608 (I45975,I46252,I46413);
nand I_2609 (I45960,I46269,I46413);
nor I_2610 (I45969,I46015,I46396);
DFFARX1 I_2611 (I46396,I2067,I45989,I45978,);
not I_2612 (I46516,I2074);
DFFARX1 I_2613 (I144316,I2067,I46516,I46542,);
nand I_2614 (I46550,I144331,I144316);
and I_2615 (I46567,I46550,I144334);
DFFARX1 I_2616 (I46567,I2067,I46516,I46593,);
nor I_2617 (I46484,I46593,I46542);
not I_2618 (I46615,I46593);
DFFARX1 I_2619 (I144340,I2067,I46516,I46641,);
nand I_2620 (I46649,I46641,I144322);
not I_2621 (I46666,I46649);
DFFARX1 I_2622 (I46666,I2067,I46516,I46692,);
not I_2623 (I46508,I46692);
nor I_2624 (I46714,I46542,I46649);
nor I_2625 (I46490,I46593,I46714);
DFFARX1 I_2626 (I144319,I2067,I46516,I46754,);
DFFARX1 I_2627 (I46754,I2067,I46516,I46771,);
not I_2628 (I46779,I46771);
not I_2629 (I46796,I46754);
nand I_2630 (I46493,I46796,I46615);
nand I_2631 (I46827,I144319,I144325);
and I_2632 (I46844,I46827,I144337);
DFFARX1 I_2633 (I46844,I2067,I46516,I46870,);
nor I_2634 (I46878,I46870,I46542);
DFFARX1 I_2635 (I46878,I2067,I46516,I46481,);
DFFARX1 I_2636 (I46870,I2067,I46516,I46499,);
nor I_2637 (I46923,I144328,I144325);
not I_2638 (I46940,I46923);
nor I_2639 (I46502,I46779,I46940);
nand I_2640 (I46487,I46796,I46940);
nor I_2641 (I46496,I46542,I46923);
DFFARX1 I_2642 (I46923,I2067,I46516,I46505,);
not I_2643 (I47043,I2074);
DFFARX1 I_2644 (I156812,I2067,I47043,I47069,);
nand I_2645 (I47077,I156794,I156818);
and I_2646 (I47094,I47077,I156809);
DFFARX1 I_2647 (I47094,I2067,I47043,I47120,);
nor I_2648 (I47011,I47120,I47069);
not I_2649 (I47142,I47120);
DFFARX1 I_2650 (I156815,I2067,I47043,I47168,);
nand I_2651 (I47176,I47168,I156803);
not I_2652 (I47193,I47176);
DFFARX1 I_2653 (I47193,I2067,I47043,I47219,);
not I_2654 (I47035,I47219);
nor I_2655 (I47241,I47069,I47176);
nor I_2656 (I47017,I47120,I47241);
DFFARX1 I_2657 (I156794,I2067,I47043,I47281,);
DFFARX1 I_2658 (I47281,I2067,I47043,I47298,);
not I_2659 (I47306,I47298);
not I_2660 (I47323,I47281);
nand I_2661 (I47020,I47323,I47142);
nand I_2662 (I47354,I156800,I156797);
and I_2663 (I47371,I47354,I156806);
DFFARX1 I_2664 (I47371,I2067,I47043,I47397,);
nor I_2665 (I47405,I47397,I47069);
DFFARX1 I_2666 (I47405,I2067,I47043,I47008,);
DFFARX1 I_2667 (I47397,I2067,I47043,I47026,);
nor I_2668 (I47450,I156797,I156797);
not I_2669 (I47467,I47450);
nor I_2670 (I47029,I47306,I47467);
nand I_2671 (I47014,I47323,I47467);
nor I_2672 (I47023,I47069,I47450);
DFFARX1 I_2673 (I47450,I2067,I47043,I47032,);
not I_2674 (I47570,I2074);
DFFARX1 I_2675 (I27458,I2067,I47570,I47596,);
nand I_2676 (I47604,I27458,I27464);
and I_2677 (I47621,I47604,I27482);
DFFARX1 I_2678 (I47621,I2067,I47570,I47647,);
nor I_2679 (I47538,I47647,I47596);
not I_2680 (I47669,I47647);
DFFARX1 I_2681 (I27470,I2067,I47570,I47695,);
nand I_2682 (I47703,I47695,I27467);
not I_2683 (I47720,I47703);
DFFARX1 I_2684 (I47720,I2067,I47570,I47746,);
not I_2685 (I47562,I47746);
nor I_2686 (I47768,I47596,I47703);
nor I_2687 (I47544,I47647,I47768);
DFFARX1 I_2688 (I27476,I2067,I47570,I47808,);
DFFARX1 I_2689 (I47808,I2067,I47570,I47825,);
not I_2690 (I47833,I47825);
not I_2691 (I47850,I47808);
nand I_2692 (I47547,I47850,I47669);
nand I_2693 (I47881,I27461,I27461);
and I_2694 (I47898,I47881,I27473);
DFFARX1 I_2695 (I47898,I2067,I47570,I47924,);
nor I_2696 (I47932,I47924,I47596);
DFFARX1 I_2697 (I47932,I2067,I47570,I47535,);
DFFARX1 I_2698 (I47924,I2067,I47570,I47553,);
nor I_2699 (I47977,I27479,I27461);
not I_2700 (I47994,I47977);
nor I_2701 (I47556,I47833,I47994);
nand I_2702 (I47541,I47850,I47994);
nor I_2703 (I47550,I47596,I47977);
DFFARX1 I_2704 (I47977,I2067,I47570,I47559,);
not I_2705 (I48097,I2074);
DFFARX1 I_2706 (I162929,I2067,I48097,I48123,);
nand I_2707 (I48131,I162926,I162917);
and I_2708 (I48148,I48131,I162914);
DFFARX1 I_2709 (I48148,I2067,I48097,I48174,);
nor I_2710 (I48065,I48174,I48123);
not I_2711 (I48196,I48174);
DFFARX1 I_2712 (I162923,I2067,I48097,I48222,);
nand I_2713 (I48230,I48222,I162932);
not I_2714 (I48247,I48230);
DFFARX1 I_2715 (I48247,I2067,I48097,I48273,);
not I_2716 (I48089,I48273);
nor I_2717 (I48295,I48123,I48230);
nor I_2718 (I48071,I48174,I48295);
DFFARX1 I_2719 (I162935,I2067,I48097,I48335,);
DFFARX1 I_2720 (I48335,I2067,I48097,I48352,);
not I_2721 (I48360,I48352);
not I_2722 (I48377,I48335);
nand I_2723 (I48074,I48377,I48196);
nand I_2724 (I48408,I162914,I162920);
and I_2725 (I48425,I48408,I162938);
DFFARX1 I_2726 (I48425,I2067,I48097,I48451,);
nor I_2727 (I48459,I48451,I48123);
DFFARX1 I_2728 (I48459,I2067,I48097,I48062,);
DFFARX1 I_2729 (I48451,I2067,I48097,I48080,);
nor I_2730 (I48504,I162917,I162920);
not I_2731 (I48521,I48504);
nor I_2732 (I48083,I48360,I48521);
nand I_2733 (I48068,I48377,I48521);
nor I_2734 (I48077,I48123,I48504);
DFFARX1 I_2735 (I48504,I2067,I48097,I48086,);
not I_2736 (I48624,I2074);
DFFARX1 I_2737 (I149518,I2067,I48624,I48650,);
nand I_2738 (I48658,I149533,I149518);
and I_2739 (I48675,I48658,I149536);
DFFARX1 I_2740 (I48675,I2067,I48624,I48701,);
nor I_2741 (I48592,I48701,I48650);
not I_2742 (I48723,I48701);
DFFARX1 I_2743 (I149542,I2067,I48624,I48749,);
nand I_2744 (I48757,I48749,I149524);
not I_2745 (I48774,I48757);
DFFARX1 I_2746 (I48774,I2067,I48624,I48800,);
not I_2747 (I48616,I48800);
nor I_2748 (I48822,I48650,I48757);
nor I_2749 (I48598,I48701,I48822);
DFFARX1 I_2750 (I149521,I2067,I48624,I48862,);
DFFARX1 I_2751 (I48862,I2067,I48624,I48879,);
not I_2752 (I48887,I48879);
not I_2753 (I48904,I48862);
nand I_2754 (I48601,I48904,I48723);
nand I_2755 (I48935,I149521,I149527);
and I_2756 (I48952,I48935,I149539);
DFFARX1 I_2757 (I48952,I2067,I48624,I48978,);
nor I_2758 (I48986,I48978,I48650);
DFFARX1 I_2759 (I48986,I2067,I48624,I48589,);
DFFARX1 I_2760 (I48978,I2067,I48624,I48607,);
nor I_2761 (I49031,I149530,I149527);
not I_2762 (I49048,I49031);
nor I_2763 (I48610,I48887,I49048);
nand I_2764 (I48595,I48904,I49048);
nor I_2765 (I48604,I48650,I49031);
DFFARX1 I_2766 (I49031,I2067,I48624,I48613,);
not I_2767 (I49151,I2074);
DFFARX1 I_2768 (I130634,I2067,I49151,I49177,);
nand I_2769 (I49185,I130631,I130634);
and I_2770 (I49202,I49185,I130643);
DFFARX1 I_2771 (I49202,I2067,I49151,I49228,);
nor I_2772 (I49119,I49228,I49177);
not I_2773 (I49250,I49228);
DFFARX1 I_2774 (I130631,I2067,I49151,I49276,);
nand I_2775 (I49284,I49276,I130649);
not I_2776 (I49301,I49284);
DFFARX1 I_2777 (I49301,I2067,I49151,I49327,);
not I_2778 (I49143,I49327);
nor I_2779 (I49349,I49177,I49284);
nor I_2780 (I49125,I49228,I49349);
DFFARX1 I_2781 (I130637,I2067,I49151,I49389,);
DFFARX1 I_2782 (I49389,I2067,I49151,I49406,);
not I_2783 (I49414,I49406);
not I_2784 (I49431,I49389);
nand I_2785 (I49128,I49431,I49250);
nand I_2786 (I49462,I130646,I130652);
and I_2787 (I49479,I49462,I130637);
DFFARX1 I_2788 (I49479,I2067,I49151,I49505,);
nor I_2789 (I49513,I49505,I49177);
DFFARX1 I_2790 (I49513,I2067,I49151,I49116,);
DFFARX1 I_2791 (I49505,I2067,I49151,I49134,);
nor I_2792 (I49558,I130640,I130652);
not I_2793 (I49575,I49558);
nor I_2794 (I49137,I49414,I49575);
nand I_2795 (I49122,I49431,I49575);
nor I_2796 (I49131,I49177,I49558);
DFFARX1 I_2797 (I49558,I2067,I49151,I49140,);
not I_2798 (I49678,I2074);
DFFARX1 I_2799 (I108653,I2067,I49678,I49704,);
nand I_2800 (I49712,I108656,I108650);
and I_2801 (I49729,I49712,I108662);
DFFARX1 I_2802 (I49729,I2067,I49678,I49755,);
nor I_2803 (I49646,I49755,I49704);
not I_2804 (I49777,I49755);
DFFARX1 I_2805 (I108665,I2067,I49678,I49803,);
nand I_2806 (I49811,I49803,I108656);
not I_2807 (I49828,I49811);
DFFARX1 I_2808 (I49828,I2067,I49678,I49854,);
not I_2809 (I49670,I49854);
nor I_2810 (I49876,I49704,I49811);
nor I_2811 (I49652,I49755,I49876);
DFFARX1 I_2812 (I108668,I2067,I49678,I49916,);
DFFARX1 I_2813 (I49916,I2067,I49678,I49933,);
not I_2814 (I49941,I49933);
not I_2815 (I49958,I49916);
nand I_2816 (I49655,I49958,I49777);
nand I_2817 (I49989,I108650,I108659);
and I_2818 (I50006,I49989,I108653);
DFFARX1 I_2819 (I50006,I2067,I49678,I50032,);
nor I_2820 (I50040,I50032,I49704);
DFFARX1 I_2821 (I50040,I2067,I49678,I49643,);
DFFARX1 I_2822 (I50032,I2067,I49678,I49661,);
nor I_2823 (I50085,I108671,I108659);
not I_2824 (I50102,I50085);
nor I_2825 (I49664,I49941,I50102);
nand I_2826 (I49649,I49958,I50102);
nor I_2827 (I49658,I49704,I50085);
DFFARX1 I_2828 (I50085,I2067,I49678,I49667,);
not I_2829 (I50205,I2074);
DFFARX1 I_2830 (I171690,I2067,I50205,I50231,);
nand I_2831 (I50239,I171669,I171669);
and I_2832 (I50256,I50239,I171696);
DFFARX1 I_2833 (I50256,I2067,I50205,I50282,);
nor I_2834 (I50173,I50282,I50231);
not I_2835 (I50304,I50282);
DFFARX1 I_2836 (I171684,I2067,I50205,I50330,);
nand I_2837 (I50338,I50330,I171687);
not I_2838 (I50355,I50338);
DFFARX1 I_2839 (I50355,I2067,I50205,I50381,);
not I_2840 (I50197,I50381);
nor I_2841 (I50403,I50231,I50338);
nor I_2842 (I50179,I50282,I50403);
DFFARX1 I_2843 (I171678,I2067,I50205,I50443,);
DFFARX1 I_2844 (I50443,I2067,I50205,I50460,);
not I_2845 (I50468,I50460);
not I_2846 (I50485,I50443);
nand I_2847 (I50182,I50485,I50304);
nand I_2848 (I50516,I171675,I171672);
and I_2849 (I50533,I50516,I171693);
DFFARX1 I_2850 (I50533,I2067,I50205,I50559,);
nor I_2851 (I50567,I50559,I50231);
DFFARX1 I_2852 (I50567,I2067,I50205,I50170,);
DFFARX1 I_2853 (I50559,I2067,I50205,I50188,);
nor I_2854 (I50612,I171681,I171672);
not I_2855 (I50629,I50612);
nor I_2856 (I50191,I50468,I50629);
nand I_2857 (I50176,I50485,I50629);
nor I_2858 (I50185,I50231,I50612);
DFFARX1 I_2859 (I50612,I2067,I50205,I50194,);
not I_2860 (I50732,I2074);
DFFARX1 I_2861 (I109707,I2067,I50732,I50758,);
nand I_2862 (I50766,I109710,I109704);
and I_2863 (I50783,I50766,I109716);
DFFARX1 I_2864 (I50783,I2067,I50732,I50809,);
nor I_2865 (I50700,I50809,I50758);
not I_2866 (I50831,I50809);
DFFARX1 I_2867 (I109719,I2067,I50732,I50857,);
nand I_2868 (I50865,I50857,I109710);
not I_2869 (I50882,I50865);
DFFARX1 I_2870 (I50882,I2067,I50732,I50908,);
not I_2871 (I50724,I50908);
nor I_2872 (I50930,I50758,I50865);
nor I_2873 (I50706,I50809,I50930);
DFFARX1 I_2874 (I109722,I2067,I50732,I50970,);
DFFARX1 I_2875 (I50970,I2067,I50732,I50987,);
not I_2876 (I50995,I50987);
not I_2877 (I51012,I50970);
nand I_2878 (I50709,I51012,I50831);
nand I_2879 (I51043,I109704,I109713);
and I_2880 (I51060,I51043,I109707);
DFFARX1 I_2881 (I51060,I2067,I50732,I51086,);
nor I_2882 (I51094,I51086,I50758);
DFFARX1 I_2883 (I51094,I2067,I50732,I50697,);
DFFARX1 I_2884 (I51086,I2067,I50732,I50715,);
nor I_2885 (I51139,I109725,I109713);
not I_2886 (I51156,I51139);
nor I_2887 (I50718,I50995,I51156);
nand I_2888 (I50703,I51012,I51156);
nor I_2889 (I50712,I50758,I51139);
DFFARX1 I_2890 (I51139,I2067,I50732,I50721,);
not I_2891 (I51259,I2074);
DFFARX1 I_2892 (I28053,I2067,I51259,I51285,);
nand I_2893 (I51293,I28053,I28059);
and I_2894 (I51310,I51293,I28077);
DFFARX1 I_2895 (I51310,I2067,I51259,I51336,);
nor I_2896 (I51227,I51336,I51285);
not I_2897 (I51358,I51336);
DFFARX1 I_2898 (I28065,I2067,I51259,I51384,);
nand I_2899 (I51392,I51384,I28062);
not I_2900 (I51409,I51392);
DFFARX1 I_2901 (I51409,I2067,I51259,I51435,);
not I_2902 (I51251,I51435);
nor I_2903 (I51457,I51285,I51392);
nor I_2904 (I51233,I51336,I51457);
DFFARX1 I_2905 (I28071,I2067,I51259,I51497,);
DFFARX1 I_2906 (I51497,I2067,I51259,I51514,);
not I_2907 (I51522,I51514);
not I_2908 (I51539,I51497);
nand I_2909 (I51236,I51539,I51358);
nand I_2910 (I51570,I28056,I28056);
and I_2911 (I51587,I51570,I28068);
DFFARX1 I_2912 (I51587,I2067,I51259,I51613,);
nor I_2913 (I51621,I51613,I51285);
DFFARX1 I_2914 (I51621,I2067,I51259,I51224,);
DFFARX1 I_2915 (I51613,I2067,I51259,I51242,);
nor I_2916 (I51666,I28074,I28056);
not I_2917 (I51683,I51666);
nor I_2918 (I51245,I51522,I51683);
nand I_2919 (I51230,I51539,I51683);
nor I_2920 (I51239,I51285,I51666);
DFFARX1 I_2921 (I51666,I2067,I51259,I51248,);
not I_2922 (I51786,I2074);
DFFARX1 I_2923 (I84219,I2067,I51786,I51812,);
nand I_2924 (I51820,I84204,I84207);
and I_2925 (I51837,I51820,I84222);
DFFARX1 I_2926 (I51837,I2067,I51786,I51863,);
nor I_2927 (I51754,I51863,I51812);
not I_2928 (I51885,I51863);
DFFARX1 I_2929 (I84216,I2067,I51786,I51911,);
nand I_2930 (I51919,I51911,I84207);
not I_2931 (I51936,I51919);
DFFARX1 I_2932 (I51936,I2067,I51786,I51962,);
not I_2933 (I51778,I51962);
nor I_2934 (I51984,I51812,I51919);
nor I_2935 (I51760,I51863,I51984);
DFFARX1 I_2936 (I84213,I2067,I51786,I52024,);
DFFARX1 I_2937 (I52024,I2067,I51786,I52041,);
not I_2938 (I52049,I52041);
not I_2939 (I52066,I52024);
nand I_2940 (I51763,I52066,I51885);
nand I_2941 (I52097,I84228,I84204);
and I_2942 (I52114,I52097,I84225);
DFFARX1 I_2943 (I52114,I2067,I51786,I52140,);
nor I_2944 (I52148,I52140,I51812);
DFFARX1 I_2945 (I52148,I2067,I51786,I51751,);
DFFARX1 I_2946 (I52140,I2067,I51786,I51769,);
nor I_2947 (I52193,I84210,I84204);
not I_2948 (I52210,I52193);
nor I_2949 (I51772,I52049,I52210);
nand I_2950 (I51757,I52066,I52210);
nor I_2951 (I51766,I51812,I52193);
DFFARX1 I_2952 (I52193,I2067,I51786,I51775,);
not I_2953 (I52313,I2074);
DFFARX1 I_2954 (I113923,I2067,I52313,I52339,);
nand I_2955 (I52347,I113920,I113938);
and I_2956 (I52364,I52347,I113929);
DFFARX1 I_2957 (I52364,I2067,I52313,I52390,);
nor I_2958 (I52281,I52390,I52339);
not I_2959 (I52412,I52390);
DFFARX1 I_2960 (I113944,I2067,I52313,I52438,);
nand I_2961 (I52446,I52438,I113926);
not I_2962 (I52463,I52446);
DFFARX1 I_2963 (I52463,I2067,I52313,I52489,);
not I_2964 (I52305,I52489);
nor I_2965 (I52511,I52339,I52446);
nor I_2966 (I52287,I52390,I52511);
DFFARX1 I_2967 (I113932,I2067,I52313,I52551,);
DFFARX1 I_2968 (I52551,I2067,I52313,I52568,);
not I_2969 (I52576,I52568);
not I_2970 (I52593,I52551);
nand I_2971 (I52290,I52593,I52412);
nand I_2972 (I52624,I113920,I113947);
and I_2973 (I52641,I52624,I113935);
DFFARX1 I_2974 (I52641,I2067,I52313,I52667,);
nor I_2975 (I52675,I52667,I52339);
DFFARX1 I_2976 (I52675,I2067,I52313,I52278,);
DFFARX1 I_2977 (I52667,I2067,I52313,I52296,);
nor I_2978 (I52720,I113941,I113947);
not I_2979 (I52737,I52720);
nor I_2980 (I52299,I52576,I52737);
nand I_2981 (I52284,I52593,I52737);
nor I_2982 (I52293,I52339,I52720);
DFFARX1 I_2983 (I52720,I2067,I52313,I52302,);
not I_2984 (I52840,I2074);
DFFARX1 I_2985 (I106545,I2067,I52840,I52866,);
nand I_2986 (I52874,I106548,I106542);
and I_2987 (I52891,I52874,I106554);
DFFARX1 I_2988 (I52891,I2067,I52840,I52917,);
nor I_2989 (I52808,I52917,I52866);
not I_2990 (I52939,I52917);
DFFARX1 I_2991 (I106557,I2067,I52840,I52965,);
nand I_2992 (I52973,I52965,I106548);
not I_2993 (I52990,I52973);
DFFARX1 I_2994 (I52990,I2067,I52840,I53016,);
not I_2995 (I52832,I53016);
nor I_2996 (I53038,I52866,I52973);
nor I_2997 (I52814,I52917,I53038);
DFFARX1 I_2998 (I106560,I2067,I52840,I53078,);
DFFARX1 I_2999 (I53078,I2067,I52840,I53095,);
not I_3000 (I53103,I53095);
not I_3001 (I53120,I53078);
nand I_3002 (I52817,I53120,I52939);
nand I_3003 (I53151,I106542,I106551);
and I_3004 (I53168,I53151,I106545);
DFFARX1 I_3005 (I53168,I2067,I52840,I53194,);
nor I_3006 (I53202,I53194,I52866);
DFFARX1 I_3007 (I53202,I2067,I52840,I52805,);
DFFARX1 I_3008 (I53194,I2067,I52840,I52823,);
nor I_3009 (I53247,I106563,I106551);
not I_3010 (I53264,I53247);
nor I_3011 (I52826,I53103,I53264);
nand I_3012 (I52811,I53120,I53264);
nor I_3013 (I52820,I52866,I53247);
DFFARX1 I_3014 (I53247,I2067,I52840,I52829,);
not I_3015 (I53367,I2074);
DFFARX1 I_3016 (I165819,I2067,I53367,I53393,);
nand I_3017 (I53401,I165816,I165807);
and I_3018 (I53418,I53401,I165804);
DFFARX1 I_3019 (I53418,I2067,I53367,I53444,);
nor I_3020 (I53335,I53444,I53393);
not I_3021 (I53466,I53444);
DFFARX1 I_3022 (I165813,I2067,I53367,I53492,);
nand I_3023 (I53500,I53492,I165822);
not I_3024 (I53517,I53500);
DFFARX1 I_3025 (I53517,I2067,I53367,I53543,);
not I_3026 (I53359,I53543);
nor I_3027 (I53565,I53393,I53500);
nor I_3028 (I53341,I53444,I53565);
DFFARX1 I_3029 (I165825,I2067,I53367,I53605,);
DFFARX1 I_3030 (I53605,I2067,I53367,I53622,);
not I_3031 (I53630,I53622);
not I_3032 (I53647,I53605);
nand I_3033 (I53344,I53647,I53466);
nand I_3034 (I53678,I165804,I165810);
and I_3035 (I53695,I53678,I165828);
DFFARX1 I_3036 (I53695,I2067,I53367,I53721,);
nor I_3037 (I53729,I53721,I53393);
DFFARX1 I_3038 (I53729,I2067,I53367,I53332,);
DFFARX1 I_3039 (I53721,I2067,I53367,I53350,);
nor I_3040 (I53774,I165807,I165810);
not I_3041 (I53791,I53774);
nor I_3042 (I53353,I53630,I53791);
nand I_3043 (I53338,I53647,I53791);
nor I_3044 (I53347,I53393,I53774);
DFFARX1 I_3045 (I53774,I2067,I53367,I53356,);
not I_3046 (I53894,I2074);
DFFARX1 I_3047 (I24483,I2067,I53894,I53920,);
nand I_3048 (I53928,I24483,I24489);
and I_3049 (I53945,I53928,I24507);
DFFARX1 I_3050 (I53945,I2067,I53894,I53971,);
nor I_3051 (I53862,I53971,I53920);
not I_3052 (I53993,I53971);
DFFARX1 I_3053 (I24495,I2067,I53894,I54019,);
nand I_3054 (I54027,I54019,I24492);
not I_3055 (I54044,I54027);
DFFARX1 I_3056 (I54044,I2067,I53894,I54070,);
not I_3057 (I53886,I54070);
nor I_3058 (I54092,I53920,I54027);
nor I_3059 (I53868,I53971,I54092);
DFFARX1 I_3060 (I24501,I2067,I53894,I54132,);
DFFARX1 I_3061 (I54132,I2067,I53894,I54149,);
not I_3062 (I54157,I54149);
not I_3063 (I54174,I54132);
nand I_3064 (I53871,I54174,I53993);
nand I_3065 (I54205,I24486,I24486);
and I_3066 (I54222,I54205,I24498);
DFFARX1 I_3067 (I54222,I2067,I53894,I54248,);
nor I_3068 (I54256,I54248,I53920);
DFFARX1 I_3069 (I54256,I2067,I53894,I53859,);
DFFARX1 I_3070 (I54248,I2067,I53894,I53877,);
nor I_3071 (I54301,I24504,I24486);
not I_3072 (I54318,I54301);
nor I_3073 (I53880,I54157,I54318);
nand I_3074 (I53865,I54174,I54318);
nor I_3075 (I53874,I53920,I54301);
DFFARX1 I_3076 (I54301,I2067,I53894,I53883,);
not I_3077 (I54421,I2074);
DFFARX1 I_3078 (I39358,I2067,I54421,I54447,);
nand I_3079 (I54455,I39358,I39364);
and I_3080 (I54472,I54455,I39382);
DFFARX1 I_3081 (I54472,I2067,I54421,I54498,);
nor I_3082 (I54389,I54498,I54447);
not I_3083 (I54520,I54498);
DFFARX1 I_3084 (I39370,I2067,I54421,I54546,);
nand I_3085 (I54554,I54546,I39367);
not I_3086 (I54571,I54554);
DFFARX1 I_3087 (I54571,I2067,I54421,I54597,);
not I_3088 (I54413,I54597);
nor I_3089 (I54619,I54447,I54554);
nor I_3090 (I54395,I54498,I54619);
DFFARX1 I_3091 (I39376,I2067,I54421,I54659,);
DFFARX1 I_3092 (I54659,I2067,I54421,I54676,);
not I_3093 (I54684,I54676);
not I_3094 (I54701,I54659);
nand I_3095 (I54398,I54701,I54520);
nand I_3096 (I54732,I39361,I39361);
and I_3097 (I54749,I54732,I39373);
DFFARX1 I_3098 (I54749,I2067,I54421,I54775,);
nor I_3099 (I54783,I54775,I54447);
DFFARX1 I_3100 (I54783,I2067,I54421,I54386,);
DFFARX1 I_3101 (I54775,I2067,I54421,I54404,);
nor I_3102 (I54828,I39379,I39361);
not I_3103 (I54845,I54828);
nor I_3104 (I54407,I54684,I54845);
nand I_3105 (I54392,I54701,I54845);
nor I_3106 (I54401,I54447,I54828);
DFFARX1 I_3107 (I54828,I2067,I54421,I54410,);
not I_3108 (I54948,I2074);
DFFARX1 I_3109 (I177045,I2067,I54948,I54974,);
nand I_3110 (I54982,I177024,I177024);
and I_3111 (I54999,I54982,I177051);
DFFARX1 I_3112 (I54999,I2067,I54948,I55025,);
nor I_3113 (I54916,I55025,I54974);
not I_3114 (I55047,I55025);
DFFARX1 I_3115 (I177039,I2067,I54948,I55073,);
nand I_3116 (I55081,I55073,I177042);
not I_3117 (I55098,I55081);
DFFARX1 I_3118 (I55098,I2067,I54948,I55124,);
not I_3119 (I54940,I55124);
nor I_3120 (I55146,I54974,I55081);
nor I_3121 (I54922,I55025,I55146);
DFFARX1 I_3122 (I177033,I2067,I54948,I55186,);
DFFARX1 I_3123 (I55186,I2067,I54948,I55203,);
not I_3124 (I55211,I55203);
not I_3125 (I55228,I55186);
nand I_3126 (I54925,I55228,I55047);
nand I_3127 (I55259,I177030,I177027);
and I_3128 (I55276,I55259,I177048);
DFFARX1 I_3129 (I55276,I2067,I54948,I55302,);
nor I_3130 (I55310,I55302,I54974);
DFFARX1 I_3131 (I55310,I2067,I54948,I54913,);
DFFARX1 I_3132 (I55302,I2067,I54948,I54931,);
nor I_3133 (I55355,I177036,I177027);
not I_3134 (I55372,I55355);
nor I_3135 (I54934,I55211,I55372);
nand I_3136 (I54919,I55228,I55372);
nor I_3137 (I54928,I54974,I55355);
DFFARX1 I_3138 (I55355,I2067,I54948,I54937,);
not I_3139 (I55475,I2074);
DFFARX1 I_3140 (I78439,I2067,I55475,I55501,);
nand I_3141 (I55509,I78424,I78427);
and I_3142 (I55526,I55509,I78442);
DFFARX1 I_3143 (I55526,I2067,I55475,I55552,);
nor I_3144 (I55443,I55552,I55501);
not I_3145 (I55574,I55552);
DFFARX1 I_3146 (I78436,I2067,I55475,I55600,);
nand I_3147 (I55608,I55600,I78427);
not I_3148 (I55625,I55608);
DFFARX1 I_3149 (I55625,I2067,I55475,I55651,);
not I_3150 (I55467,I55651);
nor I_3151 (I55673,I55501,I55608);
nor I_3152 (I55449,I55552,I55673);
DFFARX1 I_3153 (I78433,I2067,I55475,I55713,);
DFFARX1 I_3154 (I55713,I2067,I55475,I55730,);
not I_3155 (I55738,I55730);
not I_3156 (I55755,I55713);
nand I_3157 (I55452,I55755,I55574);
nand I_3158 (I55786,I78448,I78424);
and I_3159 (I55803,I55786,I78445);
DFFARX1 I_3160 (I55803,I2067,I55475,I55829,);
nor I_3161 (I55837,I55829,I55501);
DFFARX1 I_3162 (I55837,I2067,I55475,I55440,);
DFFARX1 I_3163 (I55829,I2067,I55475,I55458,);
nor I_3164 (I55882,I78430,I78424);
not I_3165 (I55899,I55882);
nor I_3166 (I55461,I55738,I55899);
nand I_3167 (I55446,I55755,I55899);
nor I_3168 (I55455,I55501,I55882);
DFFARX1 I_3169 (I55882,I2067,I55475,I55464,);
not I_3170 (I56002,I2074);
DFFARX1 I_3171 (I68924,I2067,I56002,I56028,);
nand I_3172 (I56036,I68924,I68936);
and I_3173 (I56053,I56036,I68921);
DFFARX1 I_3174 (I56053,I2067,I56002,I56079,);
nor I_3175 (I55970,I56079,I56028);
not I_3176 (I56101,I56079);
DFFARX1 I_3177 (I68945,I2067,I56002,I56127,);
nand I_3178 (I56135,I56127,I68942);
not I_3179 (I56152,I56135);
DFFARX1 I_3180 (I56152,I2067,I56002,I56178,);
not I_3181 (I55994,I56178);
nor I_3182 (I56200,I56028,I56135);
nor I_3183 (I55976,I56079,I56200);
DFFARX1 I_3184 (I68933,I2067,I56002,I56240,);
DFFARX1 I_3185 (I56240,I2067,I56002,I56257,);
not I_3186 (I56265,I56257);
not I_3187 (I56282,I56240);
nand I_3188 (I55979,I56282,I56101);
nand I_3189 (I56313,I68921,I68930);
and I_3190 (I56330,I56313,I68939);
DFFARX1 I_3191 (I56330,I2067,I56002,I56356,);
nor I_3192 (I56364,I56356,I56028);
DFFARX1 I_3193 (I56364,I2067,I56002,I55967,);
DFFARX1 I_3194 (I56356,I2067,I56002,I55985,);
nor I_3195 (I56409,I68927,I68930);
not I_3196 (I56426,I56409);
nor I_3197 (I55988,I56265,I56426);
nand I_3198 (I55973,I56282,I56426);
nor I_3199 (I55982,I56028,I56409);
DFFARX1 I_3200 (I56409,I2067,I56002,I55991,);
not I_3201 (I56529,I2074);
DFFARX1 I_3202 (I4848,I2067,I56529,I56555,);
nand I_3203 (I56563,I4872,I4851);
and I_3204 (I56580,I56563,I4848);
DFFARX1 I_3205 (I56580,I2067,I56529,I56606,);
nor I_3206 (I56497,I56606,I56555);
not I_3207 (I56628,I56606);
DFFARX1 I_3208 (I4854,I2067,I56529,I56654,);
nand I_3209 (I56662,I56654,I4863);
not I_3210 (I56679,I56662);
DFFARX1 I_3211 (I56679,I2067,I56529,I56705,);
not I_3212 (I56521,I56705);
nor I_3213 (I56727,I56555,I56662);
nor I_3214 (I56503,I56606,I56727);
DFFARX1 I_3215 (I4857,I2067,I56529,I56767,);
DFFARX1 I_3216 (I56767,I2067,I56529,I56784,);
not I_3217 (I56792,I56784);
not I_3218 (I56809,I56767);
nand I_3219 (I56506,I56809,I56628);
nand I_3220 (I56840,I4869,I4851);
and I_3221 (I56857,I56840,I4860);
DFFARX1 I_3222 (I56857,I2067,I56529,I56883,);
nor I_3223 (I56891,I56883,I56555);
DFFARX1 I_3224 (I56891,I2067,I56529,I56494,);
DFFARX1 I_3225 (I56883,I2067,I56529,I56512,);
nor I_3226 (I56936,I4866,I4851);
not I_3227 (I56953,I56936);
nor I_3228 (I56515,I56792,I56953);
nand I_3229 (I56500,I56809,I56953);
nor I_3230 (I56509,I56555,I56936);
DFFARX1 I_3231 (I56936,I2067,I56529,I56518,);
not I_3232 (I57056,I2074);
DFFARX1 I_3233 (I118445,I2067,I57056,I57082,);
nand I_3234 (I57090,I118442,I118460);
and I_3235 (I57107,I57090,I118451);
DFFARX1 I_3236 (I57107,I2067,I57056,I57133,);
nor I_3237 (I57024,I57133,I57082);
not I_3238 (I57155,I57133);
DFFARX1 I_3239 (I118466,I2067,I57056,I57181,);
nand I_3240 (I57189,I57181,I118448);
not I_3241 (I57206,I57189);
DFFARX1 I_3242 (I57206,I2067,I57056,I57232,);
not I_3243 (I57048,I57232);
nor I_3244 (I57254,I57082,I57189);
nor I_3245 (I57030,I57133,I57254);
DFFARX1 I_3246 (I118454,I2067,I57056,I57294,);
DFFARX1 I_3247 (I57294,I2067,I57056,I57311,);
not I_3248 (I57319,I57311);
not I_3249 (I57336,I57294);
nand I_3250 (I57033,I57336,I57155);
nand I_3251 (I57367,I118442,I118469);
and I_3252 (I57384,I57367,I118457);
DFFARX1 I_3253 (I57384,I2067,I57056,I57410,);
nor I_3254 (I57418,I57410,I57082);
DFFARX1 I_3255 (I57418,I2067,I57056,I57021,);
DFFARX1 I_3256 (I57410,I2067,I57056,I57039,);
nor I_3257 (I57463,I118463,I118469);
not I_3258 (I57480,I57463);
nor I_3259 (I57042,I57319,I57480);
nand I_3260 (I57027,I57336,I57480);
nor I_3261 (I57036,I57082,I57463);
DFFARX1 I_3262 (I57463,I2067,I57056,I57045,);
not I_3263 (I57583,I2074);
DFFARX1 I_3264 (I38763,I2067,I57583,I57609,);
nand I_3265 (I57617,I38763,I38769);
and I_3266 (I57634,I57617,I38787);
DFFARX1 I_3267 (I57634,I2067,I57583,I57660,);
nor I_3268 (I57551,I57660,I57609);
not I_3269 (I57682,I57660);
DFFARX1 I_3270 (I38775,I2067,I57583,I57708,);
nand I_3271 (I57716,I57708,I38772);
not I_3272 (I57733,I57716);
DFFARX1 I_3273 (I57733,I2067,I57583,I57759,);
not I_3274 (I57575,I57759);
nor I_3275 (I57781,I57609,I57716);
nor I_3276 (I57557,I57660,I57781);
DFFARX1 I_3277 (I38781,I2067,I57583,I57821,);
DFFARX1 I_3278 (I57821,I2067,I57583,I57838,);
not I_3279 (I57846,I57838);
not I_3280 (I57863,I57821);
nand I_3281 (I57560,I57863,I57682);
nand I_3282 (I57894,I38766,I38766);
and I_3283 (I57911,I57894,I38778);
DFFARX1 I_3284 (I57911,I2067,I57583,I57937,);
nor I_3285 (I57945,I57937,I57609);
DFFARX1 I_3286 (I57945,I2067,I57583,I57548,);
DFFARX1 I_3287 (I57937,I2067,I57583,I57566,);
nor I_3288 (I57990,I38784,I38766);
not I_3289 (I58007,I57990);
nor I_3290 (I57569,I57846,I58007);
nand I_3291 (I57554,I57863,I58007);
nor I_3292 (I57563,I57609,I57990);
DFFARX1 I_3293 (I57990,I2067,I57583,I57572,);
not I_3294 (I58110,I2074);
DFFARX1 I_3295 (I117153,I2067,I58110,I58136,);
nand I_3296 (I58144,I117150,I117168);
and I_3297 (I58161,I58144,I117159);
DFFARX1 I_3298 (I58161,I2067,I58110,I58187,);
nor I_3299 (I58078,I58187,I58136);
not I_3300 (I58209,I58187);
DFFARX1 I_3301 (I117174,I2067,I58110,I58235,);
nand I_3302 (I58243,I58235,I117156);
not I_3303 (I58260,I58243);
DFFARX1 I_3304 (I58260,I2067,I58110,I58286,);
not I_3305 (I58102,I58286);
nor I_3306 (I58308,I58136,I58243);
nor I_3307 (I58084,I58187,I58308);
DFFARX1 I_3308 (I117162,I2067,I58110,I58348,);
DFFARX1 I_3309 (I58348,I2067,I58110,I58365,);
not I_3310 (I58373,I58365);
not I_3311 (I58390,I58348);
nand I_3312 (I58087,I58390,I58209);
nand I_3313 (I58421,I117150,I117177);
and I_3314 (I58438,I58421,I117165);
DFFARX1 I_3315 (I58438,I2067,I58110,I58464,);
nor I_3316 (I58472,I58464,I58136);
DFFARX1 I_3317 (I58472,I2067,I58110,I58075,);
DFFARX1 I_3318 (I58464,I2067,I58110,I58093,);
nor I_3319 (I58517,I117171,I117177);
not I_3320 (I58534,I58517);
nor I_3321 (I58096,I58373,I58534);
nand I_3322 (I58081,I58390,I58534);
nor I_3323 (I58090,I58136,I58517);
DFFARX1 I_3324 (I58517,I2067,I58110,I58099,);
not I_3325 (I58637,I2074);
DFFARX1 I_3326 (I62949,I2067,I58637,I58663,);
nand I_3327 (I58671,I62961,I62940);
and I_3328 (I58688,I58671,I62964);
DFFARX1 I_3329 (I58688,I2067,I58637,I58714,);
nor I_3330 (I58605,I58714,I58663);
not I_3331 (I58736,I58714);
DFFARX1 I_3332 (I62955,I2067,I58637,I58762,);
nand I_3333 (I58770,I58762,I62937);
not I_3334 (I58787,I58770);
DFFARX1 I_3335 (I58787,I2067,I58637,I58813,);
not I_3336 (I58629,I58813);
nor I_3337 (I58835,I58663,I58770);
nor I_3338 (I58611,I58714,I58835);
DFFARX1 I_3339 (I62952,I2067,I58637,I58875,);
DFFARX1 I_3340 (I58875,I2067,I58637,I58892,);
not I_3341 (I58900,I58892);
not I_3342 (I58917,I58875);
nand I_3343 (I58614,I58917,I58736);
nand I_3344 (I58948,I62937,I62943);
and I_3345 (I58965,I58948,I62946);
DFFARX1 I_3346 (I58965,I2067,I58637,I58991,);
nor I_3347 (I58999,I58991,I58663);
DFFARX1 I_3348 (I58999,I2067,I58637,I58602,);
DFFARX1 I_3349 (I58991,I2067,I58637,I58620,);
nor I_3350 (I59044,I62958,I62943);
not I_3351 (I59061,I59044);
nor I_3352 (I58623,I58900,I59061);
nand I_3353 (I58608,I58917,I59061);
nor I_3354 (I58617,I58663,I59044);
DFFARX1 I_3355 (I59044,I2067,I58637,I58626,);
not I_3356 (I59164,I2074);
DFFARX1 I_3357 (I138539,I2067,I59164,I59190,);
DFFARX1 I_3358 (I59190,I2067,I59164,I59207,);
not I_3359 (I59156,I59207);
not I_3360 (I59229,I59190);
nand I_3361 (I59246,I138551,I138539);
and I_3362 (I59263,I59246,I138542);
DFFARX1 I_3363 (I59263,I2067,I59164,I59289,);
not I_3364 (I59297,I59289);
DFFARX1 I_3365 (I138560,I2067,I59164,I59323,);
and I_3366 (I59331,I59323,I138536);
nand I_3367 (I59348,I59323,I138536);
nand I_3368 (I59135,I59297,I59348);
DFFARX1 I_3369 (I138554,I2067,I59164,I59388,);
nor I_3370 (I59396,I59388,I59331);
DFFARX1 I_3371 (I59396,I2067,I59164,I59129,);
nor I_3372 (I59144,I59388,I59289);
nand I_3373 (I59441,I138548,I138545);
and I_3374 (I59458,I59441,I138557);
DFFARX1 I_3375 (I59458,I2067,I59164,I59484,);
nor I_3376 (I59132,I59484,I59388);
not I_3377 (I59506,I59484);
nor I_3378 (I59523,I59506,I59297);
nor I_3379 (I59540,I59229,I59523);
DFFARX1 I_3380 (I59540,I2067,I59164,I59147,);
nor I_3381 (I59571,I59506,I59388);
nor I_3382 (I59588,I138536,I138545);
nor I_3383 (I59138,I59588,I59571);
not I_3384 (I59619,I59588);
nand I_3385 (I59141,I59348,I59619);
DFFARX1 I_3386 (I59588,I2067,I59164,I59153,);
DFFARX1 I_3387 (I59588,I2067,I59164,I59150,);
not I_3388 (I59708,I2074);
DFFARX1 I_3389 (I58096,I2067,I59708,I59734,);
DFFARX1 I_3390 (I59734,I2067,I59708,I59751,);
not I_3391 (I59700,I59751);
not I_3392 (I59773,I59734);
nand I_3393 (I59790,I58075,I58099);
and I_3394 (I59807,I59790,I58102);
DFFARX1 I_3395 (I59807,I2067,I59708,I59833,);
not I_3396 (I59841,I59833);
DFFARX1 I_3397 (I58084,I2067,I59708,I59867,);
and I_3398 (I59875,I59867,I58090);
nand I_3399 (I59892,I59867,I58090);
nand I_3400 (I59679,I59841,I59892);
DFFARX1 I_3401 (I58078,I2067,I59708,I59932,);
nor I_3402 (I59940,I59932,I59875);
DFFARX1 I_3403 (I59940,I2067,I59708,I59673,);
nor I_3404 (I59688,I59932,I59833);
nand I_3405 (I59985,I58087,I58075);
and I_3406 (I60002,I59985,I58081);
DFFARX1 I_3407 (I60002,I2067,I59708,I60028,);
nor I_3408 (I59676,I60028,I59932);
not I_3409 (I60050,I60028);
nor I_3410 (I60067,I60050,I59841);
nor I_3411 (I60084,I59773,I60067);
DFFARX1 I_3412 (I60084,I2067,I59708,I59691,);
nor I_3413 (I60115,I60050,I59932);
nor I_3414 (I60132,I58093,I58075);
nor I_3415 (I59682,I60132,I60115);
not I_3416 (I60163,I60132);
nand I_3417 (I59685,I59892,I60163);
DFFARX1 I_3418 (I60132,I2067,I59708,I59697,);
DFFARX1 I_3419 (I60132,I2067,I59708,I59694,);
not I_3420 (I60252,I2074);
DFFARX1 I_3421 (I100969,I2067,I60252,I60278,);
DFFARX1 I_3422 (I60278,I2067,I60252,I60295,);
not I_3423 (I60244,I60295);
not I_3424 (I60317,I60278);
nand I_3425 (I60334,I100990,I100981);
and I_3426 (I60351,I60334,I100969);
DFFARX1 I_3427 (I60351,I2067,I60252,I60377,);
not I_3428 (I60385,I60377);
DFFARX1 I_3429 (I100975,I2067,I60252,I60411,);
and I_3430 (I60419,I60411,I100972);
nand I_3431 (I60436,I60411,I100972);
nand I_3432 (I60223,I60385,I60436);
DFFARX1 I_3433 (I100966,I2067,I60252,I60476,);
nor I_3434 (I60484,I60476,I60419);
DFFARX1 I_3435 (I60484,I2067,I60252,I60217,);
nor I_3436 (I60232,I60476,I60377);
nand I_3437 (I60529,I100966,I100978);
and I_3438 (I60546,I60529,I100987);
DFFARX1 I_3439 (I60546,I2067,I60252,I60572,);
nor I_3440 (I60220,I60572,I60476);
not I_3441 (I60594,I60572);
nor I_3442 (I60611,I60594,I60385);
nor I_3443 (I60628,I60317,I60611);
DFFARX1 I_3444 (I60628,I2067,I60252,I60235,);
nor I_3445 (I60659,I60594,I60476);
nor I_3446 (I60676,I100984,I100978);
nor I_3447 (I60226,I60676,I60659);
not I_3448 (I60707,I60676);
nand I_3449 (I60229,I60436,I60707);
DFFARX1 I_3450 (I60676,I2067,I60252,I60241,);
DFFARX1 I_3451 (I60676,I2067,I60252,I60238,);
not I_3452 (I60796,I2074);
DFFARX1 I_3453 (I155709,I2067,I60796,I60822,);
DFFARX1 I_3454 (I60822,I2067,I60796,I60839,);
not I_3455 (I60788,I60839);
not I_3456 (I60861,I60822);
nand I_3457 (I60878,I155721,I155724);
and I_3458 (I60895,I60878,I155727);
DFFARX1 I_3459 (I60895,I2067,I60796,I60921,);
not I_3460 (I60929,I60921);
DFFARX1 I_3461 (I155712,I2067,I60796,I60955,);
and I_3462 (I60963,I60955,I155718);
nand I_3463 (I60980,I60955,I155718);
nand I_3464 (I60767,I60929,I60980);
DFFARX1 I_3465 (I155706,I2067,I60796,I61020,);
nor I_3466 (I61028,I61020,I60963);
DFFARX1 I_3467 (I61028,I2067,I60796,I60761,);
nor I_3468 (I60776,I61020,I60921);
nand I_3469 (I61073,I155709,I155730);
and I_3470 (I61090,I61073,I155715);
DFFARX1 I_3471 (I61090,I2067,I60796,I61116,);
nor I_3472 (I60764,I61116,I61020);
not I_3473 (I61138,I61116);
nor I_3474 (I61155,I61138,I60929);
nor I_3475 (I61172,I60861,I61155);
DFFARX1 I_3476 (I61172,I2067,I60796,I60779,);
nor I_3477 (I61203,I61138,I61020);
nor I_3478 (I61220,I155706,I155730);
nor I_3479 (I60770,I61220,I61203);
not I_3480 (I61251,I61220);
nand I_3481 (I60773,I60980,I61251);
DFFARX1 I_3482 (I61220,I2067,I60796,I60785,);
DFFARX1 I_3483 (I61220,I2067,I60796,I60782,);
not I_3484 (I61340,I2074);
DFFARX1 I_3485 (I143163,I2067,I61340,I61366,);
DFFARX1 I_3486 (I61366,I2067,I61340,I61383,);
not I_3487 (I61332,I61383);
not I_3488 (I61405,I61366);
nand I_3489 (I61422,I143175,I143163);
and I_3490 (I61439,I61422,I143166);
DFFARX1 I_3491 (I61439,I2067,I61340,I61465,);
not I_3492 (I61473,I61465);
DFFARX1 I_3493 (I143184,I2067,I61340,I61499,);
and I_3494 (I61507,I61499,I143160);
nand I_3495 (I61524,I61499,I143160);
nand I_3496 (I61311,I61473,I61524);
DFFARX1 I_3497 (I143178,I2067,I61340,I61564,);
nor I_3498 (I61572,I61564,I61507);
DFFARX1 I_3499 (I61572,I2067,I61340,I61305,);
nor I_3500 (I61320,I61564,I61465);
nand I_3501 (I61617,I143172,I143169);
and I_3502 (I61634,I61617,I143181);
DFFARX1 I_3503 (I61634,I2067,I61340,I61660,);
nor I_3504 (I61308,I61660,I61564);
not I_3505 (I61682,I61660);
nor I_3506 (I61699,I61682,I61473);
nor I_3507 (I61716,I61405,I61699);
DFFARX1 I_3508 (I61716,I2067,I61340,I61323,);
nor I_3509 (I61747,I61682,I61564);
nor I_3510 (I61764,I143160,I143169);
nor I_3511 (I61314,I61764,I61747);
not I_3512 (I61795,I61764);
nand I_3513 (I61317,I61524,I61795);
DFFARX1 I_3514 (I61764,I2067,I61340,I61329,);
DFFARX1 I_3515 (I61764,I2067,I61340,I61326,);
not I_3516 (I61884,I2074);
DFFARX1 I_3517 (I142585,I2067,I61884,I61910,);
DFFARX1 I_3518 (I61910,I2067,I61884,I61927,);
not I_3519 (I61876,I61927);
not I_3520 (I61949,I61910);
nand I_3521 (I61966,I142597,I142585);
and I_3522 (I61983,I61966,I142588);
DFFARX1 I_3523 (I61983,I2067,I61884,I62009,);
not I_3524 (I62017,I62009);
DFFARX1 I_3525 (I142606,I2067,I61884,I62043,);
and I_3526 (I62051,I62043,I142582);
nand I_3527 (I62068,I62043,I142582);
nand I_3528 (I61855,I62017,I62068);
DFFARX1 I_3529 (I142600,I2067,I61884,I62108,);
nor I_3530 (I62116,I62108,I62051);
DFFARX1 I_3531 (I62116,I2067,I61884,I61849,);
nor I_3532 (I61864,I62108,I62009);
nand I_3533 (I62161,I142594,I142591);
and I_3534 (I62178,I62161,I142603);
DFFARX1 I_3535 (I62178,I2067,I61884,I62204,);
nor I_3536 (I61852,I62204,I62108);
not I_3537 (I62226,I62204);
nor I_3538 (I62243,I62226,I62017);
nor I_3539 (I62260,I61949,I62243);
DFFARX1 I_3540 (I62260,I2067,I61884,I61867,);
nor I_3541 (I62291,I62226,I62108);
nor I_3542 (I62308,I142582,I142591);
nor I_3543 (I61858,I62308,I62291);
not I_3544 (I62339,I62308);
nand I_3545 (I61861,I62068,I62339);
DFFARX1 I_3546 (I62308,I2067,I61884,I61873,);
DFFARX1 I_3547 (I62308,I2067,I61884,I61870,);
not I_3548 (I62428,I2074);
DFFARX1 I_3549 (I51772,I2067,I62428,I62454,);
DFFARX1 I_3550 (I62454,I2067,I62428,I62471,);
not I_3551 (I62420,I62471);
not I_3552 (I62493,I62454);
nand I_3553 (I62510,I51751,I51775);
and I_3554 (I62527,I62510,I51778);
DFFARX1 I_3555 (I62527,I2067,I62428,I62553,);
not I_3556 (I62561,I62553);
DFFARX1 I_3557 (I51760,I2067,I62428,I62587,);
and I_3558 (I62595,I62587,I51766);
nand I_3559 (I62612,I62587,I51766);
nand I_3560 (I62399,I62561,I62612);
DFFARX1 I_3561 (I51754,I2067,I62428,I62652,);
nor I_3562 (I62660,I62652,I62595);
DFFARX1 I_3563 (I62660,I2067,I62428,I62393,);
nor I_3564 (I62408,I62652,I62553);
nand I_3565 (I62705,I51763,I51751);
and I_3566 (I62722,I62705,I51757);
DFFARX1 I_3567 (I62722,I2067,I62428,I62748,);
nor I_3568 (I62396,I62748,I62652);
not I_3569 (I62770,I62748);
nor I_3570 (I62787,I62770,I62561);
nor I_3571 (I62804,I62493,I62787);
DFFARX1 I_3572 (I62804,I2067,I62428,I62411,);
nor I_3573 (I62835,I62770,I62652);
nor I_3574 (I62852,I51769,I51751);
nor I_3575 (I62402,I62852,I62835);
not I_3576 (I62883,I62852);
nand I_3577 (I62405,I62612,I62883);
DFFARX1 I_3578 (I62852,I2067,I62428,I62417,);
DFFARX1 I_3579 (I62852,I2067,I62428,I62414,);
not I_3580 (I62972,I2074);
DFFARX1 I_3581 (I107081,I2067,I62972,I62998,);
DFFARX1 I_3582 (I62998,I2067,I62972,I63015,);
not I_3583 (I62964,I63015);
not I_3584 (I63037,I62998);
nand I_3585 (I63054,I107075,I107072);
and I_3586 (I63071,I63054,I107087);
DFFARX1 I_3587 (I63071,I2067,I62972,I63097,);
not I_3588 (I63105,I63097);
DFFARX1 I_3589 (I107075,I2067,I62972,I63131,);
and I_3590 (I63139,I63131,I107069);
nand I_3591 (I63156,I63131,I107069);
nand I_3592 (I62943,I63105,I63156);
DFFARX1 I_3593 (I107069,I2067,I62972,I63196,);
nor I_3594 (I63204,I63196,I63139);
DFFARX1 I_3595 (I63204,I2067,I62972,I62937,);
nor I_3596 (I62952,I63196,I63097);
nand I_3597 (I63249,I107084,I107078);
and I_3598 (I63266,I63249,I107072);
DFFARX1 I_3599 (I63266,I2067,I62972,I63292,);
nor I_3600 (I62940,I63292,I63196);
not I_3601 (I63314,I63292);
nor I_3602 (I63331,I63314,I63105);
nor I_3603 (I63348,I63037,I63331);
DFFARX1 I_3604 (I63348,I2067,I62972,I62955,);
nor I_3605 (I63379,I63314,I63196);
nor I_3606 (I63396,I107090,I107078);
nor I_3607 (I62946,I63396,I63379);
not I_3608 (I63427,I63396);
nand I_3609 (I62949,I63156,I63427);
DFFARX1 I_3610 (I63396,I2067,I62972,I62961,);
DFFARX1 I_3611 (I63396,I2067,I62972,I62958,);
not I_3612 (I63516,I2074);
DFFARX1 I_3613 (I41152,I2067,I63516,I63542,);
DFFARX1 I_3614 (I63542,I2067,I63516,I63559,);
not I_3615 (I63508,I63559);
not I_3616 (I63581,I63542);
nand I_3617 (I63598,I41164,I41143);
and I_3618 (I63615,I63598,I41146);
DFFARX1 I_3619 (I63615,I2067,I63516,I63641,);
not I_3620 (I63649,I63641);
DFFARX1 I_3621 (I41155,I2067,I63516,I63675,);
and I_3622 (I63683,I63675,I41167);
nand I_3623 (I63700,I63675,I41167);
nand I_3624 (I63487,I63649,I63700);
DFFARX1 I_3625 (I41161,I2067,I63516,I63740,);
nor I_3626 (I63748,I63740,I63683);
DFFARX1 I_3627 (I63748,I2067,I63516,I63481,);
nor I_3628 (I63496,I63740,I63641);
nand I_3629 (I63793,I41149,I41146);
and I_3630 (I63810,I63793,I41158);
DFFARX1 I_3631 (I63810,I2067,I63516,I63836,);
nor I_3632 (I63484,I63836,I63740);
not I_3633 (I63858,I63836);
nor I_3634 (I63875,I63858,I63649);
nor I_3635 (I63892,I63581,I63875);
DFFARX1 I_3636 (I63892,I2067,I63516,I63499,);
nor I_3637 (I63923,I63858,I63740);
nor I_3638 (I63940,I41143,I41146);
nor I_3639 (I63490,I63940,I63923);
not I_3640 (I63971,I63940);
nand I_3641 (I63493,I63700,I63971);
DFFARX1 I_3642 (I63940,I2067,I63516,I63505,);
DFFARX1 I_3643 (I63940,I2067,I63516,I63502,);
not I_3644 (I64060,I2074);
DFFARX1 I_3645 (I1460,I2067,I64060,I64086,);
DFFARX1 I_3646 (I64086,I2067,I64060,I64103,);
not I_3647 (I64052,I64103);
not I_3648 (I64125,I64086);
nand I_3649 (I64142,I2004,I1500);
and I_3650 (I64159,I64142,I1860);
DFFARX1 I_3651 (I64159,I2067,I64060,I64185,);
not I_3652 (I64193,I64185);
DFFARX1 I_3653 (I1412,I2067,I64060,I64219,);
and I_3654 (I64227,I64219,I1452);
nand I_3655 (I64244,I64219,I1452);
nand I_3656 (I64031,I64193,I64244);
DFFARX1 I_3657 (I1996,I2067,I64060,I64284,);
nor I_3658 (I64292,I64284,I64227);
DFFARX1 I_3659 (I64292,I2067,I64060,I64025,);
nor I_3660 (I64040,I64284,I64185);
nand I_3661 (I64337,I1468,I1604);
and I_3662 (I64354,I64337,I1508);
DFFARX1 I_3663 (I64354,I2067,I64060,I64380,);
nor I_3664 (I64028,I64380,I64284);
not I_3665 (I64402,I64380);
nor I_3666 (I64419,I64402,I64193);
nor I_3667 (I64436,I64125,I64419);
DFFARX1 I_3668 (I64436,I2067,I64060,I64043,);
nor I_3669 (I64467,I64402,I64284);
nor I_3670 (I64484,I1428,I1604);
nor I_3671 (I64034,I64484,I64467);
not I_3672 (I64515,I64484);
nand I_3673 (I64037,I64244,I64515);
DFFARX1 I_3674 (I64484,I2067,I64060,I64049,);
DFFARX1 I_3675 (I64484,I2067,I64060,I64046,);
not I_3676 (I64604,I2074);
DFFARX1 I_3677 (I5387,I2067,I64604,I64630,);
DFFARX1 I_3678 (I64630,I2067,I64604,I64647,);
not I_3679 (I64596,I64647);
not I_3680 (I64669,I64630);
nand I_3681 (I64686,I5375,I5390);
and I_3682 (I64703,I64686,I5378);
DFFARX1 I_3683 (I64703,I2067,I64604,I64729,);
not I_3684 (I64737,I64729);
DFFARX1 I_3685 (I5399,I2067,I64604,I64763,);
and I_3686 (I64771,I64763,I5393);
nand I_3687 (I64788,I64763,I5393);
nand I_3688 (I64575,I64737,I64788);
DFFARX1 I_3689 (I5396,I2067,I64604,I64828,);
nor I_3690 (I64836,I64828,I64771);
DFFARX1 I_3691 (I64836,I2067,I64604,I64569,);
nor I_3692 (I64584,I64828,I64729);
nand I_3693 (I64881,I5375,I5378);
and I_3694 (I64898,I64881,I5381);
DFFARX1 I_3695 (I64898,I2067,I64604,I64924,);
nor I_3696 (I64572,I64924,I64828);
not I_3697 (I64946,I64924);
nor I_3698 (I64963,I64946,I64737);
nor I_3699 (I64980,I64669,I64963);
DFFARX1 I_3700 (I64980,I2067,I64604,I64587,);
nor I_3701 (I65011,I64946,I64828);
nor I_3702 (I65028,I5384,I5378);
nor I_3703 (I64578,I65028,I65011);
not I_3704 (I65059,I65028);
nand I_3705 (I64581,I64788,I65059);
DFFARX1 I_3706 (I65028,I2067,I64604,I64593,);
DFFARX1 I_3707 (I65028,I2067,I64604,I64590,);
not I_3708 (I65148,I2074);
DFFARX1 I_3709 (I45448,I2067,I65148,I65174,);
DFFARX1 I_3710 (I65174,I2067,I65148,I65191,);
not I_3711 (I65140,I65191);
not I_3712 (I65213,I65174);
nand I_3713 (I65230,I45427,I45451);
and I_3714 (I65247,I65230,I45454);
DFFARX1 I_3715 (I65247,I2067,I65148,I65273,);
not I_3716 (I65281,I65273);
DFFARX1 I_3717 (I45436,I2067,I65148,I65307,);
and I_3718 (I65315,I65307,I45442);
nand I_3719 (I65332,I65307,I45442);
nand I_3720 (I65119,I65281,I65332);
DFFARX1 I_3721 (I45430,I2067,I65148,I65372,);
nor I_3722 (I65380,I65372,I65315);
DFFARX1 I_3723 (I65380,I2067,I65148,I65113,);
nor I_3724 (I65128,I65372,I65273);
nand I_3725 (I65425,I45439,I45427);
and I_3726 (I65442,I65425,I45433);
DFFARX1 I_3727 (I65442,I2067,I65148,I65468,);
nor I_3728 (I65116,I65468,I65372);
not I_3729 (I65490,I65468);
nor I_3730 (I65507,I65490,I65281);
nor I_3731 (I65524,I65213,I65507);
DFFARX1 I_3732 (I65524,I2067,I65148,I65131,);
nor I_3733 (I65555,I65490,I65372);
nor I_3734 (I65572,I45445,I45427);
nor I_3735 (I65122,I65572,I65555);
not I_3736 (I65603,I65572);
nand I_3737 (I65125,I65332,I65603);
DFFARX1 I_3738 (I65572,I2067,I65148,I65137,);
DFFARX1 I_3739 (I65572,I2067,I65148,I65134,);
not I_3740 (I65692,I2074);
DFFARX1 I_3741 (I48083,I2067,I65692,I65718,);
DFFARX1 I_3742 (I65718,I2067,I65692,I65735,);
not I_3743 (I65684,I65735);
not I_3744 (I65757,I65718);
nand I_3745 (I65774,I48062,I48086);
and I_3746 (I65791,I65774,I48089);
DFFARX1 I_3747 (I65791,I2067,I65692,I65817,);
not I_3748 (I65825,I65817);
DFFARX1 I_3749 (I48071,I2067,I65692,I65851,);
and I_3750 (I65859,I65851,I48077);
nand I_3751 (I65876,I65851,I48077);
nand I_3752 (I65663,I65825,I65876);
DFFARX1 I_3753 (I48065,I2067,I65692,I65916,);
nor I_3754 (I65924,I65916,I65859);
DFFARX1 I_3755 (I65924,I2067,I65692,I65657,);
nor I_3756 (I65672,I65916,I65817);
nand I_3757 (I65969,I48074,I48062);
and I_3758 (I65986,I65969,I48068);
DFFARX1 I_3759 (I65986,I2067,I65692,I66012,);
nor I_3760 (I65660,I66012,I65916);
not I_3761 (I66034,I66012);
nor I_3762 (I66051,I66034,I65825);
nor I_3763 (I66068,I65757,I66051);
DFFARX1 I_3764 (I66068,I2067,I65692,I65675,);
nor I_3765 (I66099,I66034,I65916);
nor I_3766 (I66116,I48080,I48062);
nor I_3767 (I65666,I66116,I66099);
not I_3768 (I66147,I66116);
nand I_3769 (I65669,I65876,I66147);
DFFARX1 I_3770 (I66116,I2067,I65692,I65681,);
DFFARX1 I_3771 (I66116,I2067,I65692,I65678,);
not I_3772 (I66236,I2074);
DFFARX1 I_3773 (I127492,I2067,I66236,I66262,);
DFFARX1 I_3774 (I66262,I2067,I66236,I66279,);
not I_3775 (I66228,I66279);
not I_3776 (I66301,I66262);
nand I_3777 (I66318,I127507,I127495);
and I_3778 (I66335,I66318,I127486);
DFFARX1 I_3779 (I66335,I2067,I66236,I66361,);
not I_3780 (I66369,I66361);
DFFARX1 I_3781 (I127498,I2067,I66236,I66395,);
and I_3782 (I66403,I66395,I127489);
nand I_3783 (I66420,I66395,I127489);
nand I_3784 (I66207,I66369,I66420);
DFFARX1 I_3785 (I127504,I2067,I66236,I66460,);
nor I_3786 (I66468,I66460,I66403);
DFFARX1 I_3787 (I66468,I2067,I66236,I66201,);
nor I_3788 (I66216,I66460,I66361);
nand I_3789 (I66513,I127513,I127501);
and I_3790 (I66530,I66513,I127510);
DFFARX1 I_3791 (I66530,I2067,I66236,I66556,);
nor I_3792 (I66204,I66556,I66460);
not I_3793 (I66578,I66556);
nor I_3794 (I66595,I66578,I66369);
nor I_3795 (I66612,I66301,I66595);
DFFARX1 I_3796 (I66612,I2067,I66236,I66219,);
nor I_3797 (I66643,I66578,I66460);
nor I_3798 (I66660,I127486,I127501);
nor I_3799 (I66210,I66660,I66643);
not I_3800 (I66691,I66660);
nand I_3801 (I66213,I66420,I66691);
DFFARX1 I_3802 (I66660,I2067,I66236,I66225,);
DFFARX1 I_3803 (I66660,I2067,I66236,I66222,);
not I_3804 (I66780,I2074);
DFFARX1 I_3805 (I147209,I2067,I66780,I66806,);
DFFARX1 I_3806 (I66806,I2067,I66780,I66823,);
not I_3807 (I66772,I66823);
not I_3808 (I66845,I66806);
nand I_3809 (I66862,I147221,I147209);
and I_3810 (I66879,I66862,I147212);
DFFARX1 I_3811 (I66879,I2067,I66780,I66905,);
not I_3812 (I66913,I66905);
DFFARX1 I_3813 (I147230,I2067,I66780,I66939,);
and I_3814 (I66947,I66939,I147206);
nand I_3815 (I66964,I66939,I147206);
nand I_3816 (I66751,I66913,I66964);
DFFARX1 I_3817 (I147224,I2067,I66780,I67004,);
nor I_3818 (I67012,I67004,I66947);
DFFARX1 I_3819 (I67012,I2067,I66780,I66745,);
nor I_3820 (I66760,I67004,I66905);
nand I_3821 (I67057,I147218,I147215);
and I_3822 (I67074,I67057,I147227);
DFFARX1 I_3823 (I67074,I2067,I66780,I67100,);
nor I_3824 (I66748,I67100,I67004);
not I_3825 (I67122,I67100);
nor I_3826 (I67139,I67122,I66913);
nor I_3827 (I67156,I66845,I67139);
DFFARX1 I_3828 (I67156,I2067,I66780,I66763,);
nor I_3829 (I67187,I67122,I67004);
nor I_3830 (I67204,I147206,I147215);
nor I_3831 (I66754,I67204,I67187);
not I_3832 (I67235,I67204);
nand I_3833 (I66757,I66964,I67235);
DFFARX1 I_3834 (I67204,I2067,I66780,I66769,);
DFFARX1 I_3835 (I67204,I2067,I66780,I66766,);
not I_3836 (I67324,I2074);
DFFARX1 I_3837 (I115864,I2067,I67324,I67350,);
DFFARX1 I_3838 (I67350,I2067,I67324,I67367,);
not I_3839 (I67316,I67367);
not I_3840 (I67389,I67350);
nand I_3841 (I67406,I115879,I115867);
and I_3842 (I67423,I67406,I115858);
DFFARX1 I_3843 (I67423,I2067,I67324,I67449,);
not I_3844 (I67457,I67449);
DFFARX1 I_3845 (I115870,I2067,I67324,I67483,);
and I_3846 (I67491,I67483,I115861);
nand I_3847 (I67508,I67483,I115861);
nand I_3848 (I67295,I67457,I67508);
DFFARX1 I_3849 (I115876,I2067,I67324,I67548,);
nor I_3850 (I67556,I67548,I67491);
DFFARX1 I_3851 (I67556,I2067,I67324,I67289,);
nor I_3852 (I67304,I67548,I67449);
nand I_3853 (I67601,I115885,I115873);
and I_3854 (I67618,I67601,I115882);
DFFARX1 I_3855 (I67618,I2067,I67324,I67644,);
nor I_3856 (I67292,I67644,I67548);
not I_3857 (I67666,I67644);
nor I_3858 (I67683,I67666,I67457);
nor I_3859 (I67700,I67389,I67683);
DFFARX1 I_3860 (I67700,I2067,I67324,I67307,);
nor I_3861 (I67731,I67666,I67548);
nor I_3862 (I67748,I115858,I115873);
nor I_3863 (I67298,I67748,I67731);
not I_3864 (I67779,I67748);
nand I_3865 (I67301,I67508,I67779);
DFFARX1 I_3866 (I67748,I2067,I67324,I67313,);
DFFARX1 I_3867 (I67748,I2067,I67324,I67310,);
not I_3868 (I67868,I2074);
DFFARX1 I_3869 (I36392,I2067,I67868,I67894,);
DFFARX1 I_3870 (I67894,I2067,I67868,I67911,);
not I_3871 (I67860,I67911);
not I_3872 (I67933,I67894);
nand I_3873 (I67950,I36404,I36383);
and I_3874 (I67967,I67950,I36386);
DFFARX1 I_3875 (I67967,I2067,I67868,I67993,);
not I_3876 (I68001,I67993);
DFFARX1 I_3877 (I36395,I2067,I67868,I68027,);
and I_3878 (I68035,I68027,I36407);
nand I_3879 (I68052,I68027,I36407);
nand I_3880 (I67839,I68001,I68052);
DFFARX1 I_3881 (I36401,I2067,I67868,I68092,);
nor I_3882 (I68100,I68092,I68035);
DFFARX1 I_3883 (I68100,I2067,I67868,I67833,);
nor I_3884 (I67848,I68092,I67993);
nand I_3885 (I68145,I36389,I36386);
and I_3886 (I68162,I68145,I36398);
DFFARX1 I_3887 (I68162,I2067,I67868,I68188,);
nor I_3888 (I67836,I68188,I68092);
not I_3889 (I68210,I68188);
nor I_3890 (I68227,I68210,I68001);
nor I_3891 (I68244,I67933,I68227);
DFFARX1 I_3892 (I68244,I2067,I67868,I67851,);
nor I_3893 (I68275,I68210,I68092);
nor I_3894 (I68292,I36383,I36386);
nor I_3895 (I67842,I68292,I68275);
not I_3896 (I68323,I68292);
nand I_3897 (I67845,I68052,I68323);
DFFARX1 I_3898 (I68292,I2067,I67868,I67857,);
DFFARX1 I_3899 (I68292,I2067,I67868,I67854,);
not I_3900 (I68412,I2074);
DFFARX1 I_3901 (I58623,I2067,I68412,I68438,);
DFFARX1 I_3902 (I68438,I2067,I68412,I68455,);
not I_3903 (I68404,I68455);
not I_3904 (I68477,I68438);
nand I_3905 (I68494,I58602,I58626);
and I_3906 (I68511,I68494,I58629);
DFFARX1 I_3907 (I68511,I2067,I68412,I68537,);
not I_3908 (I68545,I68537);
DFFARX1 I_3909 (I58611,I2067,I68412,I68571,);
and I_3910 (I68579,I68571,I58617);
nand I_3911 (I68596,I68571,I58617);
nand I_3912 (I68383,I68545,I68596);
DFFARX1 I_3913 (I58605,I2067,I68412,I68636,);
nor I_3914 (I68644,I68636,I68579);
DFFARX1 I_3915 (I68644,I2067,I68412,I68377,);
nor I_3916 (I68392,I68636,I68537);
nand I_3917 (I68689,I58614,I58602);
and I_3918 (I68706,I68689,I58608);
DFFARX1 I_3919 (I68706,I2067,I68412,I68732,);
nor I_3920 (I68380,I68732,I68636);
not I_3921 (I68754,I68732);
nor I_3922 (I68771,I68754,I68545);
nor I_3923 (I68788,I68477,I68771);
DFFARX1 I_3924 (I68788,I2067,I68412,I68395,);
nor I_3925 (I68819,I68754,I68636);
nor I_3926 (I68836,I58620,I58602);
nor I_3927 (I68386,I68836,I68819);
not I_3928 (I68867,I68836);
nand I_3929 (I68389,I68596,I68867);
DFFARX1 I_3930 (I68836,I2067,I68412,I68401,);
DFFARX1 I_3931 (I68836,I2067,I68412,I68398,);
not I_3932 (I68953,I2074);
DFFARX1 I_3933 (I110240,I2067,I68953,I68979,);
DFFARX1 I_3934 (I68979,I2067,I68953,I68996,);
not I_3935 (I68945,I68996);
DFFARX1 I_3936 (I110237,I2067,I68953,I69027,);
not I_3937 (I69035,I110237);
nor I_3938 (I69052,I68979,I69035);
not I_3939 (I69069,I110234);
not I_3940 (I69086,I110249);
nand I_3941 (I69103,I69086,I110234);
nor I_3942 (I69120,I69035,I69103);
nor I_3943 (I69137,I69027,I69120);
DFFARX1 I_3944 (I69086,I2067,I68953,I68942,);
nor I_3945 (I69168,I110249,I110243);
nand I_3946 (I69185,I69168,I110231);
nor I_3947 (I69202,I69185,I69069);
nand I_3948 (I68927,I69202,I110237);
DFFARX1 I_3949 (I69185,I2067,I68953,I68939,);
nand I_3950 (I69247,I69069,I110249);
nor I_3951 (I69264,I69069,I110249);
nand I_3952 (I68933,I69052,I69264);
not I_3953 (I69295,I110252);
nor I_3954 (I69312,I69295,I69247);
DFFARX1 I_3955 (I69312,I2067,I68953,I68921,);
nor I_3956 (I69343,I69295,I110231);
and I_3957 (I69360,I69343,I110246);
or I_3958 (I69377,I69360,I110234);
DFFARX1 I_3959 (I69377,I2067,I68953,I69403,);
nor I_3960 (I69411,I69403,I69027);
nor I_3961 (I68930,I68979,I69411);
not I_3962 (I69442,I69403);
nor I_3963 (I69459,I69442,I69137);
DFFARX1 I_3964 (I69459,I2067,I68953,I68936,);
nand I_3965 (I69490,I69442,I69069);
nor I_3966 (I68924,I69295,I69490);
not I_3967 (I69548,I2074);
DFFARX1 I_3968 (I65113,I2067,I69548,I69574,);
DFFARX1 I_3969 (I69574,I2067,I69548,I69591,);
not I_3970 (I69540,I69591);
DFFARX1 I_3971 (I65137,I2067,I69548,I69622,);
not I_3972 (I69630,I65116);
nor I_3973 (I69647,I69574,I69630);
not I_3974 (I69664,I65122);
not I_3975 (I69681,I65128);
nand I_3976 (I69698,I69681,I65122);
nor I_3977 (I69715,I69630,I69698);
nor I_3978 (I69732,I69622,I69715);
DFFARX1 I_3979 (I69681,I2067,I69548,I69537,);
nor I_3980 (I69763,I65128,I65140);
nand I_3981 (I69780,I69763,I65134);
nor I_3982 (I69797,I69780,I69664);
nand I_3983 (I69522,I69797,I65116);
DFFARX1 I_3984 (I69780,I2067,I69548,I69534,);
nand I_3985 (I69842,I69664,I65128);
nor I_3986 (I69859,I69664,I65128);
nand I_3987 (I69528,I69647,I69859);
not I_3988 (I69890,I65119);
nor I_3989 (I69907,I69890,I69842);
DFFARX1 I_3990 (I69907,I2067,I69548,I69516,);
nor I_3991 (I69938,I69890,I65113);
and I_3992 (I69955,I69938,I65131);
or I_3993 (I69972,I69955,I65125);
DFFARX1 I_3994 (I69972,I2067,I69548,I69998,);
nor I_3995 (I70006,I69998,I69622);
nor I_3996 (I69525,I69574,I70006);
not I_3997 (I70037,I69998);
nor I_3998 (I70054,I70037,I69732);
DFFARX1 I_3999 (I70054,I2067,I69548,I69531,);
nand I_4000 (I70085,I70037,I69664);
nor I_4001 (I69519,I69890,I70085);
not I_4002 (I70143,I2074);
DFFARX1 I_4003 (I64025,I2067,I70143,I70169,);
DFFARX1 I_4004 (I70169,I2067,I70143,I70186,);
not I_4005 (I70135,I70186);
DFFARX1 I_4006 (I64049,I2067,I70143,I70217,);
not I_4007 (I70225,I64028);
nor I_4008 (I70242,I70169,I70225);
not I_4009 (I70259,I64034);
not I_4010 (I70276,I64040);
nand I_4011 (I70293,I70276,I64034);
nor I_4012 (I70310,I70225,I70293);
nor I_4013 (I70327,I70217,I70310);
DFFARX1 I_4014 (I70276,I2067,I70143,I70132,);
nor I_4015 (I70358,I64040,I64052);
nand I_4016 (I70375,I70358,I64046);
nor I_4017 (I70392,I70375,I70259);
nand I_4018 (I70117,I70392,I64028);
DFFARX1 I_4019 (I70375,I2067,I70143,I70129,);
nand I_4020 (I70437,I70259,I64040);
nor I_4021 (I70454,I70259,I64040);
nand I_4022 (I70123,I70242,I70454);
not I_4023 (I70485,I64031);
nor I_4024 (I70502,I70485,I70437);
DFFARX1 I_4025 (I70502,I2067,I70143,I70111,);
nor I_4026 (I70533,I70485,I64025);
and I_4027 (I70550,I70533,I64043);
or I_4028 (I70567,I70550,I64037);
DFFARX1 I_4029 (I70567,I2067,I70143,I70593,);
nor I_4030 (I70601,I70593,I70217);
nor I_4031 (I70120,I70169,I70601);
not I_4032 (I70632,I70593);
nor I_4033 (I70649,I70632,I70327);
DFFARX1 I_4034 (I70649,I2067,I70143,I70126,);
nand I_4035 (I70680,I70632,I70259);
nor I_4036 (I70114,I70485,I70680);
not I_4037 (I70738,I2074);
DFFARX1 I_4038 (I16978,I2067,I70738,I70764,);
DFFARX1 I_4039 (I70764,I2067,I70738,I70781,);
not I_4040 (I70730,I70781);
DFFARX1 I_4041 (I16990,I2067,I70738,I70812,);
not I_4042 (I70820,I16981);
nor I_4043 (I70837,I70764,I70820);
not I_4044 (I70854,I16972);
not I_4045 (I70871,I16969);
nand I_4046 (I70888,I70871,I16972);
nor I_4047 (I70905,I70820,I70888);
nor I_4048 (I70922,I70812,I70905);
DFFARX1 I_4049 (I70871,I2067,I70738,I70727,);
nor I_4050 (I70953,I16969,I16969);
nand I_4051 (I70970,I70953,I16987);
nor I_4052 (I70987,I70970,I70854);
nand I_4053 (I70712,I70987,I16981);
DFFARX1 I_4054 (I70970,I2067,I70738,I70724,);
nand I_4055 (I71032,I70854,I16969);
nor I_4056 (I71049,I70854,I16969);
nand I_4057 (I70718,I70837,I71049);
not I_4058 (I71080,I16993);
nor I_4059 (I71097,I71080,I71032);
DFFARX1 I_4060 (I71097,I2067,I70738,I70706,);
nor I_4061 (I71128,I71080,I16972);
and I_4062 (I71145,I71128,I16975);
or I_4063 (I71162,I71145,I16984);
DFFARX1 I_4064 (I71162,I2067,I70738,I71188,);
nor I_4065 (I71196,I71188,I70812);
nor I_4066 (I70715,I70764,I71196);
not I_4067 (I71227,I71188);
nor I_4068 (I71244,I71227,I70922);
DFFARX1 I_4069 (I71244,I2067,I70738,I70721,);
nand I_4070 (I71275,I71227,I70854);
nor I_4071 (I70709,I71080,I71275);
not I_4072 (I71333,I2074);
DFFARX1 I_4073 (I80739,I2067,I71333,I71359,);
DFFARX1 I_4074 (I71359,I2067,I71333,I71376,);
not I_4075 (I71325,I71376);
DFFARX1 I_4076 (I80751,I2067,I71333,I71407,);
not I_4077 (I71415,I80736);
nor I_4078 (I71432,I71359,I71415);
not I_4079 (I71449,I80754);
not I_4080 (I71466,I80745);
nand I_4081 (I71483,I71466,I80754);
nor I_4082 (I71500,I71415,I71483);
nor I_4083 (I71517,I71407,I71500);
DFFARX1 I_4084 (I71466,I2067,I71333,I71322,);
nor I_4085 (I71548,I80745,I80757);
nand I_4086 (I71565,I71548,I80760);
nor I_4087 (I71582,I71565,I71449);
nand I_4088 (I71307,I71582,I80736);
DFFARX1 I_4089 (I71565,I2067,I71333,I71319,);
nand I_4090 (I71627,I71449,I80745);
nor I_4091 (I71644,I71449,I80745);
nand I_4092 (I71313,I71432,I71644);
not I_4093 (I71675,I80736);
nor I_4094 (I71692,I71675,I71627);
DFFARX1 I_4095 (I71692,I2067,I71333,I71301,);
nor I_4096 (I71723,I71675,I80748);
and I_4097 (I71740,I71723,I80742);
or I_4098 (I71757,I71740,I80739);
DFFARX1 I_4099 (I71757,I2067,I71333,I71783,);
nor I_4100 (I71791,I71783,I71407);
nor I_4101 (I71310,I71359,I71791);
not I_4102 (I71822,I71783);
nor I_4103 (I71839,I71822,I71517);
DFFARX1 I_4104 (I71839,I2067,I71333,I71316,);
nand I_4105 (I71870,I71822,I71449);
nor I_4106 (I71304,I71675,I71870);
not I_4107 (I71928,I2074);
DFFARX1 I_4108 (I35788,I2067,I71928,I71954,);
DFFARX1 I_4109 (I71954,I2067,I71928,I71971,);
not I_4110 (I71920,I71971);
DFFARX1 I_4111 (I35812,I2067,I71928,I72002,);
not I_4112 (I72010,I35806);
nor I_4113 (I72027,I71954,I72010);
not I_4114 (I72044,I35800);
not I_4115 (I72061,I35797);
nand I_4116 (I72078,I72061,I35800);
nor I_4117 (I72095,I72010,I72078);
nor I_4118 (I72112,I72002,I72095);
DFFARX1 I_4119 (I72061,I2067,I71928,I71917,);
nor I_4120 (I72143,I35797,I35791);
nand I_4121 (I72160,I72143,I35809);
nor I_4122 (I72177,I72160,I72044);
nand I_4123 (I71902,I72177,I35806);
DFFARX1 I_4124 (I72160,I2067,I71928,I71914,);
nand I_4125 (I72222,I72044,I35797);
nor I_4126 (I72239,I72044,I35797);
nand I_4127 (I71908,I72027,I72239);
not I_4128 (I72270,I35803);
nor I_4129 (I72287,I72270,I72222);
DFFARX1 I_4130 (I72287,I2067,I71928,I71896,);
nor I_4131 (I72318,I72270,I35788);
and I_4132 (I72335,I72318,I35794);
or I_4133 (I72352,I72335,I35791);
DFFARX1 I_4134 (I72352,I2067,I71928,I72378,);
nor I_4135 (I72386,I72378,I72002);
nor I_4136 (I71905,I71954,I72386);
not I_4137 (I72417,I72378);
nor I_4138 (I72434,I72417,I72112);
DFFARX1 I_4139 (I72434,I2067,I71928,I71911,);
nand I_4140 (I72465,I72417,I72044);
nor I_4141 (I71899,I72270,I72465);
not I_4142 (I72523,I2074);
DFFARX1 I_4143 (I135119,I2067,I72523,I72549,);
DFFARX1 I_4144 (I72549,I2067,I72523,I72566,);
not I_4145 (I72515,I72566);
DFFARX1 I_4146 (I135122,I2067,I72523,I72597,);
not I_4147 (I72605,I135125);
nor I_4148 (I72622,I72549,I72605);
not I_4149 (I72639,I135137);
not I_4150 (I72656,I135128);
nand I_4151 (I72673,I72656,I135137);
nor I_4152 (I72690,I72605,I72673);
nor I_4153 (I72707,I72597,I72690);
DFFARX1 I_4154 (I72656,I2067,I72523,I72512,);
nor I_4155 (I72738,I135128,I135134);
nand I_4156 (I72755,I72738,I135122);
nor I_4157 (I72772,I72755,I72639);
nand I_4158 (I72497,I72772,I135125);
DFFARX1 I_4159 (I72755,I2067,I72523,I72509,);
nand I_4160 (I72817,I72639,I135128);
nor I_4161 (I72834,I72639,I135128);
nand I_4162 (I72503,I72622,I72834);
not I_4163 (I72865,I135125);
nor I_4164 (I72882,I72865,I72817);
DFFARX1 I_4165 (I72882,I2067,I72523,I72491,);
nor I_4166 (I72913,I72865,I135131);
and I_4167 (I72930,I72913,I135119);
or I_4168 (I72947,I72930,I135140);
DFFARX1 I_4169 (I72947,I2067,I72523,I72973,);
nor I_4170 (I72981,I72973,I72597);
nor I_4171 (I72500,I72549,I72981);
not I_4172 (I73012,I72973);
nor I_4173 (I73029,I73012,I72707);
DFFARX1 I_4174 (I73029,I2067,I72523,I72506,);
nand I_4175 (I73060,I73012,I72639);
nor I_4176 (I72494,I72865,I73060);
not I_4177 (I73118,I2074);
DFFARX1 I_4178 (I66745,I2067,I73118,I73144,);
DFFARX1 I_4179 (I73144,I2067,I73118,I73161,);
not I_4180 (I73110,I73161);
DFFARX1 I_4181 (I66769,I2067,I73118,I73192,);
not I_4182 (I73200,I66748);
nor I_4183 (I73217,I73144,I73200);
not I_4184 (I73234,I66754);
not I_4185 (I73251,I66760);
nand I_4186 (I73268,I73251,I66754);
nor I_4187 (I73285,I73200,I73268);
nor I_4188 (I73302,I73192,I73285);
DFFARX1 I_4189 (I73251,I2067,I73118,I73107,);
nor I_4190 (I73333,I66760,I66772);
nand I_4191 (I73350,I73333,I66766);
nor I_4192 (I73367,I73350,I73234);
nand I_4193 (I73092,I73367,I66748);
DFFARX1 I_4194 (I73350,I2067,I73118,I73104,);
nand I_4195 (I73412,I73234,I66760);
nor I_4196 (I73429,I73234,I66760);
nand I_4197 (I73098,I73217,I73429);
not I_4198 (I73460,I66751);
nor I_4199 (I73477,I73460,I73412);
DFFARX1 I_4200 (I73477,I2067,I73118,I73086,);
nor I_4201 (I73508,I73460,I66745);
and I_4202 (I73525,I73508,I66763);
or I_4203 (I73542,I73525,I66757);
DFFARX1 I_4204 (I73542,I2067,I73118,I73568,);
nor I_4205 (I73576,I73568,I73192);
nor I_4206 (I73095,I73144,I73576);
not I_4207 (I73607,I73568);
nor I_4208 (I73624,I73607,I73302);
DFFARX1 I_4209 (I73624,I2067,I73118,I73101,);
nand I_4210 (I73655,I73607,I73234);
nor I_4211 (I73089,I73460,I73655);
not I_4212 (I73713,I2074);
DFFARX1 I_4213 (I119749,I2067,I73713,I73739,);
DFFARX1 I_4214 (I73739,I2067,I73713,I73756,);
not I_4215 (I73705,I73756);
DFFARX1 I_4216 (I119737,I2067,I73713,I73787,);
not I_4217 (I73795,I119734);
nor I_4218 (I73812,I73739,I73795);
not I_4219 (I73829,I119746);
not I_4220 (I73846,I119743);
nand I_4221 (I73863,I73846,I119746);
nor I_4222 (I73880,I73795,I73863);
nor I_4223 (I73897,I73787,I73880);
DFFARX1 I_4224 (I73846,I2067,I73713,I73702,);
nor I_4225 (I73928,I119743,I119752);
nand I_4226 (I73945,I73928,I119755);
nor I_4227 (I73962,I73945,I73829);
nand I_4228 (I73687,I73962,I119734);
DFFARX1 I_4229 (I73945,I2067,I73713,I73699,);
nand I_4230 (I74007,I73829,I119743);
nor I_4231 (I74024,I73829,I119743);
nand I_4232 (I73693,I73812,I74024);
not I_4233 (I74055,I119758);
nor I_4234 (I74072,I74055,I74007);
DFFARX1 I_4235 (I74072,I2067,I73713,I73681,);
nor I_4236 (I74103,I74055,I119761);
and I_4237 (I74120,I74103,I119740);
or I_4238 (I74137,I74120,I119734);
DFFARX1 I_4239 (I74137,I2067,I73713,I74163,);
nor I_4240 (I74171,I74163,I73787);
nor I_4241 (I73690,I73739,I74171);
not I_4242 (I74202,I74163);
nor I_4243 (I74219,I74202,I73897);
DFFARX1 I_4244 (I74219,I2067,I73713,I73696,);
nand I_4245 (I74250,I74202,I73829);
nor I_4246 (I73684,I74055,I74250);
not I_4247 (I74308,I2074);
DFFARX1 I_4248 (I87103,I2067,I74308,I74334,);
DFFARX1 I_4249 (I74334,I2067,I74308,I74351,);
not I_4250 (I74300,I74351);
DFFARX1 I_4251 (I87097,I2067,I74308,I74382,);
not I_4252 (I74390,I87094);
nor I_4253 (I74407,I74334,I74390);
not I_4254 (I74424,I87106);
not I_4255 (I74441,I87109);
nand I_4256 (I74458,I74441,I87106);
nor I_4257 (I74475,I74390,I74458);
nor I_4258 (I74492,I74382,I74475);
DFFARX1 I_4259 (I74441,I2067,I74308,I74297,);
nor I_4260 (I74523,I87109,I87118);
nand I_4261 (I74540,I74523,I87112);
nor I_4262 (I74557,I74540,I74424);
nand I_4263 (I74282,I74557,I87094);
DFFARX1 I_4264 (I74540,I2067,I74308,I74294,);
nand I_4265 (I74602,I74424,I87109);
nor I_4266 (I74619,I74424,I87109);
nand I_4267 (I74288,I74407,I74619);
not I_4268 (I74650,I87100);
nor I_4269 (I74667,I74650,I74602);
DFFARX1 I_4270 (I74667,I2067,I74308,I74276,);
nor I_4271 (I74698,I74650,I87115);
and I_4272 (I74715,I74698,I87094);
or I_4273 (I74732,I74715,I87097);
DFFARX1 I_4274 (I74732,I2067,I74308,I74758,);
nor I_4275 (I74766,I74758,I74382);
nor I_4276 (I74285,I74334,I74766);
not I_4277 (I74797,I74758);
nor I_4278 (I74814,I74797,I74492);
DFFARX1 I_4279 (I74814,I2067,I74308,I74291,);
nand I_4280 (I74845,I74797,I74424);
nor I_4281 (I74279,I74650,I74845);
not I_4282 (I74903,I2074);
DFFARX1 I_4283 (I92883,I2067,I74903,I74929,);
DFFARX1 I_4284 (I74929,I2067,I74903,I74946,);
not I_4285 (I74895,I74946);
DFFARX1 I_4286 (I92877,I2067,I74903,I74977,);
not I_4287 (I74985,I92874);
nor I_4288 (I75002,I74929,I74985);
not I_4289 (I75019,I92886);
not I_4290 (I75036,I92889);
nand I_4291 (I75053,I75036,I92886);
nor I_4292 (I75070,I74985,I75053);
nor I_4293 (I75087,I74977,I75070);
DFFARX1 I_4294 (I75036,I2067,I74903,I74892,);
nor I_4295 (I75118,I92889,I92898);
nand I_4296 (I75135,I75118,I92892);
nor I_4297 (I75152,I75135,I75019);
nand I_4298 (I74877,I75152,I92874);
DFFARX1 I_4299 (I75135,I2067,I74903,I74889,);
nand I_4300 (I75197,I75019,I92889);
nor I_4301 (I75214,I75019,I92889);
nand I_4302 (I74883,I75002,I75214);
not I_4303 (I75245,I92880);
nor I_4304 (I75262,I75245,I75197);
DFFARX1 I_4305 (I75262,I2067,I74903,I74871,);
nor I_4306 (I75293,I75245,I92895);
and I_4307 (I75310,I75293,I92874);
or I_4308 (I75327,I75310,I92877);
DFFARX1 I_4309 (I75327,I2067,I74903,I75353,);
nor I_4310 (I75361,I75353,I74977);
nor I_4311 (I74880,I74929,I75361);
not I_4312 (I75392,I75353);
nor I_4313 (I75409,I75392,I75087);
DFFARX1 I_4314 (I75409,I2067,I74903,I74886,);
nand I_4315 (I75440,I75392,I75019);
nor I_4316 (I74874,I75245,I75440);
not I_4317 (I75498,I2074);
DFFARX1 I_4318 (I62393,I2067,I75498,I75524,);
DFFARX1 I_4319 (I75524,I2067,I75498,I75541,);
not I_4320 (I75490,I75541);
DFFARX1 I_4321 (I62417,I2067,I75498,I75572,);
not I_4322 (I75580,I62396);
nor I_4323 (I75597,I75524,I75580);
not I_4324 (I75614,I62402);
not I_4325 (I75631,I62408);
nand I_4326 (I75648,I75631,I62402);
nor I_4327 (I75665,I75580,I75648);
nor I_4328 (I75682,I75572,I75665);
DFFARX1 I_4329 (I75631,I2067,I75498,I75487,);
nor I_4330 (I75713,I62408,I62420);
nand I_4331 (I75730,I75713,I62414);
nor I_4332 (I75747,I75730,I75614);
nand I_4333 (I75472,I75747,I62396);
DFFARX1 I_4334 (I75730,I2067,I75498,I75484,);
nand I_4335 (I75792,I75614,I62408);
nor I_4336 (I75809,I75614,I62408);
nand I_4337 (I75478,I75597,I75809);
not I_4338 (I75840,I62399);
nor I_4339 (I75857,I75840,I75792);
DFFARX1 I_4340 (I75857,I2067,I75498,I75466,);
nor I_4341 (I75888,I75840,I62393);
and I_4342 (I75905,I75888,I62411);
or I_4343 (I75922,I75905,I62405);
DFFARX1 I_4344 (I75922,I2067,I75498,I75948,);
nor I_4345 (I75956,I75948,I75572);
nor I_4346 (I75475,I75524,I75956);
not I_4347 (I75987,I75948);
nor I_4348 (I76004,I75987,I75682);
DFFARX1 I_4349 (I76004,I2067,I75498,I75481,);
nand I_4350 (I76035,I75987,I75614);
nor I_4351 (I75469,I75840,I76035);
not I_4352 (I76093,I2074);
DFFARX1 I_4353 (I64569,I2067,I76093,I76119,);
DFFARX1 I_4354 (I76119,I2067,I76093,I76136,);
not I_4355 (I76085,I76136);
DFFARX1 I_4356 (I64593,I2067,I76093,I76167,);
not I_4357 (I76175,I64572);
nor I_4358 (I76192,I76119,I76175);
not I_4359 (I76209,I64578);
not I_4360 (I76226,I64584);
nand I_4361 (I76243,I76226,I64578);
nor I_4362 (I76260,I76175,I76243);
nor I_4363 (I76277,I76167,I76260);
DFFARX1 I_4364 (I76226,I2067,I76093,I76082,);
nor I_4365 (I76308,I64584,I64596);
nand I_4366 (I76325,I76308,I64590);
nor I_4367 (I76342,I76325,I76209);
nand I_4368 (I76067,I76342,I64572);
DFFARX1 I_4369 (I76325,I2067,I76093,I76079,);
nand I_4370 (I76387,I76209,I64584);
nor I_4371 (I76404,I76209,I64584);
nand I_4372 (I76073,I76192,I76404);
not I_4373 (I76435,I64575);
nor I_4374 (I76452,I76435,I76387);
DFFARX1 I_4375 (I76452,I2067,I76093,I76061,);
nor I_4376 (I76483,I76435,I64569);
and I_4377 (I76500,I76483,I64587);
or I_4378 (I76517,I76500,I64581);
DFFARX1 I_4379 (I76517,I2067,I76093,I76543,);
nor I_4380 (I76551,I76543,I76167);
nor I_4381 (I76070,I76119,I76551);
not I_4382 (I76582,I76543);
nor I_4383 (I76599,I76582,I76277);
DFFARX1 I_4384 (I76599,I2067,I76093,I76076,);
nand I_4385 (I76630,I76582,I76209);
nor I_4386 (I76064,I76435,I76630);
not I_4387 (I76688,I2074);
DFFARX1 I_4388 (I154074,I2067,I76688,I76714,);
DFFARX1 I_4389 (I76714,I2067,I76688,I76731,);
not I_4390 (I76680,I76731);
DFFARX1 I_4391 (I154089,I2067,I76688,I76762,);
not I_4392 (I76770,I154098);
nor I_4393 (I76787,I76714,I76770);
not I_4394 (I76804,I154077);
not I_4395 (I76821,I154083);
nand I_4396 (I76838,I76821,I154077);
nor I_4397 (I76855,I76770,I76838);
nor I_4398 (I76872,I76762,I76855);
DFFARX1 I_4399 (I76821,I2067,I76688,I76677,);
nor I_4400 (I76903,I154083,I154095);
nand I_4401 (I76920,I76903,I154092);
nor I_4402 (I76937,I76920,I76804);
nand I_4403 (I76662,I76937,I154098);
DFFARX1 I_4404 (I76920,I2067,I76688,I76674,);
nand I_4405 (I76982,I76804,I154083);
nor I_4406 (I76999,I76804,I154083);
nand I_4407 (I76668,I76787,I76999);
not I_4408 (I77030,I154074);
nor I_4409 (I77047,I77030,I76982);
DFFARX1 I_4410 (I77047,I2067,I76688,I76656,);
nor I_4411 (I77078,I77030,I154086);
and I_4412 (I77095,I77078,I154080);
or I_4413 (I77112,I77095,I154077);
DFFARX1 I_4414 (I77112,I2067,I76688,I77138,);
nor I_4415 (I77146,I77138,I76762);
nor I_4416 (I76665,I76714,I77146);
not I_4417 (I77177,I77138);
nor I_4418 (I77194,I77177,I76872);
DFFARX1 I_4419 (I77194,I2067,I76688,I76671,);
nand I_4420 (I77225,I77177,I76804);
nor I_4421 (I76659,I77030,I77225);
not I_4422 (I77283,I2074);
DFFARX1 I_4423 (I105497,I2067,I77283,I77309,);
DFFARX1 I_4424 (I77309,I2067,I77283,I77326,);
not I_4425 (I77275,I77326);
DFFARX1 I_4426 (I105494,I2067,I77283,I77357,);
not I_4427 (I77365,I105494);
nor I_4428 (I77382,I77309,I77365);
not I_4429 (I77399,I105491);
not I_4430 (I77416,I105506);
nand I_4431 (I77433,I77416,I105491);
nor I_4432 (I77450,I77365,I77433);
nor I_4433 (I77467,I77357,I77450);
DFFARX1 I_4434 (I77416,I2067,I77283,I77272,);
nor I_4435 (I77498,I105506,I105500);
nand I_4436 (I77515,I77498,I105488);
nor I_4437 (I77532,I77515,I77399);
nand I_4438 (I77257,I77532,I105494);
DFFARX1 I_4439 (I77515,I2067,I77283,I77269,);
nand I_4440 (I77577,I77399,I105506);
nor I_4441 (I77594,I77399,I105506);
nand I_4442 (I77263,I77382,I77594);
not I_4443 (I77625,I105509);
nor I_4444 (I77642,I77625,I77577);
DFFARX1 I_4445 (I77642,I2067,I77283,I77251,);
nor I_4446 (I77673,I77625,I105488);
and I_4447 (I77690,I77673,I105503);
or I_4448 (I77707,I77690,I105491);
DFFARX1 I_4449 (I77707,I2067,I77283,I77733,);
nor I_4450 (I77741,I77733,I77357);
nor I_4451 (I77260,I77309,I77741);
not I_4452 (I77772,I77733);
nor I_4453 (I77789,I77772,I77467);
DFFARX1 I_4454 (I77789,I2067,I77283,I77266,);
nand I_4455 (I77820,I77772,I77399);
nor I_4456 (I77254,I77625,I77820);
not I_4457 (I77878,I2074);
DFFARX1 I_4458 (I124908,I2067,I77878,I77904,);
not I_4459 (I77912,I77904);
DFFARX1 I_4460 (I124905,I2067,I77878,I77938,);
not I_4461 (I77946,I124902);
nand I_4462 (I77963,I77946,I124929);
not I_4463 (I77980,I77963);
nor I_4464 (I77997,I77980,I124917);
nor I_4465 (I78014,I77912,I77997);
DFFARX1 I_4466 (I78014,I2067,I77878,I77864,);
not I_4467 (I78045,I124917);
nand I_4468 (I78062,I78045,I77980);
and I_4469 (I78079,I78045,I124923);
nand I_4470 (I78096,I78079,I124914);
nor I_4471 (I77861,I78096,I78045);
and I_4472 (I77852,I77938,I78096);
not I_4473 (I78141,I78096);
nand I_4474 (I77855,I77938,I78141);
nor I_4475 (I77849,I77904,I78096);
not I_4476 (I78186,I124911);
nor I_4477 (I78203,I78186,I124923);
nand I_4478 (I78220,I78203,I78045);
nor I_4479 (I77858,I77963,I78220);
nor I_4480 (I78251,I78186,I124926);
and I_4481 (I78268,I78251,I124920);
or I_4482 (I78285,I78268,I124902);
DFFARX1 I_4483 (I78285,I2067,I77878,I78311,);
nor I_4484 (I78319,I78311,I78062);
DFFARX1 I_4485 (I78319,I2067,I77878,I77846,);
DFFARX1 I_4486 (I78311,I2067,I77878,I77870,);
not I_4487 (I78364,I78311);
nor I_4488 (I78381,I78364,I77938);
nor I_4489 (I78398,I78203,I78381);
DFFARX1 I_4490 (I78398,I2067,I77878,I77867,);
not I_4491 (I78456,I2074);
DFFARX1 I_4492 (I76064,I2067,I78456,I78482,);
not I_4493 (I78490,I78482);
DFFARX1 I_4494 (I76076,I2067,I78456,I78516,);
not I_4495 (I78524,I76082);
nand I_4496 (I78541,I78524,I76073);
not I_4497 (I78558,I78541);
nor I_4498 (I78575,I78558,I76079);
nor I_4499 (I78592,I78490,I78575);
DFFARX1 I_4500 (I78592,I2067,I78456,I78442,);
not I_4501 (I78623,I76079);
nand I_4502 (I78640,I78623,I78558);
and I_4503 (I78657,I78623,I76070);
nand I_4504 (I78674,I78657,I76061);
nor I_4505 (I78439,I78674,I78623);
and I_4506 (I78430,I78516,I78674);
not I_4507 (I78719,I78674);
nand I_4508 (I78433,I78516,I78719);
nor I_4509 (I78427,I78482,I78674);
not I_4510 (I78764,I76067);
nor I_4511 (I78781,I78764,I76070);
nand I_4512 (I78798,I78781,I78623);
nor I_4513 (I78436,I78541,I78798);
nor I_4514 (I78829,I78764,I76064);
and I_4515 (I78846,I78829,I76061);
or I_4516 (I78863,I78846,I76085);
DFFARX1 I_4517 (I78863,I2067,I78456,I78889,);
nor I_4518 (I78897,I78889,I78640);
DFFARX1 I_4519 (I78897,I2067,I78456,I78424,);
DFFARX1 I_4520 (I78889,I2067,I78456,I78448,);
not I_4521 (I78942,I78889);
nor I_4522 (I78959,I78942,I78516);
nor I_4523 (I78976,I78781,I78959);
DFFARX1 I_4524 (I78976,I2067,I78456,I78445,);
not I_4525 (I79034,I2074);
DFFARX1 I_4526 (I60229,I2067,I79034,I79060,);
not I_4527 (I79068,I79060);
DFFARX1 I_4528 (I60241,I2067,I79034,I79094,);
not I_4529 (I79102,I60217);
nand I_4530 (I79119,I79102,I60244);
not I_4531 (I79136,I79119);
nor I_4532 (I79153,I79136,I60232);
nor I_4533 (I79170,I79068,I79153);
DFFARX1 I_4534 (I79170,I2067,I79034,I79020,);
not I_4535 (I79201,I60232);
nand I_4536 (I79218,I79201,I79136);
and I_4537 (I79235,I79201,I60217);
nand I_4538 (I79252,I79235,I60220);
nor I_4539 (I79017,I79252,I79201);
and I_4540 (I79008,I79094,I79252);
not I_4541 (I79297,I79252);
nand I_4542 (I79011,I79094,I79297);
nor I_4543 (I79005,I79060,I79252);
not I_4544 (I79342,I60226);
nor I_4545 (I79359,I79342,I60217);
nand I_4546 (I79376,I79359,I79201);
nor I_4547 (I79014,I79119,I79376);
nor I_4548 (I79407,I79342,I60235);
and I_4549 (I79424,I79407,I60223);
or I_4550 (I79441,I79424,I60238);
DFFARX1 I_4551 (I79441,I2067,I79034,I79467,);
nor I_4552 (I79475,I79467,I79218);
DFFARX1 I_4553 (I79475,I2067,I79034,I79002,);
DFFARX1 I_4554 (I79467,I2067,I79034,I79026,);
not I_4555 (I79520,I79467);
nor I_4556 (I79537,I79520,I79094);
nor I_4557 (I79554,I79359,I79537);
DFFARX1 I_4558 (I79554,I2067,I79034,I79023,);
not I_4559 (I79612,I2074);
DFFARX1 I_4560 (I131774,I2067,I79612,I79638,);
not I_4561 (I79646,I79638);
DFFARX1 I_4562 (I131765,I2067,I79612,I79672,);
not I_4563 (I79680,I131759);
nand I_4564 (I79697,I79680,I131771);
not I_4565 (I79714,I79697);
nor I_4566 (I79731,I79714,I131762);
nor I_4567 (I79748,I79646,I79731);
DFFARX1 I_4568 (I79748,I2067,I79612,I79598,);
not I_4569 (I79779,I131762);
nand I_4570 (I79796,I79779,I79714);
and I_4571 (I79813,I79779,I131768);
nand I_4572 (I79830,I79813,I131753);
nor I_4573 (I79595,I79830,I79779);
and I_4574 (I79586,I79672,I79830);
not I_4575 (I79875,I79830);
nand I_4576 (I79589,I79672,I79875);
nor I_4577 (I79583,I79638,I79830);
not I_4578 (I79920,I131753);
nor I_4579 (I79937,I79920,I131768);
nand I_4580 (I79954,I79937,I79779);
nor I_4581 (I79592,I79697,I79954);
nor I_4582 (I79985,I79920,I131756);
and I_4583 (I80002,I79985,I131759);
or I_4584 (I80019,I80002,I131756);
DFFARX1 I_4585 (I80019,I2067,I79612,I80045,);
nor I_4586 (I80053,I80045,I79796);
DFFARX1 I_4587 (I80053,I2067,I79612,I79580,);
DFFARX1 I_4588 (I80045,I2067,I79612,I79604,);
not I_4589 (I80098,I80045);
nor I_4590 (I80115,I80098,I79672);
nor I_4591 (I80132,I79937,I80115);
DFFARX1 I_4592 (I80132,I2067,I79612,I79601,);
not I_4593 (I80190,I2074);
DFFARX1 I_4594 (I12250,I2067,I80190,I80216,);
not I_4595 (I80224,I80216);
DFFARX1 I_4596 (I12229,I2067,I80190,I80250,);
not I_4597 (I80258,I12226);
nand I_4598 (I80275,I80258,I12241);
not I_4599 (I80292,I80275);
nor I_4600 (I80309,I80292,I12229);
nor I_4601 (I80326,I80224,I80309);
DFFARX1 I_4602 (I80326,I2067,I80190,I80176,);
not I_4603 (I80357,I12229);
nand I_4604 (I80374,I80357,I80292);
and I_4605 (I80391,I80357,I12232);
nand I_4606 (I80408,I80391,I12247);
nor I_4607 (I80173,I80408,I80357);
and I_4608 (I80164,I80250,I80408);
not I_4609 (I80453,I80408);
nand I_4610 (I80167,I80250,I80453);
nor I_4611 (I80161,I80216,I80408);
not I_4612 (I80498,I12238);
nor I_4613 (I80515,I80498,I12232);
nand I_4614 (I80532,I80515,I80357);
nor I_4615 (I80170,I80275,I80532);
nor I_4616 (I80563,I80498,I12226);
and I_4617 (I80580,I80563,I12235);
or I_4618 (I80597,I80580,I12244);
DFFARX1 I_4619 (I80597,I2067,I80190,I80623,);
nor I_4620 (I80631,I80623,I80374);
DFFARX1 I_4621 (I80631,I2067,I80190,I80158,);
DFFARX1 I_4622 (I80623,I2067,I80190,I80182,);
not I_4623 (I80676,I80623);
nor I_4624 (I80693,I80676,I80250);
nor I_4625 (I80710,I80515,I80693);
DFFARX1 I_4626 (I80710,I2067,I80190,I80179,);
not I_4627 (I80768,I2074);
DFFARX1 I_4628 (I128138,I2067,I80768,I80794,);
not I_4629 (I80802,I80794);
DFFARX1 I_4630 (I128135,I2067,I80768,I80828,);
not I_4631 (I80836,I128132);
nand I_4632 (I80853,I80836,I128159);
not I_4633 (I80870,I80853);
nor I_4634 (I80887,I80870,I128147);
nor I_4635 (I80904,I80802,I80887);
DFFARX1 I_4636 (I80904,I2067,I80768,I80754,);
not I_4637 (I80935,I128147);
nand I_4638 (I80952,I80935,I80870);
and I_4639 (I80969,I80935,I128153);
nand I_4640 (I80986,I80969,I128144);
nor I_4641 (I80751,I80986,I80935);
and I_4642 (I80742,I80828,I80986);
not I_4643 (I81031,I80986);
nand I_4644 (I80745,I80828,I81031);
nor I_4645 (I80739,I80794,I80986);
not I_4646 (I81076,I128141);
nor I_4647 (I81093,I81076,I128153);
nand I_4648 (I81110,I81093,I80935);
nor I_4649 (I80748,I80853,I81110);
nor I_4650 (I81141,I81076,I128156);
and I_4651 (I81158,I81141,I128150);
or I_4652 (I81175,I81158,I128132);
DFFARX1 I_4653 (I81175,I2067,I80768,I81201,);
nor I_4654 (I81209,I81201,I80952);
DFFARX1 I_4655 (I81209,I2067,I80768,I80736,);
DFFARX1 I_4656 (I81201,I2067,I80768,I80760,);
not I_4657 (I81254,I81201);
nor I_4658 (I81271,I81254,I80828);
nor I_4659 (I81288,I81093,I81271);
DFFARX1 I_4660 (I81288,I2067,I80768,I80757,);
not I_4661 (I81346,I2074);
DFFARX1 I_4662 (I61861,I2067,I81346,I81372,);
not I_4663 (I81380,I81372);
DFFARX1 I_4664 (I61873,I2067,I81346,I81406,);
not I_4665 (I81414,I61849);
nand I_4666 (I81431,I81414,I61876);
not I_4667 (I81448,I81431);
nor I_4668 (I81465,I81448,I61864);
nor I_4669 (I81482,I81380,I81465);
DFFARX1 I_4670 (I81482,I2067,I81346,I81332,);
not I_4671 (I81513,I61864);
nand I_4672 (I81530,I81513,I81448);
and I_4673 (I81547,I81513,I61849);
nand I_4674 (I81564,I81547,I61852);
nor I_4675 (I81329,I81564,I81513);
and I_4676 (I81320,I81406,I81564);
not I_4677 (I81609,I81564);
nand I_4678 (I81323,I81406,I81609);
nor I_4679 (I81317,I81372,I81564);
not I_4680 (I81654,I61858);
nor I_4681 (I81671,I81654,I61849);
nand I_4682 (I81688,I81671,I81513);
nor I_4683 (I81326,I81431,I81688);
nor I_4684 (I81719,I81654,I61867);
and I_4685 (I81736,I81719,I61855);
or I_4686 (I81753,I81736,I61870);
DFFARX1 I_4687 (I81753,I2067,I81346,I81779,);
nor I_4688 (I81787,I81779,I81530);
DFFARX1 I_4689 (I81787,I2067,I81346,I81314,);
DFFARX1 I_4690 (I81779,I2067,I81346,I81338,);
not I_4691 (I81832,I81779);
nor I_4692 (I81849,I81832,I81406);
nor I_4693 (I81866,I81671,I81849);
DFFARX1 I_4694 (I81866,I2067,I81346,I81335,);
not I_4695 (I81924,I2074);
DFFARX1 I_4696 (I48595,I2067,I81924,I81950,);
not I_4697 (I81958,I81950);
DFFARX1 I_4698 (I48610,I2067,I81924,I81984,);
not I_4699 (I81992,I48613);
nand I_4700 (I82009,I81992,I48592);
not I_4701 (I82026,I82009);
nor I_4702 (I82043,I82026,I48616);
nor I_4703 (I82060,I81958,I82043);
DFFARX1 I_4704 (I82060,I2067,I81924,I81910,);
not I_4705 (I82091,I48616);
nand I_4706 (I82108,I82091,I82026);
and I_4707 (I82125,I82091,I48598);
nand I_4708 (I82142,I82125,I48589);
nor I_4709 (I81907,I82142,I82091);
and I_4710 (I81898,I81984,I82142);
not I_4711 (I82187,I82142);
nand I_4712 (I81901,I81984,I82187);
nor I_4713 (I81895,I81950,I82142);
not I_4714 (I82232,I48589);
nor I_4715 (I82249,I82232,I48598);
nand I_4716 (I82266,I82249,I82091);
nor I_4717 (I81904,I82009,I82266);
nor I_4718 (I82297,I82232,I48604);
and I_4719 (I82314,I82297,I48607);
or I_4720 (I82331,I82314,I48601);
DFFARX1 I_4721 (I82331,I2067,I81924,I82357,);
nor I_4722 (I82365,I82357,I82108);
DFFARX1 I_4723 (I82365,I2067,I81924,I81892,);
DFFARX1 I_4724 (I82357,I2067,I81924,I81916,);
not I_4725 (I82410,I82357);
nor I_4726 (I82427,I82410,I81984);
nor I_4727 (I82444,I82249,I82427);
DFFARX1 I_4728 (I82444,I2067,I81924,I81913,);
not I_4729 (I82502,I2074);
DFFARX1 I_4730 (I122970,I2067,I82502,I82528,);
not I_4731 (I82536,I82528);
DFFARX1 I_4732 (I122967,I2067,I82502,I82562,);
not I_4733 (I82570,I122964);
nand I_4734 (I82587,I82570,I122991);
not I_4735 (I82604,I82587);
nor I_4736 (I82621,I82604,I122979);
nor I_4737 (I82638,I82536,I82621);
DFFARX1 I_4738 (I82638,I2067,I82502,I82488,);
not I_4739 (I82669,I122979);
nand I_4740 (I82686,I82669,I82604);
and I_4741 (I82703,I82669,I122985);
nand I_4742 (I82720,I82703,I122976);
nor I_4743 (I82485,I82720,I82669);
and I_4744 (I82476,I82562,I82720);
not I_4745 (I82765,I82720);
nand I_4746 (I82479,I82562,I82765);
nor I_4747 (I82473,I82528,I82720);
not I_4748 (I82810,I122973);
nor I_4749 (I82827,I82810,I122985);
nand I_4750 (I82844,I82827,I82669);
nor I_4751 (I82482,I82587,I82844);
nor I_4752 (I82875,I82810,I122988);
and I_4753 (I82892,I82875,I122982);
or I_4754 (I82909,I82892,I122964);
DFFARX1 I_4755 (I82909,I2067,I82502,I82935,);
nor I_4756 (I82943,I82935,I82686);
DFFARX1 I_4757 (I82943,I2067,I82502,I82470,);
DFFARX1 I_4758 (I82935,I2067,I82502,I82494,);
not I_4759 (I82988,I82935);
nor I_4760 (I83005,I82988,I82562);
nor I_4761 (I83022,I82827,I83005);
DFFARX1 I_4762 (I83022,I2067,I82502,I82491,);
not I_4763 (I83080,I2074);
DFFARX1 I_4764 (I175239,I2067,I83080,I83106,);
not I_4765 (I83114,I83106);
DFFARX1 I_4766 (I175239,I2067,I83080,I83140,);
not I_4767 (I83148,I175263);
nand I_4768 (I83165,I83148,I175245);
not I_4769 (I83182,I83165);
nor I_4770 (I83199,I83182,I175260);
nor I_4771 (I83216,I83114,I83199);
DFFARX1 I_4772 (I83216,I2067,I83080,I83066,);
not I_4773 (I83247,I175260);
nand I_4774 (I83264,I83247,I83182);
and I_4775 (I83281,I83247,I175242);
nand I_4776 (I83298,I83281,I175251);
nor I_4777 (I83063,I83298,I83247);
and I_4778 (I83054,I83140,I83298);
not I_4779 (I83343,I83298);
nand I_4780 (I83057,I83140,I83343);
nor I_4781 (I83051,I83106,I83298);
not I_4782 (I83388,I175248);
nor I_4783 (I83405,I83388,I175242);
nand I_4784 (I83422,I83405,I83247);
nor I_4785 (I83060,I83165,I83422);
nor I_4786 (I83453,I83388,I175257);
and I_4787 (I83470,I83453,I175266);
or I_4788 (I83487,I83470,I175254);
DFFARX1 I_4789 (I83487,I2067,I83080,I83513,);
nor I_4790 (I83521,I83513,I83264);
DFFARX1 I_4791 (I83521,I2067,I83080,I83048,);
DFFARX1 I_4792 (I83513,I2067,I83080,I83072,);
not I_4793 (I83566,I83513);
nor I_4794 (I83583,I83566,I83140);
nor I_4795 (I83600,I83405,I83583);
DFFARX1 I_4796 (I83600,I2067,I83080,I83069,);
not I_4797 (I83658,I2074);
DFFARX1 I_4798 (I144894,I2067,I83658,I83684,);
not I_4799 (I83692,I83684);
DFFARX1 I_4800 (I144900,I2067,I83658,I83718,);
not I_4801 (I83726,I144894);
nand I_4802 (I83743,I83726,I144897);
not I_4803 (I83760,I83743);
nor I_4804 (I83777,I83760,I144915);
nor I_4805 (I83794,I83692,I83777);
DFFARX1 I_4806 (I83794,I2067,I83658,I83644,);
not I_4807 (I83825,I144915);
nand I_4808 (I83842,I83825,I83760);
and I_4809 (I83859,I83825,I144918);
nand I_4810 (I83876,I83859,I144897);
nor I_4811 (I83641,I83876,I83825);
and I_4812 (I83632,I83718,I83876);
not I_4813 (I83921,I83876);
nand I_4814 (I83635,I83718,I83921);
nor I_4815 (I83629,I83684,I83876);
not I_4816 (I83966,I144903);
nor I_4817 (I83983,I83966,I144918);
nand I_4818 (I84000,I83983,I83825);
nor I_4819 (I83638,I83743,I84000);
nor I_4820 (I84031,I83966,I144909);
and I_4821 (I84048,I84031,I144906);
or I_4822 (I84065,I84048,I144912);
DFFARX1 I_4823 (I84065,I2067,I83658,I84091,);
nor I_4824 (I84099,I84091,I83842);
DFFARX1 I_4825 (I84099,I2067,I83658,I83626,);
DFFARX1 I_4826 (I84091,I2067,I83658,I83650,);
not I_4827 (I84144,I84091);
nor I_4828 (I84161,I84144,I83718);
nor I_4829 (I84178,I83983,I84161);
DFFARX1 I_4830 (I84178,I2067,I83658,I83647,);
not I_4831 (I84236,I2074);
DFFARX1 I_4832 (I159532,I2067,I84236,I84262,);
not I_4833 (I84270,I84262);
DFFARX1 I_4834 (I159526,I2067,I84236,I84296,);
not I_4835 (I84304,I159535);
nand I_4836 (I84321,I84304,I159514);
not I_4837 (I84338,I84321);
nor I_4838 (I84355,I84338,I159523);
nor I_4839 (I84372,I84270,I84355);
DFFARX1 I_4840 (I84372,I2067,I84236,I84222,);
not I_4841 (I84403,I159523);
nand I_4842 (I84420,I84403,I84338);
and I_4843 (I84437,I84403,I159538);
nand I_4844 (I84454,I84437,I159517);
nor I_4845 (I84219,I84454,I84403);
and I_4846 (I84210,I84296,I84454);
not I_4847 (I84499,I84454);
nand I_4848 (I84213,I84296,I84499);
nor I_4849 (I84207,I84262,I84454);
not I_4850 (I84544,I159520);
nor I_4851 (I84561,I84544,I159538);
nand I_4852 (I84578,I84561,I84403);
nor I_4853 (I84216,I84321,I84578);
nor I_4854 (I84609,I84544,I159529);
and I_4855 (I84626,I84609,I159517);
or I_4856 (I84643,I84626,I159514);
DFFARX1 I_4857 (I84643,I2067,I84236,I84669,);
nor I_4858 (I84677,I84669,I84420);
DFFARX1 I_4859 (I84677,I2067,I84236,I84204,);
DFFARX1 I_4860 (I84669,I2067,I84236,I84228,);
not I_4861 (I84722,I84669);
nor I_4862 (I84739,I84722,I84296);
nor I_4863 (I84756,I84561,I84739);
DFFARX1 I_4864 (I84756,I2067,I84236,I84225,);
not I_4865 (I84814,I2074);
DFFARX1 I_4866 (I161770,I2067,I84814,I84840,);
not I_4867 (I84848,I84840);
DFFARX1 I_4868 (I161782,I2067,I84814,I84874,);
not I_4869 (I84882,I161773);
nand I_4870 (I84899,I84882,I161761);
not I_4871 (I84916,I84899);
nor I_4872 (I84933,I84916,I161758);
nor I_4873 (I84950,I84848,I84933);
DFFARX1 I_4874 (I84950,I2067,I84814,I84800,);
not I_4875 (I84981,I161758);
nand I_4876 (I84998,I84981,I84916);
and I_4877 (I85015,I84981,I161764);
nand I_4878 (I85032,I85015,I161761);
nor I_4879 (I84797,I85032,I84981);
and I_4880 (I84788,I84874,I85032);
not I_4881 (I85077,I85032);
nand I_4882 (I84791,I84874,I85077);
nor I_4883 (I84785,I84840,I85032);
not I_4884 (I85122,I161779);
nor I_4885 (I85139,I85122,I161764);
nand I_4886 (I85156,I85139,I84981);
nor I_4887 (I84794,I84899,I85156);
nor I_4888 (I85187,I85122,I161767);
and I_4889 (I85204,I85187,I161758);
or I_4890 (I85221,I85204,I161776);
DFFARX1 I_4891 (I85221,I2067,I84814,I85247,);
nor I_4892 (I85255,I85247,I84998);
DFFARX1 I_4893 (I85255,I2067,I84814,I84782,);
DFFARX1 I_4894 (I85247,I2067,I84814,I84806,);
not I_4895 (I85300,I85247);
nor I_4896 (I85317,I85300,I84874);
nor I_4897 (I85334,I85139,I85317);
DFFARX1 I_4898 (I85334,I2067,I84814,I84803,);
not I_4899 (I85392,I2074);
DFFARX1 I_4900 (I94608,I2067,I85392,I85418,);
not I_4901 (I85426,I85418);
DFFARX1 I_4902 (I94620,I2067,I85392,I85452,);
not I_4903 (I85460,I94611);
nand I_4904 (I85477,I85460,I94614);
not I_4905 (I85494,I85477);
nor I_4906 (I85511,I85494,I94617);
nor I_4907 (I85528,I85426,I85511);
DFFARX1 I_4908 (I85528,I2067,I85392,I85378,);
not I_4909 (I85559,I94617);
nand I_4910 (I85576,I85559,I85494);
and I_4911 (I85593,I85559,I94611);
nand I_4912 (I85610,I85593,I94623);
nor I_4913 (I85375,I85610,I85559);
and I_4914 (I85366,I85452,I85610);
not I_4915 (I85655,I85610);
nand I_4916 (I85369,I85452,I85655);
nor I_4917 (I85363,I85418,I85610);
not I_4918 (I85700,I94629);
nor I_4919 (I85717,I85700,I94611);
nand I_4920 (I85734,I85717,I85559);
nor I_4921 (I85372,I85477,I85734);
nor I_4922 (I85765,I85700,I94608);
and I_4923 (I85782,I85765,I94626);
or I_4924 (I85799,I85782,I94632);
DFFARX1 I_4925 (I85799,I2067,I85392,I85825,);
nor I_4926 (I85833,I85825,I85576);
DFFARX1 I_4927 (I85833,I2067,I85392,I85360,);
DFFARX1 I_4928 (I85825,I2067,I85392,I85384,);
not I_4929 (I85878,I85825);
nor I_4930 (I85895,I85878,I85452);
nor I_4931 (I85912,I85717,I85895);
DFFARX1 I_4932 (I85912,I2067,I85392,I85381,);
not I_4933 (I85970,I2074);
DFFARX1 I_4934 (I4324,I2067,I85970,I85996,);
not I_4935 (I86004,I85996);
DFFARX1 I_4936 (I4327,I2067,I85970,I86030,);
not I_4937 (I86038,I4321);
nand I_4938 (I86055,I86038,I4345);
not I_4939 (I86072,I86055);
nor I_4940 (I86089,I86072,I4324);
nor I_4941 (I86106,I86004,I86089);
DFFARX1 I_4942 (I86106,I2067,I85970,I85956,);
not I_4943 (I86137,I4324);
nand I_4944 (I86154,I86137,I86072);
and I_4945 (I86171,I86137,I4339);
nand I_4946 (I86188,I86171,I4333);
nor I_4947 (I85953,I86188,I86137);
and I_4948 (I85944,I86030,I86188);
not I_4949 (I86233,I86188);
nand I_4950 (I85947,I86030,I86233);
nor I_4951 (I85941,I85996,I86188);
not I_4952 (I86278,I4342);
nor I_4953 (I86295,I86278,I4339);
nand I_4954 (I86312,I86295,I86137);
nor I_4955 (I85950,I86055,I86312);
nor I_4956 (I86343,I86278,I4321);
and I_4957 (I86360,I86343,I4330);
or I_4958 (I86377,I86360,I4336);
DFFARX1 I_4959 (I86377,I2067,I85970,I86403,);
nor I_4960 (I86411,I86403,I86154);
DFFARX1 I_4961 (I86411,I2067,I85970,I85938,);
DFFARX1 I_4962 (I86403,I2067,I85970,I85962,);
not I_4963 (I86456,I86403);
nor I_4964 (I86473,I86456,I86030);
nor I_4965 (I86490,I86295,I86473);
DFFARX1 I_4966 (I86490,I2067,I85970,I85959,);
not I_4967 (I86548,I2074);
DFFARX1 I_4968 (I13810,I2067,I86548,I86574,);
not I_4969 (I86582,I86574);
nand I_4970 (I86599,I13819,I13828);
and I_4971 (I86616,I86599,I13807);
DFFARX1 I_4972 (I86616,I2067,I86548,I86642,);
not I_4973 (I86650,I13810);
DFFARX1 I_4974 (I13825,I2067,I86548,I86676,);
not I_4975 (I86684,I86676);
nor I_4976 (I86701,I86684,I86582);
and I_4977 (I86718,I86701,I13810);
nor I_4978 (I86735,I86684,I86650);
nor I_4979 (I86531,I86642,I86735);
DFFARX1 I_4980 (I13816,I2067,I86548,I86775,);
nor I_4981 (I86783,I86775,I86642);
not I_4982 (I86800,I86783);
not I_4983 (I86817,I86775);
nor I_4984 (I86834,I86817,I86718);
DFFARX1 I_4985 (I86834,I2067,I86548,I86534,);
nand I_4986 (I86865,I13831,I13807);
and I_4987 (I86882,I86865,I13813);
DFFARX1 I_4988 (I86882,I2067,I86548,I86908,);
nor I_4989 (I86916,I86908,I86775);
DFFARX1 I_4990 (I86916,I2067,I86548,I86516,);
nand I_4991 (I86947,I86908,I86817);
nand I_4992 (I86525,I86800,I86947);
not I_4993 (I86978,I86908);
nor I_4994 (I86995,I86978,I86718);
DFFARX1 I_4995 (I86995,I2067,I86548,I86537,);
nor I_4996 (I87026,I13822,I13807);
or I_4997 (I86528,I86775,I87026);
nor I_4998 (I86519,I86908,I87026);
or I_4999 (I86522,I86642,I87026);
DFFARX1 I_5000 (I87026,I2067,I86548,I86540,);
not I_5001 (I87126,I2074);
DFFARX1 I_5002 (I119112,I2067,I87126,I87152,);
not I_5003 (I87160,I87152);
nand I_5004 (I87177,I119088,I119103);
and I_5005 (I87194,I87177,I119115);
DFFARX1 I_5006 (I87194,I2067,I87126,I87220,);
not I_5007 (I87228,I119100);
DFFARX1 I_5008 (I119091,I2067,I87126,I87254,);
not I_5009 (I87262,I87254);
nor I_5010 (I87279,I87262,I87160);
and I_5011 (I87296,I87279,I119100);
nor I_5012 (I87313,I87262,I87228);
nor I_5013 (I87109,I87220,I87313);
DFFARX1 I_5014 (I119088,I2067,I87126,I87353,);
nor I_5015 (I87361,I87353,I87220);
not I_5016 (I87378,I87361);
not I_5017 (I87395,I87353);
nor I_5018 (I87412,I87395,I87296);
DFFARX1 I_5019 (I87412,I2067,I87126,I87112,);
nand I_5020 (I87443,I119106,I119097);
and I_5021 (I87460,I87443,I119109);
DFFARX1 I_5022 (I87460,I2067,I87126,I87486,);
nor I_5023 (I87494,I87486,I87353);
DFFARX1 I_5024 (I87494,I2067,I87126,I87094,);
nand I_5025 (I87525,I87486,I87395);
nand I_5026 (I87103,I87378,I87525);
not I_5027 (I87556,I87486);
nor I_5028 (I87573,I87556,I87296);
DFFARX1 I_5029 (I87573,I2067,I87126,I87115,);
nor I_5030 (I87604,I119094,I119097);
or I_5031 (I87106,I87353,I87604);
nor I_5032 (I87097,I87486,I87604);
or I_5033 (I87100,I87220,I87604);
DFFARX1 I_5034 (I87604,I2067,I87126,I87118,);
not I_5035 (I87704,I2074);
DFFARX1 I_5036 (I166397,I2067,I87704,I87730,);
not I_5037 (I87738,I87730);
nand I_5038 (I87755,I166385,I166403);
and I_5039 (I87772,I87755,I166394);
DFFARX1 I_5040 (I87772,I2067,I87704,I87798,);
not I_5041 (I87806,I166409);
DFFARX1 I_5042 (I166406,I2067,I87704,I87832,);
not I_5043 (I87840,I87832);
nor I_5044 (I87857,I87840,I87738);
and I_5045 (I87874,I87857,I166409);
nor I_5046 (I87891,I87840,I87806);
nor I_5047 (I87687,I87798,I87891);
DFFARX1 I_5048 (I166388,I2067,I87704,I87931,);
nor I_5049 (I87939,I87931,I87798);
not I_5050 (I87956,I87939);
not I_5051 (I87973,I87931);
nor I_5052 (I87990,I87973,I87874);
DFFARX1 I_5053 (I87990,I2067,I87704,I87690,);
nand I_5054 (I88021,I166382,I166382);
and I_5055 (I88038,I88021,I166391);
DFFARX1 I_5056 (I88038,I2067,I87704,I88064,);
nor I_5057 (I88072,I88064,I87931);
DFFARX1 I_5058 (I88072,I2067,I87704,I87672,);
nand I_5059 (I88103,I88064,I87973);
nand I_5060 (I87681,I87956,I88103);
not I_5061 (I88134,I88064);
nor I_5062 (I88151,I88134,I87874);
DFFARX1 I_5063 (I88151,I2067,I87704,I87693,);
nor I_5064 (I88182,I166400,I166382);
or I_5065 (I87684,I87931,I88182);
nor I_5066 (I87675,I88064,I88182);
or I_5067 (I87678,I87798,I88182);
DFFARX1 I_5068 (I88182,I2067,I87704,I87696,);
not I_5069 (I88282,I2074);
DFFARX1 I_5070 (I121696,I2067,I88282,I88308,);
not I_5071 (I88316,I88308);
nand I_5072 (I88333,I121672,I121687);
and I_5073 (I88350,I88333,I121699);
DFFARX1 I_5074 (I88350,I2067,I88282,I88376,);
not I_5075 (I88384,I121684);
DFFARX1 I_5076 (I121675,I2067,I88282,I88410,);
not I_5077 (I88418,I88410);
nor I_5078 (I88435,I88418,I88316);
and I_5079 (I88452,I88435,I121684);
nor I_5080 (I88469,I88418,I88384);
nor I_5081 (I88265,I88376,I88469);
DFFARX1 I_5082 (I121672,I2067,I88282,I88509,);
nor I_5083 (I88517,I88509,I88376);
not I_5084 (I88534,I88517);
not I_5085 (I88551,I88509);
nor I_5086 (I88568,I88551,I88452);
DFFARX1 I_5087 (I88568,I2067,I88282,I88268,);
nand I_5088 (I88599,I121690,I121681);
and I_5089 (I88616,I88599,I121693);
DFFARX1 I_5090 (I88616,I2067,I88282,I88642,);
nor I_5091 (I88650,I88642,I88509);
DFFARX1 I_5092 (I88650,I2067,I88282,I88250,);
nand I_5093 (I88681,I88642,I88551);
nand I_5094 (I88259,I88534,I88681);
not I_5095 (I88712,I88642);
nor I_5096 (I88729,I88712,I88452);
DFFARX1 I_5097 (I88729,I2067,I88282,I88271,);
nor I_5098 (I88760,I121678,I121681);
or I_5099 (I88262,I88509,I88760);
nor I_5100 (I88253,I88642,I88760);
or I_5101 (I88256,I88376,I88760);
DFFARX1 I_5102 (I88760,I2067,I88282,I88274,);
not I_5103 (I88860,I2074);
DFFARX1 I_5104 (I122342,I2067,I88860,I88886,);
not I_5105 (I88894,I88886);
nand I_5106 (I88911,I122318,I122333);
and I_5107 (I88928,I88911,I122345);
DFFARX1 I_5108 (I88928,I2067,I88860,I88954,);
not I_5109 (I88962,I122330);
DFFARX1 I_5110 (I122321,I2067,I88860,I88988,);
not I_5111 (I88996,I88988);
nor I_5112 (I89013,I88996,I88894);
and I_5113 (I89030,I89013,I122330);
nor I_5114 (I89047,I88996,I88962);
nor I_5115 (I88843,I88954,I89047);
DFFARX1 I_5116 (I122318,I2067,I88860,I89087,);
nor I_5117 (I89095,I89087,I88954);
not I_5118 (I89112,I89095);
not I_5119 (I89129,I89087);
nor I_5120 (I89146,I89129,I89030);
DFFARX1 I_5121 (I89146,I2067,I88860,I88846,);
nand I_5122 (I89177,I122336,I122327);
and I_5123 (I89194,I89177,I122339);
DFFARX1 I_5124 (I89194,I2067,I88860,I89220,);
nor I_5125 (I89228,I89220,I89087);
DFFARX1 I_5126 (I89228,I2067,I88860,I88828,);
nand I_5127 (I89259,I89220,I89129);
nand I_5128 (I88837,I89112,I89259);
not I_5129 (I89290,I89220);
nor I_5130 (I89307,I89290,I89030);
DFFARX1 I_5131 (I89307,I2067,I88860,I88849,);
nor I_5132 (I89338,I122324,I122327);
or I_5133 (I88840,I89087,I89338);
nor I_5134 (I88831,I89220,I89338);
or I_5135 (I88834,I88954,I89338);
DFFARX1 I_5136 (I89338,I2067,I88860,I88852,);
not I_5137 (I89438,I2074);
DFFARX1 I_5138 (I44924,I2067,I89438,I89464,);
not I_5139 (I89472,I89464);
nand I_5140 (I89489,I44927,I44903);
and I_5141 (I89506,I89489,I44900);
DFFARX1 I_5142 (I89506,I2067,I89438,I89532,);
not I_5143 (I89540,I44906);
DFFARX1 I_5144 (I44900,I2067,I89438,I89566,);
not I_5145 (I89574,I89566);
nor I_5146 (I89591,I89574,I89472);
and I_5147 (I89608,I89591,I44906);
nor I_5148 (I89625,I89574,I89540);
nor I_5149 (I89421,I89532,I89625);
DFFARX1 I_5150 (I44909,I2067,I89438,I89665,);
nor I_5151 (I89673,I89665,I89532);
not I_5152 (I89690,I89673);
not I_5153 (I89707,I89665);
nor I_5154 (I89724,I89707,I89608);
DFFARX1 I_5155 (I89724,I2067,I89438,I89424,);
nand I_5156 (I89755,I44912,I44921);
and I_5157 (I89772,I89755,I44918);
DFFARX1 I_5158 (I89772,I2067,I89438,I89798,);
nor I_5159 (I89806,I89798,I89665);
DFFARX1 I_5160 (I89806,I2067,I89438,I89406,);
nand I_5161 (I89837,I89798,I89707);
nand I_5162 (I89415,I89690,I89837);
not I_5163 (I89868,I89798);
nor I_5164 (I89885,I89868,I89608);
DFFARX1 I_5165 (I89885,I2067,I89438,I89427,);
nor I_5166 (I89916,I44915,I44921);
or I_5167 (I89418,I89665,I89916);
nor I_5168 (I89409,I89798,I89916);
or I_5169 (I89412,I89532,I89916);
DFFARX1 I_5170 (I89916,I2067,I89438,I89430,);
not I_5171 (I90016,I2074);
DFFARX1 I_5172 (I77251,I2067,I90016,I90042,);
not I_5173 (I90050,I90042);
nand I_5174 (I90067,I77266,I77251);
and I_5175 (I90084,I90067,I77254);
DFFARX1 I_5176 (I90084,I2067,I90016,I90110,);
not I_5177 (I90118,I77254);
DFFARX1 I_5178 (I77263,I2067,I90016,I90144,);
not I_5179 (I90152,I90144);
nor I_5180 (I90169,I90152,I90050);
and I_5181 (I90186,I90169,I77254);
nor I_5182 (I90203,I90152,I90118);
nor I_5183 (I89999,I90110,I90203);
DFFARX1 I_5184 (I77257,I2067,I90016,I90243,);
nor I_5185 (I90251,I90243,I90110);
not I_5186 (I90268,I90251);
not I_5187 (I90285,I90243);
nor I_5188 (I90302,I90285,I90186);
DFFARX1 I_5189 (I90302,I2067,I90016,I90002,);
nand I_5190 (I90333,I77260,I77269);
and I_5191 (I90350,I90333,I77275);
DFFARX1 I_5192 (I90350,I2067,I90016,I90376,);
nor I_5193 (I90384,I90376,I90243);
DFFARX1 I_5194 (I90384,I2067,I90016,I89984,);
nand I_5195 (I90415,I90376,I90285);
nand I_5196 (I89993,I90268,I90415);
not I_5197 (I90446,I90376);
nor I_5198 (I90463,I90446,I90186);
DFFARX1 I_5199 (I90463,I2067,I90016,I90005,);
nor I_5200 (I90494,I77272,I77269);
or I_5201 (I89996,I90243,I90494);
nor I_5202 (I89987,I90376,I90494);
or I_5203 (I89990,I90110,I90494);
DFFARX1 I_5204 (I90494,I2067,I90016,I90008,);
not I_5205 (I90594,I2074);
DFFARX1 I_5206 (I31623,I2067,I90594,I90620,);
not I_5207 (I90628,I90620);
nand I_5208 (I90645,I31626,I31647);
and I_5209 (I90662,I90645,I31635);
DFFARX1 I_5210 (I90662,I2067,I90594,I90688,);
not I_5211 (I90696,I31632);
DFFARX1 I_5212 (I31623,I2067,I90594,I90722,);
not I_5213 (I90730,I90722);
nor I_5214 (I90747,I90730,I90628);
and I_5215 (I90764,I90747,I31632);
nor I_5216 (I90781,I90730,I90696);
nor I_5217 (I90577,I90688,I90781);
DFFARX1 I_5218 (I31641,I2067,I90594,I90821,);
nor I_5219 (I90829,I90821,I90688);
not I_5220 (I90846,I90829);
not I_5221 (I90863,I90821);
nor I_5222 (I90880,I90863,I90764);
DFFARX1 I_5223 (I90880,I2067,I90594,I90580,);
nand I_5224 (I90911,I31626,I31629);
and I_5225 (I90928,I90911,I31638);
DFFARX1 I_5226 (I90928,I2067,I90594,I90954,);
nor I_5227 (I90962,I90954,I90821);
DFFARX1 I_5228 (I90962,I2067,I90594,I90562,);
nand I_5229 (I90993,I90954,I90863);
nand I_5230 (I90571,I90846,I90993);
not I_5231 (I91024,I90954);
nor I_5232 (I91041,I91024,I90764);
DFFARX1 I_5233 (I91041,I2067,I90594,I90583,);
nor I_5234 (I91072,I31644,I31629);
or I_5235 (I90574,I90821,I91072);
nor I_5236 (I90565,I90954,I91072);
or I_5237 (I90568,I90688,I91072);
DFFARX1 I_5238 (I91072,I2067,I90594,I90586,);
not I_5239 (I91172,I2074);
DFFARX1 I_5240 (I42289,I2067,I91172,I91198,);
not I_5241 (I91206,I91198);
nand I_5242 (I91223,I42292,I42268);
and I_5243 (I91240,I91223,I42265);
DFFARX1 I_5244 (I91240,I2067,I91172,I91266,);
not I_5245 (I91274,I42271);
DFFARX1 I_5246 (I42265,I2067,I91172,I91300,);
not I_5247 (I91308,I91300);
nor I_5248 (I91325,I91308,I91206);
and I_5249 (I91342,I91325,I42271);
nor I_5250 (I91359,I91308,I91274);
nor I_5251 (I91155,I91266,I91359);
DFFARX1 I_5252 (I42274,I2067,I91172,I91399,);
nor I_5253 (I91407,I91399,I91266);
not I_5254 (I91424,I91407);
not I_5255 (I91441,I91399);
nor I_5256 (I91458,I91441,I91342);
DFFARX1 I_5257 (I91458,I2067,I91172,I91158,);
nand I_5258 (I91489,I42277,I42286);
and I_5259 (I91506,I91489,I42283);
DFFARX1 I_5260 (I91506,I2067,I91172,I91532,);
nor I_5261 (I91540,I91532,I91399);
DFFARX1 I_5262 (I91540,I2067,I91172,I91140,);
nand I_5263 (I91571,I91532,I91441);
nand I_5264 (I91149,I91424,I91571);
not I_5265 (I91602,I91532);
nor I_5266 (I91619,I91602,I91342);
DFFARX1 I_5267 (I91619,I2067,I91172,I91161,);
nor I_5268 (I91650,I42280,I42286);
or I_5269 (I91152,I91399,I91650);
nor I_5270 (I91143,I91532,I91650);
or I_5271 (I91146,I91266,I91650);
DFFARX1 I_5272 (I91650,I2067,I91172,I91164,);
not I_5273 (I91750,I2074);
DFFARX1 I_5274 (I132881,I2067,I91750,I91776,);
not I_5275 (I91784,I91776);
nand I_5276 (I91801,I132878,I132896);
and I_5277 (I91818,I91801,I132893);
DFFARX1 I_5278 (I91818,I2067,I91750,I91844,);
not I_5279 (I91852,I132875);
DFFARX1 I_5280 (I132878,I2067,I91750,I91878,);
not I_5281 (I91886,I91878);
nor I_5282 (I91903,I91886,I91784);
and I_5283 (I91920,I91903,I132875);
nor I_5284 (I91937,I91886,I91852);
nor I_5285 (I91733,I91844,I91937);
DFFARX1 I_5286 (I132887,I2067,I91750,I91977,);
nor I_5287 (I91985,I91977,I91844);
not I_5288 (I92002,I91985);
not I_5289 (I92019,I91977);
nor I_5290 (I92036,I92019,I91920);
DFFARX1 I_5291 (I92036,I2067,I91750,I91736,);
nand I_5292 (I92067,I132890,I132875);
and I_5293 (I92084,I92067,I132881);
DFFARX1 I_5294 (I92084,I2067,I91750,I92110,);
nor I_5295 (I92118,I92110,I91977);
DFFARX1 I_5296 (I92118,I2067,I91750,I91718,);
nand I_5297 (I92149,I92110,I92019);
nand I_5298 (I91727,I92002,I92149);
not I_5299 (I92180,I92110);
nor I_5300 (I92197,I92180,I91920);
DFFARX1 I_5301 (I92197,I2067,I91750,I91739,);
nor I_5302 (I92228,I132884,I132875);
or I_5303 (I91730,I91977,I92228);
nor I_5304 (I91721,I92110,I92228);
or I_5305 (I91724,I91844,I92228);
DFFARX1 I_5306 (I92228,I2067,I91750,I91742,);
not I_5307 (I92328,I2074);
DFFARX1 I_5308 (I20661,I2067,I92328,I92354,);
not I_5309 (I92362,I92354);
nand I_5310 (I92379,I20670,I20679);
and I_5311 (I92396,I92379,I20658);
DFFARX1 I_5312 (I92396,I2067,I92328,I92422,);
not I_5313 (I92430,I20661);
DFFARX1 I_5314 (I20676,I2067,I92328,I92456,);
not I_5315 (I92464,I92456);
nor I_5316 (I92481,I92464,I92362);
and I_5317 (I92498,I92481,I20661);
nor I_5318 (I92515,I92464,I92430);
nor I_5319 (I92311,I92422,I92515);
DFFARX1 I_5320 (I20667,I2067,I92328,I92555,);
nor I_5321 (I92563,I92555,I92422);
not I_5322 (I92580,I92563);
not I_5323 (I92597,I92555);
nor I_5324 (I92614,I92597,I92498);
DFFARX1 I_5325 (I92614,I2067,I92328,I92314,);
nand I_5326 (I92645,I20682,I20658);
and I_5327 (I92662,I92645,I20664);
DFFARX1 I_5328 (I92662,I2067,I92328,I92688,);
nor I_5329 (I92696,I92688,I92555);
DFFARX1 I_5330 (I92696,I2067,I92328,I92296,);
nand I_5331 (I92727,I92688,I92597);
nand I_5332 (I92305,I92580,I92727);
not I_5333 (I92758,I92688);
nor I_5334 (I92775,I92758,I92498);
DFFARX1 I_5335 (I92775,I2067,I92328,I92317,);
nor I_5336 (I92806,I20673,I20658);
or I_5337 (I92308,I92555,I92806);
nor I_5338 (I92299,I92688,I92806);
or I_5339 (I92302,I92422,I92806);
DFFARX1 I_5340 (I92806,I2067,I92328,I92320,);
not I_5341 (I92906,I2074);
DFFARX1 I_5342 (I116528,I2067,I92906,I92932,);
not I_5343 (I92940,I92932);
nand I_5344 (I92957,I116504,I116519);
and I_5345 (I92974,I92957,I116531);
DFFARX1 I_5346 (I92974,I2067,I92906,I93000,);
not I_5347 (I93008,I116516);
DFFARX1 I_5348 (I116507,I2067,I92906,I93034,);
not I_5349 (I93042,I93034);
nor I_5350 (I93059,I93042,I92940);
and I_5351 (I93076,I93059,I116516);
nor I_5352 (I93093,I93042,I93008);
nor I_5353 (I92889,I93000,I93093);
DFFARX1 I_5354 (I116504,I2067,I92906,I93133,);
nor I_5355 (I93141,I93133,I93000);
not I_5356 (I93158,I93141);
not I_5357 (I93175,I93133);
nor I_5358 (I93192,I93175,I93076);
DFFARX1 I_5359 (I93192,I2067,I92906,I92892,);
nand I_5360 (I93223,I116522,I116513);
and I_5361 (I93240,I93223,I116525);
DFFARX1 I_5362 (I93240,I2067,I92906,I93266,);
nor I_5363 (I93274,I93266,I93133);
DFFARX1 I_5364 (I93274,I2067,I92906,I92874,);
nand I_5365 (I93305,I93266,I93175);
nand I_5366 (I92883,I93158,I93305);
not I_5367 (I93336,I93266);
nor I_5368 (I93353,I93336,I93076);
DFFARX1 I_5369 (I93353,I2067,I92906,I92895,);
nor I_5370 (I93384,I116510,I116513);
or I_5371 (I92886,I93133,I93384);
nor I_5372 (I92877,I93266,I93384);
or I_5373 (I92880,I93000,I93384);
DFFARX1 I_5374 (I93384,I2067,I92906,I92898,);
not I_5375 (I93484,I2074);
DFFARX1 I_5376 (I129448,I2067,I93484,I93510,);
not I_5377 (I93518,I93510);
nand I_5378 (I93535,I129424,I129439);
and I_5379 (I93552,I93535,I129451);
DFFARX1 I_5380 (I93552,I2067,I93484,I93578,);
not I_5381 (I93586,I129436);
DFFARX1 I_5382 (I129427,I2067,I93484,I93612,);
not I_5383 (I93620,I93612);
nor I_5384 (I93637,I93620,I93518);
and I_5385 (I93654,I93637,I129436);
nor I_5386 (I93671,I93620,I93586);
nor I_5387 (I93467,I93578,I93671);
DFFARX1 I_5388 (I129424,I2067,I93484,I93711,);
nor I_5389 (I93719,I93711,I93578);
not I_5390 (I93736,I93719);
not I_5391 (I93753,I93711);
nor I_5392 (I93770,I93753,I93654);
DFFARX1 I_5393 (I93770,I2067,I93484,I93470,);
nand I_5394 (I93801,I129442,I129433);
and I_5395 (I93818,I93801,I129445);
DFFARX1 I_5396 (I93818,I2067,I93484,I93844,);
nor I_5397 (I93852,I93844,I93711);
DFFARX1 I_5398 (I93852,I2067,I93484,I93452,);
nand I_5399 (I93883,I93844,I93753);
nand I_5400 (I93461,I93736,I93883);
not I_5401 (I93914,I93844);
nor I_5402 (I93931,I93914,I93654);
DFFARX1 I_5403 (I93931,I2067,I93484,I93473,);
nor I_5404 (I93962,I129430,I129433);
or I_5405 (I93464,I93711,I93962);
nor I_5406 (I93455,I93844,I93962);
or I_5407 (I93458,I93578,I93962);
DFFARX1 I_5408 (I93962,I2067,I93484,I93476,);
not I_5409 (I94062,I2074);
DFFARX1 I_5410 (I29838,I2067,I94062,I94088,);
not I_5411 (I94096,I94088);
nand I_5412 (I94113,I29841,I29862);
and I_5413 (I94130,I94113,I29850);
DFFARX1 I_5414 (I94130,I2067,I94062,I94156,);
not I_5415 (I94164,I29847);
DFFARX1 I_5416 (I29838,I2067,I94062,I94190,);
not I_5417 (I94198,I94190);
nor I_5418 (I94215,I94198,I94096);
and I_5419 (I94232,I94215,I29847);
nor I_5420 (I94249,I94198,I94164);
nor I_5421 (I94045,I94156,I94249);
DFFARX1 I_5422 (I29856,I2067,I94062,I94289,);
nor I_5423 (I94297,I94289,I94156);
not I_5424 (I94314,I94297);
not I_5425 (I94331,I94289);
nor I_5426 (I94348,I94331,I94232);
DFFARX1 I_5427 (I94348,I2067,I94062,I94048,);
nand I_5428 (I94379,I29841,I29844);
and I_5429 (I94396,I94379,I29853);
DFFARX1 I_5430 (I94396,I2067,I94062,I94422,);
nor I_5431 (I94430,I94422,I94289);
DFFARX1 I_5432 (I94430,I2067,I94062,I94030,);
nand I_5433 (I94461,I94422,I94331);
nand I_5434 (I94039,I94314,I94461);
not I_5435 (I94492,I94422);
nor I_5436 (I94509,I94492,I94232);
DFFARX1 I_5437 (I94509,I2067,I94062,I94051,);
nor I_5438 (I94540,I29859,I29844);
or I_5439 (I94042,I94289,I94540);
nor I_5440 (I94033,I94422,I94540);
or I_5441 (I94036,I94156,I94540);
DFFARX1 I_5442 (I94540,I2067,I94062,I94054,);
not I_5443 (I94640,I2074);
DFFARX1 I_5444 (I148958,I2067,I94640,I94666,);
not I_5445 (I94674,I94666);
nand I_5446 (I94691,I148940,I148952);
and I_5447 (I94708,I94691,I148955);
DFFARX1 I_5448 (I94708,I2067,I94640,I94734,);
not I_5449 (I94742,I148949);
DFFARX1 I_5450 (I148946,I2067,I94640,I94768,);
not I_5451 (I94776,I94768);
nor I_5452 (I94793,I94776,I94674);
and I_5453 (I94810,I94793,I148949);
nor I_5454 (I94827,I94776,I94742);
nor I_5455 (I94623,I94734,I94827);
DFFARX1 I_5456 (I148964,I2067,I94640,I94867,);
nor I_5457 (I94875,I94867,I94734);
not I_5458 (I94892,I94875);
not I_5459 (I94909,I94867);
nor I_5460 (I94926,I94909,I94810);
DFFARX1 I_5461 (I94926,I2067,I94640,I94626,);
nand I_5462 (I94957,I148943,I148943);
and I_5463 (I94974,I94957,I148940);
DFFARX1 I_5464 (I94974,I2067,I94640,I95000,);
nor I_5465 (I95008,I95000,I94867);
DFFARX1 I_5466 (I95008,I2067,I94640,I94608,);
nand I_5467 (I95039,I95000,I94909);
nand I_5468 (I94617,I94892,I95039);
not I_5469 (I95070,I95000);
nor I_5470 (I95087,I95070,I94810);
DFFARX1 I_5471 (I95087,I2067,I94640,I94629,);
nor I_5472 (I95118,I148961,I148943);
or I_5473 (I94620,I94867,I95118);
nor I_5474 (I94611,I95000,I95118);
or I_5475 (I94614,I94734,I95118);
DFFARX1 I_5476 (I95118,I2067,I94640,I94632,);
not I_5477 (I95218,I2074);
DFFARX1 I_5478 (I71301,I2067,I95218,I95244,);
not I_5479 (I95252,I95244);
nand I_5480 (I95269,I71316,I71301);
and I_5481 (I95286,I95269,I71304);
DFFARX1 I_5482 (I95286,I2067,I95218,I95312,);
not I_5483 (I95320,I71304);
DFFARX1 I_5484 (I71313,I2067,I95218,I95346,);
not I_5485 (I95354,I95346);
nor I_5486 (I95371,I95354,I95252);
and I_5487 (I95388,I95371,I71304);
nor I_5488 (I95405,I95354,I95320);
nor I_5489 (I95201,I95312,I95405);
DFFARX1 I_5490 (I71307,I2067,I95218,I95445,);
nor I_5491 (I95453,I95445,I95312);
not I_5492 (I95470,I95453);
not I_5493 (I95487,I95445);
nor I_5494 (I95504,I95487,I95388);
DFFARX1 I_5495 (I95504,I2067,I95218,I95204,);
nand I_5496 (I95535,I71310,I71319);
and I_5497 (I95552,I95535,I71325);
DFFARX1 I_5498 (I95552,I2067,I95218,I95578,);
nor I_5499 (I95586,I95578,I95445);
DFFARX1 I_5500 (I95586,I2067,I95218,I95186,);
nand I_5501 (I95617,I95578,I95487);
nand I_5502 (I95195,I95470,I95617);
not I_5503 (I95648,I95578);
nor I_5504 (I95665,I95648,I95388);
DFFARX1 I_5505 (I95665,I2067,I95218,I95207,);
nor I_5506 (I95696,I71322,I71319);
or I_5507 (I95198,I95445,I95696);
nor I_5508 (I95189,I95578,I95696);
or I_5509 (I95192,I95312,I95696);
DFFARX1 I_5510 (I95696,I2067,I95218,I95210,);
not I_5511 (I95796,I2074);
DFFARX1 I_5512 (I177646,I2067,I95796,I95822,);
not I_5513 (I95830,I95822);
nand I_5514 (I95847,I177631,I177619);
and I_5515 (I95864,I95847,I177634);
DFFARX1 I_5516 (I95864,I2067,I95796,I95890,);
not I_5517 (I95898,I177619);
DFFARX1 I_5518 (I177637,I2067,I95796,I95924,);
not I_5519 (I95932,I95924);
nor I_5520 (I95949,I95932,I95830);
and I_5521 (I95966,I95949,I177619);
nor I_5522 (I95983,I95932,I95898);
nor I_5523 (I95779,I95890,I95983);
DFFARX1 I_5524 (I177625,I2067,I95796,I96023,);
nor I_5525 (I96031,I96023,I95890);
not I_5526 (I96048,I96031);
not I_5527 (I96065,I96023);
nor I_5528 (I96082,I96065,I95966);
DFFARX1 I_5529 (I96082,I2067,I95796,I95782,);
nand I_5530 (I96113,I177622,I177628);
and I_5531 (I96130,I96113,I177643);
DFFARX1 I_5532 (I96130,I2067,I95796,I96156,);
nor I_5533 (I96164,I96156,I96023);
DFFARX1 I_5534 (I96164,I2067,I95796,I95764,);
nand I_5535 (I96195,I96156,I96065);
nand I_5536 (I95773,I96048,I96195);
not I_5537 (I96226,I96156);
nor I_5538 (I96243,I96226,I95966);
DFFARX1 I_5539 (I96243,I2067,I95796,I95785,);
nor I_5540 (I96274,I177640,I177628);
or I_5541 (I95776,I96023,I96274);
nor I_5542 (I95767,I96156,I96274);
or I_5543 (I95770,I95890,I96274);
DFFARX1 I_5544 (I96274,I2067,I95796,I95788,);
not I_5545 (I96374,I2074);
DFFARX1 I_5546 (I52829,I2067,I96374,I96400,);
not I_5547 (I96408,I96400);
nand I_5548 (I96425,I52832,I52808);
and I_5549 (I96442,I96425,I52805);
DFFARX1 I_5550 (I96442,I2067,I96374,I96468,);
not I_5551 (I96476,I52811);
DFFARX1 I_5552 (I52805,I2067,I96374,I96502,);
not I_5553 (I96510,I96502);
nor I_5554 (I96527,I96510,I96408);
and I_5555 (I96544,I96527,I52811);
nor I_5556 (I96561,I96510,I96476);
nor I_5557 (I96357,I96468,I96561);
DFFARX1 I_5558 (I52814,I2067,I96374,I96601,);
nor I_5559 (I96609,I96601,I96468);
not I_5560 (I96626,I96609);
not I_5561 (I96643,I96601);
nor I_5562 (I96660,I96643,I96544);
DFFARX1 I_5563 (I96660,I2067,I96374,I96360,);
nand I_5564 (I96691,I52817,I52826);
and I_5565 (I96708,I96691,I52823);
DFFARX1 I_5566 (I96708,I2067,I96374,I96734,);
nor I_5567 (I96742,I96734,I96601);
DFFARX1 I_5568 (I96742,I2067,I96374,I96342,);
nand I_5569 (I96773,I96734,I96643);
nand I_5570 (I96351,I96626,I96773);
not I_5571 (I96804,I96734);
nor I_5572 (I96821,I96804,I96544);
DFFARX1 I_5573 (I96821,I2067,I96374,I96363,);
nor I_5574 (I96852,I52820,I52826);
or I_5575 (I96354,I96601,I96852);
nor I_5576 (I96345,I96734,I96852);
or I_5577 (I96348,I96468,I96852);
DFFARX1 I_5578 (I96852,I2067,I96374,I96366,);
not I_5579 (I96952,I2074);
DFFARX1 I_5580 (I51248,I2067,I96952,I96978,);
not I_5581 (I96986,I96978);
nand I_5582 (I97003,I51251,I51227);
and I_5583 (I97020,I97003,I51224);
DFFARX1 I_5584 (I97020,I2067,I96952,I97046,);
not I_5585 (I97054,I51230);
DFFARX1 I_5586 (I51224,I2067,I96952,I97080,);
not I_5587 (I97088,I97080);
nor I_5588 (I97105,I97088,I96986);
and I_5589 (I97122,I97105,I51230);
nor I_5590 (I97139,I97088,I97054);
nor I_5591 (I96935,I97046,I97139);
DFFARX1 I_5592 (I51233,I2067,I96952,I97179,);
nor I_5593 (I97187,I97179,I97046);
not I_5594 (I97204,I97187);
not I_5595 (I97221,I97179);
nor I_5596 (I97238,I97221,I97122);
DFFARX1 I_5597 (I97238,I2067,I96952,I96938,);
nand I_5598 (I97269,I51236,I51245);
and I_5599 (I97286,I97269,I51242);
DFFARX1 I_5600 (I97286,I2067,I96952,I97312,);
nor I_5601 (I97320,I97312,I97179);
DFFARX1 I_5602 (I97320,I2067,I96952,I96920,);
nand I_5603 (I97351,I97312,I97221);
nand I_5604 (I96929,I97204,I97351);
not I_5605 (I97382,I97312);
nor I_5606 (I97399,I97382,I97122);
DFFARX1 I_5607 (I97399,I2067,I96952,I96941,);
nor I_5608 (I97430,I51239,I51245);
or I_5609 (I96932,I97179,I97430);
nor I_5610 (I96923,I97312,I97430);
or I_5611 (I96926,I97046,I97430);
DFFARX1 I_5612 (I97430,I2067,I96952,I96944,);
not I_5613 (I97530,I2074);
DFFARX1 I_5614 (I133442,I2067,I97530,I97556,);
not I_5615 (I97564,I97556);
nand I_5616 (I97581,I133439,I133457);
and I_5617 (I97598,I97581,I133454);
DFFARX1 I_5618 (I97598,I2067,I97530,I97624,);
not I_5619 (I97632,I133436);
DFFARX1 I_5620 (I133439,I2067,I97530,I97658,);
not I_5621 (I97666,I97658);
nor I_5622 (I97683,I97666,I97564);
and I_5623 (I97700,I97683,I133436);
nor I_5624 (I97717,I97666,I97632);
nor I_5625 (I97513,I97624,I97717);
DFFARX1 I_5626 (I133448,I2067,I97530,I97757,);
nor I_5627 (I97765,I97757,I97624);
not I_5628 (I97782,I97765);
not I_5629 (I97799,I97757);
nor I_5630 (I97816,I97799,I97700);
DFFARX1 I_5631 (I97816,I2067,I97530,I97516,);
nand I_5632 (I97847,I133451,I133436);
and I_5633 (I97864,I97847,I133442);
DFFARX1 I_5634 (I97864,I2067,I97530,I97890,);
nor I_5635 (I97898,I97890,I97757);
DFFARX1 I_5636 (I97898,I2067,I97530,I97498,);
nand I_5637 (I97929,I97890,I97799);
nand I_5638 (I97507,I97782,I97929);
not I_5639 (I97960,I97890);
nor I_5640 (I97977,I97960,I97700);
DFFARX1 I_5641 (I97977,I2067,I97530,I97519,);
nor I_5642 (I98008,I133445,I133436);
or I_5643 (I97510,I97757,I98008);
nor I_5644 (I97501,I97890,I98008);
or I_5645 (I97504,I97624,I98008);
DFFARX1 I_5646 (I98008,I2067,I97530,I97522,);
not I_5647 (I98108,I2074);
DFFARX1 I_5648 (I126218,I2067,I98108,I98134,);
not I_5649 (I98142,I98134);
nand I_5650 (I98159,I126194,I126209);
and I_5651 (I98176,I98159,I126221);
DFFARX1 I_5652 (I98176,I2067,I98108,I98202,);
not I_5653 (I98210,I126206);
DFFARX1 I_5654 (I126197,I2067,I98108,I98236,);
not I_5655 (I98244,I98236);
nor I_5656 (I98261,I98244,I98142);
and I_5657 (I98278,I98261,I126206);
nor I_5658 (I98295,I98244,I98210);
nor I_5659 (I98091,I98202,I98295);
DFFARX1 I_5660 (I126194,I2067,I98108,I98335,);
nor I_5661 (I98343,I98335,I98202);
not I_5662 (I98360,I98343);
not I_5663 (I98377,I98335);
nor I_5664 (I98394,I98377,I98278);
DFFARX1 I_5665 (I98394,I2067,I98108,I98094,);
nand I_5666 (I98425,I126212,I126203);
and I_5667 (I98442,I98425,I126215);
DFFARX1 I_5668 (I98442,I2067,I98108,I98468,);
nor I_5669 (I98476,I98468,I98335);
DFFARX1 I_5670 (I98476,I2067,I98108,I98076,);
nand I_5671 (I98507,I98468,I98377);
nand I_5672 (I98085,I98360,I98507);
not I_5673 (I98538,I98468);
nor I_5674 (I98555,I98538,I98278);
DFFARX1 I_5675 (I98555,I2067,I98108,I98097,);
nor I_5676 (I98586,I126200,I126203);
or I_5677 (I98088,I98335,I98586);
nor I_5678 (I98079,I98468,I98586);
or I_5679 (I98082,I98202,I98586);
DFFARX1 I_5680 (I98586,I2067,I98108,I98100,);
not I_5681 (I98686,I2074);
DFFARX1 I_5682 (I14864,I2067,I98686,I98712,);
not I_5683 (I98720,I98712);
nand I_5684 (I98737,I14873,I14882);
and I_5685 (I98754,I98737,I14861);
DFFARX1 I_5686 (I98754,I2067,I98686,I98780,);
not I_5687 (I98788,I14864);
DFFARX1 I_5688 (I14879,I2067,I98686,I98814,);
not I_5689 (I98822,I98814);
nor I_5690 (I98839,I98822,I98720);
and I_5691 (I98856,I98839,I14864);
nor I_5692 (I98873,I98822,I98788);
nor I_5693 (I98669,I98780,I98873);
DFFARX1 I_5694 (I14870,I2067,I98686,I98913,);
nor I_5695 (I98921,I98913,I98780);
not I_5696 (I98938,I98921);
not I_5697 (I98955,I98913);
nor I_5698 (I98972,I98955,I98856);
DFFARX1 I_5699 (I98972,I2067,I98686,I98672,);
nand I_5700 (I99003,I14885,I14861);
and I_5701 (I99020,I99003,I14867);
DFFARX1 I_5702 (I99020,I2067,I98686,I99046,);
nor I_5703 (I99054,I99046,I98913);
DFFARX1 I_5704 (I99054,I2067,I98686,I98654,);
nand I_5705 (I99085,I99046,I98955);
nand I_5706 (I98663,I98938,I99085);
not I_5707 (I99116,I99046);
nor I_5708 (I99133,I99116,I98856);
DFFARX1 I_5709 (I99133,I2067,I98686,I98675,);
nor I_5710 (I99164,I14876,I14861);
or I_5711 (I98666,I98913,I99164);
nor I_5712 (I98657,I99046,I99164);
or I_5713 (I98660,I98780,I99164);
DFFARX1 I_5714 (I99164,I2067,I98686,I98678,);
not I_5715 (I99264,I2074);
DFFARX1 I_5716 (I137976,I2067,I99264,I99290,);
not I_5717 (I99298,I99290);
nand I_5718 (I99315,I137958,I137970);
and I_5719 (I99332,I99315,I137973);
DFFARX1 I_5720 (I99332,I2067,I99264,I99358,);
not I_5721 (I99366,I137967);
DFFARX1 I_5722 (I137964,I2067,I99264,I99392,);
not I_5723 (I99400,I99392);
nor I_5724 (I99417,I99400,I99298);
and I_5725 (I99434,I99417,I137967);
nor I_5726 (I99451,I99400,I99366);
nor I_5727 (I99247,I99358,I99451);
DFFARX1 I_5728 (I137982,I2067,I99264,I99491,);
nor I_5729 (I99499,I99491,I99358);
not I_5730 (I99516,I99499);
not I_5731 (I99533,I99491);
nor I_5732 (I99550,I99533,I99434);
DFFARX1 I_5733 (I99550,I2067,I99264,I99250,);
nand I_5734 (I99581,I137961,I137961);
and I_5735 (I99598,I99581,I137958);
DFFARX1 I_5736 (I99598,I2067,I99264,I99624,);
nor I_5737 (I99632,I99624,I99491);
DFFARX1 I_5738 (I99632,I2067,I99264,I99232,);
nand I_5739 (I99663,I99624,I99533);
nand I_5740 (I99241,I99516,I99663);
not I_5741 (I99694,I99624);
nor I_5742 (I99711,I99694,I99434);
DFFARX1 I_5743 (I99711,I2067,I99264,I99253,);
nor I_5744 (I99742,I137979,I137961);
or I_5745 (I99244,I99491,I99742);
nor I_5746 (I99235,I99624,I99742);
or I_5747 (I99238,I99358,I99742);
DFFARX1 I_5748 (I99742,I2067,I99264,I99256,);
not I_5749 (I99842,I2074);
DFFARX1 I_5750 (I158970,I2067,I99842,I99868,);
not I_5751 (I99876,I99868);
nand I_5752 (I99893,I158973,I158982);
and I_5753 (I99910,I99893,I158985);
DFFARX1 I_5754 (I99910,I2067,I99842,I99936,);
not I_5755 (I99944,I158994);
DFFARX1 I_5756 (I158976,I2067,I99842,I99970,);
not I_5757 (I99978,I99970);
nor I_5758 (I99995,I99978,I99876);
and I_5759 (I100012,I99995,I158994);
nor I_5760 (I100029,I99978,I99944);
nor I_5761 (I99825,I99936,I100029);
DFFARX1 I_5762 (I158973,I2067,I99842,I100069,);
nor I_5763 (I100077,I100069,I99936);
not I_5764 (I100094,I100077);
not I_5765 (I100111,I100069);
nor I_5766 (I100128,I100111,I100012);
DFFARX1 I_5767 (I100128,I2067,I99842,I99828,);
nand I_5768 (I100159,I158991,I158970);
and I_5769 (I100176,I100159,I158988);
DFFARX1 I_5770 (I100176,I2067,I99842,I100202,);
nor I_5771 (I100210,I100202,I100069);
DFFARX1 I_5772 (I100210,I2067,I99842,I99810,);
nand I_5773 (I100241,I100202,I100111);
nand I_5774 (I99819,I100094,I100241);
not I_5775 (I100272,I100202);
nor I_5776 (I100289,I100272,I100012);
DFFARX1 I_5777 (I100289,I2067,I99842,I99831,);
nor I_5778 (I100320,I158979,I158970);
or I_5779 (I99822,I100069,I100320);
nor I_5780 (I99813,I100202,I100320);
or I_5781 (I99816,I99936,I100320);
DFFARX1 I_5782 (I100320,I2067,I99842,I99834,);
not I_5783 (I100420,I2074);
DFFARX1 I_5784 (I111300,I2067,I100420,I100446,);
not I_5785 (I100454,I100446);
nand I_5786 (I100471,I111288,I111306);
and I_5787 (I100488,I100471,I111303);
DFFARX1 I_5788 (I100488,I2067,I100420,I100514,);
not I_5789 (I100522,I111294);
DFFARX1 I_5790 (I111291,I2067,I100420,I100548,);
not I_5791 (I100556,I100548);
nor I_5792 (I100573,I100556,I100454);
and I_5793 (I100590,I100573,I111294);
nor I_5794 (I100607,I100556,I100522);
nor I_5795 (I100403,I100514,I100607);
DFFARX1 I_5796 (I111285,I2067,I100420,I100647,);
nor I_5797 (I100655,I100647,I100514);
not I_5798 (I100672,I100655);
not I_5799 (I100689,I100647);
nor I_5800 (I100706,I100689,I100590);
DFFARX1 I_5801 (I100706,I2067,I100420,I100406,);
nand I_5802 (I100737,I111285,I111288);
and I_5803 (I100754,I100737,I111291);
DFFARX1 I_5804 (I100754,I2067,I100420,I100780,);
nor I_5805 (I100788,I100780,I100647);
DFFARX1 I_5806 (I100788,I2067,I100420,I100388,);
nand I_5807 (I100819,I100780,I100689);
nand I_5808 (I100397,I100672,I100819);
not I_5809 (I100850,I100780);
nor I_5810 (I100867,I100850,I100590);
DFFARX1 I_5811 (I100867,I2067,I100420,I100409,);
nor I_5812 (I100898,I111297,I111288);
or I_5813 (I100400,I100647,I100898);
nor I_5814 (I100391,I100780,I100898);
or I_5815 (I100394,I100514,I100898);
DFFARX1 I_5816 (I100898,I2067,I100420,I100412,);
not I_5817 (I100998,I2074);
DFFARX1 I_5818 (I167531,I2067,I100998,I101024,);
not I_5819 (I101032,I101024);
nand I_5820 (I101049,I167516,I167504);
and I_5821 (I101066,I101049,I167519);
DFFARX1 I_5822 (I101066,I2067,I100998,I101092,);
not I_5823 (I101100,I167504);
DFFARX1 I_5824 (I167522,I2067,I100998,I101126,);
not I_5825 (I101134,I101126);
nor I_5826 (I101151,I101134,I101032);
and I_5827 (I101168,I101151,I167504);
nor I_5828 (I101185,I101134,I101100);
nor I_5829 (I100981,I101092,I101185);
DFFARX1 I_5830 (I167510,I2067,I100998,I101225,);
nor I_5831 (I101233,I101225,I101092);
not I_5832 (I101250,I101233);
not I_5833 (I101267,I101225);
nor I_5834 (I101284,I101267,I101168);
DFFARX1 I_5835 (I101284,I2067,I100998,I100984,);
nand I_5836 (I101315,I167507,I167513);
and I_5837 (I101332,I101315,I167528);
DFFARX1 I_5838 (I101332,I2067,I100998,I101358,);
nor I_5839 (I101366,I101358,I101225);
DFFARX1 I_5840 (I101366,I2067,I100998,I100966,);
nand I_5841 (I101397,I101358,I101267);
nand I_5842 (I100975,I101250,I101397);
not I_5843 (I101428,I101358);
nor I_5844 (I101445,I101428,I101168);
DFFARX1 I_5845 (I101445,I2067,I100998,I100987,);
nor I_5846 (I101476,I167525,I167513);
or I_5847 (I100978,I101225,I101476);
nor I_5848 (I100969,I101358,I101476);
or I_5849 (I100972,I101092,I101476);
DFFARX1 I_5850 (I101476,I2067,I100998,I100990,);
not I_5851 (I101576,I2074);
DFFARX1 I_5852 (I150114,I2067,I101576,I101602,);
not I_5853 (I101610,I101602);
nand I_5854 (I101627,I150096,I150108);
and I_5855 (I101644,I101627,I150111);
DFFARX1 I_5856 (I101644,I2067,I101576,I101670,);
not I_5857 (I101678,I150105);
DFFARX1 I_5858 (I150102,I2067,I101576,I101704,);
not I_5859 (I101712,I101704);
nor I_5860 (I101729,I101712,I101610);
and I_5861 (I101746,I101729,I150105);
nor I_5862 (I101763,I101712,I101678);
nor I_5863 (I101559,I101670,I101763);
DFFARX1 I_5864 (I150120,I2067,I101576,I101803,);
nor I_5865 (I101811,I101803,I101670);
not I_5866 (I101828,I101811);
not I_5867 (I101845,I101803);
nor I_5868 (I101862,I101845,I101746);
DFFARX1 I_5869 (I101862,I2067,I101576,I101562,);
nand I_5870 (I101893,I150099,I150099);
and I_5871 (I101910,I101893,I150096);
DFFARX1 I_5872 (I101910,I2067,I101576,I101936,);
nor I_5873 (I101944,I101936,I101803);
DFFARX1 I_5874 (I101944,I2067,I101576,I101544,);
nand I_5875 (I101975,I101936,I101845);
nand I_5876 (I101553,I101828,I101975);
not I_5877 (I102006,I101936);
nor I_5878 (I102023,I102006,I101746);
DFFARX1 I_5879 (I102023,I2067,I101576,I101565,);
nor I_5880 (I102054,I150117,I150099);
or I_5881 (I101556,I101803,I102054);
nor I_5882 (I101547,I101936,I102054);
or I_5883 (I101550,I101670,I102054);
DFFARX1 I_5884 (I102054,I2067,I101576,I101568,);
not I_5885 (I102154,I2074);
DFFARX1 I_5886 (I150692,I2067,I102154,I102180,);
not I_5887 (I102188,I102180);
nand I_5888 (I102205,I150674,I150686);
and I_5889 (I102222,I102205,I150689);
DFFARX1 I_5890 (I102222,I2067,I102154,I102248,);
not I_5891 (I102256,I150683);
DFFARX1 I_5892 (I150680,I2067,I102154,I102282,);
not I_5893 (I102290,I102282);
nor I_5894 (I102307,I102290,I102188);
and I_5895 (I102324,I102307,I150683);
nor I_5896 (I102341,I102290,I102256);
nor I_5897 (I102137,I102248,I102341);
DFFARX1 I_5898 (I150698,I2067,I102154,I102381,);
nor I_5899 (I102389,I102381,I102248);
not I_5900 (I102406,I102389);
not I_5901 (I102423,I102381);
nor I_5902 (I102440,I102423,I102324);
DFFARX1 I_5903 (I102440,I2067,I102154,I102140,);
nand I_5904 (I102471,I150677,I150677);
and I_5905 (I102488,I102471,I150674);
DFFARX1 I_5906 (I102488,I2067,I102154,I102514,);
nor I_5907 (I102522,I102514,I102381);
DFFARX1 I_5908 (I102522,I2067,I102154,I102122,);
nand I_5909 (I102553,I102514,I102423);
nand I_5910 (I102131,I102406,I102553);
not I_5911 (I102584,I102514);
nor I_5912 (I102601,I102584,I102324);
DFFARX1 I_5913 (I102601,I2067,I102154,I102143,);
nor I_5914 (I102632,I150695,I150677);
or I_5915 (I102134,I102381,I102632);
nor I_5916 (I102125,I102514,I102632);
or I_5917 (I102128,I102248,I102632);
DFFARX1 I_5918 (I102632,I2067,I102154,I102146,);
not I_5919 (I102732,I2074);
DFFARX1 I_5920 (I54937,I2067,I102732,I102758,);
not I_5921 (I102766,I102758);
nand I_5922 (I102783,I54940,I54916);
and I_5923 (I102800,I102783,I54913);
DFFARX1 I_5924 (I102800,I2067,I102732,I102826,);
not I_5925 (I102834,I54919);
DFFARX1 I_5926 (I54913,I2067,I102732,I102860,);
not I_5927 (I102868,I102860);
nor I_5928 (I102885,I102868,I102766);
and I_5929 (I102902,I102885,I54919);
nor I_5930 (I102919,I102868,I102834);
nor I_5931 (I102715,I102826,I102919);
DFFARX1 I_5932 (I54922,I2067,I102732,I102959,);
nor I_5933 (I102967,I102959,I102826);
not I_5934 (I102984,I102967);
not I_5935 (I103001,I102959);
nor I_5936 (I103018,I103001,I102902);
DFFARX1 I_5937 (I103018,I2067,I102732,I102718,);
nand I_5938 (I103049,I54925,I54934);
and I_5939 (I103066,I103049,I54931);
DFFARX1 I_5940 (I103066,I2067,I102732,I103092,);
nor I_5941 (I103100,I103092,I102959);
DFFARX1 I_5942 (I103100,I2067,I102732,I102700,);
nand I_5943 (I103131,I103092,I103001);
nand I_5944 (I102709,I102984,I103131);
not I_5945 (I103162,I103092);
nor I_5946 (I103179,I103162,I102902);
DFFARX1 I_5947 (I103179,I2067,I102732,I102721,);
nor I_5948 (I103210,I54928,I54934);
or I_5949 (I102712,I102959,I103210);
nor I_5950 (I102703,I103092,I103210);
or I_5951 (I102706,I102826,I103210);
DFFARX1 I_5952 (I103210,I2067,I102732,I102724,);
not I_5953 (I103310,I2074);
DFFARX1 I_5954 (I28648,I2067,I103310,I103336,);
not I_5955 (I103344,I103336);
nand I_5956 (I103361,I28651,I28672);
and I_5957 (I103378,I103361,I28660);
DFFARX1 I_5958 (I103378,I2067,I103310,I103404,);
not I_5959 (I103412,I28657);
DFFARX1 I_5960 (I28648,I2067,I103310,I103438,);
not I_5961 (I103446,I103438);
nor I_5962 (I103463,I103446,I103344);
and I_5963 (I103480,I103463,I28657);
nor I_5964 (I103497,I103446,I103412);
nor I_5965 (I103293,I103404,I103497);
DFFARX1 I_5966 (I28666,I2067,I103310,I103537,);
nor I_5967 (I103545,I103537,I103404);
not I_5968 (I103562,I103545);
not I_5969 (I103579,I103537);
nor I_5970 (I103596,I103579,I103480);
DFFARX1 I_5971 (I103596,I2067,I103310,I103296,);
nand I_5972 (I103627,I28651,I28654);
and I_5973 (I103644,I103627,I28663);
DFFARX1 I_5974 (I103644,I2067,I103310,I103670,);
nor I_5975 (I103678,I103670,I103537);
DFFARX1 I_5976 (I103678,I2067,I103310,I103278,);
nand I_5977 (I103709,I103670,I103579);
nand I_5978 (I103287,I103562,I103709);
not I_5979 (I103740,I103670);
nor I_5980 (I103757,I103740,I103480);
DFFARX1 I_5981 (I103757,I2067,I103310,I103299,);
nor I_5982 (I103788,I28669,I28654);
or I_5983 (I103290,I103537,I103788);
nor I_5984 (I103281,I103670,I103788);
or I_5985 (I103284,I103404,I103788);
DFFARX1 I_5986 (I103788,I2067,I103310,I103302,);
not I_5987 (I103888,I2074);
DFFARX1 I_5988 (I172291,I2067,I103888,I103914,);
not I_5989 (I103922,I103914);
nand I_5990 (I103939,I172276,I172264);
and I_5991 (I103956,I103939,I172279);
DFFARX1 I_5992 (I103956,I2067,I103888,I103982,);
not I_5993 (I103990,I172264);
DFFARX1 I_5994 (I172282,I2067,I103888,I104016,);
not I_5995 (I104024,I104016);
nor I_5996 (I104041,I104024,I103922);
and I_5997 (I104058,I104041,I172264);
nor I_5998 (I104075,I104024,I103990);
nor I_5999 (I103871,I103982,I104075);
DFFARX1 I_6000 (I172270,I2067,I103888,I104115,);
nor I_6001 (I104123,I104115,I103982);
not I_6002 (I104140,I104123);
not I_6003 (I104157,I104115);
nor I_6004 (I104174,I104157,I104058);
DFFARX1 I_6005 (I104174,I2067,I103888,I103874,);
nand I_6006 (I104205,I172267,I172273);
and I_6007 (I104222,I104205,I172288);
DFFARX1 I_6008 (I104222,I2067,I103888,I104248,);
nor I_6009 (I104256,I104248,I104115);
DFFARX1 I_6010 (I104256,I2067,I103888,I103856,);
nand I_6011 (I104287,I104248,I104157);
nand I_6012 (I103865,I104140,I104287);
not I_6013 (I104318,I104248);
nor I_6014 (I104335,I104318,I104058);
DFFARX1 I_6015 (I104335,I2067,I103888,I103877,);
nor I_6016 (I104366,I172285,I172273);
or I_6017 (I103868,I104115,I104366);
nor I_6018 (I103859,I104248,I104366);
or I_6019 (I103862,I103982,I104366);
DFFARX1 I_6020 (I104366,I2067,I103888,I103880,);
not I_6021 (I104463,I2074);
DFFARX1 I_6022 (I3803,I2067,I104463,I104489,);
not I_6023 (I104497,I104489);
nand I_6024 (I104514,I3815,I3818);
and I_6025 (I104531,I104514,I3794);
DFFARX1 I_6026 (I104531,I2067,I104463,I104557,);
DFFARX1 I_6027 (I104557,I2067,I104463,I104452,);
DFFARX1 I_6028 (I3812,I2067,I104463,I104588,);
nand I_6029 (I104596,I104588,I3800);
not I_6030 (I104613,I104596);
DFFARX1 I_6031 (I104613,I2067,I104463,I104639,);
not I_6032 (I104647,I104639);
nor I_6033 (I104455,I104497,I104647);
DFFARX1 I_6034 (I3797,I2067,I104463,I104687,);
nor I_6035 (I104446,I104687,I104557);
nor I_6036 (I104437,I104687,I104613);
nand I_6037 (I104723,I3806,I3797);
and I_6038 (I104740,I104723,I3794);
DFFARX1 I_6039 (I104740,I2067,I104463,I104766,);
not I_6040 (I104774,I104766);
nand I_6041 (I104791,I104774,I104687);
nand I_6042 (I104440,I104774,I104596);
nor I_6043 (I104822,I3809,I3797);
and I_6044 (I104839,I104687,I104822);
nor I_6045 (I104856,I104774,I104839);
DFFARX1 I_6046 (I104856,I2067,I104463,I104449,);
nor I_6047 (I104887,I104489,I104822);
DFFARX1 I_6048 (I104887,I2067,I104463,I104434,);
nor I_6049 (I104918,I104766,I104822);
not I_6050 (I104935,I104918);
nand I_6051 (I104443,I104935,I104791);
not I_6052 (I104990,I2074);
DFFARX1 I_6053 (I171089,I2067,I104990,I105016,);
not I_6054 (I105024,I105016);
nand I_6055 (I105041,I171086,I171095);
and I_6056 (I105058,I105041,I171074);
DFFARX1 I_6057 (I105058,I2067,I104990,I105084,);
DFFARX1 I_6058 (I105084,I2067,I104990,I104979,);
DFFARX1 I_6059 (I171077,I2067,I104990,I105115,);
nand I_6060 (I105123,I105115,I171092);
not I_6061 (I105140,I105123);
DFFARX1 I_6062 (I105140,I2067,I104990,I105166,);
not I_6063 (I105174,I105166);
nor I_6064 (I104982,I105024,I105174);
DFFARX1 I_6065 (I171098,I2067,I104990,I105214,);
nor I_6066 (I104973,I105214,I105084);
nor I_6067 (I104964,I105214,I105140);
nand I_6068 (I105250,I171080,I171101);
and I_6069 (I105267,I105250,I171083);
DFFARX1 I_6070 (I105267,I2067,I104990,I105293,);
not I_6071 (I105301,I105293);
nand I_6072 (I105318,I105301,I105214);
nand I_6073 (I104967,I105301,I105123);
nor I_6074 (I105349,I171074,I171101);
and I_6075 (I105366,I105214,I105349);
nor I_6076 (I105383,I105301,I105366);
DFFARX1 I_6077 (I105383,I2067,I104990,I104976,);
nor I_6078 (I105414,I105016,I105349);
DFFARX1 I_6079 (I105414,I2067,I104990,I104961,);
nor I_6080 (I105445,I105293,I105349);
not I_6081 (I105462,I105445);
nand I_6082 (I104970,I105462,I105318);
not I_6083 (I105517,I2074);
DFFARX1 I_6084 (I18574,I2067,I105517,I105543,);
not I_6085 (I105551,I105543);
nand I_6086 (I105568,I18550,I18559);
and I_6087 (I105585,I105568,I18553);
DFFARX1 I_6088 (I105585,I2067,I105517,I105611,);
DFFARX1 I_6089 (I105611,I2067,I105517,I105506,);
DFFARX1 I_6090 (I18571,I2067,I105517,I105642,);
nand I_6091 (I105650,I105642,I18562);
not I_6092 (I105667,I105650);
DFFARX1 I_6093 (I105667,I2067,I105517,I105693,);
not I_6094 (I105701,I105693);
nor I_6095 (I105509,I105551,I105701);
DFFARX1 I_6096 (I18556,I2067,I105517,I105741,);
nor I_6097 (I105500,I105741,I105611);
nor I_6098 (I105491,I105741,I105667);
nand I_6099 (I105777,I18568,I18565);
and I_6100 (I105794,I105777,I18553);
DFFARX1 I_6101 (I105794,I2067,I105517,I105820,);
not I_6102 (I105828,I105820);
nand I_6103 (I105845,I105828,I105741);
nand I_6104 (I105494,I105828,I105650);
nor I_6105 (I105876,I18550,I18565);
and I_6106 (I105893,I105741,I105876);
nor I_6107 (I105910,I105828,I105893);
DFFARX1 I_6108 (I105910,I2067,I105517,I105503,);
nor I_6109 (I105941,I105543,I105876);
DFFARX1 I_6110 (I105941,I2067,I105517,I105488,);
nor I_6111 (I105972,I105820,I105876);
not I_6112 (I105989,I105972);
nand I_6113 (I105497,I105989,I105845);
not I_6114 (I106044,I2074);
DFFARX1 I_6115 (I169304,I2067,I106044,I106070,);
not I_6116 (I106078,I106070);
nand I_6117 (I106095,I169301,I169310);
and I_6118 (I106112,I106095,I169289);
DFFARX1 I_6119 (I106112,I2067,I106044,I106138,);
DFFARX1 I_6120 (I106138,I2067,I106044,I106033,);
DFFARX1 I_6121 (I169292,I2067,I106044,I106169,);
nand I_6122 (I106177,I106169,I169307);
not I_6123 (I106194,I106177);
DFFARX1 I_6124 (I106194,I2067,I106044,I106220,);
not I_6125 (I106228,I106220);
nor I_6126 (I106036,I106078,I106228);
DFFARX1 I_6127 (I169313,I2067,I106044,I106268,);
nor I_6128 (I106027,I106268,I106138);
nor I_6129 (I106018,I106268,I106194);
nand I_6130 (I106304,I169295,I169316);
and I_6131 (I106321,I106304,I169298);
DFFARX1 I_6132 (I106321,I2067,I106044,I106347,);
not I_6133 (I106355,I106347);
nand I_6134 (I106372,I106355,I106268);
nand I_6135 (I106021,I106355,I106177);
nor I_6136 (I106403,I169289,I169316);
and I_6137 (I106420,I106268,I106403);
nor I_6138 (I106437,I106355,I106420);
DFFARX1 I_6139 (I106437,I2067,I106044,I106030,);
nor I_6140 (I106468,I106070,I106403);
DFFARX1 I_6141 (I106468,I2067,I106044,I106015,);
nor I_6142 (I106499,I106347,I106403);
not I_6143 (I106516,I106499);
nand I_6144 (I106024,I106516,I106372);
not I_6145 (I106571,I2074);
DFFARX1 I_6146 (I168709,I2067,I106571,I106597,);
not I_6147 (I106605,I106597);
nand I_6148 (I106622,I168706,I168715);
and I_6149 (I106639,I106622,I168694);
DFFARX1 I_6150 (I106639,I2067,I106571,I106665,);
DFFARX1 I_6151 (I106665,I2067,I106571,I106560,);
DFFARX1 I_6152 (I168697,I2067,I106571,I106696,);
nand I_6153 (I106704,I106696,I168712);
not I_6154 (I106721,I106704);
DFFARX1 I_6155 (I106721,I2067,I106571,I106747,);
not I_6156 (I106755,I106747);
nor I_6157 (I106563,I106605,I106755);
DFFARX1 I_6158 (I168718,I2067,I106571,I106795,);
nor I_6159 (I106554,I106795,I106665);
nor I_6160 (I106545,I106795,I106721);
nand I_6161 (I106831,I168700,I168721);
and I_6162 (I106848,I106831,I168703);
DFFARX1 I_6163 (I106848,I2067,I106571,I106874,);
not I_6164 (I106882,I106874);
nand I_6165 (I106899,I106882,I106795);
nand I_6166 (I106548,I106882,I106704);
nor I_6167 (I106930,I168694,I168721);
and I_6168 (I106947,I106795,I106930);
nor I_6169 (I106964,I106882,I106947);
DFFARX1 I_6170 (I106964,I2067,I106571,I106557,);
nor I_6171 (I106995,I106597,I106930);
DFFARX1 I_6172 (I106995,I2067,I106571,I106542,);
nor I_6173 (I107026,I106874,I106930);
not I_6174 (I107043,I107026);
nand I_6175 (I106551,I107043,I106899);
not I_6176 (I107098,I2074);
DFFARX1 I_6177 (I143756,I2067,I107098,I107124,);
not I_6178 (I107132,I107124);
nand I_6179 (I107149,I143738,I143738);
and I_6180 (I107166,I107149,I143744);
DFFARX1 I_6181 (I107166,I2067,I107098,I107192,);
DFFARX1 I_6182 (I107192,I2067,I107098,I107087,);
DFFARX1 I_6183 (I143741,I2067,I107098,I107223,);
nand I_6184 (I107231,I107223,I143750);
not I_6185 (I107248,I107231);
DFFARX1 I_6186 (I107248,I2067,I107098,I107274,);
not I_6187 (I107282,I107274);
nor I_6188 (I107090,I107132,I107282);
DFFARX1 I_6189 (I143762,I2067,I107098,I107322,);
nor I_6190 (I107081,I107322,I107192);
nor I_6191 (I107072,I107322,I107248);
nand I_6192 (I107358,I143753,I143747);
and I_6193 (I107375,I107358,I143741);
DFFARX1 I_6194 (I107375,I2067,I107098,I107401,);
not I_6195 (I107409,I107401);
nand I_6196 (I107426,I107409,I107322);
nand I_6197 (I107075,I107409,I107231);
nor I_6198 (I107457,I143759,I143747);
and I_6199 (I107474,I107322,I107457);
nor I_6200 (I107491,I107409,I107474);
DFFARX1 I_6201 (I107491,I2067,I107098,I107084,);
nor I_6202 (I107522,I107124,I107457);
DFFARX1 I_6203 (I107522,I2067,I107098,I107069,);
nor I_6204 (I107553,I107401,I107457);
not I_6205 (I107570,I107553);
nand I_6206 (I107078,I107570,I107426);
not I_6207 (I107625,I2074);
DFFARX1 I_6208 (I59135,I2067,I107625,I107651,);
not I_6209 (I107659,I107651);
nand I_6210 (I107676,I59132,I59141);
and I_6211 (I107693,I107676,I59150);
DFFARX1 I_6212 (I107693,I2067,I107625,I107719,);
DFFARX1 I_6213 (I107719,I2067,I107625,I107614,);
DFFARX1 I_6214 (I59153,I2067,I107625,I107750,);
nand I_6215 (I107758,I107750,I59156);
not I_6216 (I107775,I107758);
DFFARX1 I_6217 (I107775,I2067,I107625,I107801,);
not I_6218 (I107809,I107801);
nor I_6219 (I107617,I107659,I107809);
DFFARX1 I_6220 (I59129,I2067,I107625,I107849,);
nor I_6221 (I107608,I107849,I107719);
nor I_6222 (I107599,I107849,I107775);
nand I_6223 (I107885,I59144,I59147);
and I_6224 (I107902,I107885,I59138);
DFFARX1 I_6225 (I107902,I2067,I107625,I107928,);
not I_6226 (I107936,I107928);
nand I_6227 (I107953,I107936,I107849);
nand I_6228 (I107602,I107936,I107758);
nor I_6229 (I107984,I59129,I59147);
and I_6230 (I108001,I107849,I107984);
nor I_6231 (I108018,I107936,I108001);
DFFARX1 I_6232 (I108018,I2067,I107625,I107611,);
nor I_6233 (I108049,I107651,I107984);
DFFARX1 I_6234 (I108049,I2067,I107625,I107596,);
nor I_6235 (I108080,I107928,I107984);
not I_6236 (I108097,I108080);
nand I_6237 (I107605,I108097,I107953);
not I_6238 (I108152,I2074);
DFFARX1 I_6239 (I102122,I2067,I108152,I108178,);
not I_6240 (I108186,I108178);
nand I_6241 (I108203,I102125,I102122);
and I_6242 (I108220,I108203,I102134);
DFFARX1 I_6243 (I108220,I2067,I108152,I108246,);
DFFARX1 I_6244 (I108246,I2067,I108152,I108141,);
DFFARX1 I_6245 (I102131,I2067,I108152,I108277,);
nand I_6246 (I108285,I108277,I102137);
not I_6247 (I108302,I108285);
DFFARX1 I_6248 (I108302,I2067,I108152,I108328,);
not I_6249 (I108336,I108328);
nor I_6250 (I108144,I108186,I108336);
DFFARX1 I_6251 (I102146,I2067,I108152,I108376,);
nor I_6252 (I108135,I108376,I108246);
nor I_6253 (I108126,I108376,I108302);
nand I_6254 (I108412,I102140,I102128);
and I_6255 (I108429,I108412,I102125);
DFFARX1 I_6256 (I108429,I2067,I108152,I108455,);
not I_6257 (I108463,I108455);
nand I_6258 (I108480,I108463,I108376);
nand I_6259 (I108129,I108463,I108285);
nor I_6260 (I108511,I102143,I102128);
and I_6261 (I108528,I108376,I108511);
nor I_6262 (I108545,I108463,I108528);
DFFARX1 I_6263 (I108545,I2067,I108152,I108138,);
nor I_6264 (I108576,I108178,I108511);
DFFARX1 I_6265 (I108576,I2067,I108152,I108123,);
nor I_6266 (I108607,I108455,I108511);
not I_6267 (I108624,I108607);
nand I_6268 (I108132,I108624,I108480);
not I_6269 (I108679,I2074);
DFFARX1 I_6270 (I21736,I2067,I108679,I108705,);
not I_6271 (I108713,I108705);
nand I_6272 (I108730,I21712,I21721);
and I_6273 (I108747,I108730,I21715);
DFFARX1 I_6274 (I108747,I2067,I108679,I108773,);
DFFARX1 I_6275 (I108773,I2067,I108679,I108668,);
DFFARX1 I_6276 (I21733,I2067,I108679,I108804,);
nand I_6277 (I108812,I108804,I21724);
not I_6278 (I108829,I108812);
DFFARX1 I_6279 (I108829,I2067,I108679,I108855,);
not I_6280 (I108863,I108855);
nor I_6281 (I108671,I108713,I108863);
DFFARX1 I_6282 (I21718,I2067,I108679,I108903,);
nor I_6283 (I108662,I108903,I108773);
nor I_6284 (I108653,I108903,I108829);
nand I_6285 (I108939,I21730,I21727);
and I_6286 (I108956,I108939,I21715);
DFFARX1 I_6287 (I108956,I2067,I108679,I108982,);
not I_6288 (I108990,I108982);
nand I_6289 (I109007,I108990,I108903);
nand I_6290 (I108656,I108990,I108812);
nor I_6291 (I109038,I21712,I21727);
and I_6292 (I109055,I108903,I109038);
nor I_6293 (I109072,I108990,I109055);
DFFARX1 I_6294 (I109072,I2067,I108679,I108665,);
nor I_6295 (I109103,I108705,I109038);
DFFARX1 I_6296 (I109103,I2067,I108679,I108650,);
nor I_6297 (I109134,I108982,I109038);
not I_6298 (I109151,I109134);
nand I_6299 (I108659,I109151,I109007);
not I_6300 (I109206,I2074);
DFFARX1 I_6301 (I11723,I2067,I109206,I109232,);
not I_6302 (I109240,I109232);
nand I_6303 (I109257,I11699,I11708);
and I_6304 (I109274,I109257,I11702);
DFFARX1 I_6305 (I109274,I2067,I109206,I109300,);
DFFARX1 I_6306 (I109300,I2067,I109206,I109195,);
DFFARX1 I_6307 (I11720,I2067,I109206,I109331,);
nand I_6308 (I109339,I109331,I11711);
not I_6309 (I109356,I109339);
DFFARX1 I_6310 (I109356,I2067,I109206,I109382,);
not I_6311 (I109390,I109382);
nor I_6312 (I109198,I109240,I109390);
DFFARX1 I_6313 (I11705,I2067,I109206,I109430,);
nor I_6314 (I109189,I109430,I109300);
nor I_6315 (I109180,I109430,I109356);
nand I_6316 (I109466,I11717,I11714);
and I_6317 (I109483,I109466,I11702);
DFFARX1 I_6318 (I109483,I2067,I109206,I109509,);
not I_6319 (I109517,I109509);
nand I_6320 (I109534,I109517,I109430);
nand I_6321 (I109183,I109517,I109339);
nor I_6322 (I109565,I11699,I11714);
and I_6323 (I109582,I109430,I109565);
nor I_6324 (I109599,I109517,I109582);
DFFARX1 I_6325 (I109599,I2067,I109206,I109192,);
nor I_6326 (I109630,I109232,I109565);
DFFARX1 I_6327 (I109630,I2067,I109206,I109177,);
nor I_6328 (I109661,I109509,I109565);
not I_6329 (I109678,I109661);
nand I_6330 (I109186,I109678,I109534);
not I_6331 (I109733,I2074);
DFFARX1 I_6332 (I76662,I2067,I109733,I109759,);
not I_6333 (I109767,I109759);
nand I_6334 (I109784,I76680,I76671);
and I_6335 (I109801,I109784,I76674);
DFFARX1 I_6336 (I109801,I2067,I109733,I109827,);
DFFARX1 I_6337 (I109827,I2067,I109733,I109722,);
DFFARX1 I_6338 (I76668,I2067,I109733,I109858,);
nand I_6339 (I109866,I109858,I76659);
not I_6340 (I109883,I109866);
DFFARX1 I_6341 (I109883,I2067,I109733,I109909,);
not I_6342 (I109917,I109909);
nor I_6343 (I109725,I109767,I109917);
DFFARX1 I_6344 (I76665,I2067,I109733,I109957,);
nor I_6345 (I109716,I109957,I109827);
nor I_6346 (I109707,I109957,I109883);
nand I_6347 (I109993,I76659,I76656);
and I_6348 (I110010,I109993,I76677);
DFFARX1 I_6349 (I110010,I2067,I109733,I110036,);
not I_6350 (I110044,I110036);
nand I_6351 (I110061,I110044,I109957);
nand I_6352 (I109710,I110044,I109866);
nor I_6353 (I110092,I76656,I76656);
and I_6354 (I110109,I109957,I110092);
nor I_6355 (I110126,I110044,I110109);
DFFARX1 I_6356 (I110126,I2067,I109733,I109719,);
nor I_6357 (I110157,I109759,I110092);
DFFARX1 I_6358 (I110157,I2067,I109733,I109704,);
nor I_6359 (I110188,I110036,I110092);
not I_6360 (I110205,I110188);
nand I_6361 (I109713,I110205,I110061);
not I_6362 (I110260,I2074);
DFFARX1 I_6363 (I172874,I2067,I110260,I110286,);
not I_6364 (I110294,I110286);
nand I_6365 (I110311,I172871,I172880);
and I_6366 (I110328,I110311,I172859);
DFFARX1 I_6367 (I110328,I2067,I110260,I110354,);
DFFARX1 I_6368 (I110354,I2067,I110260,I110249,);
DFFARX1 I_6369 (I172862,I2067,I110260,I110385,);
nand I_6370 (I110393,I110385,I172877);
not I_6371 (I110410,I110393);
DFFARX1 I_6372 (I110410,I2067,I110260,I110436,);
not I_6373 (I110444,I110436);
nor I_6374 (I110252,I110294,I110444);
DFFARX1 I_6375 (I172883,I2067,I110260,I110484,);
nor I_6376 (I110243,I110484,I110354);
nor I_6377 (I110234,I110484,I110410);
nand I_6378 (I110520,I172865,I172886);
and I_6379 (I110537,I110520,I172868);
DFFARX1 I_6380 (I110537,I2067,I110260,I110563,);
not I_6381 (I110571,I110563);
nand I_6382 (I110588,I110571,I110484);
nand I_6383 (I110237,I110571,I110393);
nor I_6384 (I110619,I172859,I172886);
and I_6385 (I110636,I110484,I110619);
nor I_6386 (I110653,I110571,I110636);
DFFARX1 I_6387 (I110653,I2067,I110260,I110246,);
nor I_6388 (I110684,I110286,I110619);
DFFARX1 I_6389 (I110684,I2067,I110260,I110231,);
nor I_6390 (I110715,I110563,I110619);
not I_6391 (I110732,I110715);
nand I_6392 (I110240,I110732,I110588);
not I_6393 (I110787,I2074);
DFFARX1 I_6394 (I169899,I2067,I110787,I110813,);
not I_6395 (I110821,I110813);
nand I_6396 (I110838,I169896,I169905);
and I_6397 (I110855,I110838,I169884);
DFFARX1 I_6398 (I110855,I2067,I110787,I110881,);
DFFARX1 I_6399 (I110881,I2067,I110787,I110776,);
DFFARX1 I_6400 (I169887,I2067,I110787,I110912,);
nand I_6401 (I110920,I110912,I169902);
not I_6402 (I110937,I110920);
DFFARX1 I_6403 (I110937,I2067,I110787,I110963,);
not I_6404 (I110971,I110963);
nor I_6405 (I110779,I110821,I110971);
DFFARX1 I_6406 (I169908,I2067,I110787,I111011,);
nor I_6407 (I110770,I111011,I110881);
nor I_6408 (I110761,I111011,I110937);
nand I_6409 (I111047,I169890,I169911);
and I_6410 (I111064,I111047,I169893);
DFFARX1 I_6411 (I111064,I2067,I110787,I111090,);
not I_6412 (I111098,I111090);
nand I_6413 (I111115,I111098,I111011);
nand I_6414 (I110764,I111098,I110920);
nor I_6415 (I111146,I169884,I169911);
and I_6416 (I111163,I111011,I111146);
nor I_6417 (I111180,I111098,I111163);
DFFARX1 I_6418 (I111180,I2067,I110787,I110773,);
nor I_6419 (I111211,I110813,I111146);
DFFARX1 I_6420 (I111211,I2067,I110787,I110758,);
nor I_6421 (I111242,I111090,I111146);
not I_6422 (I111259,I111242);
nand I_6423 (I110767,I111259,I111115);
not I_6424 (I111314,I2074);
DFFARX1 I_6425 (I9615,I2067,I111314,I111340,);
not I_6426 (I111348,I111340);
nand I_6427 (I111365,I9591,I9600);
and I_6428 (I111382,I111365,I9594);
DFFARX1 I_6429 (I111382,I2067,I111314,I111408,);
DFFARX1 I_6430 (I111408,I2067,I111314,I111303,);
DFFARX1 I_6431 (I9612,I2067,I111314,I111439,);
nand I_6432 (I111447,I111439,I9603);
not I_6433 (I111464,I111447);
DFFARX1 I_6434 (I111464,I2067,I111314,I111490,);
not I_6435 (I111498,I111490);
nor I_6436 (I111306,I111348,I111498);
DFFARX1 I_6437 (I9597,I2067,I111314,I111538,);
nor I_6438 (I111297,I111538,I111408);
nor I_6439 (I111288,I111538,I111464);
nand I_6440 (I111574,I9609,I9606);
and I_6441 (I111591,I111574,I9594);
DFFARX1 I_6442 (I111591,I2067,I111314,I111617,);
not I_6443 (I111625,I111617);
nand I_6444 (I111642,I111625,I111538);
nand I_6445 (I111291,I111625,I111447);
nor I_6446 (I111673,I9591,I9606);
and I_6447 (I111690,I111538,I111673);
nor I_6448 (I111707,I111625,I111690);
DFFARX1 I_6449 (I111707,I2067,I111314,I111300,);
nor I_6450 (I111738,I111340,I111673);
DFFARX1 I_6451 (I111738,I2067,I111314,I111285,);
nor I_6452 (I111769,I111617,I111673);
not I_6453 (I111786,I111769);
nand I_6454 (I111294,I111786,I111642);
not I_6455 (I111841,I2074);
DFFARX1 I_6456 (I73092,I2067,I111841,I111867,);
not I_6457 (I111875,I111867);
nand I_6458 (I111892,I73110,I73101);
and I_6459 (I111909,I111892,I73104);
DFFARX1 I_6460 (I111909,I2067,I111841,I111935,);
DFFARX1 I_6461 (I111935,I2067,I111841,I111830,);
DFFARX1 I_6462 (I73098,I2067,I111841,I111966,);
nand I_6463 (I111974,I111966,I73089);
not I_6464 (I111991,I111974);
DFFARX1 I_6465 (I111991,I2067,I111841,I112017,);
not I_6466 (I112025,I112017);
nor I_6467 (I111833,I111875,I112025);
DFFARX1 I_6468 (I73095,I2067,I111841,I112065,);
nor I_6469 (I111824,I112065,I111935);
nor I_6470 (I111815,I112065,I111991);
nand I_6471 (I112101,I73089,I73086);
and I_6472 (I112118,I112101,I73107);
DFFARX1 I_6473 (I112118,I2067,I111841,I112144,);
not I_6474 (I112152,I112144);
nand I_6475 (I112169,I112152,I112065);
nand I_6476 (I111818,I112152,I111974);
nor I_6477 (I112200,I73086,I73086);
and I_6478 (I112217,I112065,I112200);
nor I_6479 (I112234,I112152,I112217);
DFFARX1 I_6480 (I112234,I2067,I111841,I111827,);
nor I_6481 (I112265,I111867,I112200);
DFFARX1 I_6482 (I112265,I2067,I111841,I111812,);
nor I_6483 (I112296,I112144,I112200);
not I_6484 (I112313,I112296);
nand I_6485 (I111821,I112313,I112169);
not I_6486 (I112368,I2074);
DFFARX1 I_6487 (I137398,I2067,I112368,I112394,);
not I_6488 (I112402,I112394);
nand I_6489 (I112419,I137380,I137380);
and I_6490 (I112436,I112419,I137386);
DFFARX1 I_6491 (I112436,I2067,I112368,I112462,);
DFFARX1 I_6492 (I112462,I2067,I112368,I112357,);
DFFARX1 I_6493 (I137383,I2067,I112368,I112493,);
nand I_6494 (I112501,I112493,I137392);
not I_6495 (I112518,I112501);
DFFARX1 I_6496 (I112518,I2067,I112368,I112544,);
not I_6497 (I112552,I112544);
nor I_6498 (I112360,I112402,I112552);
DFFARX1 I_6499 (I137404,I2067,I112368,I112592,);
nor I_6500 (I112351,I112592,I112462);
nor I_6501 (I112342,I112592,I112518);
nand I_6502 (I112628,I137395,I137389);
and I_6503 (I112645,I112628,I137383);
DFFARX1 I_6504 (I112645,I2067,I112368,I112671,);
not I_6505 (I112679,I112671);
nand I_6506 (I112696,I112679,I112592);
nand I_6507 (I112345,I112679,I112501);
nor I_6508 (I112727,I137401,I137389);
and I_6509 (I112744,I112592,I112727);
nor I_6510 (I112761,I112679,I112744);
DFFARX1 I_6511 (I112761,I2067,I112368,I112354,);
nor I_6512 (I112792,I112394,I112727);
DFFARX1 I_6513 (I112792,I2067,I112368,I112339,);
nor I_6514 (I112823,I112671,I112727);
not I_6515 (I112840,I112823);
nand I_6516 (I112348,I112840,I112696);
not I_6517 (I112895,I2074);
DFFARX1 I_6518 (I146646,I2067,I112895,I112921,);
not I_6519 (I112929,I112921);
nand I_6520 (I112946,I146628,I146628);
and I_6521 (I112963,I112946,I146634);
DFFARX1 I_6522 (I112963,I2067,I112895,I112989,);
DFFARX1 I_6523 (I112989,I2067,I112895,I112884,);
DFFARX1 I_6524 (I146631,I2067,I112895,I113020,);
nand I_6525 (I113028,I113020,I146640);
not I_6526 (I113045,I113028);
DFFARX1 I_6527 (I113045,I2067,I112895,I113071,);
not I_6528 (I113079,I113071);
nor I_6529 (I112887,I112929,I113079);
DFFARX1 I_6530 (I146652,I2067,I112895,I113119,);
nor I_6531 (I112878,I113119,I112989);
nor I_6532 (I112869,I113119,I113045);
nand I_6533 (I113155,I146643,I146637);
and I_6534 (I113172,I113155,I146631);
DFFARX1 I_6535 (I113172,I2067,I112895,I113198,);
not I_6536 (I113206,I113198);
nand I_6537 (I113223,I113206,I113119);
nand I_6538 (I112872,I113206,I113028);
nor I_6539 (I113254,I146649,I146637);
and I_6540 (I113271,I113119,I113254);
nor I_6541 (I113288,I113206,I113271);
DFFARX1 I_6542 (I113288,I2067,I112895,I112881,);
nor I_6543 (I113319,I112921,I113254);
DFFARX1 I_6544 (I113319,I2067,I112895,I112866,);
nor I_6545 (I113350,I113198,I113254);
not I_6546 (I113367,I113350);
nand I_6547 (I112875,I113367,I113223);
not I_6548 (I113422,I2074);
DFFARX1 I_6549 (I160070,I2067,I113422,I113448,);
not I_6550 (I113456,I113448);
nand I_6551 (I113473,I160076,I160058);
and I_6552 (I113490,I113473,I160067);
DFFARX1 I_6553 (I113490,I2067,I113422,I113516,);
DFFARX1 I_6554 (I113516,I2067,I113422,I113411,);
DFFARX1 I_6555 (I160073,I2067,I113422,I113547,);
nand I_6556 (I113555,I113547,I160061);
not I_6557 (I113572,I113555);
DFFARX1 I_6558 (I113572,I2067,I113422,I113598,);
not I_6559 (I113606,I113598);
nor I_6560 (I113414,I113456,I113606);
DFFARX1 I_6561 (I160079,I2067,I113422,I113646,);
nor I_6562 (I113405,I113646,I113516);
nor I_6563 (I113396,I113646,I113572);
nand I_6564 (I113682,I160058,I160064);
and I_6565 (I113699,I113682,I160082);
DFFARX1 I_6566 (I113699,I2067,I113422,I113725,);
not I_6567 (I113733,I113725);
nand I_6568 (I113750,I113733,I113646);
nand I_6569 (I113399,I113733,I113555);
nor I_6570 (I113781,I160061,I160064);
and I_6571 (I113798,I113646,I113781);
nor I_6572 (I113815,I113733,I113798);
DFFARX1 I_6573 (I113815,I2067,I113422,I113408,);
nor I_6574 (I113846,I113448,I113781);
DFFARX1 I_6575 (I113846,I2067,I113422,I113393,);
nor I_6576 (I113877,I113725,I113781);
not I_6577 (I113894,I113877);
nand I_6578 (I113402,I113894,I113750);
not I_6579 (I113955,I2074);
DFFARX1 I_6580 (I13280,I2067,I113955,I113981,);
DFFARX1 I_6581 (I13286,I2067,I113955,I113998,);
not I_6582 (I114006,I113998);
not I_6583 (I114023,I13304);
nor I_6584 (I114040,I114023,I13283);
not I_6585 (I114057,I13289);
nor I_6586 (I114074,I114040,I13295);
nor I_6587 (I114091,I113998,I114074);
DFFARX1 I_6588 (I114091,I2067,I113955,I113941,);
nor I_6589 (I114122,I13295,I13283);
nand I_6590 (I114139,I114122,I13304);
DFFARX1 I_6591 (I114139,I2067,I113955,I113944,);
nor I_6592 (I114170,I114057,I13295);
nand I_6593 (I114187,I114170,I13301);
nor I_6594 (I114204,I113981,I114187);
DFFARX1 I_6595 (I114204,I2067,I113955,I113920,);
not I_6596 (I114235,I114187);
nand I_6597 (I113932,I113998,I114235);
DFFARX1 I_6598 (I114187,I2067,I113955,I114275,);
not I_6599 (I114283,I114275);
not I_6600 (I114300,I13295);
not I_6601 (I114317,I13283);
nor I_6602 (I114334,I114317,I13289);
nor I_6603 (I113947,I114283,I114334);
nor I_6604 (I114365,I114317,I13292);
and I_6605 (I114382,I114365,I13280);
or I_6606 (I114399,I114382,I13298);
DFFARX1 I_6607 (I114399,I2067,I113955,I114425,);
nor I_6608 (I113935,I114425,I113981);
not I_6609 (I114447,I114425);
and I_6610 (I114464,I114447,I113981);
nor I_6611 (I113929,I114006,I114464);
nand I_6612 (I114495,I114447,I114057);
nor I_6613 (I113923,I114317,I114495);
nand I_6614 (I113926,I114447,I114235);
nand I_6615 (I114540,I114057,I13283);
nor I_6616 (I113938,I114300,I114540);
not I_6617 (I114601,I2074);
DFFARX1 I_6618 (I55440,I2067,I114601,I114627,);
DFFARX1 I_6619 (I55446,I2067,I114601,I114644,);
not I_6620 (I114652,I114644);
not I_6621 (I114669,I55467);
nor I_6622 (I114686,I114669,I55455);
not I_6623 (I114703,I55464);
nor I_6624 (I114720,I114686,I55449);
nor I_6625 (I114737,I114644,I114720);
DFFARX1 I_6626 (I114737,I2067,I114601,I114587,);
nor I_6627 (I114768,I55449,I55455);
nand I_6628 (I114785,I114768,I55467);
DFFARX1 I_6629 (I114785,I2067,I114601,I114590,);
nor I_6630 (I114816,I114703,I55449);
nand I_6631 (I114833,I114816,I55440);
nor I_6632 (I114850,I114627,I114833);
DFFARX1 I_6633 (I114850,I2067,I114601,I114566,);
not I_6634 (I114881,I114833);
nand I_6635 (I114578,I114644,I114881);
DFFARX1 I_6636 (I114833,I2067,I114601,I114921,);
not I_6637 (I114929,I114921);
not I_6638 (I114946,I55449);
not I_6639 (I114963,I55452);
nor I_6640 (I114980,I114963,I55464);
nor I_6641 (I114593,I114929,I114980);
nor I_6642 (I115011,I114963,I55461);
and I_6643 (I115028,I115011,I55443);
or I_6644 (I115045,I115028,I55458);
DFFARX1 I_6645 (I115045,I2067,I114601,I115071,);
nor I_6646 (I114581,I115071,I114627);
not I_6647 (I115093,I115071);
and I_6648 (I115110,I115093,I114627);
nor I_6649 (I114575,I114652,I115110);
nand I_6650 (I115141,I115093,I114703);
nor I_6651 (I114569,I114963,I115141);
nand I_6652 (I114572,I115093,I114881);
nand I_6653 (I115186,I114703,I55452);
nor I_6654 (I114584,I114946,I115186);
not I_6655 (I115247,I2074);
DFFARX1 I_6656 (I31034,I2067,I115247,I115273,);
DFFARX1 I_6657 (I31046,I2067,I115247,I115290,);
not I_6658 (I115298,I115290);
not I_6659 (I115315,I31052);
nor I_6660 (I115332,I115315,I31037);
not I_6661 (I115349,I31028);
nor I_6662 (I115366,I115332,I31049);
nor I_6663 (I115383,I115290,I115366);
DFFARX1 I_6664 (I115383,I2067,I115247,I115233,);
nor I_6665 (I115414,I31049,I31037);
nand I_6666 (I115431,I115414,I31052);
DFFARX1 I_6667 (I115431,I2067,I115247,I115236,);
nor I_6668 (I115462,I115349,I31049);
nand I_6669 (I115479,I115462,I31031);
nor I_6670 (I115496,I115273,I115479);
DFFARX1 I_6671 (I115496,I2067,I115247,I115212,);
not I_6672 (I115527,I115479);
nand I_6673 (I115224,I115290,I115527);
DFFARX1 I_6674 (I115479,I2067,I115247,I115567,);
not I_6675 (I115575,I115567);
not I_6676 (I115592,I31049);
not I_6677 (I115609,I31040);
nor I_6678 (I115626,I115609,I31028);
nor I_6679 (I115239,I115575,I115626);
nor I_6680 (I115657,I115609,I31043);
and I_6681 (I115674,I115657,I31031);
or I_6682 (I115691,I115674,I31028);
DFFARX1 I_6683 (I115691,I2067,I115247,I115717,);
nor I_6684 (I115227,I115717,I115273);
not I_6685 (I115739,I115717);
and I_6686 (I115756,I115739,I115273);
nor I_6687 (I115221,I115298,I115756);
nand I_6688 (I115787,I115739,I115349);
nor I_6689 (I115215,I115609,I115787);
nand I_6690 (I115218,I115739,I115527);
nand I_6691 (I115832,I115349,I31040);
nor I_6692 (I115230,I115592,I115832);
not I_6693 (I115893,I2074);
DFFARX1 I_6694 (I26274,I2067,I115893,I115919,);
DFFARX1 I_6695 (I26286,I2067,I115893,I115936,);
not I_6696 (I115944,I115936);
not I_6697 (I115961,I26292);
nor I_6698 (I115978,I115961,I26277);
not I_6699 (I115995,I26268);
nor I_6700 (I116012,I115978,I26289);
nor I_6701 (I116029,I115936,I116012);
DFFARX1 I_6702 (I116029,I2067,I115893,I115879,);
nor I_6703 (I116060,I26289,I26277);
nand I_6704 (I116077,I116060,I26292);
DFFARX1 I_6705 (I116077,I2067,I115893,I115882,);
nor I_6706 (I116108,I115995,I26289);
nand I_6707 (I116125,I116108,I26271);
nor I_6708 (I116142,I115919,I116125);
DFFARX1 I_6709 (I116142,I2067,I115893,I115858,);
not I_6710 (I116173,I116125);
nand I_6711 (I115870,I115936,I116173);
DFFARX1 I_6712 (I116125,I2067,I115893,I116213,);
not I_6713 (I116221,I116213);
not I_6714 (I116238,I26289);
not I_6715 (I116255,I26280);
nor I_6716 (I116272,I116255,I26268);
nor I_6717 (I115885,I116221,I116272);
nor I_6718 (I116303,I116255,I26283);
and I_6719 (I116320,I116303,I26271);
or I_6720 (I116337,I116320,I26268);
DFFARX1 I_6721 (I116337,I2067,I115893,I116363,);
nor I_6722 (I115873,I116363,I115919);
not I_6723 (I116385,I116363);
and I_6724 (I116402,I116385,I115919);
nor I_6725 (I115867,I115944,I116402);
nand I_6726 (I116433,I116385,I115995);
nor I_6727 (I115861,I116255,I116433);
nand I_6728 (I115864,I116385,I116173);
nand I_6729 (I116478,I115995,I26280);
nor I_6730 (I115876,I116238,I116478);
not I_6731 (I116539,I2074);
DFFARX1 I_6732 (I77849,I2067,I116539,I116565,);
DFFARX1 I_6733 (I77861,I2067,I116539,I116582,);
not I_6734 (I116590,I116582);
not I_6735 (I116607,I77870);
nor I_6736 (I116624,I116607,I77846);
not I_6737 (I116641,I77864);
nor I_6738 (I116658,I116624,I77858);
nor I_6739 (I116675,I116582,I116658);
DFFARX1 I_6740 (I116675,I2067,I116539,I116525,);
nor I_6741 (I116706,I77858,I77846);
nand I_6742 (I116723,I116706,I77870);
DFFARX1 I_6743 (I116723,I2067,I116539,I116528,);
nor I_6744 (I116754,I116641,I77858);
nand I_6745 (I116771,I116754,I77852);
nor I_6746 (I116788,I116565,I116771);
DFFARX1 I_6747 (I116788,I2067,I116539,I116504,);
not I_6748 (I116819,I116771);
nand I_6749 (I116516,I116582,I116819);
DFFARX1 I_6750 (I116771,I2067,I116539,I116859,);
not I_6751 (I116867,I116859);
not I_6752 (I116884,I77858);
not I_6753 (I116901,I77867);
nor I_6754 (I116918,I116901,I77864);
nor I_6755 (I116531,I116867,I116918);
nor I_6756 (I116949,I116901,I77849);
and I_6757 (I116966,I116949,I77846);
or I_6758 (I116983,I116966,I77855);
DFFARX1 I_6759 (I116983,I2067,I116539,I117009,);
nor I_6760 (I116519,I117009,I116565);
not I_6761 (I117031,I117009);
and I_6762 (I117048,I117031,I116565);
nor I_6763 (I116513,I116590,I117048);
nand I_6764 (I117079,I117031,I116641);
nor I_6765 (I116507,I116901,I117079);
nand I_6766 (I116510,I117031,I116819);
nand I_6767 (I117124,I116641,I77867);
nor I_6768 (I116522,I116884,I117124);
not I_6769 (I117185,I2074);
DFFARX1 I_6770 (I15388,I2067,I117185,I117211,);
DFFARX1 I_6771 (I15394,I2067,I117185,I117228,);
not I_6772 (I117236,I117228);
not I_6773 (I117253,I15412);
nor I_6774 (I117270,I117253,I15391);
not I_6775 (I117287,I15397);
nor I_6776 (I117304,I117270,I15403);
nor I_6777 (I117321,I117228,I117304);
DFFARX1 I_6778 (I117321,I2067,I117185,I117171,);
nor I_6779 (I117352,I15403,I15391);
nand I_6780 (I117369,I117352,I15412);
DFFARX1 I_6781 (I117369,I2067,I117185,I117174,);
nor I_6782 (I117400,I117287,I15403);
nand I_6783 (I117417,I117400,I15409);
nor I_6784 (I117434,I117211,I117417);
DFFARX1 I_6785 (I117434,I2067,I117185,I117150,);
not I_6786 (I117465,I117417);
nand I_6787 (I117162,I117228,I117465);
DFFARX1 I_6788 (I117417,I2067,I117185,I117505,);
not I_6789 (I117513,I117505);
not I_6790 (I117530,I15403);
not I_6791 (I117547,I15391);
nor I_6792 (I117564,I117547,I15397);
nor I_6793 (I117177,I117513,I117564);
nor I_6794 (I117595,I117547,I15400);
and I_6795 (I117612,I117595,I15388);
or I_6796 (I117629,I117612,I15406);
DFFARX1 I_6797 (I117629,I2067,I117185,I117655,);
nor I_6798 (I117165,I117655,I117211);
not I_6799 (I117677,I117655);
and I_6800 (I117694,I117677,I117211);
nor I_6801 (I117159,I117236,I117694);
nand I_6802 (I117725,I117677,I117287);
nor I_6803 (I117153,I117547,I117725);
nand I_6804 (I117156,I117677,I117465);
nand I_6805 (I117770,I117287,I15391);
nor I_6806 (I117168,I117530,I117770);
not I_6807 (I117831,I2074);
DFFARX1 I_6808 (I157356,I2067,I117831,I117857,);
DFFARX1 I_6809 (I157362,I2067,I117831,I117874,);
not I_6810 (I117882,I117874);
not I_6811 (I117899,I157359);
nor I_6812 (I117916,I117899,I157338);
not I_6813 (I117933,I157341);
nor I_6814 (I117950,I117916,I157347);
nor I_6815 (I117967,I117874,I117950);
DFFARX1 I_6816 (I117967,I2067,I117831,I117817,);
nor I_6817 (I117998,I157347,I157338);
nand I_6818 (I118015,I117998,I157359);
DFFARX1 I_6819 (I118015,I2067,I117831,I117820,);
nor I_6820 (I118046,I117933,I157347);
nand I_6821 (I118063,I118046,I157341);
nor I_6822 (I118080,I117857,I118063);
DFFARX1 I_6823 (I118080,I2067,I117831,I117796,);
not I_6824 (I118111,I118063);
nand I_6825 (I117808,I117874,I118111);
DFFARX1 I_6826 (I118063,I2067,I117831,I118151,);
not I_6827 (I118159,I118151);
not I_6828 (I118176,I157347);
not I_6829 (I118193,I157350);
nor I_6830 (I118210,I118193,I157341);
nor I_6831 (I117823,I118159,I118210);
nor I_6832 (I118241,I118193,I157338);
and I_6833 (I118258,I118241,I157344);
or I_6834 (I118275,I118258,I157353);
DFFARX1 I_6835 (I118275,I2067,I117831,I118301,);
nor I_6836 (I117811,I118301,I117857);
not I_6837 (I118323,I118301);
and I_6838 (I118340,I118323,I117857);
nor I_6839 (I117805,I117882,I118340);
nand I_6840 (I118371,I118323,I117933);
nor I_6841 (I117799,I118193,I118371);
nand I_6842 (I117802,I118323,I118111);
nand I_6843 (I118416,I117933,I157350);
nor I_6844 (I117814,I118176,I118416);
not I_6845 (I118477,I2074);
DFFARX1 I_6846 (I37579,I2067,I118477,I118503,);
DFFARX1 I_6847 (I37591,I2067,I118477,I118520,);
not I_6848 (I118528,I118520);
not I_6849 (I118545,I37597);
nor I_6850 (I118562,I118545,I37582);
not I_6851 (I118579,I37573);
nor I_6852 (I118596,I118562,I37594);
nor I_6853 (I118613,I118520,I118596);
DFFARX1 I_6854 (I118613,I2067,I118477,I118463,);
nor I_6855 (I118644,I37594,I37582);
nand I_6856 (I118661,I118644,I37597);
DFFARX1 I_6857 (I118661,I2067,I118477,I118466,);
nor I_6858 (I118692,I118579,I37594);
nand I_6859 (I118709,I118692,I37576);
nor I_6860 (I118726,I118503,I118709);
DFFARX1 I_6861 (I118726,I2067,I118477,I118442,);
not I_6862 (I118757,I118709);
nand I_6863 (I118454,I118520,I118757);
DFFARX1 I_6864 (I118709,I2067,I118477,I118797,);
not I_6865 (I118805,I118797);
not I_6866 (I118822,I37594);
not I_6867 (I118839,I37585);
nor I_6868 (I118856,I118839,I37573);
nor I_6869 (I118469,I118805,I118856);
nor I_6870 (I118887,I118839,I37588);
and I_6871 (I118904,I118887,I37576);
or I_6872 (I118921,I118904,I37573);
DFFARX1 I_6873 (I118921,I2067,I118477,I118947,);
nor I_6874 (I118457,I118947,I118503);
not I_6875 (I118969,I118947);
and I_6876 (I118986,I118969,I118503);
nor I_6877 (I118451,I118528,I118986);
nand I_6878 (I119017,I118969,I118579);
nor I_6879 (I118445,I118839,I119017);
nand I_6880 (I118448,I118969,I118757);
nand I_6881 (I119062,I118579,I37585);
nor I_6882 (I118460,I118822,I119062);
not I_6883 (I119123,I2074);
DFFARX1 I_6884 (I65663,I2067,I119123,I119149,);
DFFARX1 I_6885 (I65660,I2067,I119123,I119166,);
not I_6886 (I119174,I119166);
not I_6887 (I119191,I65675);
nor I_6888 (I119208,I119191,I65678);
not I_6889 (I119225,I65666);
nor I_6890 (I119242,I119208,I65672);
nor I_6891 (I119259,I119166,I119242);
DFFARX1 I_6892 (I119259,I2067,I119123,I119109,);
nor I_6893 (I119290,I65672,I65678);
nand I_6894 (I119307,I119290,I65675);
DFFARX1 I_6895 (I119307,I2067,I119123,I119112,);
nor I_6896 (I119338,I119225,I65672);
nand I_6897 (I119355,I119338,I65684);
nor I_6898 (I119372,I119149,I119355);
DFFARX1 I_6899 (I119372,I2067,I119123,I119088,);
not I_6900 (I119403,I119355);
nand I_6901 (I119100,I119166,I119403);
DFFARX1 I_6902 (I119355,I2067,I119123,I119443,);
not I_6903 (I119451,I119443);
not I_6904 (I119468,I65672);
not I_6905 (I119485,I65657);
nor I_6906 (I119502,I119485,I65666);
nor I_6907 (I119115,I119451,I119502);
nor I_6908 (I119533,I119485,I65669);
and I_6909 (I119550,I119533,I65657);
or I_6910 (I119567,I119550,I65681);
DFFARX1 I_6911 (I119567,I2067,I119123,I119593,);
nor I_6912 (I119103,I119593,I119149);
not I_6913 (I119615,I119593);
and I_6914 (I119632,I119615,I119149);
nor I_6915 (I119097,I119174,I119632);
nand I_6916 (I119663,I119615,I119225);
nor I_6917 (I119091,I119485,I119663);
nand I_6918 (I119094,I119615,I119403);
nand I_6919 (I119708,I119225,I65657);
nor I_6920 (I119106,I119468,I119708);
not I_6921 (I119769,I2074);
DFFARX1 I_6922 (I23311,I2067,I119769,I119795,);
DFFARX1 I_6923 (I23314,I2067,I119769,I119812,);
not I_6924 (I119820,I119812);
not I_6925 (I119837,I23299);
nor I_6926 (I119854,I119837,I23293);
not I_6927 (I119871,I23302);
nor I_6928 (I119888,I119854,I23317);
nor I_6929 (I119905,I119812,I119888);
DFFARX1 I_6930 (I119905,I2067,I119769,I119755,);
nor I_6931 (I119936,I23317,I23293);
nand I_6932 (I119953,I119936,I23299);
DFFARX1 I_6933 (I119953,I2067,I119769,I119758,);
nor I_6934 (I119984,I119871,I23317);
nand I_6935 (I120001,I119984,I23320);
nor I_6936 (I120018,I119795,I120001);
DFFARX1 I_6937 (I120018,I2067,I119769,I119734,);
not I_6938 (I120049,I120001);
nand I_6939 (I119746,I119812,I120049);
DFFARX1 I_6940 (I120001,I2067,I119769,I120089,);
not I_6941 (I120097,I120089);
not I_6942 (I120114,I23317);
not I_6943 (I120131,I23296);
nor I_6944 (I120148,I120131,I23302);
nor I_6945 (I119761,I120097,I120148);
nor I_6946 (I120179,I120131,I23305);
and I_6947 (I120196,I120179,I23293);
or I_6948 (I120213,I120196,I23308);
DFFARX1 I_6949 (I120213,I2067,I119769,I120239,);
nor I_6950 (I119749,I120239,I119795);
not I_6951 (I120261,I120239);
and I_6952 (I120278,I120261,I119795);
nor I_6953 (I119743,I119820,I120278);
nand I_6954 (I120309,I120261,I119871);
nor I_6955 (I119737,I120131,I120309);
nand I_6956 (I119740,I120261,I120049);
nand I_6957 (I120354,I119871,I23296);
nor I_6958 (I119752,I120114,I120354);
not I_6959 (I120415,I2074);
DFFARX1 I_6960 (I176429,I2067,I120415,I120441,);
DFFARX1 I_6961 (I176453,I2067,I120415,I120458,);
not I_6962 (I120466,I120458);
not I_6963 (I120483,I176435);
nor I_6964 (I120500,I120483,I176444);
not I_6965 (I120517,I176429);
nor I_6966 (I120534,I120500,I176450);
nor I_6967 (I120551,I120458,I120534);
DFFARX1 I_6968 (I120551,I2067,I120415,I120401,);
nor I_6969 (I120582,I176450,I176444);
nand I_6970 (I120599,I120582,I176435);
DFFARX1 I_6971 (I120599,I2067,I120415,I120404,);
nor I_6972 (I120630,I120517,I176450);
nand I_6973 (I120647,I120630,I176447);
nor I_6974 (I120664,I120441,I120647);
DFFARX1 I_6975 (I120664,I2067,I120415,I120380,);
not I_6976 (I120695,I120647);
nand I_6977 (I120392,I120458,I120695);
DFFARX1 I_6978 (I120647,I2067,I120415,I120735,);
not I_6979 (I120743,I120735);
not I_6980 (I120760,I176450);
not I_6981 (I120777,I176441);
nor I_6982 (I120794,I120777,I176429);
nor I_6983 (I120407,I120743,I120794);
nor I_6984 (I120825,I120777,I176432);
and I_6985 (I120842,I120825,I176456);
or I_6986 (I120859,I120842,I176438);
DFFARX1 I_6987 (I120859,I2067,I120415,I120885,);
nor I_6988 (I120395,I120885,I120441);
not I_6989 (I120907,I120885);
and I_6990 (I120924,I120907,I120441);
nor I_6991 (I120389,I120466,I120924);
nand I_6992 (I120955,I120907,I120517);
nor I_6993 (I120383,I120777,I120955);
nand I_6994 (I120386,I120907,I120695);
nand I_6995 (I121000,I120517,I176441);
nor I_6996 (I120398,I120760,I121000);
not I_6997 (I121061,I2074);
DFFARX1 I_6998 (I57021,I2067,I121061,I121087,);
DFFARX1 I_6999 (I57027,I2067,I121061,I121104,);
not I_7000 (I121112,I121104);
not I_7001 (I121129,I57048);
nor I_7002 (I121146,I121129,I57036);
not I_7003 (I121163,I57045);
nor I_7004 (I121180,I121146,I57030);
nor I_7005 (I121197,I121104,I121180);
DFFARX1 I_7006 (I121197,I2067,I121061,I121047,);
nor I_7007 (I121228,I57030,I57036);
nand I_7008 (I121245,I121228,I57048);
DFFARX1 I_7009 (I121245,I2067,I121061,I121050,);
nor I_7010 (I121276,I121163,I57030);
nand I_7011 (I121293,I121276,I57021);
nor I_7012 (I121310,I121087,I121293);
DFFARX1 I_7013 (I121310,I2067,I121061,I121026,);
not I_7014 (I121341,I121293);
nand I_7015 (I121038,I121104,I121341);
DFFARX1 I_7016 (I121293,I2067,I121061,I121381,);
not I_7017 (I121389,I121381);
not I_7018 (I121406,I57030);
not I_7019 (I121423,I57033);
nor I_7020 (I121440,I121423,I57045);
nor I_7021 (I121053,I121389,I121440);
nor I_7022 (I121471,I121423,I57042);
and I_7023 (I121488,I121471,I57024);
or I_7024 (I121505,I121488,I57039);
DFFARX1 I_7025 (I121505,I2067,I121061,I121531,);
nor I_7026 (I121041,I121531,I121087);
not I_7027 (I121553,I121531);
and I_7028 (I121570,I121553,I121087);
nor I_7029 (I121035,I121112,I121570);
nand I_7030 (I121601,I121553,I121163);
nor I_7031 (I121029,I121423,I121601);
nand I_7032 (I121032,I121553,I121341);
nand I_7033 (I121646,I121163,I57033);
nor I_7034 (I121044,I121406,I121646);
not I_7035 (I121707,I2074);
DFFARX1 I_7036 (I40554,I2067,I121707,I121733,);
DFFARX1 I_7037 (I40566,I2067,I121707,I121750,);
not I_7038 (I121758,I121750);
not I_7039 (I121775,I40572);
nor I_7040 (I121792,I121775,I40557);
not I_7041 (I121809,I40548);
nor I_7042 (I121826,I121792,I40569);
nor I_7043 (I121843,I121750,I121826);
DFFARX1 I_7044 (I121843,I2067,I121707,I121693,);
nor I_7045 (I121874,I40569,I40557);
nand I_7046 (I121891,I121874,I40572);
DFFARX1 I_7047 (I121891,I2067,I121707,I121696,);
nor I_7048 (I121922,I121809,I40569);
nand I_7049 (I121939,I121922,I40551);
nor I_7050 (I121956,I121733,I121939);
DFFARX1 I_7051 (I121956,I2067,I121707,I121672,);
not I_7052 (I121987,I121939);
nand I_7053 (I121684,I121750,I121987);
DFFARX1 I_7054 (I121939,I2067,I121707,I122027,);
not I_7055 (I122035,I122027);
not I_7056 (I122052,I40569);
not I_7057 (I122069,I40560);
nor I_7058 (I122086,I122069,I40548);
nor I_7059 (I121699,I122035,I122086);
nor I_7060 (I122117,I122069,I40563);
and I_7061 (I122134,I122117,I40551);
or I_7062 (I122151,I122134,I40548);
DFFARX1 I_7063 (I122151,I2067,I121707,I122177,);
nor I_7064 (I121687,I122177,I121733);
not I_7065 (I122199,I122177);
and I_7066 (I122216,I122199,I121733);
nor I_7067 (I121681,I121758,I122216);
nand I_7068 (I122247,I122199,I121809);
nor I_7069 (I121675,I122069,I122247);
nand I_7070 (I121678,I122199,I121987);
nand I_7071 (I122292,I121809,I40560);
nor I_7072 (I121690,I122052,I122292);
not I_7073 (I122353,I2074);
DFFARX1 I_7074 (I111818,I2067,I122353,I122379,);
DFFARX1 I_7075 (I111815,I2067,I122353,I122396,);
not I_7076 (I122404,I122396);
not I_7077 (I122421,I111815);
nor I_7078 (I122438,I122421,I111818);
not I_7079 (I122455,I111830);
nor I_7080 (I122472,I122438,I111824);
nor I_7081 (I122489,I122396,I122472);
DFFARX1 I_7082 (I122489,I2067,I122353,I122339,);
nor I_7083 (I122520,I111824,I111818);
nand I_7084 (I122537,I122520,I111815);
DFFARX1 I_7085 (I122537,I2067,I122353,I122342,);
nor I_7086 (I122568,I122455,I111824);
nand I_7087 (I122585,I122568,I111812);
nor I_7088 (I122602,I122379,I122585);
DFFARX1 I_7089 (I122602,I2067,I122353,I122318,);
not I_7090 (I122633,I122585);
nand I_7091 (I122330,I122396,I122633);
DFFARX1 I_7092 (I122585,I2067,I122353,I122673,);
not I_7093 (I122681,I122673);
not I_7094 (I122698,I111824);
not I_7095 (I122715,I111821);
nor I_7096 (I122732,I122715,I111830);
nor I_7097 (I122345,I122681,I122732);
nor I_7098 (I122763,I122715,I111827);
and I_7099 (I122780,I122763,I111833);
or I_7100 (I122797,I122780,I111812);
DFFARX1 I_7101 (I122797,I2067,I122353,I122823,);
nor I_7102 (I122333,I122823,I122379);
not I_7103 (I122845,I122823);
and I_7104 (I122862,I122845,I122379);
nor I_7105 (I122327,I122404,I122862);
nand I_7106 (I122893,I122845,I122455);
nor I_7107 (I122321,I122715,I122893);
nand I_7108 (I122324,I122845,I122633);
nand I_7109 (I122938,I122455,I111821);
nor I_7110 (I122336,I122698,I122938);
not I_7111 (I122999,I2074);
DFFARX1 I_7112 (I8537,I2067,I122999,I123025,);
DFFARX1 I_7113 (I8543,I2067,I122999,I123042,);
not I_7114 (I123050,I123042);
not I_7115 (I123067,I8537);
nor I_7116 (I123084,I123067,I8549);
not I_7117 (I123101,I8561);
nor I_7118 (I123118,I123084,I8555);
nor I_7119 (I123135,I123042,I123118);
DFFARX1 I_7120 (I123135,I2067,I122999,I122985,);
nor I_7121 (I123166,I8555,I8549);
nand I_7122 (I123183,I123166,I8537);
DFFARX1 I_7123 (I123183,I2067,I122999,I122988,);
nor I_7124 (I123214,I123101,I8555);
nand I_7125 (I123231,I123214,I8540);
nor I_7126 (I123248,I123025,I123231);
DFFARX1 I_7127 (I123248,I2067,I122999,I122964,);
not I_7128 (I123279,I123231);
nand I_7129 (I122976,I123042,I123279);
DFFARX1 I_7130 (I123231,I2067,I122999,I123319,);
not I_7131 (I123327,I123319);
not I_7132 (I123344,I8555);
not I_7133 (I123361,I8540);
nor I_7134 (I123378,I123361,I8561);
nor I_7135 (I122991,I123327,I123378);
nor I_7136 (I123409,I123361,I8558);
and I_7137 (I123426,I123409,I8552);
or I_7138 (I123443,I123426,I8546);
DFFARX1 I_7139 (I123443,I2067,I122999,I123469,);
nor I_7140 (I122979,I123469,I123025);
not I_7141 (I123491,I123469);
and I_7142 (I123508,I123491,I123025);
nor I_7143 (I122973,I123050,I123508);
nand I_7144 (I123539,I123491,I123101);
nor I_7145 (I122967,I123361,I123539);
nand I_7146 (I122970,I123491,I123279);
nand I_7147 (I123584,I123101,I8540);
nor I_7148 (I122982,I123344,I123584);
not I_7149 (I123645,I2074);
DFFARX1 I_7150 (I94036,I2067,I123645,I123671,);
DFFARX1 I_7151 (I94030,I2067,I123645,I123688,);
not I_7152 (I123696,I123688);
not I_7153 (I123713,I94045);
nor I_7154 (I123730,I123713,I94030);
not I_7155 (I123747,I94039);
nor I_7156 (I123764,I123730,I94048);
nor I_7157 (I123781,I123688,I123764);
DFFARX1 I_7158 (I123781,I2067,I123645,I123631,);
nor I_7159 (I123812,I94048,I94030);
nand I_7160 (I123829,I123812,I94045);
DFFARX1 I_7161 (I123829,I2067,I123645,I123634,);
nor I_7162 (I123860,I123747,I94048);
nand I_7163 (I123877,I123860,I94033);
nor I_7164 (I123894,I123671,I123877);
DFFARX1 I_7165 (I123894,I2067,I123645,I123610,);
not I_7166 (I123925,I123877);
nand I_7167 (I123622,I123688,I123925);
DFFARX1 I_7168 (I123877,I2067,I123645,I123965,);
not I_7169 (I123973,I123965);
not I_7170 (I123990,I94048);
not I_7171 (I124007,I94042);
nor I_7172 (I124024,I124007,I94039);
nor I_7173 (I123637,I123973,I124024);
nor I_7174 (I124055,I124007,I94051);
and I_7175 (I124072,I124055,I94054);
or I_7176 (I124089,I124072,I94033);
DFFARX1 I_7177 (I124089,I2067,I123645,I124115,);
nor I_7178 (I123625,I124115,I123671);
not I_7179 (I124137,I124115);
and I_7180 (I124154,I124137,I123671);
nor I_7181 (I123619,I123696,I124154);
nand I_7182 (I124185,I124137,I123747);
nor I_7183 (I123613,I124007,I124185);
nand I_7184 (I123616,I124137,I123925);
nand I_7185 (I124230,I123747,I94042);
nor I_7186 (I123628,I123990,I124230);
not I_7187 (I124291,I2074);
DFFARX1 I_7188 (I141444,I2067,I124291,I124317,);
DFFARX1 I_7189 (I141426,I2067,I124291,I124334,);
not I_7190 (I124342,I124334);
not I_7191 (I124359,I141435);
nor I_7192 (I124376,I124359,I141447);
not I_7193 (I124393,I141429);
nor I_7194 (I124410,I124376,I141438);
nor I_7195 (I124427,I124334,I124410);
DFFARX1 I_7196 (I124427,I2067,I124291,I124277,);
nor I_7197 (I124458,I141438,I141447);
nand I_7198 (I124475,I124458,I141435);
DFFARX1 I_7199 (I124475,I2067,I124291,I124280,);
nor I_7200 (I124506,I124393,I141438);
nand I_7201 (I124523,I124506,I141450);
nor I_7202 (I124540,I124317,I124523);
DFFARX1 I_7203 (I124540,I2067,I124291,I124256,);
not I_7204 (I124571,I124523);
nand I_7205 (I124268,I124334,I124571);
DFFARX1 I_7206 (I124523,I2067,I124291,I124611,);
not I_7207 (I124619,I124611);
not I_7208 (I124636,I141438);
not I_7209 (I124653,I141426);
nor I_7210 (I124670,I124653,I141429);
nor I_7211 (I124283,I124619,I124670);
nor I_7212 (I124701,I124653,I141432);
and I_7213 (I124718,I124701,I141441);
or I_7214 (I124735,I124718,I141429);
DFFARX1 I_7215 (I124735,I2067,I124291,I124761,);
nor I_7216 (I124271,I124761,I124317);
not I_7217 (I124783,I124761);
and I_7218 (I124800,I124783,I124317);
nor I_7219 (I124265,I124342,I124800);
nand I_7220 (I124831,I124783,I124393);
nor I_7221 (I124259,I124653,I124831);
nand I_7222 (I124262,I124783,I124571);
nand I_7223 (I124876,I124393,I141426);
nor I_7224 (I124274,I124636,I124876);
not I_7225 (I124937,I2074);
DFFARX1 I_7226 (I63487,I2067,I124937,I124963,);
DFFARX1 I_7227 (I63484,I2067,I124937,I124980,);
not I_7228 (I124988,I124980);
not I_7229 (I125005,I63499);
nor I_7230 (I125022,I125005,I63502);
not I_7231 (I125039,I63490);
nor I_7232 (I125056,I125022,I63496);
nor I_7233 (I125073,I124980,I125056);
DFFARX1 I_7234 (I125073,I2067,I124937,I124923,);
nor I_7235 (I125104,I63496,I63502);
nand I_7236 (I125121,I125104,I63499);
DFFARX1 I_7237 (I125121,I2067,I124937,I124926,);
nor I_7238 (I125152,I125039,I63496);
nand I_7239 (I125169,I125152,I63508);
nor I_7240 (I125186,I124963,I125169);
DFFARX1 I_7241 (I125186,I2067,I124937,I124902,);
not I_7242 (I125217,I125169);
nand I_7243 (I124914,I124980,I125217);
DFFARX1 I_7244 (I125169,I2067,I124937,I125257,);
not I_7245 (I125265,I125257);
not I_7246 (I125282,I63496);
not I_7247 (I125299,I63481);
nor I_7248 (I125316,I125299,I63490);
nor I_7249 (I124929,I125265,I125316);
nor I_7250 (I125347,I125299,I63493);
and I_7251 (I125364,I125347,I63481);
or I_7252 (I125381,I125364,I63505);
DFFARX1 I_7253 (I125381,I2067,I124937,I125407,);
nor I_7254 (I124917,I125407,I124963);
not I_7255 (I125429,I125407);
and I_7256 (I125446,I125429,I124963);
nor I_7257 (I124911,I124988,I125446);
nand I_7258 (I125477,I125429,I125039);
nor I_7259 (I124905,I125299,I125477);
nand I_7260 (I124908,I125429,I125217);
nand I_7261 (I125522,I125039,I63481);
nor I_7262 (I124920,I125282,I125522);
not I_7263 (I125583,I2074);
DFFARX1 I_7264 (I88834,I2067,I125583,I125609,);
DFFARX1 I_7265 (I88828,I2067,I125583,I125626,);
not I_7266 (I125634,I125626);
not I_7267 (I125651,I88843);
nor I_7268 (I125668,I125651,I88828);
not I_7269 (I125685,I88837);
nor I_7270 (I125702,I125668,I88846);
nor I_7271 (I125719,I125626,I125702);
DFFARX1 I_7272 (I125719,I2067,I125583,I125569,);
nor I_7273 (I125750,I88846,I88828);
nand I_7274 (I125767,I125750,I88843);
DFFARX1 I_7275 (I125767,I2067,I125583,I125572,);
nor I_7276 (I125798,I125685,I88846);
nand I_7277 (I125815,I125798,I88831);
nor I_7278 (I125832,I125609,I125815);
DFFARX1 I_7279 (I125832,I2067,I125583,I125548,);
not I_7280 (I125863,I125815);
nand I_7281 (I125560,I125626,I125863);
DFFARX1 I_7282 (I125815,I2067,I125583,I125903,);
not I_7283 (I125911,I125903);
not I_7284 (I125928,I88846);
not I_7285 (I125945,I88840);
nor I_7286 (I125962,I125945,I88837);
nor I_7287 (I125575,I125911,I125962);
nor I_7288 (I125993,I125945,I88849);
and I_7289 (I126010,I125993,I88852);
or I_7290 (I126027,I126010,I88831);
DFFARX1 I_7291 (I126027,I2067,I125583,I126053,);
nor I_7292 (I125563,I126053,I125609);
not I_7293 (I126075,I126053);
and I_7294 (I126092,I126075,I125609);
nor I_7295 (I125557,I125634,I126092);
nand I_7296 (I126123,I126075,I125685);
nor I_7297 (I125551,I125945,I126123);
nand I_7298 (I125554,I126075,I125863);
nand I_7299 (I126168,I125685,I88840);
nor I_7300 (I125566,I125928,I126168);
not I_7301 (I126229,I2074);
DFFARX1 I_7302 (I19077,I2067,I126229,I126255,);
DFFARX1 I_7303 (I19083,I2067,I126229,I126272,);
not I_7304 (I126280,I126272);
not I_7305 (I126297,I19101);
nor I_7306 (I126314,I126297,I19080);
not I_7307 (I126331,I19086);
nor I_7308 (I126348,I126314,I19092);
nor I_7309 (I126365,I126272,I126348);
DFFARX1 I_7310 (I126365,I2067,I126229,I126215,);
nor I_7311 (I126396,I19092,I19080);
nand I_7312 (I126413,I126396,I19101);
DFFARX1 I_7313 (I126413,I2067,I126229,I126218,);
nor I_7314 (I126444,I126331,I19092);
nand I_7315 (I126461,I126444,I19098);
nor I_7316 (I126478,I126255,I126461);
DFFARX1 I_7317 (I126478,I2067,I126229,I126194,);
not I_7318 (I126509,I126461);
nand I_7319 (I126206,I126272,I126509);
DFFARX1 I_7320 (I126461,I2067,I126229,I126549,);
not I_7321 (I126557,I126549);
not I_7322 (I126574,I19092);
not I_7323 (I126591,I19080);
nor I_7324 (I126608,I126591,I19086);
nor I_7325 (I126221,I126557,I126608);
nor I_7326 (I126639,I126591,I19089);
and I_7327 (I126656,I126639,I19077);
or I_7328 (I126673,I126656,I19095);
DFFARX1 I_7329 (I126673,I2067,I126229,I126699,);
nor I_7330 (I126209,I126699,I126255);
not I_7331 (I126721,I126699);
and I_7332 (I126738,I126721,I126255);
nor I_7333 (I126203,I126280,I126738);
nand I_7334 (I126769,I126721,I126331);
nor I_7335 (I126197,I126591,I126769);
nand I_7336 (I126200,I126721,I126509);
nand I_7337 (I126814,I126331,I19080);
nor I_7338 (I126212,I126574,I126814);
not I_7339 (I126875,I2074);
DFFARX1 I_7340 (I72494,I2067,I126875,I126901,);
DFFARX1 I_7341 (I72506,I2067,I126875,I126918,);
not I_7342 (I126926,I126918);
not I_7343 (I126943,I72491);
nor I_7344 (I126960,I126943,I72509);
not I_7345 (I126977,I72515);
nor I_7346 (I126994,I126960,I72497);
nor I_7347 (I127011,I126918,I126994);
DFFARX1 I_7348 (I127011,I2067,I126875,I126861,);
nor I_7349 (I127042,I72497,I72509);
nand I_7350 (I127059,I127042,I72491);
DFFARX1 I_7351 (I127059,I2067,I126875,I126864,);
nor I_7352 (I127090,I126977,I72497);
nand I_7353 (I127107,I127090,I72500);
nor I_7354 (I127124,I126901,I127107);
DFFARX1 I_7355 (I127124,I2067,I126875,I126840,);
not I_7356 (I127155,I127107);
nand I_7357 (I126852,I126918,I127155);
DFFARX1 I_7358 (I127107,I2067,I126875,I127195,);
not I_7359 (I127203,I127195);
not I_7360 (I127220,I72497);
not I_7361 (I127237,I72503);
nor I_7362 (I127254,I127237,I72515);
nor I_7363 (I126867,I127203,I127254);
nor I_7364 (I127285,I127237,I72512);
and I_7365 (I127302,I127285,I72491);
or I_7366 (I127319,I127302,I72494);
DFFARX1 I_7367 (I127319,I2067,I126875,I127345,);
nor I_7368 (I126855,I127345,I126901);
not I_7369 (I127367,I127345);
and I_7370 (I127384,I127367,I126901);
nor I_7371 (I126849,I126926,I127384);
nand I_7372 (I127415,I127367,I126977);
nor I_7373 (I126843,I127237,I127415);
nand I_7374 (I126846,I127367,I127155);
nand I_7375 (I127460,I126977,I72503);
nor I_7376 (I126858,I127220,I127460);
not I_7377 (I127521,I2074);
DFFARX1 I_7378 (I134558,I2067,I127521,I127547,);
DFFARX1 I_7379 (I134561,I2067,I127521,I127564,);
not I_7380 (I127572,I127564);
not I_7381 (I127589,I134558);
nor I_7382 (I127606,I127589,I134570);
not I_7383 (I127623,I134579);
nor I_7384 (I127640,I127606,I134567);
nor I_7385 (I127657,I127564,I127640);
DFFARX1 I_7386 (I127657,I2067,I127521,I127507,);
nor I_7387 (I127688,I134567,I134570);
nand I_7388 (I127705,I127688,I134558);
DFFARX1 I_7389 (I127705,I2067,I127521,I127510,);
nor I_7390 (I127736,I127623,I134567);
nand I_7391 (I127753,I127736,I134573);
nor I_7392 (I127770,I127547,I127753);
DFFARX1 I_7393 (I127770,I2067,I127521,I127486,);
not I_7394 (I127801,I127753);
nand I_7395 (I127498,I127564,I127801);
DFFARX1 I_7396 (I127753,I2067,I127521,I127841,);
not I_7397 (I127849,I127841);
not I_7398 (I127866,I134567);
not I_7399 (I127883,I134564);
nor I_7400 (I127900,I127883,I134579);
nor I_7401 (I127513,I127849,I127900);
nor I_7402 (I127931,I127883,I134576);
and I_7403 (I127948,I127931,I134564);
or I_7404 (I127965,I127948,I134561);
DFFARX1 I_7405 (I127965,I2067,I127521,I127991,);
nor I_7406 (I127501,I127991,I127547);
not I_7407 (I128013,I127991);
and I_7408 (I128030,I128013,I127547);
nor I_7409 (I127495,I127572,I128030);
nand I_7410 (I128061,I128013,I127623);
nor I_7411 (I127489,I127883,I128061);
nand I_7412 (I127492,I128013,I127801);
nand I_7413 (I128106,I127623,I134564);
nor I_7414 (I127504,I127866,I128106);
not I_7415 (I128167,I2074);
DFFARX1 I_7416 (I79005,I2067,I128167,I128193,);
DFFARX1 I_7417 (I79017,I2067,I128167,I128210,);
not I_7418 (I128218,I128210);
not I_7419 (I128235,I79026);
nor I_7420 (I128252,I128235,I79002);
not I_7421 (I128269,I79020);
nor I_7422 (I128286,I128252,I79014);
nor I_7423 (I128303,I128210,I128286);
DFFARX1 I_7424 (I128303,I2067,I128167,I128153,);
nor I_7425 (I128334,I79014,I79002);
nand I_7426 (I128351,I128334,I79026);
DFFARX1 I_7427 (I128351,I2067,I128167,I128156,);
nor I_7428 (I128382,I128269,I79014);
nand I_7429 (I128399,I128382,I79008);
nor I_7430 (I128416,I128193,I128399);
DFFARX1 I_7431 (I128416,I2067,I128167,I128132,);
not I_7432 (I128447,I128399);
nand I_7433 (I128144,I128210,I128447);
DFFARX1 I_7434 (I128399,I2067,I128167,I128487,);
not I_7435 (I128495,I128487);
not I_7436 (I128512,I79014);
not I_7437 (I128529,I79023);
nor I_7438 (I128546,I128529,I79020);
nor I_7439 (I128159,I128495,I128546);
nor I_7440 (I128577,I128529,I79005);
and I_7441 (I128594,I128577,I79002);
or I_7442 (I128611,I128594,I79011);
DFFARX1 I_7443 (I128611,I2067,I128167,I128637,);
nor I_7444 (I128147,I128637,I128193);
not I_7445 (I128659,I128637);
and I_7446 (I128676,I128659,I128193);
nor I_7447 (I128141,I128218,I128676);
nand I_7448 (I128707,I128659,I128269);
nor I_7449 (I128135,I128529,I128707);
nand I_7450 (I128138,I128659,I128447);
nand I_7451 (I128752,I128269,I79023);
nor I_7452 (I128150,I128512,I128752);
not I_7453 (I128813,I2074);
DFFARX1 I_7454 (I41738,I2067,I128813,I128839,);
DFFARX1 I_7455 (I41744,I2067,I128813,I128856,);
not I_7456 (I128864,I128856);
not I_7457 (I128881,I41765);
nor I_7458 (I128898,I128881,I41753);
not I_7459 (I128915,I41762);
nor I_7460 (I128932,I128898,I41747);
nor I_7461 (I128949,I128856,I128932);
DFFARX1 I_7462 (I128949,I2067,I128813,I128799,);
nor I_7463 (I128980,I41747,I41753);
nand I_7464 (I128997,I128980,I41765);
DFFARX1 I_7465 (I128997,I2067,I128813,I128802,);
nor I_7466 (I129028,I128915,I41747);
nand I_7467 (I129045,I129028,I41738);
nor I_7468 (I129062,I128839,I129045);
DFFARX1 I_7469 (I129062,I2067,I128813,I128778,);
not I_7470 (I129093,I129045);
nand I_7471 (I128790,I128856,I129093);
DFFARX1 I_7472 (I129045,I2067,I128813,I129133,);
not I_7473 (I129141,I129133);
not I_7474 (I129158,I41747);
not I_7475 (I129175,I41750);
nor I_7476 (I129192,I129175,I41762);
nor I_7477 (I128805,I129141,I129192);
nor I_7478 (I129223,I129175,I41759);
and I_7479 (I129240,I129223,I41741);
or I_7480 (I129257,I129240,I41756);
DFFARX1 I_7481 (I129257,I2067,I128813,I129283,);
nor I_7482 (I128793,I129283,I128839);
not I_7483 (I129305,I129283);
and I_7484 (I129322,I129305,I128839);
nor I_7485 (I128787,I128864,I129322);
nand I_7486 (I129353,I129305,I128915);
nor I_7487 (I128781,I129175,I129353);
nand I_7488 (I128784,I129305,I129093);
nand I_7489 (I129398,I128915,I41750);
nor I_7490 (I128796,I129158,I129398);
not I_7491 (I129459,I2074);
DFFARX1 I_7492 (I136820,I2067,I129459,I129485,);
DFFARX1 I_7493 (I136802,I2067,I129459,I129502,);
not I_7494 (I129510,I129502);
not I_7495 (I129527,I136811);
nor I_7496 (I129544,I129527,I136823);
not I_7497 (I129561,I136805);
nor I_7498 (I129578,I129544,I136814);
nor I_7499 (I129595,I129502,I129578);
DFFARX1 I_7500 (I129595,I2067,I129459,I129445,);
nor I_7501 (I129626,I136814,I136823);
nand I_7502 (I129643,I129626,I136811);
DFFARX1 I_7503 (I129643,I2067,I129459,I129448,);
nor I_7504 (I129674,I129561,I136814);
nand I_7505 (I129691,I129674,I136826);
nor I_7506 (I129708,I129485,I129691);
DFFARX1 I_7507 (I129708,I2067,I129459,I129424,);
not I_7508 (I129739,I129691);
nand I_7509 (I129436,I129502,I129739);
DFFARX1 I_7510 (I129691,I2067,I129459,I129779,);
not I_7511 (I129787,I129779);
not I_7512 (I129804,I136814);
not I_7513 (I129821,I136802);
nor I_7514 (I129838,I129821,I136805);
nor I_7515 (I129451,I129787,I129838);
nor I_7516 (I129869,I129821,I136808);
and I_7517 (I129886,I129869,I136817);
or I_7518 (I129903,I129886,I136805);
DFFARX1 I_7519 (I129903,I2067,I129459,I129929,);
nor I_7520 (I129439,I129929,I129485);
not I_7521 (I129951,I129929);
and I_7522 (I129968,I129951,I129485);
nor I_7523 (I129433,I129510,I129968);
nand I_7524 (I129999,I129951,I129561);
nor I_7525 (I129427,I129821,I129999);
nand I_7526 (I129430,I129951,I129739);
nand I_7527 (I130044,I129561,I136802);
nor I_7528 (I129442,I129804,I130044);
not I_7529 (I130099,I2074);
DFFARX1 I_7530 (I20143,I2067,I130099,I130125,);
DFFARX1 I_7531 (I130125,I2067,I130099,I130142,);
not I_7532 (I130091,I130142);
not I_7533 (I130164,I130125);
DFFARX1 I_7534 (I20131,I2067,I130099,I130190,);
nand I_7535 (I130198,I130190,I20146);
not I_7536 (I130215,I20146);
not I_7537 (I130232,I20134);
nand I_7538 (I130249,I20155,I20149);
and I_7539 (I130266,I20155,I20149);
not I_7540 (I130283,I20137);
nand I_7541 (I130300,I130283,I130232);
nor I_7542 (I130073,I130300,I130198);
nor I_7543 (I130331,I130215,I130300);
nand I_7544 (I130076,I130266,I130331);
not I_7545 (I130362,I20140);
nor I_7546 (I130379,I130362,I20155);
nor I_7547 (I130396,I130379,I20137);
nor I_7548 (I130413,I130164,I130396);
DFFARX1 I_7549 (I130413,I2067,I130099,I130085,);
not I_7550 (I130444,I130379);
DFFARX1 I_7551 (I130444,I2067,I130099,I130088,);
and I_7552 (I130082,I130190,I130379);
nor I_7553 (I130489,I130362,I20134);
and I_7554 (I130506,I130489,I20131);
or I_7555 (I130523,I130506,I20152);
DFFARX1 I_7556 (I130523,I2067,I130099,I130549,);
nor I_7557 (I130557,I130549,I130283);
DFFARX1 I_7558 (I130557,I2067,I130099,I130070,);
nand I_7559 (I130588,I130549,I130190);
nand I_7560 (I130605,I130283,I130588);
nor I_7561 (I130079,I130605,I130249);
not I_7562 (I130660,I2074);
DFFARX1 I_7563 (I152992,I2067,I130660,I130686,);
DFFARX1 I_7564 (I130686,I2067,I130660,I130703,);
not I_7565 (I130652,I130703);
not I_7566 (I130725,I130686);
DFFARX1 I_7567 (I152998,I2067,I130660,I130751,);
nand I_7568 (I130759,I130751,I153007);
not I_7569 (I130776,I153007);
not I_7570 (I130793,I152986);
nand I_7571 (I130810,I152989,I152989);
and I_7572 (I130827,I152989,I152989);
not I_7573 (I130844,I153001);
nand I_7574 (I130861,I130844,I130793);
nor I_7575 (I130634,I130861,I130759);
nor I_7576 (I130892,I130776,I130861);
nand I_7577 (I130637,I130827,I130892);
not I_7578 (I130923,I152995);
nor I_7579 (I130940,I130923,I152989);
nor I_7580 (I130957,I130940,I153001);
nor I_7581 (I130974,I130725,I130957);
DFFARX1 I_7582 (I130974,I2067,I130660,I130646,);
not I_7583 (I131005,I130940);
DFFARX1 I_7584 (I131005,I2067,I130660,I130649,);
and I_7585 (I130643,I130751,I130940);
nor I_7586 (I131050,I130923,I153010);
and I_7587 (I131067,I131050,I152986);
or I_7588 (I131084,I131067,I153004);
DFFARX1 I_7589 (I131084,I2067,I130660,I131110,);
nor I_7590 (I131118,I131110,I130844);
DFFARX1 I_7591 (I131118,I2067,I130660,I130631,);
nand I_7592 (I131149,I131110,I130751);
nand I_7593 (I131166,I130844,I131149);
nor I_7594 (I130640,I131166,I130810);
not I_7595 (I131221,I2074);
DFFARX1 I_7596 (I153536,I2067,I131221,I131247,);
DFFARX1 I_7597 (I131247,I2067,I131221,I131264,);
not I_7598 (I131213,I131264);
not I_7599 (I131286,I131247);
DFFARX1 I_7600 (I153542,I2067,I131221,I131312,);
nand I_7601 (I131320,I131312,I153551);
not I_7602 (I131337,I153551);
not I_7603 (I131354,I153530);
nand I_7604 (I131371,I153533,I153533);
and I_7605 (I131388,I153533,I153533);
not I_7606 (I131405,I153545);
nand I_7607 (I131422,I131405,I131354);
nor I_7608 (I131195,I131422,I131320);
nor I_7609 (I131453,I131337,I131422);
nand I_7610 (I131198,I131388,I131453);
not I_7611 (I131484,I153539);
nor I_7612 (I131501,I131484,I153533);
nor I_7613 (I131518,I131501,I153545);
nor I_7614 (I131535,I131286,I131518);
DFFARX1 I_7615 (I131535,I2067,I131221,I131207,);
not I_7616 (I131566,I131501);
DFFARX1 I_7617 (I131566,I2067,I131221,I131210,);
and I_7618 (I131204,I131312,I131501);
nor I_7619 (I131611,I131484,I153554);
and I_7620 (I131628,I131611,I153530);
or I_7621 (I131645,I131628,I153548);
DFFARX1 I_7622 (I131645,I2067,I131221,I131671,);
nor I_7623 (I131679,I131671,I131405);
DFFARX1 I_7624 (I131679,I2067,I131221,I131192,);
nand I_7625 (I131710,I131671,I131312);
nand I_7626 (I131727,I131405,I131710);
nor I_7627 (I131201,I131727,I131371);
not I_7628 (I131782,I2074);
DFFARX1 I_7629 (I99235,I2067,I131782,I131808,);
DFFARX1 I_7630 (I131808,I2067,I131782,I131825,);
not I_7631 (I131774,I131825);
not I_7632 (I131847,I131808);
DFFARX1 I_7633 (I99247,I2067,I131782,I131873,);
nand I_7634 (I131881,I131873,I99256);
not I_7635 (I131898,I99256);
not I_7636 (I131915,I99238);
nand I_7637 (I131932,I99241,I99232);
and I_7638 (I131949,I99241,I99232);
not I_7639 (I131966,I99250);
nand I_7640 (I131983,I131966,I131915);
nor I_7641 (I131756,I131983,I131881);
nor I_7642 (I132014,I131898,I131983);
nand I_7643 (I131759,I131949,I132014);
not I_7644 (I132045,I99253);
nor I_7645 (I132062,I132045,I99241);
nor I_7646 (I132079,I132062,I99250);
nor I_7647 (I132096,I131847,I132079);
DFFARX1 I_7648 (I132096,I2067,I131782,I131768,);
not I_7649 (I132127,I132062);
DFFARX1 I_7650 (I132127,I2067,I131782,I131771,);
and I_7651 (I131765,I131873,I132062);
nor I_7652 (I132172,I132045,I99232);
and I_7653 (I132189,I132172,I99244);
or I_7654 (I132206,I132189,I99235);
DFFARX1 I_7655 (I132206,I2067,I131782,I132232,);
nor I_7656 (I132240,I132232,I131966);
DFFARX1 I_7657 (I132240,I2067,I131782,I131753,);
nand I_7658 (I132271,I132232,I131873);
nand I_7659 (I132288,I131966,I132271);
nor I_7660 (I131762,I132288,I131932);
not I_7661 (I132343,I2074);
DFFARX1 I_7662 (I1972,I2067,I132343,I132369,);
DFFARX1 I_7663 (I132369,I2067,I132343,I132386,);
not I_7664 (I132335,I132386);
not I_7665 (I132408,I132369);
DFFARX1 I_7666 (I1652,I2067,I132343,I132434,);
nand I_7667 (I132442,I132434,I1612);
not I_7668 (I132459,I1612);
not I_7669 (I132476,I2036);
nand I_7670 (I132493,I1876,I1892);
and I_7671 (I132510,I1876,I1892);
not I_7672 (I132527,I1684);
nand I_7673 (I132544,I132527,I132476);
nor I_7674 (I132317,I132544,I132442);
nor I_7675 (I132575,I132459,I132544);
nand I_7676 (I132320,I132510,I132575);
not I_7677 (I132606,I1724);
nor I_7678 (I132623,I132606,I1876);
nor I_7679 (I132640,I132623,I1684);
nor I_7680 (I132657,I132408,I132640);
DFFARX1 I_7681 (I132657,I2067,I132343,I132329,);
not I_7682 (I132688,I132623);
DFFARX1 I_7683 (I132688,I2067,I132343,I132332,);
and I_7684 (I132326,I132434,I132623);
nor I_7685 (I132733,I132606,I1484);
and I_7686 (I132750,I132733,I1564);
or I_7687 (I132767,I132750,I1772);
DFFARX1 I_7688 (I132767,I2067,I132343,I132793,);
nor I_7689 (I132801,I132793,I132527);
DFFARX1 I_7690 (I132801,I2067,I132343,I132314,);
nand I_7691 (I132832,I132793,I132434);
nand I_7692 (I132849,I132527,I132832);
nor I_7693 (I132323,I132849,I132493);
not I_7694 (I132904,I2074);
DFFARX1 I_7695 (I117796,I2067,I132904,I132930,);
DFFARX1 I_7696 (I132930,I2067,I132904,I132947,);
not I_7697 (I132896,I132947);
not I_7698 (I132969,I132930);
DFFARX1 I_7699 (I117823,I2067,I132904,I132995,);
nand I_7700 (I133003,I132995,I117814);
not I_7701 (I133020,I117814);
not I_7702 (I133037,I117796);
nand I_7703 (I133054,I117808,I117811);
and I_7704 (I133071,I117808,I117811);
not I_7705 (I133088,I117820);
nand I_7706 (I133105,I133088,I133037);
nor I_7707 (I132878,I133105,I133003);
nor I_7708 (I133136,I133020,I133105);
nand I_7709 (I132881,I133071,I133136);
not I_7710 (I133167,I117805);
nor I_7711 (I133184,I133167,I117808);
nor I_7712 (I133201,I133184,I117820);
nor I_7713 (I133218,I132969,I133201);
DFFARX1 I_7714 (I133218,I2067,I132904,I132890,);
not I_7715 (I133249,I133184);
DFFARX1 I_7716 (I133249,I2067,I132904,I132893,);
and I_7717 (I132887,I132995,I133184);
nor I_7718 (I133294,I133167,I117799);
and I_7719 (I133311,I133294,I117802);
or I_7720 (I133328,I133311,I117817);
DFFARX1 I_7721 (I133328,I2067,I132904,I133354,);
nor I_7722 (I133362,I133354,I133088);
DFFARX1 I_7723 (I133362,I2067,I132904,I132875,);
nand I_7724 (I133393,I133354,I132995);
nand I_7725 (I133410,I133088,I133393);
nor I_7726 (I132884,I133410,I133054);
not I_7727 (I133465,I2074);
DFFARX1 I_7728 (I121026,I2067,I133465,I133491,);
DFFARX1 I_7729 (I133491,I2067,I133465,I133508,);
not I_7730 (I133457,I133508);
not I_7731 (I133530,I133491);
DFFARX1 I_7732 (I121053,I2067,I133465,I133556,);
nand I_7733 (I133564,I133556,I121044);
not I_7734 (I133581,I121044);
not I_7735 (I133598,I121026);
nand I_7736 (I133615,I121038,I121041);
and I_7737 (I133632,I121038,I121041);
not I_7738 (I133649,I121050);
nand I_7739 (I133666,I133649,I133598);
nor I_7740 (I133439,I133666,I133564);
nor I_7741 (I133697,I133581,I133666);
nand I_7742 (I133442,I133632,I133697);
not I_7743 (I133728,I121035);
nor I_7744 (I133745,I133728,I121038);
nor I_7745 (I133762,I133745,I121050);
nor I_7746 (I133779,I133530,I133762);
DFFARX1 I_7747 (I133779,I2067,I133465,I133451,);
not I_7748 (I133810,I133745);
DFFARX1 I_7749 (I133810,I2067,I133465,I133454,);
and I_7750 (I133448,I133556,I133745);
nor I_7751 (I133855,I133728,I121029);
and I_7752 (I133872,I133855,I121032);
or I_7753 (I133889,I133872,I121047);
DFFARX1 I_7754 (I133889,I2067,I133465,I133915,);
nor I_7755 (I133923,I133915,I133649);
DFFARX1 I_7756 (I133923,I2067,I133465,I133436,);
nand I_7757 (I133954,I133915,I133556);
nand I_7758 (I133971,I133649,I133954);
nor I_7759 (I133445,I133971,I133615);
not I_7760 (I134026,I2074);
DFFARX1 I_7761 (I142019,I2067,I134026,I134052,);
DFFARX1 I_7762 (I134052,I2067,I134026,I134069,);
not I_7763 (I134018,I134069);
not I_7764 (I134091,I134052);
DFFARX1 I_7765 (I142010,I2067,I134026,I134117,);
nand I_7766 (I134125,I134117,I142007);
not I_7767 (I134142,I142007);
not I_7768 (I134159,I142016);
nand I_7769 (I134176,I142025,I142007);
and I_7770 (I134193,I142025,I142007);
not I_7771 (I134210,I142004);
nand I_7772 (I134227,I134210,I134159);
nor I_7773 (I134000,I134227,I134125);
nor I_7774 (I134258,I134142,I134227);
nand I_7775 (I134003,I134193,I134258);
not I_7776 (I134289,I142013);
nor I_7777 (I134306,I134289,I142025);
nor I_7778 (I134323,I134306,I142004);
nor I_7779 (I134340,I134091,I134323);
DFFARX1 I_7780 (I134340,I2067,I134026,I134012,);
not I_7781 (I134371,I134306);
DFFARX1 I_7782 (I134371,I2067,I134026,I134015,);
and I_7783 (I134009,I134117,I134306);
nor I_7784 (I134416,I134289,I142028);
and I_7785 (I134433,I134416,I142004);
or I_7786 (I134450,I134433,I142022);
DFFARX1 I_7787 (I134450,I2067,I134026,I134476,);
nor I_7788 (I134484,I134476,I134210);
DFFARX1 I_7789 (I134484,I2067,I134026,I133997,);
nand I_7790 (I134515,I134476,I134117);
nand I_7791 (I134532,I134210,I134515);
nor I_7792 (I134006,I134532,I134176);
not I_7793 (I134587,I2074);
DFFARX1 I_7794 (I165229,I2067,I134587,I134613,);
DFFARX1 I_7795 (I134613,I2067,I134587,I134630,);
not I_7796 (I134579,I134630);
not I_7797 (I134652,I134613);
DFFARX1 I_7798 (I165226,I2067,I134587,I134678,);
nand I_7799 (I134686,I134678,I165232);
not I_7800 (I134703,I165232);
not I_7801 (I134720,I165241);
nand I_7802 (I134737,I165235,I165229);
and I_7803 (I134754,I165235,I165229);
not I_7804 (I134771,I165247);
nand I_7805 (I134788,I134771,I134720);
nor I_7806 (I134561,I134788,I134686);
nor I_7807 (I134819,I134703,I134788);
nand I_7808 (I134564,I134754,I134819);
not I_7809 (I134850,I165244);
nor I_7810 (I134867,I134850,I165235);
nor I_7811 (I134884,I134867,I165247);
nor I_7812 (I134901,I134652,I134884);
DFFARX1 I_7813 (I134901,I2067,I134587,I134573,);
not I_7814 (I134932,I134867);
DFFARX1 I_7815 (I134932,I2067,I134587,I134576,);
and I_7816 (I134570,I134678,I134867);
nor I_7817 (I134977,I134850,I165238);
and I_7818 (I134994,I134977,I165250);
or I_7819 (I135011,I134994,I165226);
DFFARX1 I_7820 (I135011,I2067,I134587,I135037,);
nor I_7821 (I135045,I135037,I134771);
DFFARX1 I_7822 (I135045,I2067,I134587,I134558,);
nand I_7823 (I135076,I135037,I134678);
nand I_7824 (I135093,I134771,I135076);
nor I_7825 (I134567,I135093,I134737);
not I_7826 (I135148,I2074);
DFFARX1 I_7827 (I91143,I2067,I135148,I135174,);
DFFARX1 I_7828 (I135174,I2067,I135148,I135191,);
not I_7829 (I135140,I135191);
not I_7830 (I135213,I135174);
DFFARX1 I_7831 (I91155,I2067,I135148,I135239,);
nand I_7832 (I135247,I135239,I91164);
not I_7833 (I135264,I91164);
not I_7834 (I135281,I91146);
nand I_7835 (I135298,I91149,I91140);
and I_7836 (I135315,I91149,I91140);
not I_7837 (I135332,I91158);
nand I_7838 (I135349,I135332,I135281);
nor I_7839 (I135122,I135349,I135247);
nor I_7840 (I135380,I135264,I135349);
nand I_7841 (I135125,I135315,I135380);
not I_7842 (I135411,I91161);
nor I_7843 (I135428,I135411,I91149);
nor I_7844 (I135445,I135428,I91158);
nor I_7845 (I135462,I135213,I135445);
DFFARX1 I_7846 (I135462,I2067,I135148,I135134,);
not I_7847 (I135493,I135428);
DFFARX1 I_7848 (I135493,I2067,I135148,I135137,);
and I_7849 (I135131,I135239,I135428);
nor I_7850 (I135538,I135411,I91140);
and I_7851 (I135555,I135538,I91152);
or I_7852 (I135572,I135555,I91143);
DFFARX1 I_7853 (I135572,I2067,I135148,I135598,);
nor I_7854 (I135606,I135598,I135332);
DFFARX1 I_7855 (I135606,I2067,I135148,I135119,);
nand I_7856 (I135637,I135598,I135239);
nand I_7857 (I135654,I135332,I135637);
nor I_7858 (I135128,I135654,I135298);
not I_7859 (I135709,I2074);
DFFARX1 I_7860 (I166964,I2067,I135709,I135735,);
DFFARX1 I_7861 (I135735,I2067,I135709,I135752,);
not I_7862 (I135701,I135752);
not I_7863 (I135774,I135735);
DFFARX1 I_7864 (I166949,I2067,I135709,I135800,);
nand I_7865 (I135808,I135800,I166958);
not I_7866 (I135825,I166958);
not I_7867 (I135842,I166952);
nand I_7868 (I135859,I166970,I166967);
and I_7869 (I135876,I166970,I166967);
not I_7870 (I135893,I166943);
nand I_7871 (I135910,I135893,I135842);
nor I_7872 (I135683,I135910,I135808);
nor I_7873 (I135941,I135825,I135910);
nand I_7874 (I135686,I135876,I135941);
not I_7875 (I135972,I166946);
nor I_7876 (I135989,I135972,I166970);
nor I_7877 (I136006,I135989,I166943);
nor I_7878 (I136023,I135774,I136006);
DFFARX1 I_7879 (I136023,I2067,I135709,I135695,);
not I_7880 (I136054,I135989);
DFFARX1 I_7881 (I136054,I2067,I135709,I135698,);
and I_7882 (I135692,I135800,I135989);
nor I_7883 (I136099,I135972,I166943);
and I_7884 (I136116,I136099,I166961);
or I_7885 (I136133,I136116,I166955);
DFFARX1 I_7886 (I136133,I2067,I135709,I136159,);
nor I_7887 (I136167,I136159,I135893);
DFFARX1 I_7888 (I136167,I2067,I135709,I135680,);
nand I_7889 (I136198,I136159,I135800);
nand I_7890 (I136215,I135893,I136198);
nor I_7891 (I135689,I136215,I135859);
not I_7892 (I136270,I2074);
DFFARX1 I_7893 (I99813,I2067,I136270,I136296,);
DFFARX1 I_7894 (I136296,I2067,I136270,I136313,);
not I_7895 (I136262,I136313);
not I_7896 (I136335,I136296);
DFFARX1 I_7897 (I99825,I2067,I136270,I136361,);
nand I_7898 (I136369,I136361,I99834);
not I_7899 (I136386,I99834);
not I_7900 (I136403,I99816);
nand I_7901 (I136420,I99819,I99810);
and I_7902 (I136437,I99819,I99810);
not I_7903 (I136454,I99828);
nand I_7904 (I136471,I136454,I136403);
nor I_7905 (I136244,I136471,I136369);
nor I_7906 (I136502,I136386,I136471);
nand I_7907 (I136247,I136437,I136502);
not I_7908 (I136533,I99831);
nor I_7909 (I136550,I136533,I99819);
nor I_7910 (I136567,I136550,I99828);
nor I_7911 (I136584,I136335,I136567);
DFFARX1 I_7912 (I136584,I2067,I136270,I136256,);
not I_7913 (I136615,I136550);
DFFARX1 I_7914 (I136615,I2067,I136270,I136259,);
and I_7915 (I136253,I136361,I136550);
nor I_7916 (I136660,I136533,I99810);
and I_7917 (I136677,I136660,I99822);
or I_7918 (I136694,I136677,I99813);
DFFARX1 I_7919 (I136694,I2067,I136270,I136720,);
nor I_7920 (I136728,I136720,I136454);
DFFARX1 I_7921 (I136728,I2067,I136270,I136241,);
nand I_7922 (I136759,I136720,I136361);
nand I_7923 (I136776,I136454,I136759);
nor I_7924 (I136250,I136776,I136420);
not I_7925 (I136834,I2074);
DFFARX1 I_7926 (I1492,I2067,I136834,I136860,);
and I_7927 (I136868,I136860,I1796);
DFFARX1 I_7928 (I136868,I2067,I136834,I136817,);
DFFARX1 I_7929 (I1388,I2067,I136834,I136908,);
not I_7930 (I136916,I1708);
not I_7931 (I136933,I1924);
nand I_7932 (I136950,I136933,I136916);
nor I_7933 (I136805,I136908,I136950);
DFFARX1 I_7934 (I136950,I2067,I136834,I136990,);
not I_7935 (I136826,I136990);
not I_7936 (I137012,I1900);
nand I_7937 (I137029,I136933,I137012);
DFFARX1 I_7938 (I137029,I2067,I136834,I137055,);
not I_7939 (I137063,I137055);
not I_7940 (I137080,I2020);
nand I_7941 (I137097,I137080,I1884);
and I_7942 (I137114,I136916,I137097);
nor I_7943 (I137131,I137029,I137114);
DFFARX1 I_7944 (I137131,I2067,I136834,I136802,);
DFFARX1 I_7945 (I137114,I2067,I136834,I136823,);
nor I_7946 (I137176,I2020,I1812);
nor I_7947 (I136814,I137029,I137176);
or I_7948 (I137207,I2020,I1812);
nor I_7949 (I137224,I1836,I1948);
DFFARX1 I_7950 (I137224,I2067,I136834,I137250,);
not I_7951 (I137258,I137250);
nor I_7952 (I136820,I137258,I137063);
nand I_7953 (I137289,I137258,I136908);
not I_7954 (I137306,I1836);
nand I_7955 (I137323,I137306,I137012);
nand I_7956 (I137340,I137258,I137323);
nand I_7957 (I136811,I137340,I137289);
nand I_7958 (I136808,I137323,I137207);
not I_7959 (I137412,I2074);
DFFARX1 I_7960 (I80173,I2067,I137412,I137438,);
and I_7961 (I137446,I137438,I80161);
DFFARX1 I_7962 (I137446,I2067,I137412,I137395,);
DFFARX1 I_7963 (I80176,I2067,I137412,I137486,);
not I_7964 (I137494,I80167);
not I_7965 (I137511,I80158);
nand I_7966 (I137528,I137511,I137494);
nor I_7967 (I137383,I137486,I137528);
DFFARX1 I_7968 (I137528,I2067,I137412,I137568,);
not I_7969 (I137404,I137568);
not I_7970 (I137590,I80164);
nand I_7971 (I137607,I137511,I137590);
DFFARX1 I_7972 (I137607,I2067,I137412,I137633,);
not I_7973 (I137641,I137633);
not I_7974 (I137658,I80179);
nand I_7975 (I137675,I137658,I80182);
and I_7976 (I137692,I137494,I137675);
nor I_7977 (I137709,I137607,I137692);
DFFARX1 I_7978 (I137709,I2067,I137412,I137380,);
DFFARX1 I_7979 (I137692,I2067,I137412,I137401,);
nor I_7980 (I137754,I80179,I80158);
nor I_7981 (I137392,I137607,I137754);
or I_7982 (I137785,I80179,I80158);
nor I_7983 (I137802,I80170,I80161);
DFFARX1 I_7984 (I137802,I2067,I137412,I137828,);
not I_7985 (I137836,I137828);
nor I_7986 (I137398,I137836,I137641);
nand I_7987 (I137867,I137836,I137486);
not I_7988 (I137884,I80170);
nand I_7989 (I137901,I137884,I137590);
nand I_7990 (I137918,I137836,I137901);
nand I_7991 (I137389,I137918,I137867);
nand I_7992 (I137386,I137901,I137785);
not I_7993 (I137990,I2074);
DFFARX1 I_7994 (I120386,I2067,I137990,I138016,);
and I_7995 (I138024,I138016,I120380);
DFFARX1 I_7996 (I138024,I2067,I137990,I137973,);
DFFARX1 I_7997 (I120398,I2067,I137990,I138064,);
not I_7998 (I138072,I120389);
not I_7999 (I138089,I120401);
nand I_8000 (I138106,I138089,I138072);
nor I_8001 (I137961,I138064,I138106);
DFFARX1 I_8002 (I138106,I2067,I137990,I138146,);
not I_8003 (I137982,I138146);
not I_8004 (I138168,I120407);
nand I_8005 (I138185,I138089,I138168);
DFFARX1 I_8006 (I138185,I2067,I137990,I138211,);
not I_8007 (I138219,I138211);
not I_8008 (I138236,I120383);
nand I_8009 (I138253,I138236,I120404);
and I_8010 (I138270,I138072,I138253);
nor I_8011 (I138287,I138185,I138270);
DFFARX1 I_8012 (I138287,I2067,I137990,I137958,);
DFFARX1 I_8013 (I138270,I2067,I137990,I137979,);
nor I_8014 (I138332,I120383,I120395);
nor I_8015 (I137970,I138185,I138332);
or I_8016 (I138363,I120383,I120395);
nor I_8017 (I138380,I120380,I120392);
DFFARX1 I_8018 (I138380,I2067,I137990,I138406,);
not I_8019 (I138414,I138406);
nor I_8020 (I137976,I138414,I138219);
nand I_8021 (I138445,I138414,I138064);
not I_8022 (I138462,I120380);
nand I_8023 (I138479,I138462,I138168);
nand I_8024 (I138496,I138414,I138479);
nand I_8025 (I137967,I138496,I138445);
nand I_8026 (I137964,I138479,I138363);
not I_8027 (I138568,I2074);
DFFARX1 I_8028 (I83063,I2067,I138568,I138594,);
and I_8029 (I138602,I138594,I83051);
DFFARX1 I_8030 (I138602,I2067,I138568,I138551,);
DFFARX1 I_8031 (I83066,I2067,I138568,I138642,);
not I_8032 (I138650,I83057);
not I_8033 (I138667,I83048);
nand I_8034 (I138684,I138667,I138650);
nor I_8035 (I138539,I138642,I138684);
DFFARX1 I_8036 (I138684,I2067,I138568,I138724,);
not I_8037 (I138560,I138724);
not I_8038 (I138746,I83054);
nand I_8039 (I138763,I138667,I138746);
DFFARX1 I_8040 (I138763,I2067,I138568,I138789,);
not I_8041 (I138797,I138789);
not I_8042 (I138814,I83069);
nand I_8043 (I138831,I138814,I83072);
and I_8044 (I138848,I138650,I138831);
nor I_8045 (I138865,I138763,I138848);
DFFARX1 I_8046 (I138865,I2067,I138568,I138536,);
DFFARX1 I_8047 (I138848,I2067,I138568,I138557,);
nor I_8048 (I138910,I83069,I83048);
nor I_8049 (I138548,I138763,I138910);
or I_8050 (I138941,I83069,I83048);
nor I_8051 (I138958,I83060,I83051);
DFFARX1 I_8052 (I138958,I2067,I138568,I138984,);
not I_8053 (I138992,I138984);
nor I_8054 (I138554,I138992,I138797);
nand I_8055 (I139023,I138992,I138642);
not I_8056 (I139040,I83060);
nand I_8057 (I139057,I139040,I138746);
nand I_8058 (I139074,I138992,I139057);
nand I_8059 (I138545,I139074,I139023);
nand I_8060 (I138542,I139057,I138941);
not I_8061 (I139146,I2074);
DFFARX1 I_8062 (I70114,I2067,I139146,I139172,);
and I_8063 (I139180,I139172,I70129);
DFFARX1 I_8064 (I139180,I2067,I139146,I139129,);
DFFARX1 I_8065 (I70120,I2067,I139146,I139220,);
not I_8066 (I139228,I70114);
not I_8067 (I139245,I70132);
nand I_8068 (I139262,I139245,I139228);
nor I_8069 (I139117,I139220,I139262);
DFFARX1 I_8070 (I139262,I2067,I139146,I139302,);
not I_8071 (I139138,I139302);
not I_8072 (I139324,I70123);
nand I_8073 (I139341,I139245,I139324);
DFFARX1 I_8074 (I139341,I2067,I139146,I139367,);
not I_8075 (I139375,I139367);
not I_8076 (I139392,I70135);
nand I_8077 (I139409,I139392,I70111);
and I_8078 (I139426,I139228,I139409);
nor I_8079 (I139443,I139341,I139426);
DFFARX1 I_8080 (I139443,I2067,I139146,I139114,);
DFFARX1 I_8081 (I139426,I2067,I139146,I139135,);
nor I_8082 (I139488,I70135,I70111);
nor I_8083 (I139126,I139341,I139488);
or I_8084 (I139519,I70135,I70111);
nor I_8085 (I139536,I70117,I70126);
DFFARX1 I_8086 (I139536,I2067,I139146,I139562,);
not I_8087 (I139570,I139562);
nor I_8088 (I139132,I139570,I139375);
nand I_8089 (I139601,I139570,I139220);
not I_8090 (I139618,I70117);
nand I_8091 (I139635,I139618,I139324);
nand I_8092 (I139652,I139570,I139635);
nand I_8093 (I139123,I139652,I139601);
nand I_8094 (I139120,I139635,I139519);
not I_8095 (I139724,I2074);
DFFARX1 I_8096 (I60761,I2067,I139724,I139750,);
and I_8097 (I139758,I139750,I60776);
DFFARX1 I_8098 (I139758,I2067,I139724,I139707,);
DFFARX1 I_8099 (I60779,I2067,I139724,I139798,);
not I_8100 (I139806,I60773);
not I_8101 (I139823,I60788);
nand I_8102 (I139840,I139823,I139806);
nor I_8103 (I139695,I139798,I139840);
DFFARX1 I_8104 (I139840,I2067,I139724,I139880,);
not I_8105 (I139716,I139880);
not I_8106 (I139902,I60764);
nand I_8107 (I139919,I139823,I139902);
DFFARX1 I_8108 (I139919,I2067,I139724,I139945,);
not I_8109 (I139953,I139945);
not I_8110 (I139970,I60767);
nand I_8111 (I139987,I139970,I60761);
and I_8112 (I140004,I139806,I139987);
nor I_8113 (I140021,I139919,I140004);
DFFARX1 I_8114 (I140021,I2067,I139724,I139692,);
DFFARX1 I_8115 (I140004,I2067,I139724,I139713,);
nor I_8116 (I140066,I60767,I60770);
nor I_8117 (I139704,I139919,I140066);
or I_8118 (I140097,I60767,I60770);
nor I_8119 (I140114,I60785,I60782);
DFFARX1 I_8120 (I140114,I2067,I139724,I140140,);
not I_8121 (I140148,I140140);
nor I_8122 (I139710,I140148,I139953);
nand I_8123 (I140179,I140148,I139798);
not I_8124 (I140196,I60785);
nand I_8125 (I140213,I140196,I139902);
nand I_8126 (I140230,I140148,I140213);
nand I_8127 (I139701,I140230,I140179);
nand I_8128 (I139698,I140213,I140097);
not I_8129 (I140302,I2074);
DFFARX1 I_8130 (I81907,I2067,I140302,I140328,);
and I_8131 (I140336,I140328,I81895);
DFFARX1 I_8132 (I140336,I2067,I140302,I140285,);
DFFARX1 I_8133 (I81910,I2067,I140302,I140376,);
not I_8134 (I140384,I81901);
not I_8135 (I140401,I81892);
nand I_8136 (I140418,I140401,I140384);
nor I_8137 (I140273,I140376,I140418);
DFFARX1 I_8138 (I140418,I2067,I140302,I140458,);
not I_8139 (I140294,I140458);
not I_8140 (I140480,I81898);
nand I_8141 (I140497,I140401,I140480);
DFFARX1 I_8142 (I140497,I2067,I140302,I140523,);
not I_8143 (I140531,I140523);
not I_8144 (I140548,I81913);
nand I_8145 (I140565,I140548,I81916);
and I_8146 (I140582,I140384,I140565);
nor I_8147 (I140599,I140497,I140582);
DFFARX1 I_8148 (I140599,I2067,I140302,I140270,);
DFFARX1 I_8149 (I140582,I2067,I140302,I140291,);
nor I_8150 (I140644,I81913,I81892);
nor I_8151 (I140282,I140497,I140644);
or I_8152 (I140675,I81913,I81892);
nor I_8153 (I140692,I81904,I81895);
DFFARX1 I_8154 (I140692,I2067,I140302,I140718,);
not I_8155 (I140726,I140718);
nor I_8156 (I140288,I140726,I140531);
nand I_8157 (I140757,I140726,I140376);
not I_8158 (I140774,I81904);
nand I_8159 (I140791,I140774,I140480);
nand I_8160 (I140808,I140726,I140791);
nand I_8161 (I140279,I140808,I140757);
nand I_8162 (I140276,I140791,I140675);
not I_8163 (I140880,I2074);
DFFARX1 I_8164 (I43346,I2067,I140880,I140906,);
and I_8165 (I140914,I140906,I43331);
DFFARX1 I_8166 (I140914,I2067,I140880,I140863,);
DFFARX1 I_8167 (I43337,I2067,I140880,I140954,);
not I_8168 (I140962,I43319);
not I_8169 (I140979,I43340);
nand I_8170 (I140996,I140979,I140962);
nor I_8171 (I140851,I140954,I140996);
DFFARX1 I_8172 (I140996,I2067,I140880,I141036,);
not I_8173 (I140872,I141036);
not I_8174 (I141058,I43343);
nand I_8175 (I141075,I140979,I141058);
DFFARX1 I_8176 (I141075,I2067,I140880,I141101,);
not I_8177 (I141109,I141101);
not I_8178 (I141126,I43334);
nand I_8179 (I141143,I141126,I43322);
and I_8180 (I141160,I140962,I141143);
nor I_8181 (I141177,I141075,I141160);
DFFARX1 I_8182 (I141177,I2067,I140880,I140848,);
DFFARX1 I_8183 (I141160,I2067,I140880,I140869,);
nor I_8184 (I141222,I43334,I43328);
nor I_8185 (I140860,I141075,I141222);
or I_8186 (I141253,I43334,I43328);
nor I_8187 (I141270,I43325,I43319);
DFFARX1 I_8188 (I141270,I2067,I140880,I141296,);
not I_8189 (I141304,I141296);
nor I_8190 (I140866,I141304,I141109);
nand I_8191 (I141335,I141304,I140954);
not I_8192 (I141352,I43325);
nand I_8193 (I141369,I141352,I141058);
nand I_8194 (I141386,I141304,I141369);
nand I_8195 (I140857,I141386,I141335);
nand I_8196 (I140854,I141369,I141253);
not I_8197 (I141458,I2074);
DFFARX1 I_8198 (I134000,I2067,I141458,I141484,);
and I_8199 (I141492,I141484,I133997);
DFFARX1 I_8200 (I141492,I2067,I141458,I141441,);
DFFARX1 I_8201 (I134003,I2067,I141458,I141532,);
not I_8202 (I141540,I134006);
not I_8203 (I141557,I134000);
nand I_8204 (I141574,I141557,I141540);
nor I_8205 (I141429,I141532,I141574);
DFFARX1 I_8206 (I141574,I2067,I141458,I141614,);
not I_8207 (I141450,I141614);
not I_8208 (I141636,I134015);
nand I_8209 (I141653,I141557,I141636);
DFFARX1 I_8210 (I141653,I2067,I141458,I141679,);
not I_8211 (I141687,I141679);
not I_8212 (I141704,I134012);
nand I_8213 (I141721,I141704,I134018);
and I_8214 (I141738,I141540,I141721);
nor I_8215 (I141755,I141653,I141738);
DFFARX1 I_8216 (I141755,I2067,I141458,I141426,);
DFFARX1 I_8217 (I141738,I2067,I141458,I141447,);
nor I_8218 (I141800,I134012,I133997);
nor I_8219 (I141438,I141653,I141800);
or I_8220 (I141831,I134012,I133997);
nor I_8221 (I141848,I134009,I134003);
DFFARX1 I_8222 (I141848,I2067,I141458,I141874,);
not I_8223 (I141882,I141874);
nor I_8224 (I141444,I141882,I141687);
nand I_8225 (I141913,I141882,I141532);
not I_8226 (I141930,I134009);
nand I_8227 (I141947,I141930,I141636);
nand I_8228 (I141964,I141882,I141947);
nand I_8229 (I141435,I141964,I141913);
nand I_8230 (I141432,I141947,I141831);
not I_8231 (I142036,I2074);
DFFARX1 I_8232 (I113396,I2067,I142036,I142062,);
and I_8233 (I142070,I142062,I113402);
DFFARX1 I_8234 (I142070,I2067,I142036,I142019,);
DFFARX1 I_8235 (I113408,I2067,I142036,I142110,);
not I_8236 (I142118,I113393);
not I_8237 (I142135,I113393);
nand I_8238 (I142152,I142135,I142118);
nor I_8239 (I142007,I142110,I142152);
DFFARX1 I_8240 (I142152,I2067,I142036,I142192,);
not I_8241 (I142028,I142192);
not I_8242 (I142214,I113411);
nand I_8243 (I142231,I142135,I142214);
DFFARX1 I_8244 (I142231,I2067,I142036,I142257,);
not I_8245 (I142265,I142257);
not I_8246 (I142282,I113405);
nand I_8247 (I142299,I142282,I113396);
and I_8248 (I142316,I142118,I142299);
nor I_8249 (I142333,I142231,I142316);
DFFARX1 I_8250 (I142333,I2067,I142036,I142004,);
DFFARX1 I_8251 (I142316,I2067,I142036,I142025,);
nor I_8252 (I142378,I113405,I113414);
nor I_8253 (I142016,I142231,I142378);
or I_8254 (I142409,I113405,I113414);
nor I_8255 (I142426,I113399,I113399);
DFFARX1 I_8256 (I142426,I2067,I142036,I142452,);
not I_8257 (I142460,I142452);
nor I_8258 (I142022,I142460,I142265);
nand I_8259 (I142491,I142460,I142110);
not I_8260 (I142508,I113399);
nand I_8261 (I142525,I142508,I142214);
nand I_8262 (I142542,I142460,I142525);
nand I_8263 (I142013,I142542,I142491);
nand I_8264 (I142010,I142525,I142409);
not I_8265 (I142614,I2074);
DFFARX1 I_8266 (I114572,I2067,I142614,I142640,);
and I_8267 (I142648,I142640,I114566);
DFFARX1 I_8268 (I142648,I2067,I142614,I142597,);
DFFARX1 I_8269 (I114584,I2067,I142614,I142688,);
not I_8270 (I142696,I114575);
not I_8271 (I142713,I114587);
nand I_8272 (I142730,I142713,I142696);
nor I_8273 (I142585,I142688,I142730);
DFFARX1 I_8274 (I142730,I2067,I142614,I142770,);
not I_8275 (I142606,I142770);
not I_8276 (I142792,I114593);
nand I_8277 (I142809,I142713,I142792);
DFFARX1 I_8278 (I142809,I2067,I142614,I142835,);
not I_8279 (I142843,I142835);
not I_8280 (I142860,I114569);
nand I_8281 (I142877,I142860,I114590);
and I_8282 (I142894,I142696,I142877);
nor I_8283 (I142911,I142809,I142894);
DFFARX1 I_8284 (I142911,I2067,I142614,I142582,);
DFFARX1 I_8285 (I142894,I2067,I142614,I142603,);
nor I_8286 (I142956,I114569,I114581);
nor I_8287 (I142594,I142809,I142956);
or I_8288 (I142987,I114569,I114581);
nor I_8289 (I143004,I114566,I114578);
DFFARX1 I_8290 (I143004,I2067,I142614,I143030,);
not I_8291 (I143038,I143030);
nor I_8292 (I142600,I143038,I142843);
nand I_8293 (I143069,I143038,I142688);
not I_8294 (I143086,I114566);
nand I_8295 (I143103,I143086,I142792);
nand I_8296 (I143120,I143038,I143103);
nand I_8297 (I142591,I143120,I143069);
nand I_8298 (I142588,I143103,I142987);
not I_8299 (I143192,I2074);
DFFARX1 I_8300 (I59673,I2067,I143192,I143218,);
and I_8301 (I143226,I143218,I59688);
DFFARX1 I_8302 (I143226,I2067,I143192,I143175,);
DFFARX1 I_8303 (I59691,I2067,I143192,I143266,);
not I_8304 (I143274,I59685);
not I_8305 (I143291,I59700);
nand I_8306 (I143308,I143291,I143274);
nor I_8307 (I143163,I143266,I143308);
DFFARX1 I_8308 (I143308,I2067,I143192,I143348,);
not I_8309 (I143184,I143348);
not I_8310 (I143370,I59676);
nand I_8311 (I143387,I143291,I143370);
DFFARX1 I_8312 (I143387,I2067,I143192,I143413,);
not I_8313 (I143421,I143413);
not I_8314 (I143438,I59679);
nand I_8315 (I143455,I143438,I59673);
and I_8316 (I143472,I143274,I143455);
nor I_8317 (I143489,I143387,I143472);
DFFARX1 I_8318 (I143489,I2067,I143192,I143160,);
DFFARX1 I_8319 (I143472,I2067,I143192,I143181,);
nor I_8320 (I143534,I59679,I59682);
nor I_8321 (I143172,I143387,I143534);
or I_8322 (I143565,I59679,I59682);
nor I_8323 (I143582,I59697,I59694);
DFFARX1 I_8324 (I143582,I2067,I143192,I143608,);
not I_8325 (I143616,I143608);
nor I_8326 (I143178,I143616,I143421);
nand I_8327 (I143647,I143616,I143266);
not I_8328 (I143664,I59697);
nand I_8329 (I143681,I143664,I143370);
nand I_8330 (I143698,I143616,I143681);
nand I_8331 (I143169,I143698,I143647);
nand I_8332 (I143166,I143681,I143565);
not I_8333 (I143770,I2074);
DFFARX1 I_8334 (I107599,I2067,I143770,I143796,);
and I_8335 (I143804,I143796,I107605);
DFFARX1 I_8336 (I143804,I2067,I143770,I143753,);
DFFARX1 I_8337 (I107611,I2067,I143770,I143844,);
not I_8338 (I143852,I107596);
not I_8339 (I143869,I107596);
nand I_8340 (I143886,I143869,I143852);
nor I_8341 (I143741,I143844,I143886);
DFFARX1 I_8342 (I143886,I2067,I143770,I143926,);
not I_8343 (I143762,I143926);
not I_8344 (I143948,I107614);
nand I_8345 (I143965,I143869,I143948);
DFFARX1 I_8346 (I143965,I2067,I143770,I143991,);
not I_8347 (I143999,I143991);
not I_8348 (I144016,I107608);
nand I_8349 (I144033,I144016,I107599);
and I_8350 (I144050,I143852,I144033);
nor I_8351 (I144067,I143965,I144050);
DFFARX1 I_8352 (I144067,I2067,I143770,I143738,);
DFFARX1 I_8353 (I144050,I2067,I143770,I143759,);
nor I_8354 (I144112,I107608,I107617);
nor I_8355 (I143750,I143965,I144112);
or I_8356 (I144143,I107608,I107617);
nor I_8357 (I144160,I107602,I107602);
DFFARX1 I_8358 (I144160,I2067,I143770,I144186,);
not I_8359 (I144194,I144186);
nor I_8360 (I143756,I144194,I143999);
nand I_8361 (I144225,I144194,I143844);
not I_8362 (I144242,I107602);
nand I_8363 (I144259,I144242,I143948);
nand I_8364 (I144276,I144194,I144259);
nand I_8365 (I143747,I144276,I144225);
nand I_8366 (I143744,I144259,I144143);
not I_8367 (I144348,I2074);
DFFARX1 I_8368 (I130073,I2067,I144348,I144374,);
and I_8369 (I144382,I144374,I130070);
DFFARX1 I_8370 (I144382,I2067,I144348,I144331,);
DFFARX1 I_8371 (I130076,I2067,I144348,I144422,);
not I_8372 (I144430,I130079);
not I_8373 (I144447,I130073);
nand I_8374 (I144464,I144447,I144430);
nor I_8375 (I144319,I144422,I144464);
DFFARX1 I_8376 (I144464,I2067,I144348,I144504,);
not I_8377 (I144340,I144504);
not I_8378 (I144526,I130088);
nand I_8379 (I144543,I144447,I144526);
DFFARX1 I_8380 (I144543,I2067,I144348,I144569,);
not I_8381 (I144577,I144569);
not I_8382 (I144594,I130085);
nand I_8383 (I144611,I144594,I130091);
and I_8384 (I144628,I144430,I144611);
nor I_8385 (I144645,I144543,I144628);
DFFARX1 I_8386 (I144645,I2067,I144348,I144316,);
DFFARX1 I_8387 (I144628,I2067,I144348,I144337,);
nor I_8388 (I144690,I130085,I130070);
nor I_8389 (I144328,I144543,I144690);
or I_8390 (I144721,I130085,I130070);
nor I_8391 (I144738,I130082,I130076);
DFFARX1 I_8392 (I144738,I2067,I144348,I144764,);
not I_8393 (I144772,I144764);
nor I_8394 (I144334,I144772,I144577);
nand I_8395 (I144803,I144772,I144422);
not I_8396 (I144820,I130082);
nand I_8397 (I144837,I144820,I144526);
nand I_8398 (I144854,I144772,I144837);
nand I_8399 (I144325,I144854,I144803);
nand I_8400 (I144322,I144837,I144721);
not I_8401 (I144926,I2074);
DFFARX1 I_8402 (I9064,I2067,I144926,I144952,);
and I_8403 (I144960,I144952,I9067);
DFFARX1 I_8404 (I144960,I2067,I144926,I144909,);
DFFARX1 I_8405 (I9067,I2067,I144926,I145000,);
not I_8406 (I145008,I9070);
not I_8407 (I145025,I9085);
nand I_8408 (I145042,I145025,I145008);
nor I_8409 (I144897,I145000,I145042);
DFFARX1 I_8410 (I145042,I2067,I144926,I145082,);
not I_8411 (I144918,I145082);
not I_8412 (I145104,I9079);
nand I_8413 (I145121,I145025,I145104);
DFFARX1 I_8414 (I145121,I2067,I144926,I145147,);
not I_8415 (I145155,I145147);
not I_8416 (I145172,I9082);
nand I_8417 (I145189,I145172,I9064);
and I_8418 (I145206,I145008,I145189);
nor I_8419 (I145223,I145121,I145206);
DFFARX1 I_8420 (I145223,I2067,I144926,I144894,);
DFFARX1 I_8421 (I145206,I2067,I144926,I144915,);
nor I_8422 (I145268,I9082,I9076);
nor I_8423 (I144906,I145121,I145268);
or I_8424 (I145299,I9082,I9076);
nor I_8425 (I145316,I9073,I9088);
DFFARX1 I_8426 (I145316,I2067,I144926,I145342,);
not I_8427 (I145350,I145342);
nor I_8428 (I144912,I145350,I145155);
nand I_8429 (I145381,I145350,I145000);
not I_8430 (I145398,I9073);
nand I_8431 (I145415,I145398,I145104);
nand I_8432 (I145432,I145350,I145415);
nand I_8433 (I144903,I145432,I145381);
nand I_8434 (I144900,I145415,I145299);
not I_8435 (I145504,I2074);
DFFARX1 I_8436 (I1620,I2067,I145504,I145530,);
and I_8437 (I145538,I145530,I1676);
DFFARX1 I_8438 (I145538,I2067,I145504,I145487,);
DFFARX1 I_8439 (I1852,I2067,I145504,I145578,);
not I_8440 (I145586,I1444);
not I_8441 (I145603,I1844);
nand I_8442 (I145620,I145603,I145586);
nor I_8443 (I145475,I145578,I145620);
DFFARX1 I_8444 (I145620,I2067,I145504,I145660,);
not I_8445 (I145496,I145660);
not I_8446 (I145682,I1372);
nand I_8447 (I145699,I145603,I145682);
DFFARX1 I_8448 (I145699,I2067,I145504,I145725,);
not I_8449 (I145733,I145725);
not I_8450 (I145750,I1596);
nand I_8451 (I145767,I145750,I1556);
and I_8452 (I145784,I145586,I145767);
nor I_8453 (I145801,I145699,I145784);
DFFARX1 I_8454 (I145801,I2067,I145504,I145472,);
DFFARX1 I_8455 (I145784,I2067,I145504,I145493,);
nor I_8456 (I145846,I1596,I1572);
nor I_8457 (I145484,I145699,I145846);
or I_8458 (I145877,I1596,I1572);
nor I_8459 (I145894,I1716,I2012);
DFFARX1 I_8460 (I145894,I2067,I145504,I145920,);
not I_8461 (I145928,I145920);
nor I_8462 (I145490,I145928,I145733);
nand I_8463 (I145959,I145928,I145578);
not I_8464 (I145976,I1716);
nand I_8465 (I145993,I145976,I145682);
nand I_8466 (I146010,I145928,I145993);
nand I_8467 (I145481,I146010,I145959);
nand I_8468 (I145478,I145993,I145877);
not I_8469 (I146082,I2074);
DFFARX1 I_8470 (I8010,I2067,I146082,I146108,);
and I_8471 (I146116,I146108,I8013);
DFFARX1 I_8472 (I146116,I2067,I146082,I146065,);
DFFARX1 I_8473 (I8013,I2067,I146082,I146156,);
not I_8474 (I146164,I8016);
not I_8475 (I146181,I8031);
nand I_8476 (I146198,I146181,I146164);
nor I_8477 (I146053,I146156,I146198);
DFFARX1 I_8478 (I146198,I2067,I146082,I146238,);
not I_8479 (I146074,I146238);
not I_8480 (I146260,I8025);
nand I_8481 (I146277,I146181,I146260);
DFFARX1 I_8482 (I146277,I2067,I146082,I146303,);
not I_8483 (I146311,I146303);
not I_8484 (I146328,I8028);
nand I_8485 (I146345,I146328,I8010);
and I_8486 (I146362,I146164,I146345);
nor I_8487 (I146379,I146277,I146362);
DFFARX1 I_8488 (I146379,I2067,I146082,I146050,);
DFFARX1 I_8489 (I146362,I2067,I146082,I146071,);
nor I_8490 (I146424,I8028,I8022);
nor I_8491 (I146062,I146277,I146424);
or I_8492 (I146455,I8028,I8022);
nor I_8493 (I146472,I8019,I8034);
DFFARX1 I_8494 (I146472,I2067,I146082,I146498,);
not I_8495 (I146506,I146498);
nor I_8496 (I146068,I146506,I146311);
nand I_8497 (I146537,I146506,I146156);
not I_8498 (I146554,I8019);
nand I_8499 (I146571,I146554,I146260);
nand I_8500 (I146588,I146506,I146571);
nand I_8501 (I146059,I146588,I146537);
nand I_8502 (I146056,I146571,I146455);
not I_8503 (I146660,I2074);
DFFARX1 I_8504 (I2687,I2067,I146660,I146686,);
and I_8505 (I146694,I146686,I2693);
DFFARX1 I_8506 (I146694,I2067,I146660,I146643,);
DFFARX1 I_8507 (I2672,I2067,I146660,I146734,);
not I_8508 (I146742,I2678);
not I_8509 (I146759,I2684);
nand I_8510 (I146776,I146759,I146742);
nor I_8511 (I146631,I146734,I146776);
DFFARX1 I_8512 (I146776,I2067,I146660,I146816,);
not I_8513 (I146652,I146816);
not I_8514 (I146838,I2675);
nand I_8515 (I146855,I146759,I146838);
DFFARX1 I_8516 (I146855,I2067,I146660,I146881,);
not I_8517 (I146889,I146881);
not I_8518 (I146906,I2690);
nand I_8519 (I146923,I146906,I2675);
and I_8520 (I146940,I146742,I146923);
nor I_8521 (I146957,I146855,I146940);
DFFARX1 I_8522 (I146957,I2067,I146660,I146628,);
DFFARX1 I_8523 (I146940,I2067,I146660,I146649,);
nor I_8524 (I147002,I2690,I2678);
nor I_8525 (I146640,I146855,I147002);
or I_8526 (I147033,I2690,I2678);
nor I_8527 (I147050,I2681,I2672);
DFFARX1 I_8528 (I147050,I2067,I146660,I147076,);
not I_8529 (I147084,I147076);
nor I_8530 (I146646,I147084,I146889);
nand I_8531 (I147115,I147084,I146734);
not I_8532 (I147132,I2681);
nand I_8533 (I147149,I147132,I146838);
nand I_8534 (I147166,I147084,I147149);
nand I_8535 (I146637,I147166,I147115);
nand I_8536 (I146634,I147149,I147033);
not I_8537 (I147238,I2074);
DFFARX1 I_8538 (I21209,I2067,I147238,I147264,);
and I_8539 (I147272,I147264,I21185);
DFFARX1 I_8540 (I147272,I2067,I147238,I147221,);
DFFARX1 I_8541 (I21203,I2067,I147238,I147312,);
not I_8542 (I147320,I21191);
not I_8543 (I147337,I21188);
nand I_8544 (I147354,I147337,I147320);
nor I_8545 (I147209,I147312,I147354);
DFFARX1 I_8546 (I147354,I2067,I147238,I147394,);
not I_8547 (I147230,I147394);
not I_8548 (I147416,I21197);
nand I_8549 (I147433,I147337,I147416);
DFFARX1 I_8550 (I147433,I2067,I147238,I147459,);
not I_8551 (I147467,I147459);
not I_8552 (I147484,I21188);
nand I_8553 (I147501,I147484,I21206);
and I_8554 (I147518,I147320,I147501);
nor I_8555 (I147535,I147433,I147518);
DFFARX1 I_8556 (I147535,I2067,I147238,I147206,);
DFFARX1 I_8557 (I147518,I2067,I147238,I147227,);
nor I_8558 (I147580,I21188,I21200);
nor I_8559 (I147218,I147433,I147580);
or I_8560 (I147611,I21188,I21200);
nor I_8561 (I147628,I21194,I21185);
DFFARX1 I_8562 (I147628,I2067,I147238,I147654,);
not I_8563 (I147662,I147654);
nor I_8564 (I147224,I147662,I147467);
nand I_8565 (I147693,I147662,I147312);
not I_8566 (I147710,I21194);
nand I_8567 (I147727,I147710,I147416);
nand I_8568 (I147744,I147662,I147727);
nand I_8569 (I147215,I147744,I147693);
nand I_8570 (I147212,I147727,I147611);
not I_8571 (I147816,I2074);
DFFARX1 I_8572 (I66201,I2067,I147816,I147842,);
and I_8573 (I147850,I147842,I66216);
DFFARX1 I_8574 (I147850,I2067,I147816,I147799,);
DFFARX1 I_8575 (I66219,I2067,I147816,I147890,);
not I_8576 (I147898,I66213);
not I_8577 (I147915,I66228);
nand I_8578 (I147932,I147915,I147898);
nor I_8579 (I147787,I147890,I147932);
DFFARX1 I_8580 (I147932,I2067,I147816,I147972,);
not I_8581 (I147808,I147972);
not I_8582 (I147994,I66204);
nand I_8583 (I148011,I147915,I147994);
DFFARX1 I_8584 (I148011,I2067,I147816,I148037,);
not I_8585 (I148045,I148037);
not I_8586 (I148062,I66207);
nand I_8587 (I148079,I148062,I66201);
and I_8588 (I148096,I147898,I148079);
nor I_8589 (I148113,I148011,I148096);
DFFARX1 I_8590 (I148113,I2067,I147816,I147784,);
DFFARX1 I_8591 (I148096,I2067,I147816,I147805,);
nor I_8592 (I148158,I66207,I66210);
nor I_8593 (I147796,I148011,I148158);
or I_8594 (I148189,I66207,I66210);
nor I_8595 (I148206,I66225,I66222);
DFFARX1 I_8596 (I148206,I2067,I147816,I148232,);
not I_8597 (I148240,I148232);
nor I_8598 (I147802,I148240,I148045);
nand I_8599 (I148271,I148240,I147890);
not I_8600 (I148288,I66225);
nand I_8601 (I148305,I148288,I147994);
nand I_8602 (I148322,I148240,I148305);
nand I_8603 (I147793,I148322,I148271);
nand I_8604 (I147790,I148305,I148189);
not I_8605 (I148394,I2074);
DFFARX1 I_8606 (I45981,I2067,I148394,I148420,);
and I_8607 (I148428,I148420,I45966);
DFFARX1 I_8608 (I148428,I2067,I148394,I148377,);
DFFARX1 I_8609 (I45972,I2067,I148394,I148468,);
not I_8610 (I148476,I45954);
not I_8611 (I148493,I45975);
nand I_8612 (I148510,I148493,I148476);
nor I_8613 (I148365,I148468,I148510);
DFFARX1 I_8614 (I148510,I2067,I148394,I148550,);
not I_8615 (I148386,I148550);
not I_8616 (I148572,I45978);
nand I_8617 (I148589,I148493,I148572);
DFFARX1 I_8618 (I148589,I2067,I148394,I148615,);
not I_8619 (I148623,I148615);
not I_8620 (I148640,I45969);
nand I_8621 (I148657,I148640,I45957);
and I_8622 (I148674,I148476,I148657);
nor I_8623 (I148691,I148589,I148674);
DFFARX1 I_8624 (I148691,I2067,I148394,I148362,);
DFFARX1 I_8625 (I148674,I2067,I148394,I148383,);
nor I_8626 (I148736,I45969,I45963);
nor I_8627 (I148374,I148589,I148736);
or I_8628 (I148767,I45969,I45963);
nor I_8629 (I148784,I45960,I45954);
DFFARX1 I_8630 (I148784,I2067,I148394,I148810,);
not I_8631 (I148818,I148810);
nor I_8632 (I148380,I148818,I148623);
nand I_8633 (I148849,I148818,I148468);
not I_8634 (I148866,I45960);
nand I_8635 (I148883,I148866,I148572);
nand I_8636 (I148900,I148818,I148883);
nand I_8637 (I148371,I148900,I148849);
nand I_8638 (I148368,I148883,I148767);
not I_8639 (I148972,I2074);
DFFARX1 I_8640 (I85953,I2067,I148972,I148998,);
and I_8641 (I149006,I148998,I85941);
DFFARX1 I_8642 (I149006,I2067,I148972,I148955,);
DFFARX1 I_8643 (I85956,I2067,I148972,I149046,);
not I_8644 (I149054,I85947);
not I_8645 (I149071,I85938);
nand I_8646 (I149088,I149071,I149054);
nor I_8647 (I148943,I149046,I149088);
DFFARX1 I_8648 (I149088,I2067,I148972,I149128,);
not I_8649 (I148964,I149128);
not I_8650 (I149150,I85944);
nand I_8651 (I149167,I149071,I149150);
DFFARX1 I_8652 (I149167,I2067,I148972,I149193,);
not I_8653 (I149201,I149193);
not I_8654 (I149218,I85959);
nand I_8655 (I149235,I149218,I85962);
and I_8656 (I149252,I149054,I149235);
nor I_8657 (I149269,I149167,I149252);
DFFARX1 I_8658 (I149269,I2067,I148972,I148940,);
DFFARX1 I_8659 (I149252,I2067,I148972,I148961,);
nor I_8660 (I149314,I85959,I85938);
nor I_8661 (I148952,I149167,I149314);
or I_8662 (I149345,I85959,I85938);
nor I_8663 (I149362,I85950,I85941);
DFFARX1 I_8664 (I149362,I2067,I148972,I149388,);
not I_8665 (I149396,I149388);
nor I_8666 (I148958,I149396,I149201);
nand I_8667 (I149427,I149396,I149046);
not I_8668 (I149444,I85950);
nand I_8669 (I149461,I149444,I149150);
nand I_8670 (I149478,I149396,I149461);
nand I_8671 (I148949,I149478,I149427);
nand I_8672 (I148946,I149461,I149345);
not I_8673 (I149550,I2074);
DFFARX1 I_8674 (I126846,I2067,I149550,I149576,);
and I_8675 (I149584,I149576,I126840);
DFFARX1 I_8676 (I149584,I2067,I149550,I149533,);
DFFARX1 I_8677 (I126858,I2067,I149550,I149624,);
not I_8678 (I149632,I126849);
not I_8679 (I149649,I126861);
nand I_8680 (I149666,I149649,I149632);
nor I_8681 (I149521,I149624,I149666);
DFFARX1 I_8682 (I149666,I2067,I149550,I149706,);
not I_8683 (I149542,I149706);
not I_8684 (I149728,I126867);
nand I_8685 (I149745,I149649,I149728);
DFFARX1 I_8686 (I149745,I2067,I149550,I149771,);
not I_8687 (I149779,I149771);
not I_8688 (I149796,I126843);
nand I_8689 (I149813,I149796,I126864);
and I_8690 (I149830,I149632,I149813);
nor I_8691 (I149847,I149745,I149830);
DFFARX1 I_8692 (I149847,I2067,I149550,I149518,);
DFFARX1 I_8693 (I149830,I2067,I149550,I149539,);
nor I_8694 (I149892,I126843,I126855);
nor I_8695 (I149530,I149745,I149892);
or I_8696 (I149923,I126843,I126855);
nor I_8697 (I149940,I126840,I126852);
DFFARX1 I_8698 (I149940,I2067,I149550,I149966,);
not I_8699 (I149974,I149966);
nor I_8700 (I149536,I149974,I149779);
nand I_8701 (I150005,I149974,I149624);
not I_8702 (I150022,I126840);
nand I_8703 (I150039,I150022,I149728);
nand I_8704 (I150056,I149974,I150039);
nand I_8705 (I149527,I150056,I150005);
nand I_8706 (I149524,I150039,I149923);
not I_8707 (I150128,I2074);
DFFARX1 I_8708 (I32218,I2067,I150128,I150154,);
and I_8709 (I150162,I150154,I32221);
DFFARX1 I_8710 (I150162,I2067,I150128,I150111,);
DFFARX1 I_8711 (I32221,I2067,I150128,I150202,);
not I_8712 (I150210,I32236);
not I_8713 (I150227,I32242);
nand I_8714 (I150244,I150227,I150210);
nor I_8715 (I150099,I150202,I150244);
DFFARX1 I_8716 (I150244,I2067,I150128,I150284,);
not I_8717 (I150120,I150284);
not I_8718 (I150306,I32230);
nand I_8719 (I150323,I150227,I150306);
DFFARX1 I_8720 (I150323,I2067,I150128,I150349,);
not I_8721 (I150357,I150349);
not I_8722 (I150374,I32227);
nand I_8723 (I150391,I150374,I32224);
and I_8724 (I150408,I150210,I150391);
nor I_8725 (I150425,I150323,I150408);
DFFARX1 I_8726 (I150425,I2067,I150128,I150096,);
DFFARX1 I_8727 (I150408,I2067,I150128,I150117,);
nor I_8728 (I150470,I32227,I32218);
nor I_8729 (I150108,I150323,I150470);
or I_8730 (I150501,I32227,I32218);
nor I_8731 (I150518,I32233,I32239);
DFFARX1 I_8732 (I150518,I2067,I150128,I150544,);
not I_8733 (I150552,I150544);
nor I_8734 (I150114,I150552,I150357);
nand I_8735 (I150583,I150552,I150202);
not I_8736 (I150600,I32233);
nand I_8737 (I150617,I150600,I150306);
nand I_8738 (I150634,I150552,I150617);
nand I_8739 (I150105,I150634,I150583);
nand I_8740 (I150102,I150617,I150501);
not I_8741 (I150706,I2074);
DFFARX1 I_8742 (I170506,I2067,I150706,I150732,);
and I_8743 (I150740,I150732,I170488);
DFFARX1 I_8744 (I150740,I2067,I150706,I150689,);
DFFARX1 I_8745 (I170479,I2067,I150706,I150780,);
not I_8746 (I150788,I170494);
not I_8747 (I150805,I170482);
nand I_8748 (I150822,I150805,I150788);
nor I_8749 (I150677,I150780,I150822);
DFFARX1 I_8750 (I150822,I2067,I150706,I150862,);
not I_8751 (I150698,I150862);
not I_8752 (I150884,I170491);
nand I_8753 (I150901,I150805,I150884);
DFFARX1 I_8754 (I150901,I2067,I150706,I150927,);
not I_8755 (I150935,I150927);
not I_8756 (I150952,I170500);
nand I_8757 (I150969,I150952,I170479);
and I_8758 (I150986,I150788,I150969);
nor I_8759 (I151003,I150901,I150986);
DFFARX1 I_8760 (I151003,I2067,I150706,I150674,);
DFFARX1 I_8761 (I150986,I2067,I150706,I150695,);
nor I_8762 (I151048,I170500,I170503);
nor I_8763 (I150686,I150901,I151048);
or I_8764 (I151079,I170500,I170503);
nor I_8765 (I151096,I170497,I170485);
DFFARX1 I_8766 (I151096,I2067,I150706,I151122,);
not I_8767 (I151130,I151122);
nor I_8768 (I150692,I151130,I150935);
nand I_8769 (I151161,I151130,I150780);
not I_8770 (I151178,I170497);
nand I_8771 (I151195,I151178,I150884);
nand I_8772 (I151212,I151130,I151195);
nand I_8773 (I150683,I151212,I151161);
nand I_8774 (I150680,I151195,I151079);
not I_8775 (I151284,I2074);
DFFARX1 I_8776 (I73684,I2067,I151284,I151310,);
and I_8777 (I151318,I151310,I73699);
DFFARX1 I_8778 (I151318,I2067,I151284,I151267,);
DFFARX1 I_8779 (I73690,I2067,I151284,I151358,);
not I_8780 (I151366,I73684);
not I_8781 (I151383,I73702);
nand I_8782 (I151400,I151383,I151366);
nor I_8783 (I151255,I151358,I151400);
DFFARX1 I_8784 (I151400,I2067,I151284,I151440,);
not I_8785 (I151276,I151440);
not I_8786 (I151462,I73693);
nand I_8787 (I151479,I151383,I151462);
DFFARX1 I_8788 (I151479,I2067,I151284,I151505,);
not I_8789 (I151513,I151505);
not I_8790 (I151530,I73705);
nand I_8791 (I151547,I151530,I73681);
and I_8792 (I151564,I151366,I151547);
nor I_8793 (I151581,I151479,I151564);
DFFARX1 I_8794 (I151581,I2067,I151284,I151252,);
DFFARX1 I_8795 (I151564,I2067,I151284,I151273,);
nor I_8796 (I151626,I73705,I73681);
nor I_8797 (I151264,I151479,I151626);
or I_8798 (I151657,I73705,I73681);
nor I_8799 (I151674,I73687,I73696);
DFFARX1 I_8800 (I151674,I2067,I151284,I151700,);
not I_8801 (I151708,I151700);
nor I_8802 (I151270,I151708,I151513);
nand I_8803 (I151739,I151708,I151358);
not I_8804 (I151756,I73687);
nand I_8805 (I151773,I151756,I151462);
nand I_8806 (I151790,I151708,I151773);
nand I_8807 (I151261,I151790,I151739);
nand I_8808 (I151258,I151773,I151657);
not I_8809 (I151862,I2074);
DFFARX1 I_8810 (I38168,I2067,I151862,I151888,);
and I_8811 (I151896,I151888,I38171);
DFFARX1 I_8812 (I151896,I2067,I151862,I151845,);
DFFARX1 I_8813 (I38171,I2067,I151862,I151936,);
not I_8814 (I151944,I38186);
not I_8815 (I151961,I38192);
nand I_8816 (I151978,I151961,I151944);
nor I_8817 (I151833,I151936,I151978);
DFFARX1 I_8818 (I151978,I2067,I151862,I152018,);
not I_8819 (I151854,I152018);
not I_8820 (I152040,I38180);
nand I_8821 (I152057,I151961,I152040);
DFFARX1 I_8822 (I152057,I2067,I151862,I152083,);
not I_8823 (I152091,I152083);
not I_8824 (I152108,I38177);
nand I_8825 (I152125,I152108,I38174);
and I_8826 (I152142,I151944,I152125);
nor I_8827 (I152159,I152057,I152142);
DFFARX1 I_8828 (I152159,I2067,I151862,I151830,);
DFFARX1 I_8829 (I152142,I2067,I151862,I151851,);
nor I_8830 (I152204,I38177,I38168);
nor I_8831 (I151842,I152057,I152204);
or I_8832 (I152235,I38177,I38168);
nor I_8833 (I152252,I38183,I38189);
DFFARX1 I_8834 (I152252,I2067,I151862,I152278,);
not I_8835 (I152286,I152278);
nor I_8836 (I151848,I152286,I152091);
nand I_8837 (I152317,I152286,I151936);
not I_8838 (I152334,I38183);
nand I_8839 (I152351,I152334,I152040);
nand I_8840 (I152368,I152286,I152351);
nand I_8841 (I151839,I152368,I152317);
nand I_8842 (I151836,I152351,I152235);
not I_8843 (I152440,I2074);
DFFARX1 I_8844 (I158447,I2067,I152440,I152466,);
and I_8845 (I152474,I152466,I158441);
DFFARX1 I_8846 (I152474,I2067,I152440,I152423,);
DFFARX1 I_8847 (I158426,I2067,I152440,I152514,);
not I_8848 (I152522,I158432);
not I_8849 (I152539,I158444);
nand I_8850 (I152556,I152539,I152522);
nor I_8851 (I152411,I152514,I152556);
DFFARX1 I_8852 (I152556,I2067,I152440,I152596,);
not I_8853 (I152432,I152596);
not I_8854 (I152618,I158426);
nand I_8855 (I152635,I152539,I152618);
DFFARX1 I_8856 (I152635,I2067,I152440,I152661,);
not I_8857 (I152669,I152661);
not I_8858 (I152686,I158450);
nand I_8859 (I152703,I152686,I158438);
and I_8860 (I152720,I152522,I152703);
nor I_8861 (I152737,I152635,I152720);
DFFARX1 I_8862 (I152737,I2067,I152440,I152408,);
DFFARX1 I_8863 (I152720,I2067,I152440,I152429,);
nor I_8864 (I152782,I158450,I158429);
nor I_8865 (I152420,I152635,I152782);
or I_8866 (I152813,I158450,I158429);
nor I_8867 (I152830,I158435,I158429);
DFFARX1 I_8868 (I152830,I2067,I152440,I152856,);
not I_8869 (I152864,I152856);
nor I_8870 (I152426,I152864,I152669);
nand I_8871 (I152895,I152864,I152514);
not I_8872 (I152912,I158435);
nand I_8873 (I152929,I152912,I152618);
nand I_8874 (I152946,I152864,I152929);
nand I_8875 (I152417,I152946,I152895);
nand I_8876 (I152414,I152929,I152813);
not I_8877 (I153018,I2074);
DFFARX1 I_8878 (I108129,I2067,I153018,I153044,);
nand I_8879 (I153052,I153044,I108123);
DFFARX1 I_8880 (I108126,I2067,I153018,I153078,);
DFFARX1 I_8881 (I153078,I2067,I153018,I153095,);
not I_8882 (I153010,I153095);
not I_8883 (I153117,I108132);
nor I_8884 (I153134,I108132,I108126);
not I_8885 (I153151,I108135);
nand I_8886 (I153168,I153117,I153151);
nor I_8887 (I153185,I108135,I108132);
and I_8888 (I152989,I153185,I153052);
not I_8889 (I153216,I108144);
nand I_8890 (I153233,I153216,I108138);
nor I_8891 (I153250,I108144,I108141);
not I_8892 (I153267,I153250);
nand I_8893 (I152992,I153134,I153267);
DFFARX1 I_8894 (I153250,I2067,I153018,I153007,);
nor I_8895 (I153312,I108123,I108135);
nor I_8896 (I153329,I153312,I108126);
and I_8897 (I153346,I153329,I153233);
DFFARX1 I_8898 (I153346,I2067,I153018,I153004,);
nor I_8899 (I153001,I153312,I153168);
or I_8900 (I152998,I153250,I153312);
nor I_8901 (I153405,I108123,I108129);
DFFARX1 I_8902 (I153405,I2067,I153018,I153431,);
not I_8903 (I153439,I153431);
nand I_8904 (I153456,I153439,I153117);
nor I_8905 (I153473,I153456,I108126);
DFFARX1 I_8906 (I153473,I2067,I153018,I152986,);
nor I_8907 (I153504,I153439,I153168);
nor I_8908 (I152995,I153312,I153504);
not I_8909 (I153562,I2074);
DFFARX1 I_8910 (I109183,I2067,I153562,I153588,);
nand I_8911 (I153596,I153588,I109177);
DFFARX1 I_8912 (I109180,I2067,I153562,I153622,);
DFFARX1 I_8913 (I153622,I2067,I153562,I153639,);
not I_8914 (I153554,I153639);
not I_8915 (I153661,I109186);
nor I_8916 (I153678,I109186,I109180);
not I_8917 (I153695,I109189);
nand I_8918 (I153712,I153661,I153695);
nor I_8919 (I153729,I109189,I109186);
and I_8920 (I153533,I153729,I153596);
not I_8921 (I153760,I109198);
nand I_8922 (I153777,I153760,I109192);
nor I_8923 (I153794,I109198,I109195);
not I_8924 (I153811,I153794);
nand I_8925 (I153536,I153678,I153811);
DFFARX1 I_8926 (I153794,I2067,I153562,I153551,);
nor I_8927 (I153856,I109177,I109189);
nor I_8928 (I153873,I153856,I109180);
and I_8929 (I153890,I153873,I153777);
DFFARX1 I_8930 (I153890,I2067,I153562,I153548,);
nor I_8931 (I153545,I153856,I153712);
or I_8932 (I153542,I153794,I153856);
nor I_8933 (I153949,I109177,I109183);
DFFARX1 I_8934 (I153949,I2067,I153562,I153975,);
not I_8935 (I153983,I153975);
nand I_8936 (I154000,I153983,I153661);
nor I_8937 (I154017,I154000,I109180);
DFFARX1 I_8938 (I154017,I2067,I153562,I153530,);
nor I_8939 (I154048,I153983,I153712);
nor I_8940 (I153539,I153856,I154048);
not I_8941 (I154106,I2074);
DFFARX1 I_8942 (I16463,I2067,I154106,I154132,);
nand I_8943 (I154140,I154132,I16445);
DFFARX1 I_8944 (I16442,I2067,I154106,I154166,);
DFFARX1 I_8945 (I154166,I2067,I154106,I154183,);
not I_8946 (I154098,I154183);
not I_8947 (I154205,I16460);
nor I_8948 (I154222,I16460,I16454);
not I_8949 (I154239,I16442);
nand I_8950 (I154256,I154205,I154239);
nor I_8951 (I154273,I16442,I16460);
and I_8952 (I154077,I154273,I154140);
not I_8953 (I154304,I16451);
nand I_8954 (I154321,I154304,I16457);
nor I_8955 (I154338,I16451,I16445);
not I_8956 (I154355,I154338);
nand I_8957 (I154080,I154222,I154355);
DFFARX1 I_8958 (I154338,I2067,I154106,I154095,);
nor I_8959 (I154400,I16448,I16442);
nor I_8960 (I154417,I154400,I16454);
and I_8961 (I154434,I154417,I154321);
DFFARX1 I_8962 (I154434,I2067,I154106,I154092,);
nor I_8963 (I154089,I154400,I154256);
or I_8964 (I154086,I154338,I154400);
nor I_8965 (I154493,I16448,I16466);
DFFARX1 I_8966 (I154493,I2067,I154106,I154519,);
not I_8967 (I154527,I154519);
nand I_8968 (I154544,I154527,I154205);
nor I_8969 (I154561,I154544,I16454);
DFFARX1 I_8970 (I154561,I2067,I154106,I154074,);
nor I_8971 (I154592,I154527,I154256);
nor I_8972 (I154083,I154400,I154592);
not I_8973 (I154650,I2074);
DFFARX1 I_8974 (I54398,I2067,I154650,I154676,);
nand I_8975 (I154684,I154676,I54401);
DFFARX1 I_8976 (I54395,I2067,I154650,I154710,);
DFFARX1 I_8977 (I154710,I2067,I154650,I154727,);
not I_8978 (I154642,I154727);
not I_8979 (I154749,I54404);
nor I_8980 (I154766,I54404,I54389);
not I_8981 (I154783,I54413);
nand I_8982 (I154800,I154749,I154783);
nor I_8983 (I154817,I54413,I54404);
and I_8984 (I154621,I154817,I154684);
not I_8985 (I154848,I54392);
nand I_8986 (I154865,I154848,I54410);
nor I_8987 (I154882,I54392,I54386);
not I_8988 (I154899,I154882);
nand I_8989 (I154624,I154766,I154899);
DFFARX1 I_8990 (I154882,I2067,I154650,I154639,);
nor I_8991 (I154944,I54407,I54413);
nor I_8992 (I154961,I154944,I54389);
and I_8993 (I154978,I154961,I154865);
DFFARX1 I_8994 (I154978,I2067,I154650,I154636,);
nor I_8995 (I154633,I154944,I154800);
or I_8996 (I154630,I154882,I154944);
nor I_8997 (I155037,I54407,I54386);
DFFARX1 I_8998 (I155037,I2067,I154650,I155063,);
not I_8999 (I155071,I155063);
nand I_9000 (I155088,I155071,I154749);
nor I_9001 (I155105,I155088,I54389);
DFFARX1 I_9002 (I155105,I2067,I154650,I154618,);
nor I_9003 (I155136,I155071,I154800);
nor I_9004 (I154627,I154944,I155136);
not I_9005 (I155194,I2074);
DFFARX1 I_9006 (I178241,I2067,I155194,I155220,);
nand I_9007 (I155228,I155220,I178226);
DFFARX1 I_9008 (I178220,I2067,I155194,I155254,);
DFFARX1 I_9009 (I155254,I2067,I155194,I155271,);
not I_9010 (I155186,I155271);
not I_9011 (I155293,I178214);
nor I_9012 (I155310,I178214,I178235);
not I_9013 (I155327,I178223);
nand I_9014 (I155344,I155293,I155327);
nor I_9015 (I155361,I178223,I178214);
and I_9016 (I155165,I155361,I155228);
not I_9017 (I155392,I178232);
nand I_9018 (I155409,I155392,I178238);
nor I_9019 (I155426,I178232,I178229);
not I_9020 (I155443,I155426);
nand I_9021 (I155168,I155310,I155443);
DFFARX1 I_9022 (I155426,I2067,I155194,I155183,);
nor I_9023 (I155488,I178217,I178223);
nor I_9024 (I155505,I155488,I178235);
and I_9025 (I155522,I155505,I155409);
DFFARX1 I_9026 (I155522,I2067,I155194,I155180,);
nor I_9027 (I155177,I155488,I155344);
or I_9028 (I155174,I155426,I155488);
nor I_9029 (I155581,I178217,I178214);
DFFARX1 I_9030 (I155581,I2067,I155194,I155607,);
not I_9031 (I155615,I155607);
nand I_9032 (I155632,I155615,I155293);
nor I_9033 (I155649,I155632,I178235);
DFFARX1 I_9034 (I155649,I2067,I155194,I155162,);
nor I_9035 (I155680,I155615,I155344);
nor I_9036 (I155171,I155488,I155680);
not I_9037 (I155738,I2074);
DFFARX1 I_9038 (I35202,I2067,I155738,I155764,);
nand I_9039 (I155772,I155764,I35217);
DFFARX1 I_9040 (I35214,I2067,I155738,I155798,);
DFFARX1 I_9041 (I155798,I2067,I155738,I155815,);
not I_9042 (I155730,I155815);
not I_9043 (I155837,I35193);
nor I_9044 (I155854,I35193,I35199);
not I_9045 (I155871,I35205);
nand I_9046 (I155888,I155837,I155871);
nor I_9047 (I155905,I35205,I35193);
and I_9048 (I155709,I155905,I155772);
not I_9049 (I155936,I35211);
nand I_9050 (I155953,I155936,I35193);
nor I_9051 (I155970,I35211,I35196);
not I_9052 (I155987,I155970);
nand I_9053 (I155712,I155854,I155987);
DFFARX1 I_9054 (I155970,I2067,I155738,I155727,);
nor I_9055 (I156032,I35196,I35205);
nor I_9056 (I156049,I156032,I35199);
and I_9057 (I156066,I156049,I155953);
DFFARX1 I_9058 (I156066,I2067,I155738,I155724,);
nor I_9059 (I155721,I156032,I155888);
or I_9060 (I155718,I155970,I156032);
nor I_9061 (I156125,I35196,I35208);
DFFARX1 I_9062 (I156125,I2067,I155738,I156151,);
not I_9063 (I156159,I156151);
nand I_9064 (I156176,I156159,I155837);
nor I_9065 (I156193,I156176,I35199);
DFFARX1 I_9066 (I156193,I2067,I155738,I155706,);
nor I_9067 (I156224,I156159,I155888);
nor I_9068 (I155715,I156032,I156224);
not I_9069 (I156282,I2074);
DFFARX1 I_9070 (I10666,I2067,I156282,I156308,);
nand I_9071 (I156316,I156308,I10648);
DFFARX1 I_9072 (I10645,I2067,I156282,I156342,);
DFFARX1 I_9073 (I156342,I2067,I156282,I156359,);
not I_9074 (I156274,I156359);
not I_9075 (I156381,I10663);
nor I_9076 (I156398,I10663,I10657);
not I_9077 (I156415,I10645);
nand I_9078 (I156432,I156381,I156415);
nor I_9079 (I156449,I10645,I10663);
and I_9080 (I156253,I156449,I156316);
not I_9081 (I156480,I10654);
nand I_9082 (I156497,I156480,I10660);
nor I_9083 (I156514,I10654,I10648);
not I_9084 (I156531,I156514);
nand I_9085 (I156256,I156398,I156531);
DFFARX1 I_9086 (I156514,I2067,I156282,I156271,);
nor I_9087 (I156576,I10651,I10645);
nor I_9088 (I156593,I156576,I10657);
and I_9089 (I156610,I156593,I156497);
DFFARX1 I_9090 (I156610,I2067,I156282,I156268,);
nor I_9091 (I156265,I156576,I156432);
or I_9092 (I156262,I156514,I156576);
nor I_9093 (I156669,I10651,I10669);
DFFARX1 I_9094 (I156669,I2067,I156282,I156695,);
not I_9095 (I156703,I156695);
nand I_9096 (I156720,I156703,I156381);
nor I_9097 (I156737,I156720,I10657);
DFFARX1 I_9098 (I156737,I2067,I156282,I156250,);
nor I_9099 (I156768,I156703,I156432);
nor I_9100 (I156259,I156576,I156768);
not I_9101 (I156826,I2074);
DFFARX1 I_9102 (I11193,I2067,I156826,I156852,);
nand I_9103 (I156860,I156852,I11175);
DFFARX1 I_9104 (I11172,I2067,I156826,I156886,);
DFFARX1 I_9105 (I156886,I2067,I156826,I156903,);
not I_9106 (I156818,I156903);
not I_9107 (I156925,I11190);
nor I_9108 (I156942,I11190,I11184);
not I_9109 (I156959,I11172);
nand I_9110 (I156976,I156925,I156959);
nor I_9111 (I156993,I11172,I11190);
and I_9112 (I156797,I156993,I156860);
not I_9113 (I157024,I11181);
nand I_9114 (I157041,I157024,I11187);
nor I_9115 (I157058,I11181,I11175);
not I_9116 (I157075,I157058);
nand I_9117 (I156800,I156942,I157075);
DFFARX1 I_9118 (I157058,I2067,I156826,I156815,);
nor I_9119 (I157120,I11178,I11172);
nor I_9120 (I157137,I157120,I11184);
and I_9121 (I157154,I157137,I157041);
DFFARX1 I_9122 (I157154,I2067,I156826,I156812,);
nor I_9123 (I156809,I157120,I156976);
or I_9124 (I156806,I157058,I157120);
nor I_9125 (I157213,I11178,I11196);
DFFARX1 I_9126 (I157213,I2067,I156826,I157239,);
not I_9127 (I157247,I157239);
nand I_9128 (I157264,I157247,I156925);
nor I_9129 (I157281,I157264,I11184);
DFFARX1 I_9130 (I157281,I2067,I156826,I156794,);
nor I_9131 (I157312,I157247,I156976);
nor I_9132 (I156803,I157120,I157312);
not I_9133 (I157370,I2074);
DFFARX1 I_9134 (I30442,I2067,I157370,I157396,);
nand I_9135 (I157404,I157396,I30457);
DFFARX1 I_9136 (I30454,I2067,I157370,I157430,);
DFFARX1 I_9137 (I157430,I2067,I157370,I157447,);
not I_9138 (I157362,I157447);
not I_9139 (I157469,I30433);
nor I_9140 (I157486,I30433,I30439);
not I_9141 (I157503,I30445);
nand I_9142 (I157520,I157469,I157503);
nor I_9143 (I157537,I30445,I30433);
and I_9144 (I157341,I157537,I157404);
not I_9145 (I157568,I30451);
nand I_9146 (I157585,I157568,I30433);
nor I_9147 (I157602,I30451,I30436);
not I_9148 (I157619,I157602);
nand I_9149 (I157344,I157486,I157619);
DFFARX1 I_9150 (I157602,I2067,I157370,I157359,);
nor I_9151 (I157664,I30436,I30445);
nor I_9152 (I157681,I157664,I30439);
and I_9153 (I157698,I157681,I157585);
DFFARX1 I_9154 (I157698,I2067,I157370,I157356,);
nor I_9155 (I157353,I157664,I157520);
or I_9156 (I157350,I157602,I157664);
nor I_9157 (I157757,I30436,I30448);
DFFARX1 I_9158 (I157757,I2067,I157370,I157783,);
not I_9159 (I157791,I157783);
nand I_9160 (I157808,I157791,I157469);
nor I_9161 (I157825,I157808,I30439);
DFFARX1 I_9162 (I157825,I2067,I157370,I157338,);
nor I_9163 (I157856,I157791,I157520);
nor I_9164 (I157347,I157664,I157856);
not I_9165 (I157914,I2074);
DFFARX1 I_9166 (I46493,I2067,I157914,I157940,);
nand I_9167 (I157948,I157940,I46496);
DFFARX1 I_9168 (I46490,I2067,I157914,I157974,);
DFFARX1 I_9169 (I157974,I2067,I157914,I157991,);
not I_9170 (I157906,I157991);
not I_9171 (I158013,I46499);
nor I_9172 (I158030,I46499,I46484);
not I_9173 (I158047,I46508);
nand I_9174 (I158064,I158013,I158047);
nor I_9175 (I158081,I46508,I46499);
and I_9176 (I157885,I158081,I157948);
not I_9177 (I158112,I46487);
nand I_9178 (I158129,I158112,I46505);
nor I_9179 (I158146,I46487,I46481);
not I_9180 (I158163,I158146);
nand I_9181 (I157888,I158030,I158163);
DFFARX1 I_9182 (I158146,I2067,I157914,I157903,);
nor I_9183 (I158208,I46502,I46508);
nor I_9184 (I158225,I158208,I46484);
and I_9185 (I158242,I158225,I158129);
DFFARX1 I_9186 (I158242,I2067,I157914,I157900,);
nor I_9187 (I157897,I158208,I158064);
or I_9188 (I157894,I158146,I158208);
nor I_9189 (I158301,I46502,I46481);
DFFARX1 I_9190 (I158301,I2067,I157914,I158327,);
not I_9191 (I158335,I158327);
nand I_9192 (I158352,I158335,I158013);
nor I_9193 (I158369,I158352,I46484);
DFFARX1 I_9194 (I158369,I2067,I157914,I157882,);
nor I_9195 (I158400,I158335,I158064);
nor I_9196 (I157891,I158208,I158400);
not I_9197 (I158458,I2074);
DFFARX1 I_9198 (I55979,I2067,I158458,I158484,);
nand I_9199 (I158492,I158484,I55982);
DFFARX1 I_9200 (I55976,I2067,I158458,I158518,);
DFFARX1 I_9201 (I158518,I2067,I158458,I158535,);
not I_9202 (I158450,I158535);
not I_9203 (I158557,I55985);
nor I_9204 (I158574,I55985,I55970);
not I_9205 (I158591,I55994);
nand I_9206 (I158608,I158557,I158591);
nor I_9207 (I158625,I55994,I55985);
and I_9208 (I158429,I158625,I158492);
not I_9209 (I158656,I55973);
nand I_9210 (I158673,I158656,I55991);
nor I_9211 (I158690,I55973,I55967);
not I_9212 (I158707,I158690);
nand I_9213 (I158432,I158574,I158707);
DFFARX1 I_9214 (I158690,I2067,I158458,I158447,);
nor I_9215 (I158752,I55988,I55994);
nor I_9216 (I158769,I158752,I55970);
and I_9217 (I158786,I158769,I158673);
DFFARX1 I_9218 (I158786,I2067,I158458,I158444,);
nor I_9219 (I158441,I158752,I158608);
or I_9220 (I158438,I158690,I158752);
nor I_9221 (I158845,I55988,I55967);
DFFARX1 I_9222 (I158845,I2067,I158458,I158871,);
not I_9223 (I158879,I158871);
nand I_9224 (I158896,I158879,I158557);
nor I_9225 (I158913,I158896,I55970);
DFFARX1 I_9226 (I158913,I2067,I158458,I158426,);
nor I_9227 (I158944,I158879,I158608);
nor I_9228 (I158435,I158752,I158944);
not I_9229 (I159002,I2074);
DFFARX1 I_9230 (I56506,I2067,I159002,I159028,);
nand I_9231 (I159036,I159028,I56509);
DFFARX1 I_9232 (I56503,I2067,I159002,I159062,);
DFFARX1 I_9233 (I159062,I2067,I159002,I159079,);
not I_9234 (I158994,I159079);
not I_9235 (I159101,I56512);
nor I_9236 (I159118,I56512,I56497);
not I_9237 (I159135,I56521);
nand I_9238 (I159152,I159101,I159135);
nor I_9239 (I159169,I56521,I56512);
and I_9240 (I158973,I159169,I159036);
not I_9241 (I159200,I56500);
nand I_9242 (I159217,I159200,I56518);
nor I_9243 (I159234,I56500,I56494);
not I_9244 (I159251,I159234);
nand I_9245 (I158976,I159118,I159251);
DFFARX1 I_9246 (I159234,I2067,I159002,I158991,);
nor I_9247 (I159296,I56515,I56521);
nor I_9248 (I159313,I159296,I56497);
and I_9249 (I159330,I159313,I159217);
DFFARX1 I_9250 (I159330,I2067,I159002,I158988,);
nor I_9251 (I158985,I159296,I159152);
or I_9252 (I158982,I159234,I159296);
nor I_9253 (I159389,I56515,I56494);
DFFARX1 I_9254 (I159389,I2067,I159002,I159415,);
not I_9255 (I159423,I159415);
nand I_9256 (I159440,I159423,I159101);
nor I_9257 (I159457,I159440,I56497);
DFFARX1 I_9258 (I159457,I2067,I159002,I158970,);
nor I_9259 (I159488,I159423,I159152);
nor I_9260 (I158979,I159296,I159488);
not I_9261 (I159546,I2074);
DFFARX1 I_9262 (I29252,I2067,I159546,I159572,);
nand I_9263 (I159580,I159572,I29267);
DFFARX1 I_9264 (I29264,I2067,I159546,I159606,);
DFFARX1 I_9265 (I159606,I2067,I159546,I159623,);
not I_9266 (I159538,I159623);
not I_9267 (I159645,I29243);
nor I_9268 (I159662,I29243,I29249);
not I_9269 (I159679,I29255);
nand I_9270 (I159696,I159645,I159679);
nor I_9271 (I159713,I29255,I29243);
and I_9272 (I159517,I159713,I159580);
not I_9273 (I159744,I29261);
nand I_9274 (I159761,I159744,I29243);
nor I_9275 (I159778,I29261,I29246);
not I_9276 (I159795,I159778);
nand I_9277 (I159520,I159662,I159795);
DFFARX1 I_9278 (I159778,I2067,I159546,I159535,);
nor I_9279 (I159840,I29246,I29255);
nor I_9280 (I159857,I159840,I29249);
and I_9281 (I159874,I159857,I159761);
DFFARX1 I_9282 (I159874,I2067,I159546,I159532,);
nor I_9283 (I159529,I159840,I159696);
or I_9284 (I159526,I159778,I159840);
nor I_9285 (I159933,I29246,I29258);
DFFARX1 I_9286 (I159933,I2067,I159546,I159959,);
not I_9287 (I159967,I159959);
nand I_9288 (I159984,I159967,I159645);
nor I_9289 (I160001,I159984,I29249);
DFFARX1 I_9290 (I160001,I2067,I159546,I159514,);
nor I_9291 (I160032,I159967,I159696);
nor I_9292 (I159523,I159840,I160032);
not I_9293 (I160090,I2074);
DFFARX1 I_9294 (I174076,I2067,I160090,I160116,);
nand I_9295 (I160124,I160116,I174061);
DFFARX1 I_9296 (I174055,I2067,I160090,I160150,);
DFFARX1 I_9297 (I160150,I2067,I160090,I160167,);
not I_9298 (I160082,I160167);
not I_9299 (I160189,I174049);
nor I_9300 (I160206,I174049,I174070);
not I_9301 (I160223,I174058);
nand I_9302 (I160240,I160189,I160223);
nor I_9303 (I160257,I174058,I174049);
and I_9304 (I160061,I160257,I160124);
not I_9305 (I160288,I174067);
nand I_9306 (I160305,I160288,I174073);
nor I_9307 (I160322,I174067,I174064);
not I_9308 (I160339,I160322);
nand I_9309 (I160064,I160206,I160339);
DFFARX1 I_9310 (I160322,I2067,I160090,I160079,);
nor I_9311 (I160384,I174052,I174058);
nor I_9312 (I160401,I160384,I174070);
and I_9313 (I160418,I160401,I160305);
DFFARX1 I_9314 (I160418,I2067,I160090,I160076,);
nor I_9315 (I160073,I160384,I160240);
or I_9316 (I160070,I160322,I160384);
nor I_9317 (I160477,I174052,I174049);
DFFARX1 I_9318 (I160477,I2067,I160090,I160503,);
not I_9319 (I160511,I160503);
nand I_9320 (I160528,I160511,I160189);
nor I_9321 (I160545,I160528,I174070);
DFFARX1 I_9322 (I160545,I2067,I160090,I160058,);
nor I_9323 (I160576,I160511,I160240);
nor I_9324 (I160067,I160384,I160576);
not I_9325 (I160634,I2074);
DFFARX1 I_9326 (I151270,I2067,I160634,I160660,);
nand I_9327 (I160668,I160660,I151255);
not I_9328 (I160685,I160668);
DFFARX1 I_9329 (I151258,I2067,I160634,I160711,);
not I_9330 (I160719,I160711);
not I_9331 (I160736,I151273);
or I_9332 (I160753,I151276,I151273);
nor I_9333 (I160770,I151276,I151273);
or I_9334 (I160787,I151252,I151276);
DFFARX1 I_9335 (I160787,I2067,I160634,I160626,);
not I_9336 (I160818,I151264);
nand I_9337 (I160835,I160818,I151267);
nand I_9338 (I160852,I160736,I160835);
and I_9339 (I160605,I160719,I160852);
nor I_9340 (I160883,I151264,I151261);
and I_9341 (I160900,I160719,I160883);
nor I_9342 (I160611,I160685,I160900);
DFFARX1 I_9343 (I160883,I2067,I160634,I160940,);
not I_9344 (I160948,I160940);
nor I_9345 (I160620,I160719,I160948);
or I_9346 (I160979,I160787,I151252);
nor I_9347 (I160996,I151252,I151252);
nand I_9348 (I161013,I160852,I160996);
nand I_9349 (I161030,I160979,I161013);
DFFARX1 I_9350 (I161030,I2067,I160634,I160623,);
nor I_9351 (I161061,I160996,I160753);
DFFARX1 I_9352 (I161061,I2067,I160634,I160602,);
nor I_9353 (I161092,I151252,I151255);
DFFARX1 I_9354 (I161092,I2067,I160634,I161118,);
DFFARX1 I_9355 (I161118,I2067,I160634,I160617,);
not I_9356 (I161140,I161118);
nand I_9357 (I160614,I161140,I160668);
nand I_9358 (I160608,I161140,I160770);
not I_9359 (I161212,I2074);
DFFARX1 I_9360 (I96342,I2067,I161212,I161238,);
nand I_9361 (I161246,I161238,I96345);
not I_9362 (I161263,I161246);
DFFARX1 I_9363 (I96357,I2067,I161212,I161289,);
not I_9364 (I161297,I161289);
not I_9365 (I161314,I96342);
or I_9366 (I161331,I96351,I96342);
nor I_9367 (I161348,I96351,I96342);
or I_9368 (I161365,I96360,I96351);
DFFARX1 I_9369 (I161365,I2067,I161212,I161204,);
not I_9370 (I161396,I96363);
nand I_9371 (I161413,I161396,I96345);
nand I_9372 (I161430,I161314,I161413);
and I_9373 (I161183,I161297,I161430);
nor I_9374 (I161461,I96363,I96348);
and I_9375 (I161478,I161297,I161461);
nor I_9376 (I161189,I161263,I161478);
DFFARX1 I_9377 (I161461,I2067,I161212,I161518,);
not I_9378 (I161526,I161518);
nor I_9379 (I161198,I161297,I161526);
or I_9380 (I161557,I161365,I96354);
nor I_9381 (I161574,I96354,I96360);
nand I_9382 (I161591,I161430,I161574);
nand I_9383 (I161608,I161557,I161591);
DFFARX1 I_9384 (I161608,I2067,I161212,I161201,);
nor I_9385 (I161639,I161574,I161331);
DFFARX1 I_9386 (I161639,I2067,I161212,I161180,);
nor I_9387 (I161670,I96354,I96366);
DFFARX1 I_9388 (I161670,I2067,I161212,I161696,);
DFFARX1 I_9389 (I161696,I2067,I161212,I161195,);
not I_9390 (I161718,I161696);
nand I_9391 (I161192,I161718,I161246);
nand I_9392 (I161186,I161718,I161348);
not I_9393 (I161790,I2074);
DFFARX1 I_9394 (I95764,I2067,I161790,I161816,);
nand I_9395 (I161824,I161816,I95767);
not I_9396 (I161841,I161824);
DFFARX1 I_9397 (I95779,I2067,I161790,I161867,);
not I_9398 (I161875,I161867);
not I_9399 (I161892,I95764);
or I_9400 (I161909,I95773,I95764);
nor I_9401 (I161926,I95773,I95764);
or I_9402 (I161943,I95782,I95773);
DFFARX1 I_9403 (I161943,I2067,I161790,I161782,);
not I_9404 (I161974,I95785);
nand I_9405 (I161991,I161974,I95767);
nand I_9406 (I162008,I161892,I161991);
and I_9407 (I161761,I161875,I162008);
nor I_9408 (I162039,I95785,I95770);
and I_9409 (I162056,I161875,I162039);
nor I_9410 (I161767,I161841,I162056);
DFFARX1 I_9411 (I162039,I2067,I161790,I162096,);
not I_9412 (I162104,I162096);
nor I_9413 (I161776,I161875,I162104);
or I_9414 (I162135,I161943,I95776);
nor I_9415 (I162152,I95776,I95782);
nand I_9416 (I162169,I162008,I162152);
nand I_9417 (I162186,I162135,I162169);
DFFARX1 I_9418 (I162186,I2067,I161790,I161779,);
nor I_9419 (I162217,I162152,I161909);
DFFARX1 I_9420 (I162217,I2067,I161790,I161758,);
nor I_9421 (I162248,I95776,I95788);
DFFARX1 I_9422 (I162248,I2067,I161790,I162274,);
DFFARX1 I_9423 (I162274,I2067,I161790,I161773,);
not I_9424 (I162296,I162274);
nand I_9425 (I161770,I162296,I161824);
nand I_9426 (I161764,I162296,I161926);
not I_9427 (I162368,I2074);
DFFARX1 I_9428 (I88250,I2067,I162368,I162394,);
nand I_9429 (I162402,I162394,I88253);
not I_9430 (I162419,I162402);
DFFARX1 I_9431 (I88265,I2067,I162368,I162445,);
not I_9432 (I162453,I162445);
not I_9433 (I162470,I88250);
or I_9434 (I162487,I88259,I88250);
nor I_9435 (I162504,I88259,I88250);
or I_9436 (I162521,I88268,I88259);
DFFARX1 I_9437 (I162521,I2067,I162368,I162360,);
not I_9438 (I162552,I88271);
nand I_9439 (I162569,I162552,I88253);
nand I_9440 (I162586,I162470,I162569);
and I_9441 (I162339,I162453,I162586);
nor I_9442 (I162617,I88271,I88256);
and I_9443 (I162634,I162453,I162617);
nor I_9444 (I162345,I162419,I162634);
DFFARX1 I_9445 (I162617,I2067,I162368,I162674,);
not I_9446 (I162682,I162674);
nor I_9447 (I162354,I162453,I162682);
or I_9448 (I162713,I162521,I88262);
nor I_9449 (I162730,I88262,I88268);
nand I_9450 (I162747,I162586,I162730);
nand I_9451 (I162764,I162713,I162747);
DFFARX1 I_9452 (I162764,I2067,I162368,I162357,);
nor I_9453 (I162795,I162730,I162487);
DFFARX1 I_9454 (I162795,I2067,I162368,I162336,);
nor I_9455 (I162826,I88262,I88274);
DFFARX1 I_9456 (I162826,I2067,I162368,I162852,);
DFFARX1 I_9457 (I162852,I2067,I162368,I162351,);
not I_9458 (I162874,I162852);
nand I_9459 (I162348,I162874,I162402);
nand I_9460 (I162342,I162874,I162504);
not I_9461 (I162946,I2074);
DFFARX1 I_9462 (I131201,I2067,I162946,I162972,);
nand I_9463 (I162980,I162972,I131198);
not I_9464 (I162997,I162980);
DFFARX1 I_9465 (I131198,I2067,I162946,I163023,);
not I_9466 (I163031,I163023);
not I_9467 (I163048,I131195);
or I_9468 (I163065,I131204,I131195);
nor I_9469 (I163082,I131204,I131195);
or I_9470 (I163099,I131207,I131204);
DFFARX1 I_9471 (I163099,I2067,I162946,I162938,);
not I_9472 (I163130,I131195);
nand I_9473 (I163147,I163130,I131192);
nand I_9474 (I163164,I163048,I163147);
and I_9475 (I162917,I163031,I163164);
nor I_9476 (I163195,I131195,I131210);
and I_9477 (I163212,I163031,I163195);
nor I_9478 (I162923,I162997,I163212);
DFFARX1 I_9479 (I163195,I2067,I162946,I163252,);
not I_9480 (I163260,I163252);
nor I_9481 (I162932,I163031,I163260);
or I_9482 (I163291,I163099,I131213);
nor I_9483 (I163308,I131213,I131207);
nand I_9484 (I163325,I163164,I163308);
nand I_9485 (I163342,I163291,I163325);
DFFARX1 I_9486 (I163342,I2067,I162946,I162935,);
nor I_9487 (I163373,I163308,I163065);
DFFARX1 I_9488 (I163373,I2067,I162946,I162914,);
nor I_9489 (I163404,I131213,I131192);
DFFARX1 I_9490 (I163404,I2067,I162946,I163430,);
DFFARX1 I_9491 (I163430,I2067,I162946,I162929,);
not I_9492 (I163452,I163430);
nand I_9493 (I162926,I163452,I162980);
nand I_9494 (I162920,I163452,I163082);
not I_9495 (I163524,I2074);
DFFARX1 I_9496 (I93452,I2067,I163524,I163550,);
nand I_9497 (I163558,I163550,I93455);
not I_9498 (I163575,I163558);
DFFARX1 I_9499 (I93467,I2067,I163524,I163601,);
not I_9500 (I163609,I163601);
not I_9501 (I163626,I93452);
or I_9502 (I163643,I93461,I93452);
nor I_9503 (I163660,I93461,I93452);
or I_9504 (I163677,I93470,I93461);
DFFARX1 I_9505 (I163677,I2067,I163524,I163516,);
not I_9506 (I163708,I93473);
nand I_9507 (I163725,I163708,I93455);
nand I_9508 (I163742,I163626,I163725);
and I_9509 (I163495,I163609,I163742);
nor I_9510 (I163773,I93473,I93458);
and I_9511 (I163790,I163609,I163773);
nor I_9512 (I163501,I163575,I163790);
DFFARX1 I_9513 (I163773,I2067,I163524,I163830,);
not I_9514 (I163838,I163830);
nor I_9515 (I163510,I163609,I163838);
or I_9516 (I163869,I163677,I93464);
nor I_9517 (I163886,I93464,I93470);
nand I_9518 (I163903,I163742,I163886);
nand I_9519 (I163920,I163869,I163903);
DFFARX1 I_9520 (I163920,I2067,I163524,I163513,);
nor I_9521 (I163951,I163886,I163643);
DFFARX1 I_9522 (I163951,I2067,I163524,I163492,);
nor I_9523 (I163982,I93464,I93476);
DFFARX1 I_9524 (I163982,I2067,I163524,I164008,);
DFFARX1 I_9525 (I164008,I2067,I163524,I163507,);
not I_9526 (I164030,I164008);
nand I_9527 (I163504,I164030,I163558);
nand I_9528 (I163498,I164030,I163660);
not I_9529 (I164102,I2074);
DFFARX1 I_9530 (I49649,I2067,I164102,I164128,);
nand I_9531 (I164136,I164128,I49670);
not I_9532 (I164153,I164136);
DFFARX1 I_9533 (I49664,I2067,I164102,I164179,);
not I_9534 (I164187,I164179);
not I_9535 (I164204,I49652);
or I_9536 (I164221,I49667,I49652);
nor I_9537 (I164238,I49667,I49652);
or I_9538 (I164255,I49658,I49667);
DFFARX1 I_9539 (I164255,I2067,I164102,I164094,);
not I_9540 (I164286,I49646);
nand I_9541 (I164303,I164286,I49643);
nand I_9542 (I164320,I164204,I164303);
and I_9543 (I164073,I164187,I164320);
nor I_9544 (I164351,I49646,I49655);
and I_9545 (I164368,I164187,I164351);
nor I_9546 (I164079,I164153,I164368);
DFFARX1 I_9547 (I164351,I2067,I164102,I164408,);
not I_9548 (I164416,I164408);
nor I_9549 (I164088,I164187,I164416);
or I_9550 (I164447,I164255,I49661);
nor I_9551 (I164464,I49661,I49658);
nand I_9552 (I164481,I164320,I164464);
nand I_9553 (I164498,I164447,I164481);
DFFARX1 I_9554 (I164498,I2067,I164102,I164091,);
nor I_9555 (I164529,I164464,I164221);
DFFARX1 I_9556 (I164529,I2067,I164102,I164070,);
nor I_9557 (I164560,I49661,I49643);
DFFARX1 I_9558 (I164560,I2067,I164102,I164586,);
DFFARX1 I_9559 (I164586,I2067,I164102,I164085,);
not I_9560 (I164608,I164586);
nand I_9561 (I164082,I164608,I164136);
nand I_9562 (I164076,I164608,I164238);
not I_9563 (I164680,I2074);
DFFARX1 I_9564 (I103856,I2067,I164680,I164706,);
nand I_9565 (I164714,I164706,I103859);
not I_9566 (I164731,I164714);
DFFARX1 I_9567 (I103871,I2067,I164680,I164757,);
not I_9568 (I164765,I164757);
not I_9569 (I164782,I103856);
or I_9570 (I164799,I103865,I103856);
nor I_9571 (I164816,I103865,I103856);
or I_9572 (I164833,I103874,I103865);
DFFARX1 I_9573 (I164833,I2067,I164680,I164672,);
not I_9574 (I164864,I103877);
nand I_9575 (I164881,I164864,I103859);
nand I_9576 (I164898,I164782,I164881);
and I_9577 (I164651,I164765,I164898);
nor I_9578 (I164929,I103877,I103862);
and I_9579 (I164946,I164765,I164929);
nor I_9580 (I164657,I164731,I164946);
DFFARX1 I_9581 (I164929,I2067,I164680,I164986,);
not I_9582 (I164994,I164986);
nor I_9583 (I164666,I164765,I164994);
or I_9584 (I165025,I164833,I103868);
nor I_9585 (I165042,I103868,I103874);
nand I_9586 (I165059,I164898,I165042);
nand I_9587 (I165076,I165025,I165059);
DFFARX1 I_9588 (I165076,I2067,I164680,I164669,);
nor I_9589 (I165107,I165042,I164799);
DFFARX1 I_9590 (I165107,I2067,I164680,I164648,);
nor I_9591 (I165138,I103868,I103880);
DFFARX1 I_9592 (I165138,I2067,I164680,I165164,);
DFFARX1 I_9593 (I165164,I2067,I164680,I164663,);
not I_9594 (I165186,I165164);
nand I_9595 (I164660,I165186,I164714);
nand I_9596 (I164654,I165186,I164816);
not I_9597 (I165258,I2074);
DFFARX1 I_9598 (I154633,I2067,I165258,I165284,);
nand I_9599 (I165292,I165284,I154642);
not I_9600 (I165309,I165292);
DFFARX1 I_9601 (I154618,I2067,I165258,I165335,);
not I_9602 (I165343,I165335);
not I_9603 (I165360,I154621);
or I_9604 (I165377,I154618,I154621);
nor I_9605 (I165394,I154618,I154621);
or I_9606 (I165411,I154636,I154618);
DFFARX1 I_9607 (I165411,I2067,I165258,I165250,);
not I_9608 (I165442,I154624);
nand I_9609 (I165459,I165442,I154639);
nand I_9610 (I165476,I165360,I165459);
and I_9611 (I165229,I165343,I165476);
nor I_9612 (I165507,I154624,I154627);
and I_9613 (I165524,I165343,I165507);
nor I_9614 (I165235,I165309,I165524);
DFFARX1 I_9615 (I165507,I2067,I165258,I165564,);
not I_9616 (I165572,I165564);
nor I_9617 (I165244,I165343,I165572);
or I_9618 (I165603,I165411,I154630);
nor I_9619 (I165620,I154630,I154636);
nand I_9620 (I165637,I165476,I165620);
nand I_9621 (I165654,I165603,I165637);
DFFARX1 I_9622 (I165654,I2067,I165258,I165247,);
nor I_9623 (I165685,I165620,I165377);
DFFARX1 I_9624 (I165685,I2067,I165258,I165226,);
nor I_9625 (I165716,I154630,I154621);
DFFARX1 I_9626 (I165716,I2067,I165258,I165742,);
DFFARX1 I_9627 (I165742,I2067,I165258,I165241,);
not I_9628 (I165764,I165742);
nand I_9629 (I165238,I165764,I165292);
nand I_9630 (I165232,I165764,I165394);
not I_9631 (I165836,I2074);
DFFARX1 I_9632 (I98654,I2067,I165836,I165862,);
nand I_9633 (I165870,I165862,I98657);
not I_9634 (I165887,I165870);
DFFARX1 I_9635 (I98669,I2067,I165836,I165913,);
not I_9636 (I165921,I165913);
not I_9637 (I165938,I98654);
or I_9638 (I165955,I98663,I98654);
nor I_9639 (I165972,I98663,I98654);
or I_9640 (I165989,I98672,I98663);
DFFARX1 I_9641 (I165989,I2067,I165836,I165828,);
not I_9642 (I166020,I98675);
nand I_9643 (I166037,I166020,I98657);
nand I_9644 (I166054,I165938,I166037);
and I_9645 (I165807,I165921,I166054);
nor I_9646 (I166085,I98675,I98660);
and I_9647 (I166102,I165921,I166085);
nor I_9648 (I165813,I165887,I166102);
DFFARX1 I_9649 (I166085,I2067,I165836,I166142,);
not I_9650 (I166150,I166142);
nor I_9651 (I165822,I165921,I166150);
or I_9652 (I166181,I165989,I98666);
nor I_9653 (I166198,I98666,I98672);
nand I_9654 (I166215,I166054,I166198);
nand I_9655 (I166232,I166181,I166215);
DFFARX1 I_9656 (I166232,I2067,I165836,I165825,);
nor I_9657 (I166263,I166198,I165955);
DFFARX1 I_9658 (I166263,I2067,I165836,I165804,);
nor I_9659 (I166294,I98666,I98678);
DFFARX1 I_9660 (I166294,I2067,I165836,I166320,);
DFFARX1 I_9661 (I166320,I2067,I165836,I165819,);
not I_9662 (I166342,I166320);
nand I_9663 (I165816,I166342,I165870);
nand I_9664 (I165810,I166342,I165972);
not I_9665 (I166417,I2074);
DFFARX1 I_9666 (I18047,I2067,I166417,I166443,);
nand I_9667 (I166451,I166443,I18038);
not I_9668 (I166468,I166451);
DFFARX1 I_9669 (I18026,I2067,I166417,I166494,);
not I_9670 (I166502,I166494);
nor I_9671 (I166519,I18029,I18026);
not I_9672 (I166536,I166519);
DFFARX1 I_9673 (I166536,I2067,I166417,I166403,);
or I_9674 (I166567,I18023,I18029);
DFFARX1 I_9675 (I166567,I2067,I166417,I166406,);
not I_9676 (I166598,I18032);
nor I_9677 (I166615,I166598,I18023);
nor I_9678 (I166632,I166615,I18026);
nor I_9679 (I166649,I18023,I18035);
nor I_9680 (I166666,I166502,I166649);
nor I_9681 (I166391,I166468,I166666);
not I_9682 (I166697,I166649);
nand I_9683 (I166394,I166697,I166451);
nand I_9684 (I166388,I166697,I166519);
nor I_9685 (I166385,I166649,I166632);
nor I_9686 (I166756,I18041,I18023);
not I_9687 (I166773,I166756);
DFFARX1 I_9688 (I166756,I2067,I166417,I166799,);
not I_9689 (I166409,I166799);
nor I_9690 (I166821,I18041,I18044);
DFFARX1 I_9691 (I166821,I2067,I166417,I166847,);
and I_9692 (I166855,I166847,I18029);
nor I_9693 (I166872,I166855,I166773);
DFFARX1 I_9694 (I166872,I2067,I166417,I166400,);
nor I_9695 (I166903,I166847,I166632);
DFFARX1 I_9696 (I166903,I2067,I166417,I166382,);
nor I_9697 (I166397,I166847,I166536);
not I_9698 (I166978,I2074);
DFFARX1 I_9699 (I71908,I2067,I166978,I167004,);
nand I_9700 (I167012,I167004,I71899);
not I_9701 (I167029,I167012);
DFFARX1 I_9702 (I71899,I2067,I166978,I167055,);
not I_9703 (I167063,I167055);
nor I_9704 (I167080,I71896,I71917);
not I_9705 (I167097,I167080);
DFFARX1 I_9706 (I167097,I2067,I166978,I166964,);
or I_9707 (I167128,I71911,I71896);
DFFARX1 I_9708 (I167128,I2067,I166978,I166967,);
not I_9709 (I167159,I71902);
nor I_9710 (I167176,I167159,I71896);
nor I_9711 (I167193,I167176,I71917);
nor I_9712 (I167210,I71896,I71905);
nor I_9713 (I167227,I167063,I167210);
nor I_9714 (I166952,I167029,I167227);
not I_9715 (I167258,I167210);
nand I_9716 (I166955,I167258,I167012);
nand I_9717 (I166949,I167258,I167080);
nor I_9718 (I166946,I167210,I167193);
nor I_9719 (I167317,I71920,I71911);
not I_9720 (I167334,I167317);
DFFARX1 I_9721 (I167317,I2067,I166978,I167360,);
not I_9722 (I166970,I167360);
nor I_9723 (I167382,I71920,I71914);
DFFARX1 I_9724 (I167382,I2067,I166978,I167408,);
and I_9725 (I167416,I167408,I71896);
nor I_9726 (I167433,I167416,I167334);
DFFARX1 I_9727 (I167433,I2067,I166978,I166961,);
nor I_9728 (I167464,I167408,I167193);
DFFARX1 I_9729 (I167464,I2067,I166978,I166943,);
nor I_9730 (I166958,I167408,I167097);
not I_9731 (I167539,I2074);
DFFARX1 I_9732 (I82491,I2067,I167539,I167565,);
DFFARX1 I_9733 (I82485,I2067,I167539,I167582,);
not I_9734 (I167590,I167582);
nor I_9735 (I167507,I167565,I167590);
DFFARX1 I_9736 (I167590,I2067,I167539,I167522,);
nor I_9737 (I167635,I82482,I82473);
and I_9738 (I167652,I167635,I82470);
nor I_9739 (I167669,I167652,I82482);
not I_9740 (I167686,I82482);
and I_9741 (I167703,I167686,I82476);
nand I_9742 (I167720,I167703,I82488);
nor I_9743 (I167737,I167686,I167720);
DFFARX1 I_9744 (I167737,I2067,I167539,I167504,);
not I_9745 (I167768,I167720);
nand I_9746 (I167785,I167590,I167768);
nand I_9747 (I167516,I167652,I167768);
DFFARX1 I_9748 (I167686,I2067,I167539,I167531,);
not I_9749 (I167830,I82494);
nor I_9750 (I167847,I167830,I82476);
nor I_9751 (I167864,I167847,I167669);
DFFARX1 I_9752 (I167864,I2067,I167539,I167528,);
not I_9753 (I167895,I167847);
DFFARX1 I_9754 (I167895,I2067,I167539,I167921,);
not I_9755 (I167929,I167921);
nor I_9756 (I167525,I167929,I167847);
nor I_9757 (I167960,I167830,I82473);
and I_9758 (I167977,I167960,I82479);
or I_9759 (I167994,I167977,I82470);
DFFARX1 I_9760 (I167994,I2067,I167539,I168020,);
not I_9761 (I168028,I168020);
nand I_9762 (I168045,I168028,I167768);
not I_9763 (I167519,I168045);
nand I_9764 (I167513,I168045,I167785);
nand I_9765 (I167510,I168028,I167652);
not I_9766 (I168134,I2074);
DFFARX1 I_9767 (I47029,I2067,I168134,I168160,);
DFFARX1 I_9768 (I47023,I2067,I168134,I168177,);
not I_9769 (I168185,I168177);
nor I_9770 (I168102,I168160,I168185);
DFFARX1 I_9771 (I168185,I2067,I168134,I168117,);
nor I_9772 (I168230,I47011,I47032);
and I_9773 (I168247,I168230,I47026);
nor I_9774 (I168264,I168247,I47011);
not I_9775 (I168281,I47011);
and I_9776 (I168298,I168281,I47008);
nand I_9777 (I168315,I168298,I47020);
nor I_9778 (I168332,I168281,I168315);
DFFARX1 I_9779 (I168332,I2067,I168134,I168099,);
not I_9780 (I168363,I168315);
nand I_9781 (I168380,I168185,I168363);
nand I_9782 (I168111,I168247,I168363);
DFFARX1 I_9783 (I168281,I2067,I168134,I168126,);
not I_9784 (I168425,I47035);
nor I_9785 (I168442,I168425,I47008);
nor I_9786 (I168459,I168442,I168264);
DFFARX1 I_9787 (I168459,I2067,I168134,I168123,);
not I_9788 (I168490,I168442);
DFFARX1 I_9789 (I168490,I2067,I168134,I168516,);
not I_9790 (I168524,I168516);
nor I_9791 (I168120,I168524,I168442);
nor I_9792 (I168555,I168425,I47017);
and I_9793 (I168572,I168555,I47014);
or I_9794 (I168589,I168572,I47008);
DFFARX1 I_9795 (I168589,I2067,I168134,I168615,);
not I_9796 (I168623,I168615);
nand I_9797 (I168640,I168623,I168363);
not I_9798 (I168114,I168640);
nand I_9799 (I168108,I168640,I168380);
nand I_9800 (I168105,I168623,I168247);
not I_9801 (I168729,I2074);
DFFARX1 I_9802 (I96941,I2067,I168729,I168755,);
DFFARX1 I_9803 (I96923,I2067,I168729,I168772,);
not I_9804 (I168780,I168772);
nor I_9805 (I168697,I168755,I168780);
DFFARX1 I_9806 (I168780,I2067,I168729,I168712,);
nor I_9807 (I168825,I96929,I96932);
and I_9808 (I168842,I168825,I96920);
nor I_9809 (I168859,I168842,I96929);
not I_9810 (I168876,I96929);
and I_9811 (I168893,I168876,I96938);
nand I_9812 (I168910,I168893,I96926);
nor I_9813 (I168927,I168876,I168910);
DFFARX1 I_9814 (I168927,I2067,I168729,I168694,);
not I_9815 (I168958,I168910);
nand I_9816 (I168975,I168780,I168958);
nand I_9817 (I168706,I168842,I168958);
DFFARX1 I_9818 (I168876,I2067,I168729,I168721,);
not I_9819 (I169020,I96923);
nor I_9820 (I169037,I169020,I96938);
nor I_9821 (I169054,I169037,I168859);
DFFARX1 I_9822 (I169054,I2067,I168729,I168718,);
not I_9823 (I169085,I169037);
DFFARX1 I_9824 (I169085,I2067,I168729,I169111,);
not I_9825 (I169119,I169111);
nor I_9826 (I168715,I169119,I169037);
nor I_9827 (I169150,I169020,I96935);
and I_9828 (I169167,I169150,I96944);
or I_9829 (I169184,I169167,I96920);
DFFARX1 I_9830 (I169184,I2067,I168729,I169210,);
not I_9831 (I169218,I169210);
nand I_9832 (I169235,I169218,I168958);
not I_9833 (I168709,I169235);
nand I_9834 (I168703,I169235,I168975);
nand I_9835 (I168700,I169218,I168842);
not I_9836 (I169324,I2074);
DFFARX1 I_9837 (I156250,I2067,I169324,I169350,);
DFFARX1 I_9838 (I156253,I2067,I169324,I169367,);
not I_9839 (I169375,I169367);
nor I_9840 (I169292,I169350,I169375);
DFFARX1 I_9841 (I169375,I2067,I169324,I169307,);
nor I_9842 (I169420,I156253,I156268);
and I_9843 (I169437,I169420,I156262);
nor I_9844 (I169454,I169437,I156253);
not I_9845 (I169471,I156253);
and I_9846 (I169488,I169471,I156271);
nand I_9847 (I169505,I169488,I156259);
nor I_9848 (I169522,I169471,I169505);
DFFARX1 I_9849 (I169522,I2067,I169324,I169289,);
not I_9850 (I169553,I169505);
nand I_9851 (I169570,I169375,I169553);
nand I_9852 (I169301,I169437,I169553);
DFFARX1 I_9853 (I169471,I2067,I169324,I169316,);
not I_9854 (I169615,I156265);
nor I_9855 (I169632,I169615,I156271);
nor I_9856 (I169649,I169632,I169454);
DFFARX1 I_9857 (I169649,I2067,I169324,I169313,);
not I_9858 (I169680,I169632);
DFFARX1 I_9859 (I169680,I2067,I169324,I169706,);
not I_9860 (I169714,I169706);
nor I_9861 (I169310,I169714,I169632);
nor I_9862 (I169745,I169615,I156250);
and I_9863 (I169762,I169745,I156274);
or I_9864 (I169779,I169762,I156256);
DFFARX1 I_9865 (I169779,I2067,I169324,I169805,);
not I_9866 (I169813,I169805);
nand I_9867 (I169830,I169813,I169553);
not I_9868 (I169304,I169830);
nand I_9869 (I169298,I169830,I169570);
nand I_9870 (I169295,I169813,I169437);
not I_9871 (I169919,I2074);
DFFARX1 I_9872 (I139695,I2067,I169919,I169945,);
DFFARX1 I_9873 (I139707,I2067,I169919,I169962,);
not I_9874 (I169970,I169962);
nor I_9875 (I169887,I169945,I169970);
DFFARX1 I_9876 (I169970,I2067,I169919,I169902,);
nor I_9877 (I170015,I139704,I139698);
and I_9878 (I170032,I170015,I139692);
nor I_9879 (I170049,I170032,I139704);
not I_9880 (I170066,I139704);
and I_9881 (I170083,I170066,I139701);
nand I_9882 (I170100,I170083,I139692);
nor I_9883 (I170117,I170066,I170100);
DFFARX1 I_9884 (I170117,I2067,I169919,I169884,);
not I_9885 (I170148,I170100);
nand I_9886 (I170165,I169970,I170148);
nand I_9887 (I169896,I170032,I170148);
DFFARX1 I_9888 (I170066,I2067,I169919,I169911,);
not I_9889 (I170210,I139716);
nor I_9890 (I170227,I170210,I139701);
nor I_9891 (I170244,I170227,I170049);
DFFARX1 I_9892 (I170244,I2067,I169919,I169908,);
not I_9893 (I170275,I170227);
DFFARX1 I_9894 (I170275,I2067,I169919,I170301,);
not I_9895 (I170309,I170301);
nor I_9896 (I169905,I170309,I170227);
nor I_9897 (I170340,I170210,I139710);
and I_9898 (I170357,I170340,I139713);
or I_9899 (I170374,I170357,I139695);
DFFARX1 I_9900 (I170374,I2067,I169919,I170400,);
not I_9901 (I170408,I170400);
nand I_9902 (I170425,I170408,I170148);
not I_9903 (I169899,I170425);
nand I_9904 (I169893,I170425,I170165);
nand I_9905 (I169890,I170408,I170032);
not I_9906 (I170514,I2074);
DFFARX1 I_9907 (I81335,I2067,I170514,I170540,);
DFFARX1 I_9908 (I81329,I2067,I170514,I170557,);
not I_9909 (I170565,I170557);
nor I_9910 (I170482,I170540,I170565);
DFFARX1 I_9911 (I170565,I2067,I170514,I170497,);
nor I_9912 (I170610,I81326,I81317);
and I_9913 (I170627,I170610,I81314);
nor I_9914 (I170644,I170627,I81326);
not I_9915 (I170661,I81326);
and I_9916 (I170678,I170661,I81320);
nand I_9917 (I170695,I170678,I81332);
nor I_9918 (I170712,I170661,I170695);
DFFARX1 I_9919 (I170712,I2067,I170514,I170479,);
not I_9920 (I170743,I170695);
nand I_9921 (I170760,I170565,I170743);
nand I_9922 (I170491,I170627,I170743);
DFFARX1 I_9923 (I170661,I2067,I170514,I170506,);
not I_9924 (I170805,I81338);
nor I_9925 (I170822,I170805,I81320);
nor I_9926 (I170839,I170822,I170644);
DFFARX1 I_9927 (I170839,I2067,I170514,I170503,);
not I_9928 (I170870,I170822);
DFFARX1 I_9929 (I170870,I2067,I170514,I170896,);
not I_9930 (I170904,I170896);
nor I_9931 (I170500,I170904,I170822);
nor I_9932 (I170935,I170805,I81317);
and I_9933 (I170952,I170935,I81323);
or I_9934 (I170969,I170952,I81314);
DFFARX1 I_9935 (I170969,I2067,I170514,I170995,);
not I_9936 (I171003,I170995);
nand I_9937 (I171020,I171003,I170743);
not I_9938 (I170494,I171020);
nand I_9939 (I170488,I171020,I170760);
nand I_9940 (I170485,I171003,I170627);
not I_9941 (I171109,I2074);
DFFARX1 I_9942 (I23888,I2067,I171109,I171135,);
DFFARX1 I_9943 (I23891,I2067,I171109,I171152,);
not I_9944 (I171160,I171152);
nor I_9945 (I171077,I171135,I171160);
DFFARX1 I_9946 (I171160,I2067,I171109,I171092,);
nor I_9947 (I171205,I23897,I23891);
and I_9948 (I171222,I171205,I23894);
nor I_9949 (I171239,I171222,I23897);
not I_9950 (I171256,I23897);
and I_9951 (I171273,I171256,I23888);
nand I_9952 (I171290,I171273,I23906);
nor I_9953 (I171307,I171256,I171290);
DFFARX1 I_9954 (I171307,I2067,I171109,I171074,);
not I_9955 (I171338,I171290);
nand I_9956 (I171355,I171160,I171338);
nand I_9957 (I171086,I171222,I171338);
DFFARX1 I_9958 (I171256,I2067,I171109,I171101,);
not I_9959 (I171400,I23900);
nor I_9960 (I171417,I171400,I23888);
nor I_9961 (I171434,I171417,I171239);
DFFARX1 I_9962 (I171434,I2067,I171109,I171098,);
not I_9963 (I171465,I171417);
DFFARX1 I_9964 (I171465,I2067,I171109,I171491,);
not I_9965 (I171499,I171491);
nor I_9966 (I171095,I171499,I171417);
nor I_9967 (I171530,I171400,I23903);
and I_9968 (I171547,I171530,I23909);
or I_9969 (I171564,I171547,I23912);
DFFARX1 I_9970 (I171564,I2067,I171109,I171590,);
not I_9971 (I171598,I171590);
nand I_9972 (I171615,I171598,I171338);
not I_9973 (I171089,I171615);
nand I_9974 (I171083,I171615,I171355);
nand I_9975 (I171080,I171598,I171222);
not I_9976 (I171704,I2074);
DFFARX1 I_9977 (I157882,I2067,I171704,I171730,);
DFFARX1 I_9978 (I157885,I2067,I171704,I171747,);
not I_9979 (I171755,I171747);
nor I_9980 (I171672,I171730,I171755);
DFFARX1 I_9981 (I171755,I2067,I171704,I171687,);
nor I_9982 (I171800,I157885,I157900);
and I_9983 (I171817,I171800,I157894);
nor I_9984 (I171834,I171817,I157885);
not I_9985 (I171851,I157885);
and I_9986 (I171868,I171851,I157903);
nand I_9987 (I171885,I171868,I157891);
nor I_9988 (I171902,I171851,I171885);
DFFARX1 I_9989 (I171902,I2067,I171704,I171669,);
not I_9990 (I171933,I171885);
nand I_9991 (I171950,I171755,I171933);
nand I_9992 (I171681,I171817,I171933);
DFFARX1 I_9993 (I171851,I2067,I171704,I171696,);
not I_9994 (I171995,I157897);
nor I_9995 (I172012,I171995,I157903);
nor I_9996 (I172029,I172012,I171834);
DFFARX1 I_9997 (I172029,I2067,I171704,I171693,);
not I_9998 (I172060,I172012);
DFFARX1 I_9999 (I172060,I2067,I171704,I172086,);
not I_10000 (I172094,I172086);
nor I_10001 (I171690,I172094,I172012);
nor I_10002 (I172125,I171995,I157882);
and I_10003 (I172142,I172125,I157906);
or I_10004 (I172159,I172142,I157888);
DFFARX1 I_10005 (I172159,I2067,I171704,I172185,);
not I_10006 (I172193,I172185);
nand I_10007 (I172210,I172193,I171933);
not I_10008 (I171684,I172210);
nand I_10009 (I171678,I172210,I171950);
nand I_10010 (I171675,I172193,I171817);
not I_10011 (I172299,I2074);
DFFARX1 I_10012 (I139117,I2067,I172299,I172325,);
DFFARX1 I_10013 (I139129,I2067,I172299,I172342,);
not I_10014 (I172350,I172342);
nor I_10015 (I172267,I172325,I172350);
DFFARX1 I_10016 (I172350,I2067,I172299,I172282,);
nor I_10017 (I172395,I139126,I139120);
and I_10018 (I172412,I172395,I139114);
nor I_10019 (I172429,I172412,I139126);
not I_10020 (I172446,I139126);
and I_10021 (I172463,I172446,I139123);
nand I_10022 (I172480,I172463,I139114);
nor I_10023 (I172497,I172446,I172480);
DFFARX1 I_10024 (I172497,I2067,I172299,I172264,);
not I_10025 (I172528,I172480);
nand I_10026 (I172545,I172350,I172528);
nand I_10027 (I172276,I172412,I172528);
DFFARX1 I_10028 (I172446,I2067,I172299,I172291,);
not I_10029 (I172590,I139138);
nor I_10030 (I172607,I172590,I139123);
nor I_10031 (I172624,I172607,I172429);
DFFARX1 I_10032 (I172624,I2067,I172299,I172288,);
not I_10033 (I172655,I172607);
DFFARX1 I_10034 (I172655,I2067,I172299,I172681,);
not I_10035 (I172689,I172681);
nor I_10036 (I172285,I172689,I172607);
nor I_10037 (I172720,I172590,I139132);
and I_10038 (I172737,I172720,I139135);
or I_10039 (I172754,I172737,I139117);
DFFARX1 I_10040 (I172754,I2067,I172299,I172780,);
not I_10041 (I172788,I172780);
nand I_10042 (I172805,I172788,I172528);
not I_10043 (I172279,I172805);
nand I_10044 (I172273,I172805,I172545);
nand I_10045 (I172270,I172788,I172412);
not I_10046 (I172894,I2074);
DFFARX1 I_10047 (I95207,I2067,I172894,I172920,);
DFFARX1 I_10048 (I95189,I2067,I172894,I172937,);
not I_10049 (I172945,I172937);
nor I_10050 (I172862,I172920,I172945);
DFFARX1 I_10051 (I172945,I2067,I172894,I172877,);
nor I_10052 (I172990,I95195,I95198);
and I_10053 (I173007,I172990,I95186);
nor I_10054 (I173024,I173007,I95195);
not I_10055 (I173041,I95195);
and I_10056 (I173058,I173041,I95204);
nand I_10057 (I173075,I173058,I95192);
nor I_10058 (I173092,I173041,I173075);
DFFARX1 I_10059 (I173092,I2067,I172894,I172859,);
not I_10060 (I173123,I173075);
nand I_10061 (I173140,I172945,I173123);
nand I_10062 (I172871,I173007,I173123);
DFFARX1 I_10063 (I173041,I2067,I172894,I172886,);
not I_10064 (I173185,I95189);
nor I_10065 (I173202,I173185,I95204);
nor I_10066 (I173219,I173202,I173024);
DFFARX1 I_10067 (I173219,I2067,I172894,I172883,);
not I_10068 (I173250,I173202);
DFFARX1 I_10069 (I173250,I2067,I172894,I173276,);
not I_10070 (I173284,I173276);
nor I_10071 (I172880,I173284,I173202);
nor I_10072 (I173315,I173185,I95201);
and I_10073 (I173332,I173315,I95210);
or I_10074 (I173349,I173332,I95186);
DFFARX1 I_10075 (I173349,I2067,I172894,I173375,);
not I_10076 (I173383,I173375);
nand I_10077 (I173400,I173383,I173123);
not I_10078 (I172874,I173400);
nand I_10079 (I172868,I173400,I173140);
nand I_10080 (I172865,I173383,I173007);
not I_10081 (I173489,I2074);
DFFARX1 I_10082 (I5920,I2067,I173489,I173515,);
DFFARX1 I_10083 (I5902,I2067,I173489,I173532,);
not I_10084 (I173540,I173532);
nor I_10085 (I173457,I173515,I173540);
DFFARX1 I_10086 (I173540,I2067,I173489,I173472,);
nor I_10087 (I173585,I5902,I5917);
and I_10088 (I173602,I173585,I5911);
nor I_10089 (I173619,I173602,I5902);
not I_10090 (I173636,I5902);
and I_10091 (I173653,I173636,I5905);
nand I_10092 (I173670,I173653,I5908);
nor I_10093 (I173687,I173636,I173670);
DFFARX1 I_10094 (I173687,I2067,I173489,I173454,);
not I_10095 (I173718,I173670);
nand I_10096 (I173735,I173540,I173718);
nand I_10097 (I173466,I173602,I173718);
DFFARX1 I_10098 (I173636,I2067,I173489,I173481,);
not I_10099 (I173780,I5914);
nor I_10100 (I173797,I173780,I5905);
nor I_10101 (I173814,I173797,I173619);
DFFARX1 I_10102 (I173814,I2067,I173489,I173478,);
not I_10103 (I173845,I173797);
DFFARX1 I_10104 (I173845,I2067,I173489,I173871,);
not I_10105 (I173879,I173871);
nor I_10106 (I173475,I173879,I173797);
nor I_10107 (I173910,I173780,I5926);
and I_10108 (I173927,I173910,I5923);
or I_10109 (I173944,I173927,I5905);
DFFARX1 I_10110 (I173944,I2067,I173489,I173970,);
not I_10111 (I173978,I173970);
nand I_10112 (I173995,I173978,I173718);
not I_10113 (I173469,I173995);
nand I_10114 (I173463,I173995,I173735);
nand I_10115 (I173460,I173978,I173602);
not I_10116 (I174084,I2074);
DFFARX1 I_10117 (I86537,I2067,I174084,I174110,);
DFFARX1 I_10118 (I86519,I2067,I174084,I174127,);
not I_10119 (I174135,I174127);
nor I_10120 (I174052,I174110,I174135);
DFFARX1 I_10121 (I174135,I2067,I174084,I174067,);
nor I_10122 (I174180,I86525,I86528);
and I_10123 (I174197,I174180,I86516);
nor I_10124 (I174214,I174197,I86525);
not I_10125 (I174231,I86525);
and I_10126 (I174248,I174231,I86534);
nand I_10127 (I174265,I174248,I86522);
nor I_10128 (I174282,I174231,I174265);
DFFARX1 I_10129 (I174282,I2067,I174084,I174049,);
not I_10130 (I174313,I174265);
nand I_10131 (I174330,I174135,I174313);
nand I_10132 (I174061,I174197,I174313);
DFFARX1 I_10133 (I174231,I2067,I174084,I174076,);
not I_10134 (I174375,I86519);
nor I_10135 (I174392,I174375,I86534);
nor I_10136 (I174409,I174392,I174214);
DFFARX1 I_10137 (I174409,I2067,I174084,I174073,);
not I_10138 (I174440,I174392);
DFFARX1 I_10139 (I174440,I2067,I174084,I174466,);
not I_10140 (I174474,I174466);
nor I_10141 (I174070,I174474,I174392);
nor I_10142 (I174505,I174375,I86531);
and I_10143 (I174522,I174505,I86540);
or I_10144 (I174539,I174522,I86516);
DFFARX1 I_10145 (I174539,I2067,I174084,I174565,);
not I_10146 (I174573,I174565);
nand I_10147 (I174590,I174573,I174313);
not I_10148 (I174064,I174590);
nand I_10149 (I174058,I174590,I174330);
nand I_10150 (I174055,I174573,I174197);
not I_10151 (I174679,I2074);
DFFARX1 I_10152 (I148365,I2067,I174679,I174705,);
DFFARX1 I_10153 (I148377,I2067,I174679,I174722,);
not I_10154 (I174730,I174722);
nor I_10155 (I174647,I174705,I174730);
DFFARX1 I_10156 (I174730,I2067,I174679,I174662,);
nor I_10157 (I174775,I148374,I148368);
and I_10158 (I174792,I174775,I148362);
nor I_10159 (I174809,I174792,I148374);
not I_10160 (I174826,I148374);
and I_10161 (I174843,I174826,I148371);
nand I_10162 (I174860,I174843,I148362);
nor I_10163 (I174877,I174826,I174860);
DFFARX1 I_10164 (I174877,I2067,I174679,I174644,);
not I_10165 (I174908,I174860);
nand I_10166 (I174925,I174730,I174908);
nand I_10167 (I174656,I174792,I174908);
DFFARX1 I_10168 (I174826,I2067,I174679,I174671,);
not I_10169 (I174970,I148386);
nor I_10170 (I174987,I174970,I148371);
nor I_10171 (I175004,I174987,I174809);
DFFARX1 I_10172 (I175004,I2067,I174679,I174668,);
not I_10173 (I175035,I174987);
DFFARX1 I_10174 (I175035,I2067,I174679,I175061,);
not I_10175 (I175069,I175061);
nor I_10176 (I174665,I175069,I174987);
nor I_10177 (I175100,I174970,I148380);
and I_10178 (I175117,I175100,I148383);
or I_10179 (I175134,I175117,I148365);
DFFARX1 I_10180 (I175134,I2067,I174679,I175160,);
not I_10181 (I175168,I175160);
nand I_10182 (I175185,I175168,I174908);
not I_10183 (I174659,I175185);
nand I_10184 (I174653,I175185,I174925);
nand I_10185 (I174650,I175168,I174792);
not I_10186 (I175274,I2074);
DFFARX1 I_10187 (I110767,I2067,I175274,I175300,);
DFFARX1 I_10188 (I110764,I2067,I175274,I175317,);
not I_10189 (I175325,I175317);
nor I_10190 (I175242,I175300,I175325);
DFFARX1 I_10191 (I175325,I2067,I175274,I175257,);
nor I_10192 (I175370,I110779,I110761);
and I_10193 (I175387,I175370,I110758);
nor I_10194 (I175404,I175387,I110779);
not I_10195 (I175421,I110779);
and I_10196 (I175438,I175421,I110764);
nand I_10197 (I175455,I175438,I110776);
nor I_10198 (I175472,I175421,I175455);
DFFARX1 I_10199 (I175472,I2067,I175274,I175239,);
not I_10200 (I175503,I175455);
nand I_10201 (I175520,I175325,I175503);
nand I_10202 (I175251,I175387,I175503);
DFFARX1 I_10203 (I175421,I2067,I175274,I175266,);
not I_10204 (I175565,I110770);
nor I_10205 (I175582,I175565,I110764);
nor I_10206 (I175599,I175582,I175404);
DFFARX1 I_10207 (I175599,I2067,I175274,I175263,);
not I_10208 (I175630,I175582);
DFFARX1 I_10209 (I175630,I2067,I175274,I175656,);
not I_10210 (I175664,I175656);
nor I_10211 (I175260,I175664,I175582);
nor I_10212 (I175695,I175565,I110758);
and I_10213 (I175712,I175695,I110773);
or I_10214 (I175729,I175712,I110761);
DFFARX1 I_10215 (I175729,I2067,I175274,I175755,);
not I_10216 (I175763,I175755);
nand I_10217 (I175780,I175763,I175503);
not I_10218 (I175254,I175780);
nand I_10219 (I175248,I175780,I175520);
nand I_10220 (I175245,I175763,I175387);
not I_10221 (I175869,I2074);
DFFARX1 I_10222 (I12774,I2067,I175869,I175895,);
DFFARX1 I_10223 (I12762,I2067,I175869,I175912,);
not I_10224 (I175920,I175912);
nor I_10225 (I175837,I175895,I175920);
DFFARX1 I_10226 (I175920,I2067,I175869,I175852,);
nor I_10227 (I175965,I12753,I12777);
and I_10228 (I175982,I175965,I12756);
nor I_10229 (I175999,I175982,I12753);
not I_10230 (I176016,I12753);
and I_10231 (I176033,I176016,I12759);
nand I_10232 (I176050,I176033,I12771);
nor I_10233 (I176067,I176016,I176050);
DFFARX1 I_10234 (I176067,I2067,I175869,I175834,);
not I_10235 (I176098,I176050);
nand I_10236 (I176115,I175920,I176098);
nand I_10237 (I175846,I175982,I176098);
DFFARX1 I_10238 (I176016,I2067,I175869,I175861,);
not I_10239 (I176160,I12753);
nor I_10240 (I176177,I176160,I12759);
nor I_10241 (I176194,I176177,I175999);
DFFARX1 I_10242 (I176194,I2067,I175869,I175858,);
not I_10243 (I176225,I176177);
DFFARX1 I_10244 (I176225,I2067,I175869,I176251,);
not I_10245 (I176259,I176251);
nor I_10246 (I175855,I176259,I176177);
nor I_10247 (I176290,I176160,I12756);
and I_10248 (I176307,I176290,I12765);
or I_10249 (I176324,I176307,I12768);
DFFARX1 I_10250 (I176324,I2067,I175869,I176350,);
not I_10251 (I176358,I176350);
nand I_10252 (I176375,I176358,I176098);
not I_10253 (I175849,I176375);
nand I_10254 (I175843,I176375,I176115);
nand I_10255 (I175840,I176358,I175982);
not I_10256 (I176464,I2074);
DFFARX1 I_10257 (I155162,I2067,I176464,I176490,);
DFFARX1 I_10258 (I155165,I2067,I176464,I176507,);
not I_10259 (I176515,I176507);
nor I_10260 (I176432,I176490,I176515);
DFFARX1 I_10261 (I176515,I2067,I176464,I176447,);
nor I_10262 (I176560,I155165,I155180);
and I_10263 (I176577,I176560,I155174);
nor I_10264 (I176594,I176577,I155165);
not I_10265 (I176611,I155165);
and I_10266 (I176628,I176611,I155183);
nand I_10267 (I176645,I176628,I155171);
nor I_10268 (I176662,I176611,I176645);
DFFARX1 I_10269 (I176662,I2067,I176464,I176429,);
not I_10270 (I176693,I176645);
nand I_10271 (I176710,I176515,I176693);
nand I_10272 (I176441,I176577,I176693);
DFFARX1 I_10273 (I176611,I2067,I176464,I176456,);
not I_10274 (I176755,I155177);
nor I_10275 (I176772,I176755,I155183);
nor I_10276 (I176789,I176772,I176594);
DFFARX1 I_10277 (I176789,I2067,I176464,I176453,);
not I_10278 (I176820,I176772);
DFFARX1 I_10279 (I176820,I2067,I176464,I176846,);
not I_10280 (I176854,I176846);
nor I_10281 (I176450,I176854,I176772);
nor I_10282 (I176885,I176755,I155162);
and I_10283 (I176902,I176885,I155186);
or I_10284 (I176919,I176902,I155168);
DFFARX1 I_10285 (I176919,I2067,I176464,I176945,);
not I_10286 (I176953,I176945);
nand I_10287 (I176970,I176953,I176693);
not I_10288 (I176444,I176970);
nand I_10289 (I176438,I176970,I176710);
nand I_10290 (I176435,I176953,I176577);
not I_10291 (I177059,I2074);
DFFARX1 I_10292 (I112348,I2067,I177059,I177085,);
DFFARX1 I_10293 (I112345,I2067,I177059,I177102,);
not I_10294 (I177110,I177102);
nor I_10295 (I177027,I177085,I177110);
DFFARX1 I_10296 (I177110,I2067,I177059,I177042,);
nor I_10297 (I177155,I112360,I112342);
and I_10298 (I177172,I177155,I112339);
nor I_10299 (I177189,I177172,I112360);
not I_10300 (I177206,I112360);
and I_10301 (I177223,I177206,I112345);
nand I_10302 (I177240,I177223,I112357);
nor I_10303 (I177257,I177206,I177240);
DFFARX1 I_10304 (I177257,I2067,I177059,I177024,);
not I_10305 (I177288,I177240);
nand I_10306 (I177305,I177110,I177288);
nand I_10307 (I177036,I177172,I177288);
DFFARX1 I_10308 (I177206,I2067,I177059,I177051,);
not I_10309 (I177350,I112351);
nor I_10310 (I177367,I177350,I112345);
nor I_10311 (I177384,I177367,I177189);
DFFARX1 I_10312 (I177384,I2067,I177059,I177048,);
not I_10313 (I177415,I177367);
DFFARX1 I_10314 (I177415,I2067,I177059,I177441,);
not I_10315 (I177449,I177441);
nor I_10316 (I177045,I177449,I177367);
nor I_10317 (I177480,I177350,I112339);
and I_10318 (I177497,I177480,I112354);
or I_10319 (I177514,I177497,I112342);
DFFARX1 I_10320 (I177514,I2067,I177059,I177540,);
not I_10321 (I177548,I177540);
nand I_10322 (I177565,I177548,I177288);
not I_10323 (I177039,I177565);
nand I_10324 (I177033,I177565,I177305);
nand I_10325 (I177030,I177548,I177172);
not I_10326 (I177654,I2074);
DFFARX1 I_10327 (I123616,I2067,I177654,I177680,);
DFFARX1 I_10328 (I123634,I2067,I177654,I177697,);
not I_10329 (I177705,I177697);
nor I_10330 (I177622,I177680,I177705);
DFFARX1 I_10331 (I177705,I2067,I177654,I177637,);
nor I_10332 (I177750,I123613,I123625);
and I_10333 (I177767,I177750,I123610);
nor I_10334 (I177784,I177767,I123613);
not I_10335 (I177801,I123613);
and I_10336 (I177818,I177801,I123619);
nand I_10337 (I177835,I177818,I123631);
nor I_10338 (I177852,I177801,I177835);
DFFARX1 I_10339 (I177852,I2067,I177654,I177619,);
not I_10340 (I177883,I177835);
nand I_10341 (I177900,I177705,I177883);
nand I_10342 (I177631,I177767,I177883);
DFFARX1 I_10343 (I177801,I2067,I177654,I177646,);
not I_10344 (I177945,I123622);
nor I_10345 (I177962,I177945,I123619);
nor I_10346 (I177979,I177962,I177784);
DFFARX1 I_10347 (I177979,I2067,I177654,I177643,);
not I_10348 (I178010,I177962);
DFFARX1 I_10349 (I178010,I2067,I177654,I178036,);
not I_10350 (I178044,I178036);
nor I_10351 (I177640,I178044,I177962);
nor I_10352 (I178075,I177945,I123610);
and I_10353 (I178092,I178075,I123637);
or I_10354 (I178109,I178092,I123628);
DFFARX1 I_10355 (I178109,I2067,I177654,I178135,);
not I_10356 (I178143,I178135);
nand I_10357 (I178160,I178143,I177883);
not I_10358 (I177634,I178160);
nand I_10359 (I177628,I178160,I177900);
nand I_10360 (I177625,I178143,I177767);
not I_10361 (I178249,I2074);
DFFARX1 I_10362 (I34003,I2067,I178249,I178275,);
DFFARX1 I_10363 (I34006,I2067,I178249,I178292,);
not I_10364 (I178300,I178292);
nor I_10365 (I178217,I178275,I178300);
DFFARX1 I_10366 (I178300,I2067,I178249,I178232,);
nor I_10367 (I178345,I34012,I34006);
and I_10368 (I178362,I178345,I34009);
nor I_10369 (I178379,I178362,I34012);
not I_10370 (I178396,I34012);
and I_10371 (I178413,I178396,I34003);
nand I_10372 (I178430,I178413,I34021);
nor I_10373 (I178447,I178396,I178430);
DFFARX1 I_10374 (I178447,I2067,I178249,I178214,);
not I_10375 (I178478,I178430);
nand I_10376 (I178495,I178300,I178478);
nand I_10377 (I178226,I178362,I178478);
DFFARX1 I_10378 (I178396,I2067,I178249,I178241,);
not I_10379 (I178540,I34015);
nor I_10380 (I178557,I178540,I34003);
nor I_10381 (I178574,I178557,I178379);
DFFARX1 I_10382 (I178574,I2067,I178249,I178238,);
not I_10383 (I178605,I178557);
DFFARX1 I_10384 (I178605,I2067,I178249,I178631,);
not I_10385 (I178639,I178631);
nor I_10386 (I178235,I178639,I178557);
nor I_10387 (I178670,I178540,I34018);
and I_10388 (I178687,I178670,I34024);
or I_10389 (I178704,I178687,I34027);
DFFARX1 I_10390 (I178704,I2067,I178249,I178730,);
not I_10391 (I178738,I178730);
nand I_10392 (I178755,I178738,I178478);
not I_10393 (I178229,I178755);
nand I_10394 (I178223,I178755,I178495);
nand I_10395 (I178220,I178738,I178362);
not I_10396 (I178844,I2074);
DFFARX1 I_10397 (I36978,I2067,I178844,I178870,);
DFFARX1 I_10398 (I36981,I2067,I178844,I178887,);
not I_10399 (I178895,I178887);
nor I_10400 (I178812,I178870,I178895);
DFFARX1 I_10401 (I178895,I2067,I178844,I178827,);
nor I_10402 (I178940,I36987,I36981);
and I_10403 (I178957,I178940,I36984);
nor I_10404 (I178974,I178957,I36987);
not I_10405 (I178991,I36987);
and I_10406 (I179008,I178991,I36978);
nand I_10407 (I179025,I179008,I36996);
nor I_10408 (I179042,I178991,I179025);
DFFARX1 I_10409 (I179042,I2067,I178844,I178809,);
not I_10410 (I179073,I179025);
nand I_10411 (I179090,I178895,I179073);
nand I_10412 (I178821,I178957,I179073);
DFFARX1 I_10413 (I178991,I2067,I178844,I178836,);
not I_10414 (I179135,I36990);
nor I_10415 (I179152,I179135,I36978);
nor I_10416 (I179169,I179152,I178974);
DFFARX1 I_10417 (I179169,I2067,I178844,I178833,);
not I_10418 (I179200,I179152);
DFFARX1 I_10419 (I179200,I2067,I178844,I179226,);
not I_10420 (I179234,I179226);
nor I_10421 (I178830,I179234,I179152);
nor I_10422 (I179265,I179135,I36993);
and I_10423 (I179282,I179265,I36999);
or I_10424 (I179299,I179282,I37002);
DFFARX1 I_10425 (I179299,I2067,I178844,I179325,);
not I_10426 (I179333,I179325);
nand I_10427 (I179350,I179333,I179073);
not I_10428 (I178824,I179350);
nand I_10429 (I178818,I179350,I179090);
nand I_10430 (I178815,I179333,I178957);
endmodule


