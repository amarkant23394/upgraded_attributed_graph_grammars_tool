module test_final(IN_1_1_l_8,IN_2_1_l_8,IN_3_1_l_8,IN_1_3_l_8,IN_2_3_l_8,IN_3_3_l_8,IN_1_6_l_8,IN_2_6_l_8,IN_3_6_l_8,IN_4_6_l_8,IN_5_6_l_8,IN_1_8_l_8,IN_2_8_l_8,IN_3_8_l_8,IN_6_8_l_8,blif_clk_net_8_r_6,blif_reset_net_8_r_6,N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,N1372_10_r_6,N1508_10_r_6);
input IN_1_1_l_8,IN_2_1_l_8,IN_3_1_l_8,IN_1_3_l_8,IN_2_3_l_8,IN_3_3_l_8,IN_1_6_l_8,IN_2_6_l_8,IN_3_6_l_8,IN_4_6_l_8,IN_5_6_l_8,IN_1_8_l_8,IN_2_8_l_8,IN_3_8_l_8,IN_6_8_l_8,blif_clk_net_8_r_6,blif_reset_net_8_r_6;
output N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,N1372_10_r_6,N1508_10_r_6;
wire N1371_0_r_8,N1508_0_r_8,N1372_1_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,I_BUFF_1_9_r_8,N1372_10_r_8,N1508_10_r_8,N3_8_l_8,n53_8,n29_8,N3_8_r_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8,n38_8,n39_8,n40_8,n41_8,n42_8,n43_8,n44_8,n45_8,n46_8,n47_8,n48_8,n49_8,n50_8,n51_8,n52_8,I_BUFF_1_9_r_6,N3_8_r_6,n9_6,n30_6,n31_6,n32_6,n33_6,n34_6,n35_6,n36_6,n37_6,n38_6,n39_6,n40_6,n41_6,n42_6,n43_6,n44_6,n45_6,n46_6,n47_6,n48_6,n49_6,n50_6,n51_6,n52_6,n53_6,n54_6;
nor I_0(N1371_0_r_8,n46_8,n51_8);
not I_1(N1508_0_r_8,n46_8);
nor I_2(N1372_1_r_8,n37_8,n49_8);
and I_3(N1508_1_r_8,N1372_1_r_8,n29_8);
nor I_4(N1507_6_r_8,n47_8,n48_8);
nor I_5(N1508_6_r_8,n37_8,n38_8);
nor I_6(n_42_8_r_8,I_BUFF_1_9_r_8,n53_8);
DFFARX1 I_7(N3_8_r_8,blif_clk_net_8_r_6,n9_6,G199_8_r_8,);
nor I_8(N6147_9_r_8,n29_8,n30_8);
nor I_9(N6134_9_r_8,n30_8,n31_8);
not I_10(I_BUFF_1_9_r_8,n35_8);
nor I_11(N1372_10_r_8,n46_8,n49_8);
nor I_12(N1508_10_r_8,n40_8,n41_8);
and I_13(N3_8_l_8,IN_6_8_l_8,n36_8);
DFFARX1 I_14(N3_8_l_8,blif_clk_net_8_r_6,n9_6,n53_8,);
not I_15(n29_8,n53_8);
nor I_16(N3_8_r_8,n33_8,n34_8);
and I_17(n30_8,n32_8,n33_8);
nor I_18(n31_8,IN_1_8_l_8,IN_3_8_l_8);
nand I_19(n32_8,IN_2_6_l_8,n42_8);
or I_20(n33_8,IN_3_1_l_8,n46_8);
nor I_21(n34_8,n32_8,n35_8);
nand I_22(n35_8,IN_5_6_l_8,n44_8);
nand I_23(n36_8,IN_2_8_l_8,IN_3_8_l_8);
not I_24(n37_8,n31_8);
nand I_25(n38_8,N1508_0_r_8,n39_8);
nand I_26(n39_8,n33_8,n50_8);
and I_27(n40_8,n32_8,n35_8);
not I_28(n41_8,N1372_10_r_8);
and I_29(n42_8,IN_1_6_l_8,n43_8);
nand I_30(n43_8,n44_8,n45_8);
nand I_31(n44_8,IN_3_6_l_8,IN_4_6_l_8);
not I_32(n45_8,IN_5_6_l_8);
nand I_33(n46_8,IN_1_1_l_8,IN_2_1_l_8);
not I_34(n47_8,n39_8);
nor I_35(n48_8,n35_8,n49_8);
not I_36(n49_8,n51_8);
nand I_37(n50_8,I_BUFF_1_9_r_8,n51_8);
nor I_38(n51_8,IN_1_3_l_8,n52_8);
or I_39(n52_8,IN_2_3_l_8,IN_3_3_l_8);
nor I_40(N1371_0_r_6,n30_6,n33_6);
nor I_41(N1508_0_r_6,n33_6,n44_6);
not I_42(N1372_1_r_6,n41_6);
nor I_43(N1508_1_r_6,n40_6,n41_6);
nor I_44(N1507_6_r_6,n39_6,n45_6);
nor I_45(N1508_6_r_6,n37_6,n38_6);
nor I_46(n_42_8_r_6,n30_6,n31_6);
DFFARX1 I_47(N3_8_r_6,blif_clk_net_8_r_6,n9_6,G199_8_r_6,);
nor I_48(N6147_9_r_6,n32_6,n33_6);
nor I_49(N6134_9_r_6,I_BUFF_1_9_r_6,n35_6);
not I_50(I_BUFF_1_9_r_6,n37_6);
not I_51(N1372_10_r_6,n43_6);
nor I_52(N1508_10_r_6,n42_6,n43_6);
nor I_53(N3_8_r_6,n36_6,N6134_9_r_8);
not I_54(n9_6,blif_reset_net_8_r_6);
nor I_55(n30_6,n53_6,N1508_6_r_8);
not I_56(n31_6,n36_6);
nor I_57(n32_6,I_BUFF_1_9_r_6,n34_6);
not I_58(n33_6,N6134_9_r_8);
not I_59(n34_6,n35_6);
nand I_60(n35_6,n49_6,N1507_6_r_8);
nand I_61(n36_6,n51_6,n_42_8_r_8);
nand I_62(n37_6,n54_6,n_42_8_r_8);
or I_63(n38_6,n35_6,n39_6);
nor I_64(n39_6,n40_6,n45_6);
and I_65(n40_6,n46_6,n47_6);
nand I_66(n41_6,n30_6,n31_6);
nor I_67(n42_6,n34_6,n40_6);
nand I_68(n43_6,n30_6,N6134_9_r_8);
nor I_69(n44_6,n31_6,n40_6);
nor I_70(n45_6,n35_6,n36_6);
nor I_71(n46_6,N1508_1_r_8,N1371_0_r_8);
or I_72(n47_6,n48_6,N1508_1_r_8);
nor I_73(n48_6,N1371_0_r_8,N1508_10_r_8);
and I_74(n49_6,n50_6,G199_8_r_8);
nand I_75(n50_6,n51_6,n52_6);
nand I_76(n51_6,N1508_6_r_8,G199_8_r_8);
not I_77(n52_6,n_42_8_r_8);
nor I_78(n53_6,N1507_6_r_8,N6147_9_r_8);
or I_79(n54_6,N1507_6_r_8,N6147_9_r_8);
endmodule


