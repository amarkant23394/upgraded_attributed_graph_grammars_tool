module test_I1917(I1410,I1294,I1828,I1639,I1301,I1917);
input I1410,I1294,I1828,I1639,I1301;
output I1917;
wire I1328,I2313,I1937,I2505,I1331,I2389,I2406,I2488;
nand I_0(I1328,I1639,I1828);
nand I_1(I1917,I2406,I2505);
DFFARX1 I_2(I1331,I1294,I1937,,,I2313,);
not I_3(I1937,I1301);
nor I_4(I2505,I2313,I2488);
nor I_5(I1331,I1639,I1410);
DFFARX1 I_6(I1328,I1294,I1937,,,I2389,);
not I_7(I2406,I2389);
not I_8(I2488,I2406);
endmodule


