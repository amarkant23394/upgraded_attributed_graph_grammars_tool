module test_final(IN_1_1_l_2,IN_2_1_l_2,IN_3_1_l_2,IN_1_3_l_2,IN_2_3_l_2,IN_3_3_l_2,IN_1_4_l_2,IN_2_4_l_2,IN_3_4_l_2,IN_4_4_l_2,IN_5_4_l_2,blif_clk_net_5_r_0,blif_reset_net_5_r_0,N1371_0_r_0,N6147_2_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_547_5_r_0,N1507_6_r_0,N1508_6_r_0);
input IN_1_1_l_2,IN_2_1_l_2,IN_3_1_l_2,IN_1_3_l_2,IN_2_3_l_2,IN_3_3_l_2,IN_1_4_l_2,IN_2_4_l_2,IN_3_4_l_2,IN_4_4_l_2,IN_5_4_l_2,blif_clk_net_5_r_0,blif_reset_net_5_r_0;
output N1371_0_r_0,N6147_2_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_547_5_r_0,N1507_6_r_0,N1508_6_r_0;
wire N1371_0_r_2,N1508_0_r_2,N6147_3_r_2,n_429_or_0_5_r_2,G78_5_r_2,n_576_5_r_2,n_102_5_r_2,n_547_5_r_2,N1372_10_r_2,N1508_10_r_2,n_431_5_r_2,n21_2,n22_2,n23_2,n24_2,n25_2,n26_2,n27_2,n28_2,n29_2,n30_2,n31_2,n32_2,N1508_0_r_0,n_102_5_r_0,N3_8_l_0,n5_0,n40_0,n4_0,n23_0,n24_0,n25_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0,n37_0,n38_0,n39_0;
nor I_0(N1371_0_r_2,n23_2,n24_2);
not I_1(N1508_0_r_2,n24_2);
nor I_2(N6147_3_r_2,n22_2,n26_2);
nand I_3(n_429_or_0_5_r_2,IN_3_1_l_2,n22_2);
DFFARX1 I_4(n_431_5_r_2,blif_clk_net_5_r_0,n5_0,G78_5_r_2,);
nand I_5(n_576_5_r_2,n21_2,n22_2);
not I_6(n_102_5_r_2,n23_2);
nand I_7(n_547_5_r_2,n22_2,n24_2);
not I_8(N1372_10_r_2,n29_2);
nor I_9(N1508_10_r_2,n28_2,n29_2);
nand I_10(n_431_5_r_2,n_102_5_r_2,n25_2);
nor I_11(n21_2,IN_3_1_l_2,n23_2);
and I_12(n22_2,IN_1_1_l_2,IN_2_1_l_2);
nor I_13(n23_2,n24_2,n31_2);
nand I_14(n24_2,IN_1_4_l_2,IN_2_4_l_2);
nand I_15(n25_2,n26_2,n27_2);
nor I_16(n26_2,IN_1_3_l_2,n30_2);
not I_17(n27_2,n_429_or_0_5_r_2);
nor I_18(n28_2,n22_2,n23_2);
nand I_19(n29_2,N1508_0_r_2,n26_2);
or I_20(n30_2,IN_2_3_l_2,IN_3_3_l_2);
nor I_21(n31_2,IN_5_4_l_2,n32_2);
and I_22(n32_2,IN_3_4_l_2,IN_4_4_l_2);
nor I_23(N1371_0_r_0,n24_0,n25_0);
not I_24(N1508_0_r_0,n25_0);
nor I_25(N6147_2_r_0,n28_0,n29_0);
nand I_26(n_429_or_0_5_r_0,n4_0,n25_0);
DFFARX1 I_27(n4_0,blif_clk_net_5_r_0,n5_0,G78_5_r_0,);
nand I_28(n_576_5_r_0,n23_0,n24_0);
not I_29(n_102_5_r_0,n40_0);
nand I_30(n_547_5_r_0,n26_0,n27_0);
nor I_31(N1507_6_r_0,n_102_5_r_0,n37_0);
nor I_32(N1508_6_r_0,n25_0,n33_0);
and I_33(N3_8_l_0,n32_0,n_547_5_r_2);
not I_34(n5_0,blif_reset_net_5_r_0);
DFFARX1 I_35(N3_8_l_0,blif_clk_net_5_r_0,n5_0,n40_0,);
not I_36(n4_0,n31_0);
nor I_37(n23_0,n40_0,n25_0);
and I_38(n24_0,n4_0,n39_0);
nand I_39(n25_0,G78_5_r_2,n_576_5_r_2);
nor I_40(n26_0,n40_0,n24_0);
nor I_41(n27_0,N6147_3_r_2,N1508_10_r_2);
nor I_42(n28_0,n25_0,N6147_3_r_2);
nand I_43(n29_0,n_102_5_r_0,n30_0);
nand I_44(n30_0,n27_0,n31_0);
nand I_45(n31_0,n_576_5_r_2,N1371_0_r_2);
nand I_46(n32_0,N1371_0_r_2,N1508_10_r_2);
nand I_47(n33_0,n34_0,n35_0);
nand I_48(n34_0,n_102_5_r_0,n36_0);
not I_49(n35_0,N6147_3_r_2);
not I_50(n36_0,n27_0);
nor I_51(n37_0,n36_0,n38_0);
nand I_52(n38_0,N1508_0_r_0,n35_0);
or I_53(n39_0,n_547_5_r_2,N1372_10_r_2);
endmodule


