module test_final(IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_6_2_l_10,IN_1_3_l_10,IN_2_3_l_10,IN_4_3_l_10,IN_1_4_l_10,IN_2_4_l_10,IN_3_4_l_10,IN_6_4_l_10,blif_clk_net_1_r_15,blif_reset_net_1_r_15,G42_1_r_15,n_572_1_r_15,n_573_1_r_15,n_549_1_r_15,n_569_1_r_15,ACVQN2_3_r_15,n_266_and_0_3_r_15,G199_4_r_15,G214_4_r_15);
input IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_6_2_l_10,IN_1_3_l_10,IN_2_3_l_10,IN_4_3_l_10,IN_1_4_l_10,IN_2_4_l_10,IN_3_4_l_10,IN_6_4_l_10,blif_clk_net_1_r_15,blif_reset_net_1_r_15;
output G42_1_r_15,n_572_1_r_15,n_573_1_r_15,n_549_1_r_15,n_569_1_r_15,ACVQN2_3_r_15,n_266_and_0_3_r_15,G199_4_r_15,G214_4_r_15;
wire G42_1_r_10,n_572_1_r_10,n_573_1_r_10,n_549_1_r_10,n_452_1_r_10,n_42_2_r_10,G199_2_r_10,ACVQN2_3_r_10,n_266_and_0_3_r_10,N3_2_l_10,n25_10,n16_10,n26_10,ACVQN1_3_l_10,N1_4_l_10,G199_4_l_10,n27_10,n17_10,n4_1_r_10,N3_2_r_10,n3_10,n13_internal_10,n13_10,n18_10,n19_10,n20_10,n21_10,n22_10,n23_10,n24_10,n_452_1_r_15,n4_1_l_15,n4_15,G42_1_l_15,n15_15,n17_internal_15,n17_15,n30_15,n_572_1_l_15,n14_internal_15,n14_15,N1_4_r_15,n_573_1_l_15,n18_15,n19_15,n20_15,n21_15,n22_15,n23_15,n24_15,n25_15,n26_15,n27_15,n28_15,n29_15;
DFFARX1 I_0(n4_1_r_10,blif_clk_net_1_r_15,n4_15,G42_1_r_10,);
nor I_1(n_572_1_r_10,n26_10,n3_10);
nand I_2(n_573_1_r_10,n16_10,n18_10);
nand I_3(n_549_1_r_10,n19_10,n20_10);
nor I_4(n_452_1_r_10,n25_10,n21_10);
nor I_5(n_42_2_r_10,n26_10,G199_4_l_10);
DFFARX1 I_6(N3_2_r_10,blif_clk_net_1_r_15,n4_15,G199_2_r_10,);
DFFARX1 I_7(G199_4_l_10,blif_clk_net_1_r_15,n4_15,ACVQN2_3_r_10,);
nor I_8(n_266_and_0_3_r_10,n17_10,n13_10);
and I_9(N3_2_l_10,IN_6_2_l_10,n23_10);
DFFARX1 I_10(N3_2_l_10,blif_clk_net_1_r_15,n4_15,n25_10,);
not I_11(n16_10,n25_10);
DFFARX1 I_12(IN_1_3_l_10,blif_clk_net_1_r_15,n4_15,n26_10,);
DFFARX1 I_13(IN_2_3_l_10,blif_clk_net_1_r_15,n4_15,ACVQN1_3_l_10,);
and I_14(N1_4_l_10,IN_6_4_l_10,n24_10);
DFFARX1 I_15(N1_4_l_10,blif_clk_net_1_r_15,n4_15,G199_4_l_10,);
DFFARX1 I_16(IN_3_4_l_10,blif_clk_net_1_r_15,n4_15,n27_10,);
not I_17(n17_10,n27_10);
nor I_18(n4_1_r_10,n27_10,n21_10);
nor I_19(N3_2_r_10,n16_10,n22_10);
not I_20(n3_10,n18_10);
DFFARX1 I_21(n3_10,blif_clk_net_1_r_15,n4_15,n13_internal_10,);
not I_22(n13_10,n13_internal_10);
nand I_23(n18_10,IN_4_3_l_10,ACVQN1_3_l_10);
not I_24(n19_10,n_452_1_r_10);
nand I_25(n20_10,n16_10,n26_10);
nor I_26(n21_10,IN_1_2_l_10,IN_3_2_l_10);
and I_27(n22_10,n26_10,n21_10);
nand I_28(n23_10,IN_2_2_l_10,IN_3_2_l_10);
nand I_29(n24_10,IN_1_4_l_10,IN_2_4_l_10);
DFFARX1 I_30(n_452_1_r_15,blif_clk_net_1_r_15,n4_15,G42_1_r_15,);
and I_31(n_572_1_r_15,n17_15,n19_15);
nand I_32(n_573_1_r_15,n15_15,n18_15);
nor I_33(n_549_1_r_15,n21_15,n22_15);
nand I_34(n_569_1_r_15,n15_15,n20_15);
nor I_35(n_452_1_r_15,n23_15,n24_15);
DFFARX1 I_36(G42_1_l_15,blif_clk_net_1_r_15,n4_15,ACVQN2_3_r_15,);
nor I_37(n_266_and_0_3_r_15,n17_15,n14_15);
DFFARX1 I_38(N1_4_r_15,blif_clk_net_1_r_15,n4_15,G199_4_r_15,);
DFFARX1 I_39(n_573_1_l_15,blif_clk_net_1_r_15,n4_15,G214_4_r_15,);
nor I_40(n4_1_l_15,n_42_2_r_10,n_572_1_r_10);
not I_41(n4_15,blif_reset_net_1_r_15);
DFFARX1 I_42(n4_1_l_15,blif_clk_net_1_r_15,n4_15,G42_1_l_15,);
not I_43(n15_15,G42_1_l_15);
DFFARX1 I_44(n_549_1_r_10,blif_clk_net_1_r_15,n4_15,n17_internal_15,);
not I_45(n17_15,n17_internal_15);
DFFARX1 I_46(G42_1_r_10,blif_clk_net_1_r_15,n4_15,n30_15,);
nor I_47(n_572_1_l_15,n_572_1_r_10,n_266_and_0_3_r_10);
DFFARX1 I_48(n_572_1_l_15,blif_clk_net_1_r_15,n4_15,n14_internal_15,);
not I_49(n14_15,n14_internal_15);
nand I_50(N1_4_r_15,n25_15,n26_15);
or I_51(n_573_1_l_15,G42_1_r_10,ACVQN2_3_r_10);
nor I_52(n18_15,G42_1_r_10,n_573_1_r_10);
nand I_53(n19_15,n27_15,n28_15);
nand I_54(n20_15,n30_15,G199_2_r_10);
not I_55(n21_15,n20_15);
and I_56(n22_15,n17_15,n_572_1_l_15);
nor I_57(n23_15,n_42_2_r_10,ACVQN2_3_r_10);
or I_58(n24_15,G42_1_r_10,n_573_1_r_10);
or I_59(n25_15,n_573_1_l_15,n_42_2_r_10);
nand I_60(n26_15,n19_15,n23_15);
not I_61(n27_15,n_573_1_r_10);
nand I_62(n28_15,n29_15,n_573_1_r_10);
not I_63(n29_15,n_572_1_r_10);
endmodule


