module test_I11310_rst(I1477_rst,I11310_rst);
,I11310_rst);
input I1477_rst;
output I11310_rst;
wire ;
not I_0(I11310_rst,I1477_rst);
endmodule


