module test_I15341(I12930,I1477,I1470,I12882,I15341);
input I12930,I1477,I1470,I12882;
output I15341;
wire I12619,I12718,I14982,I10615,I12596,I13119,I10639,I15276,I12599,I12964,I14965;
not I_0(I12619,I1477);
nor I_1(I12718,I10615,I10639);
not I_2(I14982,I12596);
DFFARX1 I_3(I1470,,,I10615,);
DFFARX1 I_4(I13119,I1470,I12619,,,I12596,);
or I_5(I13119,I12718);
DFFARX1 I_6(I1470,,,I10639,);
nand I_7(I15276,I14982,I12599);
nand I_8(I12599,I12718,I12964);
nor I_9(I12964,I12930,I12882);
not I_10(I14965,I1477);
DFFARX1 I_11(I15276,I1470,I14965,,,I15341,);
endmodule


