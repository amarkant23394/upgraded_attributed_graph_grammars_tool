module test_I3168(I2815,I2668,I1911,I1301,I2022,I1294,I3168);
input I2815,I2668,I1911,I1301,I2022,I1294;
output I3168;
wire I2897,I2600,I2583,I2313,I2344,I2849,I1923,I2685,I2914,I3086,I3103,I2832,I1920;
nand I_0(I2897,I2600,I1923);
not I_1(I2600,I1911);
or I_2(I3168,I3103,I2914);
not I_3(I2583,I1301);
DFFARX1 I_4(I1294,,,I2313,);
nor I_5(I2344,I2313);
nor I_6(I2849,I2832,I2685);
nand I_7(I1923,I2022,I2344);
not I_8(I2685,I2668);
and I_9(I2914,I2897,I2849);
DFFARX1 I_10(I1920,I1294,I2583,,,I3086,);
not I_11(I3103,I3086);
DFFARX1 I_12(I2815,I1294,I2583,,,I2832,);
not I_13(I1920,I2313);
endmodule


