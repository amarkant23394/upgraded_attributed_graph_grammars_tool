module test_final(IN_1_1_l_16,IN_2_1_l_16,IN_3_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_3_3_l_16,IN_1_6_l_16,IN_2_6_l_16,IN_3_6_l_16,IN_4_6_l_16,IN_5_6_l_16,IN_1_8_l_16,IN_2_8_l_16,IN_3_8_l_16,IN_6_8_l_16,blif_clk_net_7_r_12,blif_reset_net_7_r_12,N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_549_7_r_12,n_569_7_r_12,N6147_9_r_12);
input IN_1_1_l_16,IN_2_1_l_16,IN_3_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_3_3_l_16,IN_1_6_l_16,IN_2_6_l_16,IN_3_6_l_16,IN_4_6_l_16,IN_5_6_l_16,IN_1_8_l_16,IN_2_8_l_16,IN_3_8_l_16,IN_6_8_l_16,blif_clk_net_7_r_12,blif_reset_net_7_r_12;
output N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_549_7_r_12,n_569_7_r_12,N6147_9_r_12;
wire N1371_0_r_16,N1508_0_r_16,N1372_1_r_16,N1508_1_r_16,N6147_2_r_16,N1507_6_r_16,N1508_6_r_16,G42_7_r_16,n_572_7_r_16,n_573_7_r_16,n_549_7_r_16,n_569_7_r_16,n_452_7_r_16,N3_8_l_16,n53_16,n29_16,n4_7_r_16,n30_16,n31_16,n32_16,n33_16,n34_16,n35_16,n36_16,n37_16,n38_16,n39_16,n40_16,n41_16,n42_16,n43_16,n44_16,n45_16,n46_16,n47_16,n48_16,n49_16,n50_16,n51_16,n52_16,n_573_7_r_12,n_452_7_r_12,N6134_9_r_12,I_BUFF_1_9_r_12,n1_12,n8_12,n23_12,n24_12,n25_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12,n41_12,n42_12;
nor I_0(N1371_0_r_16,n35_16,n39_16);
nor I_1(N1508_0_r_16,n39_16,n46_16);
not I_2(N1372_1_r_16,n45_16);
nor I_3(N1508_1_r_16,n53_16,n45_16);
nor I_4(N6147_2_r_16,n37_16,n38_16);
nor I_5(N1507_6_r_16,n44_16,n49_16);
nor I_6(N1508_6_r_16,n29_16,n42_16);
DFFARX1 I_7(n4_7_r_16,blif_clk_net_7_r_12,n8_12,G42_7_r_16,);
nor I_8(n_572_7_r_16,n32_16,n33_16);
nand I_9(n_573_7_r_16,n30_16,n31_16);
nand I_10(n_549_7_r_16,IN_5_6_l_16,n47_16);
nand I_11(n_569_7_r_16,n_549_7_r_16,n30_16);
nor I_12(n_452_7_r_16,n34_16,n35_16);
and I_13(N3_8_l_16,IN_6_8_l_16,n41_16);
DFFARX1 I_14(N3_8_l_16,blif_clk_net_7_r_12,n8_12,n53_16,);
not I_15(n29_16,n53_16);
nor I_16(n4_7_r_16,n35_16,n36_16);
nand I_17(n30_16,IN_1_1_l_16,IN_2_1_l_16);
not I_18(n31_16,n34_16);
nor I_19(n32_16,IN_3_1_l_16,n30_16);
not I_20(n33_16,n_549_7_r_16);
nor I_21(n34_16,IN_1_3_l_16,n48_16);
and I_22(n35_16,IN_2_6_l_16,n50_16);
not I_23(n36_16,n30_16);
nor I_24(n37_16,n31_16,n40_16);
nand I_25(n38_16,n29_16,n39_16);
not I_26(n39_16,n32_16);
nor I_27(n40_16,IN_1_8_l_16,IN_3_8_l_16);
nand I_28(n41_16,IN_2_8_l_16,IN_3_8_l_16);
nand I_29(n42_16,n35_16,n43_16);
not I_30(n43_16,n44_16);
nor I_31(n44_16,n32_16,n49_16);
nand I_32(n45_16,n36_16,n40_16);
nor I_33(n46_16,n33_16,n34_16);
nand I_34(n47_16,IN_3_6_l_16,IN_4_6_l_16);
or I_35(n48_16,IN_2_3_l_16,IN_3_3_l_16);
and I_36(n49_16,n35_16,n36_16);
and I_37(n50_16,IN_1_6_l_16,n51_16);
nand I_38(n51_16,n47_16,n52_16);
not I_39(n52_16,IN_5_6_l_16);
nor I_40(N1371_0_r_12,I_BUFF_1_9_r_12,n36_12);
nand I_41(N1508_0_r_12,n30_12,n37_12);
nor I_42(N1507_6_r_12,n25_12,n39_12);
nor I_43(N1508_6_r_12,n25_12,n29_12);
DFFARX1 I_44(n1_12,blif_clk_net_7_r_12,n8_12,G42_7_r_12,);
nor I_45(n_572_7_r_12,n23_12,n24_12);
nand I_46(n_573_7_r_12,n_452_7_r_12,n25_12);
nand I_47(n_549_7_r_12,n27_12,n28_12);
nand I_48(n_569_7_r_12,n25_12,n26_12);
nand I_49(n_452_7_r_12,N1372_1_r_16,N1507_6_r_16);
nand I_50(N6147_9_r_12,n30_12,n31_12);
nor I_51(N6134_9_r_12,n35_12,n36_12);
not I_52(I_BUFF_1_9_r_12,n_452_7_r_12);
not I_53(n1_12,n_573_7_r_12);
not I_54(n8_12,blif_reset_net_7_r_12);
not I_55(n23_12,n36_12);
nor I_56(n24_12,n_452_7_r_12,G42_7_r_16);
nand I_57(n25_12,n23_12,n40_12);
not I_58(n26_12,n35_12);
not I_59(n27_12,N6134_9_r_12);
nand I_60(n28_12,n26_12,n29_12);
not I_61(n29_12,n24_12);
nand I_62(n30_12,n33_12,n41_12);
nand I_63(n31_12,n32_12,n33_12);
nor I_64(n32_12,n26_12,n34_12);
nor I_65(n33_12,N1371_0_r_16,N1508_0_r_16);
nor I_66(n34_12,n42_12,n_569_7_r_16);
nor I_67(n35_12,n38_12,n_452_7_r_16);
nand I_68(n36_12,N1508_1_r_16,n_573_7_r_16);
nand I_69(n37_12,n23_12,n35_12);
or I_70(n38_12,N6147_2_r_16,N1508_6_r_16);
not I_71(n39_12,n30_12);
or I_72(n40_12,N1508_0_r_16,N1372_1_r_16);
nor I_73(n41_12,n34_12,n36_12);
nor I_74(n42_12,n_572_7_r_16,N1371_0_r_16);
endmodule


