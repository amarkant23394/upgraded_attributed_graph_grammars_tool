module test_I7881(I6589,I1477,I1470,I4263,I4068,I7881);
input I6589,I1477,I1470,I4263,I4068;
output I7881;
wire I6606,I6300,I3948,I7587,I6329,I6688,I6705,I6291,I3972;
DFFARX1 I_0(I6589,I1470,I6329,,,I6606,);
DFFARX1 I_1(I6606,I1470,I6329,,,I6300,);
nand I_2(I7881,I7587,I6291);
DFFARX1 I_3(I1470,,,I3948,);
not I_4(I7587,I6300);
not I_5(I6329,I1477);
DFFARX1 I_6(I3948,I1470,I6329,,,I6688,);
and I_7(I6705,I6688,I3972);
DFFARX1 I_8(I6705,I1470,I6329,,,I6291,);
or I_9(I3972,I4263,I4068);
endmodule


