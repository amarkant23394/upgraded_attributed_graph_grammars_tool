module test_I12106(I1477,I1470,I10202,I10120,I12106);
input I1477,I1470,I10202,I10120;
output I12106;
wire I10219,I10154,I10020,I10137,I10052,I10287;
DFFARX1 I_0(I10202,I1470,I10052,,,I10219,);
nand I_1(I10154,I10137,I10120);
DFFARX1 I_2(I10287,I1470,I10052,,,I10020,);
not I_3(I12106,I10020);
DFFARX1 I_4(I1470,I10052,,,I10137,);
not I_5(I10052,I1477);
and I_6(I10287,I10219,I10154);
endmodule


