module test_final(G18_1_l_14,G15_1_l_14,IN_1_1_l_14,IN_4_1_l_14,IN_5_1_l_14,IN_7_1_l_14,IN_9_1_l_14,IN_10_1_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_4_3_l_14,blif_clk_net_1_r_5,blif_reset_net_1_r_5,G42_1_r_5,n_572_1_r_5,n_573_1_r_5,n_549_1_r_5,n_569_1_r_5,n_452_1_r_5,ACVQN2_3_r_5,n_266_and_0_3_r_5,ACVQN1_5_r_5,P6_5_r_5);
input G18_1_l_14,G15_1_l_14,IN_1_1_l_14,IN_4_1_l_14,IN_5_1_l_14,IN_7_1_l_14,IN_9_1_l_14,IN_10_1_l_14,IN_1_3_l_14,IN_2_3_l_14,IN_4_3_l_14,blif_clk_net_1_r_5,blif_reset_net_1_r_5;
output G42_1_r_5,n_572_1_r_5,n_573_1_r_5,n_549_1_r_5,n_569_1_r_5,n_452_1_r_5,ACVQN2_3_r_5,n_266_and_0_3_r_5,ACVQN1_5_r_5,P6_5_r_5;
wire G42_1_r_14,n_572_1_r_14,n_573_1_r_14,n_549_1_r_14,n_569_1_r_14,n_452_1_r_14,n_42_2_r_14,G199_2_r_14,ACVQN1_5_r_14,P6_5_r_14,n4_1_l_14,n15_internal_14,n15_14,ACVQN2_3_l_14,ACVQN1_3_l_14,N3_2_r_14,n_572_1_l_14,P6_5_r_internal_14,n16_14,n17_14,n18_14,n19_14,n20_14,n21_14,n22_14,n23_14,n24_14,n25_14,n26_14,n27_14,n28_14,N3_2_l_5,n5_5,G199_2_l_5,ACVQN2_3_l_5,n13_5,ACVQN1_3_l_5,N1_4_l_5,n21_5,n15_5,n22_5,n4_1_r_5,n11_internal_5,n11_5,n_42_2_l_5,n1_5,P6_5_r_internal_5,n16_5,n17_5,n18_5,n19_5,n20_5;
DFFARX1 I_0(n_452_1_r_14,blif_clk_net_1_r_5,n5_5,G42_1_r_14,);
and I_1(n_572_1_r_14,n18_14,n19_14);
nand I_2(n_573_1_r_14,n16_14,n17_14);
nor I_3(n_549_1_r_14,n20_14,n21_14);
or I_4(n_569_1_r_14,n_572_1_l_14,n20_14);
nor I_5(n_452_1_r_14,IN_10_1_l_14,n23_14);
nor I_6(n_42_2_r_14,n20_14,n22_14);
DFFARX1 I_7(N3_2_r_14,blif_clk_net_1_r_5,n5_5,G199_2_r_14,);
DFFARX1 I_8(n_572_1_l_14,blif_clk_net_1_r_5,n5_5,ACVQN1_5_r_14,);
not I_9(P6_5_r_14,P6_5_r_internal_14);
nor I_10(n4_1_l_14,G18_1_l_14,IN_1_1_l_14);
DFFARX1 I_11(n4_1_l_14,blif_clk_net_1_r_5,n5_5,n15_internal_14,);
not I_12(n15_14,n15_internal_14);
DFFARX1 I_13(IN_1_3_l_14,blif_clk_net_1_r_5,n5_5,ACVQN2_3_l_14,);
DFFARX1 I_14(IN_2_3_l_14,blif_clk_net_1_r_5,n5_5,ACVQN1_3_l_14,);
and I_15(N3_2_r_14,n26_14,n27_14);
nor I_16(n_572_1_l_14,G15_1_l_14,IN_7_1_l_14);
DFFARX1 I_17(ACVQN2_3_l_14,blif_clk_net_1_r_5,n5_5,P6_5_r_internal_14,);
nor I_18(n16_14,IN_9_1_l_14,IN_10_1_l_14);
not I_19(n17_14,n_572_1_l_14);
nor I_20(n18_14,IN_5_1_l_14,IN_9_1_l_14);
nand I_21(n19_14,IN_4_3_l_14,ACVQN1_3_l_14);
nor I_22(n20_14,G18_1_l_14,IN_5_1_l_14);
nor I_23(n21_14,n15_14,n22_14);
nand I_24(n22_14,n24_14,n25_14);
nand I_25(n23_14,n15_14,n24_14);
not I_26(n24_14,IN_9_1_l_14);
not I_27(n25_14,IN_5_1_l_14);
nor I_28(n26_14,IN_10_1_l_14,n20_14);
nand I_29(n27_14,IN_4_1_l_14,n28_14);
not I_30(n28_14,G15_1_l_14);
DFFARX1 I_31(n4_1_r_5,blif_clk_net_1_r_5,n5_5,G42_1_r_5,);
nor I_32(n_572_1_r_5,n21_5,n22_5);
nand I_33(n_573_1_r_5,n13_5,n16_5);
nor I_34(n_549_1_r_5,n21_5,n17_5);
nand I_35(n_569_1_r_5,n13_5,n15_5);
nor I_36(n_452_1_r_5,n22_5,n_42_2_l_5);
DFFARX1 I_37(G199_2_l_5,blif_clk_net_1_r_5,n5_5,ACVQN2_3_r_5,);
nor I_38(n_266_and_0_3_r_5,n11_5,n16_5);
DFFARX1 I_39(n_42_2_l_5,blif_clk_net_1_r_5,n5_5,ACVQN1_5_r_5,);
not I_40(P6_5_r_5,P6_5_r_internal_5);
and I_41(N3_2_l_5,n19_5,n_569_1_r_14);
not I_42(n5_5,blif_reset_net_1_r_5);
DFFARX1 I_43(N3_2_l_5,blif_clk_net_1_r_5,n5_5,G199_2_l_5,);
DFFARX1 I_44(G42_1_r_14,blif_clk_net_1_r_5,n5_5,ACVQN2_3_l_5,);
not I_45(n13_5,ACVQN2_3_l_5);
DFFARX1 I_46(ACVQN1_5_r_14,blif_clk_net_1_r_5,n5_5,ACVQN1_3_l_5,);
and I_47(N1_4_l_5,n20_5,n_42_2_r_14);
DFFARX1 I_48(N1_4_l_5,blif_clk_net_1_r_5,n5_5,n21_5,);
not I_49(n15_5,n21_5);
DFFARX1 I_50(G199_2_r_14,blif_clk_net_1_r_5,n5_5,n22_5,);
nor I_51(n4_1_r_5,G199_2_l_5,n22_5);
DFFARX1 I_52(ACVQN2_3_l_5,blif_clk_net_1_r_5,n5_5,n11_internal_5,);
not I_53(n11_5,n11_internal_5);
nor I_54(n_42_2_l_5,n_572_1_r_14,n_573_1_r_14);
not I_55(n1_5,n18_5);
DFFARX1 I_56(n1_5,blif_clk_net_1_r_5,n5_5,P6_5_r_internal_5,);
not I_57(n16_5,n_42_2_l_5);
nor I_58(n17_5,n22_5,n18_5);
nand I_59(n18_5,ACVQN1_3_l_5,n_549_1_r_14);
nand I_60(n19_5,n_572_1_r_14,n_573_1_r_14);
nand I_61(n20_5,G42_1_r_14,P6_5_r_14);
endmodule


