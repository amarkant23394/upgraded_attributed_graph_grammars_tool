module test_final(IN_1_2_l_0,IN_2_2_l_0,IN_3_2_l_0,IN_4_2_l_0,IN_5_2_l_0,IN_1_4_l_0,IN_2_4_l_0,IN_3_4_l_0,IN_4_4_l_0,IN_5_4_l_0,IN_1_9_l_0,IN_2_9_l_0,IN_3_9_l_0,IN_4_9_l_0,IN_5_9_l_0,blif_clk_net_7_r_3,blif_reset_net_7_r_3,N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6134_9_r_3);
input IN_1_2_l_0,IN_2_2_l_0,IN_3_2_l_0,IN_4_2_l_0,IN_5_2_l_0,IN_1_4_l_0,IN_2_4_l_0,IN_3_4_l_0,IN_4_4_l_0,IN_5_4_l_0,IN_1_9_l_0,IN_2_9_l_0,IN_3_9_l_0,IN_4_9_l_0,IN_5_9_l_0,blif_clk_net_7_r_3,blif_reset_net_7_r_3;
output N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6134_9_r_3;
wire N1371_0_r_0,N1508_0_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_102_5_r_0,n_547_5_r_0,G42_7_r_0,n_572_7_r_0,n_573_7_r_0,n_549_7_r_0,n_569_7_r_0,n_452_7_r_0,n_431_5_r_0,n4_7_r_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0,n37_0,n38_0,n39_0,n40_0,n41_0,n42_0,n43_0,n44_0,n45_0,n_572_7_r_3,N6147_9_r_3,I_BUFF_1_9_r_3,n4_7_r_3,n10_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3,n40_3,n41_3,n42_3,n43_3,n44_3,n45_3,n46_3,n47_3,n48_3,n49_3,n50_3,n51_3;
nor I_0(N1371_0_r_0,n_102_5_r_0,n29_0);
nor I_1(N1508_0_r_0,n_102_5_r_0,n_452_7_r_0);
or I_2(n_429_or_0_5_r_0,IN_1_9_l_0,n38_0);
DFFARX1 I_3(n_431_5_r_0,blif_clk_net_7_r_3,n10_3,G78_5_r_0,);
nand I_4(n_576_5_r_0,IN_1_9_l_0,n26_0);
not I_5(n_102_5_r_0,n27_0);
nand I_6(n_547_5_r_0,n30_0,n34_0);
DFFARX1 I_7(n4_7_r_0,blif_clk_net_7_r_3,n10_3,G42_7_r_0,);
nor I_8(n_572_7_r_0,IN_1_9_l_0,n31_0);
or I_9(n_573_7_r_0,n29_0,n30_0);
nor I_10(n_549_7_r_0,n29_0,n33_0);
nand I_11(n_569_7_r_0,n28_0,n32_0);
nor I_12(n_452_7_r_0,n30_0,n31_0);
nand I_13(n_431_5_r_0,n_102_5_r_0,n35_0);
nor I_14(n4_7_r_0,n31_0,n37_0);
nor I_15(n26_0,n27_0,n28_0);
nor I_16(n27_0,n28_0,n44_0);
nand I_17(n28_0,IN_1_4_l_0,IN_2_4_l_0);
not I_18(n29_0,n32_0);
nor I_19(n30_0,IN_5_9_l_0,n39_0);
not I_20(n31_0,n38_0);
nand I_21(n32_0,n41_0,n42_0);
nor I_22(n33_0,IN_1_9_l_0,n_102_5_r_0);
nor I_23(n34_0,IN_1_9_l_0,n27_0);
nand I_24(n35_0,n29_0,n36_0);
nor I_25(n36_0,n37_0,n38_0);
not I_26(n37_0,n28_0);
nand I_27(n38_0,IN_2_9_l_0,n40_0);
nor I_28(n39_0,IN_3_9_l_0,IN_4_9_l_0);
or I_29(n40_0,IN_3_9_l_0,IN_4_9_l_0);
nor I_30(n41_0,IN_1_2_l_0,IN_2_2_l_0);
or I_31(n42_0,IN_5_2_l_0,n43_0);
nor I_32(n43_0,IN_3_2_l_0,IN_4_2_l_0);
nor I_33(n44_0,IN_5_4_l_0,n45_0);
and I_34(n45_0,IN_3_4_l_0,IN_4_4_l_0);
not I_35(N1372_1_r_3,n40_3);
nor I_36(N1508_1_r_3,N6147_9_r_3,n40_3);
nor I_37(N1507_6_r_3,n31_3,n42_3);
nor I_38(N1508_6_r_3,n30_3,n38_3);
DFFARX1 I_39(n4_7_r_3,blif_clk_net_7_r_3,n10_3,G42_7_r_3,);
nor I_40(n_572_7_r_3,I_BUFF_1_9_r_3,n35_3);
nand I_41(n_573_7_r_3,n30_3,n31_3);
nor I_42(n_549_7_r_3,N6147_9_r_3,n33_3);
nand I_43(n_569_7_r_3,n30_3,n32_3);
nor I_44(n_452_7_r_3,n35_3,n_569_7_r_0);
not I_45(N6147_9_r_3,n32_3);
nor I_46(N6134_9_r_3,n36_3,n37_3);
not I_47(I_BUFF_1_9_r_3,n45_3);
nor I_48(n4_7_r_3,I_BUFF_1_9_r_3,n_569_7_r_0);
not I_49(n10_3,blif_reset_net_7_r_3);
not I_50(n30_3,n39_3);
not I_51(n31_3,n35_3);
nand I_52(n32_3,n41_3,n_429_or_0_5_r_0);
nor I_53(n33_3,I_BUFF_1_9_r_3,n34_3);
nand I_54(n34_3,n46_3,G78_5_r_0);
nor I_55(n35_3,n43_3,n44_3);
not I_56(n36_3,n34_3);
nor I_57(n37_3,N6147_9_r_3,n_569_7_r_0);
or I_58(n38_3,n_572_7_r_3,n34_3);
nor I_59(n39_3,n44_3,n_549_7_r_0);
nand I_60(n40_3,n39_3,n_569_7_r_0);
nand I_61(n41_3,G42_7_r_0,N1371_0_r_0);
nor I_62(n42_3,n34_3,n45_3);
not I_63(n43_3,n_573_7_r_0);
nor I_64(n44_3,n_547_5_r_0,G78_5_r_0);
nand I_65(n45_3,n49_3,n50_3);
and I_66(n46_3,n47_3,n_576_5_r_0);
nand I_67(n47_3,n41_3,n48_3);
not I_68(n48_3,n_429_or_0_5_r_0);
nor I_69(n49_3,N1371_0_r_0,n_572_7_r_0);
or I_70(n50_3,n51_3,N1508_0_r_0);
nor I_71(n51_3,N1508_0_r_0,n_429_or_0_5_r_0);
endmodule


