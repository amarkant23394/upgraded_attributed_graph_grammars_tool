module test_final(IN_1_2_l_6,IN_2_2_l_6,G1_3_l_6,G2_3_l_6,IN_2_3_l_6,IN_4_3_l_6,IN_5_3_l_6,IN_7_3_l_6,IN_8_3_l_6,IN_10_3_l_6,IN_11_3_l_6,blif_clk_net_1_r_9,blif_reset_net_1_r_9,G199_1_r_9,G214_1_r_9,ACVQN1_2_r_9,P6_2_r_9,n_429_or_0_3_r_9,G78_3_r_9,n_576_3_r_9,n_102_3_r_9,n_547_3_r_9,n_42_5_r_9,G199_5_r_9);
input IN_1_2_l_6,IN_2_2_l_6,G1_3_l_6,G2_3_l_6,IN_2_3_l_6,IN_4_3_l_6,IN_5_3_l_6,IN_7_3_l_6,IN_8_3_l_6,IN_10_3_l_6,IN_11_3_l_6,blif_clk_net_1_r_9,blif_reset_net_1_r_9;
output G199_1_r_9,G214_1_r_9,ACVQN1_2_r_9,P6_2_r_9,n_429_or_0_3_r_9,G78_3_r_9,n_576_3_r_9,n_102_3_r_9,n_547_3_r_9,n_42_5_r_9,G199_5_r_9;
wire ACVQN2_0_r_6,n_266_and_0_0_r_6,ACVQN1_2_r_6,P6_2_r_6,n_429_or_0_3_r_6,G78_3_r_6,n_576_3_r_6,n_102_3_r_6,n_547_3_r_6,n_42_5_r_6,G199_5_r_6,ACVQN1_2_l_6,P6_2_l_6,P6_internal_2_l_6,n_429_or_0_3_l_6,n12_3_l_6,n_431_3_l_6,G78_3_l_6,n_576_3_l_6,n11_3_l_6,n_102_3_l_6,n_547_3_l_6,n13_3_l_6,n14_3_l_6,n15_3_l_6,n16_3_l_6,ACVQN1_0_r_6,P6_internal_2_r_6,n12_3_r_6,n_431_3_r_6,n11_3_r_6,n13_3_r_6,n14_3_r_6,n15_3_r_6,n16_3_r_6,N3_5_r_6,n3_5_r_6,n1_1_r_9,ACVQN2_0_l_9,n_266_and_0_0_l_9,ACVQN1_0_l_9,n4_4_l_9,G42_4_l_9,n_87_4_l_9,n_572_4_l_9,n_573_4_l_9,n_549_4_l_9,n7_4_l_9,n_569_4_l_9,n_452_4_l_9,N1_1_r_9,n3_1_r_9,P6_internal_2_r_9,n12_3_r_9,n_431_3_r_9,n11_3_r_9,n13_3_r_9,n14_3_r_9,n15_3_r_9,n16_3_r_9,N3_5_r_9,n3_5_r_9;
DFFARX1 I_0(G78_3_l_6,blif_clk_net_1_r_9,n1_1_r_9,ACVQN2_0_r_6,);
and I_1(n_266_and_0_0_r_6,n_429_or_0_3_l_6,ACVQN1_0_r_6);
DFFARX1 I_2(G78_3_l_6,blif_clk_net_1_r_9,n1_1_r_9,ACVQN1_2_r_6,);
not I_3(P6_2_r_6,P6_internal_2_r_6);
nand I_4(n_429_or_0_3_r_6,n_102_3_l_6,n12_3_r_6);
DFFARX1 I_5(n_431_3_r_6,blif_clk_net_1_r_9,n1_1_r_9,G78_3_r_6,);
nand I_6(n_576_3_r_6,P6_2_l_6,n11_3_r_6);
not I_7(n_102_3_r_6,ACVQN1_2_l_6);
nand I_8(n_547_3_r_6,n_576_3_l_6,n13_3_r_6);
nor I_9(n_42_5_r_6,ACVQN1_2_l_6,n_429_or_0_3_l_6);
DFFARX1 I_10(N3_5_r_6,blif_clk_net_1_r_9,n1_1_r_9,G199_5_r_6,);
DFFARX1 I_11(IN_2_2_l_6,blif_clk_net_1_r_9,n1_1_r_9,ACVQN1_2_l_6,);
not I_12(P6_2_l_6,P6_internal_2_l_6);
DFFARX1 I_13(IN_1_2_l_6,blif_clk_net_1_r_9,n1_1_r_9,P6_internal_2_l_6,);
nand I_14(n_429_or_0_3_l_6,G1_3_l_6,n12_3_l_6);
not I_15(n12_3_l_6,IN_5_3_l_6);
or I_16(n_431_3_l_6,IN_8_3_l_6,n14_3_l_6);
DFFARX1 I_17(n_431_3_l_6,blif_clk_net_1_r_9,n1_1_r_9,G78_3_l_6,);
nand I_18(n_576_3_l_6,IN_7_3_l_6,n11_3_l_6);
nor I_19(n11_3_l_6,G2_3_l_6,n12_3_l_6);
not I_20(n_102_3_l_6,G2_3_l_6);
nand I_21(n_547_3_l_6,IN_11_3_l_6,n13_3_l_6);
nor I_22(n13_3_l_6,G2_3_l_6,IN_10_3_l_6);
and I_23(n14_3_l_6,IN_2_3_l_6,n15_3_l_6);
nor I_24(n15_3_l_6,IN_4_3_l_6,n16_3_l_6);
not I_25(n16_3_l_6,G1_3_l_6);
DFFARX1 I_26(G78_3_l_6,blif_clk_net_1_r_9,n1_1_r_9,ACVQN1_0_r_6,);
DFFARX1 I_27(n_576_3_l_6,blif_clk_net_1_r_9,n1_1_r_9,P6_internal_2_r_6,);
not I_28(n12_3_r_6,P6_2_l_6);
or I_29(n_431_3_r_6,n_429_or_0_3_l_6,n14_3_r_6);
nor I_30(n11_3_r_6,ACVQN1_2_l_6,n12_3_r_6);
nor I_31(n13_3_r_6,ACVQN1_2_l_6,n_547_3_l_6);
and I_32(n14_3_r_6,ACVQN1_2_l_6,n15_3_r_6);
nor I_33(n15_3_r_6,P6_2_l_6,n16_3_r_6);
not I_34(n16_3_r_6,n_102_3_l_6);
and I_35(N3_5_r_6,n_102_3_l_6,n3_5_r_6);
nand I_36(n3_5_r_6,n_429_or_0_3_l_6,n_547_3_l_6);
DFFARX1 I_37(N1_1_r_9,blif_clk_net_1_r_9,n1_1_r_9,G199_1_r_9,);
DFFARX1 I_38(G42_4_l_9,blif_clk_net_1_r_9,n1_1_r_9,G214_1_r_9,);
DFFARX1 I_39(n_572_4_l_9,blif_clk_net_1_r_9,n1_1_r_9,ACVQN1_2_r_9,);
not I_40(P6_2_r_9,P6_internal_2_r_9);
nand I_41(n_429_or_0_3_r_9,n_572_4_l_9,n12_3_r_9);
DFFARX1 I_42(n_431_3_r_9,blif_clk_net_1_r_9,n1_1_r_9,G78_3_r_9,);
nand I_43(n_576_3_r_9,n_573_4_l_9,n11_3_r_9);
not I_44(n_102_3_r_9,n_266_and_0_0_l_9);
nand I_45(n_547_3_r_9,n_549_4_l_9,n13_3_r_9);
nor I_46(n_42_5_r_9,n_569_4_l_9,n_452_4_l_9);
DFFARX1 I_47(N3_5_r_9,blif_clk_net_1_r_9,n1_1_r_9,G199_5_r_9,);
not I_48(n1_1_r_9,blif_reset_net_1_r_9);
DFFARX1 I_49(n_429_or_0_3_r_6,blif_clk_net_1_r_9,n1_1_r_9,ACVQN2_0_l_9,);
and I_50(n_266_and_0_0_l_9,ACVQN1_0_l_9,n_102_3_r_6);
DFFARX1 I_51(P6_2_r_6,blif_clk_net_1_r_9,n1_1_r_9,ACVQN1_0_l_9,);
nor I_52(n4_4_l_9,ACVQN2_0_r_6,ACVQN1_2_r_6);
DFFARX1 I_53(n4_4_l_9,blif_clk_net_1_r_9,n1_1_r_9,G42_4_l_9,);
not I_54(n_87_4_l_9,n_266_and_0_0_r_6);
nor I_55(n_572_4_l_9,n_266_and_0_0_r_6,n_547_3_r_6);
or I_56(n_573_4_l_9,n_42_5_r_6,G199_5_r_6);
nor I_57(n_549_4_l_9,n7_4_l_9,n_576_3_r_6);
and I_58(n7_4_l_9,n_87_4_l_9,G78_3_r_6);
or I_59(n_569_4_l_9,n_576_3_r_6,n_42_5_r_6);
nor I_60(n_452_4_l_9,ACVQN1_2_r_6,G199_5_r_6);
and I_61(N1_1_r_9,n_266_and_0_0_l_9,n3_1_r_9);
nand I_62(n3_1_r_9,n_572_4_l_9,n_569_4_l_9);
DFFARX1 I_63(n_266_and_0_0_l_9,blif_clk_net_1_r_9,n1_1_r_9,P6_internal_2_r_9,);
not I_64(n12_3_r_9,G42_4_l_9);
or I_65(n_431_3_r_9,n_549_4_l_9,n14_3_r_9);
nor I_66(n11_3_r_9,ACVQN2_0_l_9,n12_3_r_9);
nor I_67(n13_3_r_9,ACVQN2_0_l_9,n_266_and_0_0_l_9);
and I_68(n14_3_r_9,n_452_4_l_9,n15_3_r_9);
nor I_69(n15_3_r_9,G42_4_l_9,n16_3_r_9);
not I_70(n16_3_r_9,n_572_4_l_9);
and I_71(N3_5_r_9,ACVQN2_0_l_9,n3_5_r_9);
nand I_72(n3_5_r_9,n_573_4_l_9,n_452_4_l_9);
endmodule


