module test_I2560(I2600,I1923,I1294,I2685,I1920,I1301,I2560);
input I2600,I1923,I1294,I2685,I1920,I1301;
output I2560;
wire I2897,I3168,I2583,I2849,I2914,I3086,I3103,I2832;
nand I_0(I2897,I2600,I1923);
or I_1(I3168,I3103,I2914);
DFFARX1 I_2(I3168,I1294,I2583,,,I2560,);
not I_3(I2583,I1301);
nor I_4(I2849,I2832,I2685);
and I_5(I2914,I2897,I2849);
DFFARX1 I_6(I1920,I1294,I2583,,,I3086,);
not I_7(I3103,I3086);
DFFARX1 I_8(I1294,I2583,,,I2832,);
endmodule


