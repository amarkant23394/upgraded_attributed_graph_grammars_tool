module test_I5731(I2167,I2173,I1477,I1470,I4578,I5731);
input I2167,I2173,I1477,I1470,I4578;
output I5731;
wire I4629,I5864,I5751,I4595,I4536,I4515,I4527,I4544,I4869,I5881,I5915;
nor I_0(I4629,I2167,I2173);
nor I_1(I5864,I4536,I4515);
not I_2(I5751,I1477);
DFFARX1 I_3(I4578,I1470,I4544,,,I4595,);
nor I_4(I4536,I4869,I4595);
not I_5(I4515,I4629);
or I_6(I4527,I4629,I4595);
not I_7(I4544,I1477);
DFFARX1 I_8(I1470,I4544,,,I4869,);
not I_9(I5881,I5864);
DFFARX1 I_10(I4527,I1470,I5751,,,I5915,);
nand I_11(I5731,I5915,I5881);
endmodule


