module test_I5740(I4515,I1477,I1470,I4530,I5740);
input I4515,I1477,I1470,I4530;
output I5740;
wire I5751,I4595,I4524,I5785,I4742,I5802,I5768;
not I_0(I5751,I1477);
DFFARX1 I_1(I1470,,,I4595,);
nor I_2(I4524,I4742,I4595);
and I_3(I5785,I5768,I4524);
DFFARX1 I_4(I1470,,,I4742,);
DFFARX1 I_5(I5785,I1470,I5751,,,I5802,);
nand I_6(I5768,I4530,I4515);
not I_7(I5740,I5802);
endmodule


