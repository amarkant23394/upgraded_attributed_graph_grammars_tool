module test_I2362(I1477,I1470,I1375,I2362);
input I1477,I1470,I1375;
output I2362;
wire I2181,I2345;
not I_0(I2362,I2345);
not I_1(I2181,I1477);
DFFARX1 I_2(I1375,I1470,I2181,,,I2345,);
endmodule


