module test_I11847(I9320,I8830,I1477,I9049,I6881,I9413,I1470,I8879,I11847);
input I9320,I8830,I1477,I9049,I6881,I9413,I1470,I8879;
output I11847;
wire I9179,I8854,I11830,I11395,I8862,I8848,I9083,I11378,I8851,I9066,I11813,I11327,I11310;
DFFARX1 I_0(I1470,I8862,,,I9179,);
nor I_1(I8854,I9179,I9320);
not I_2(I11830,I11813);
nand I_3(I11395,I11378,I8851);
nand I_4(I11847,I11830,I11395);
not I_5(I8862,I1477);
nor I_6(I8848,I9083,I9413);
nand I_7(I9083,I8879,I6881);
nor I_8(I11378,I11327,I8848);
or I_9(I8851,I9083,I9066);
DFFARX1 I_10(I9049,I1470,I8862,,,I9066,);
DFFARX1 I_11(I8854,I1470,I11310,,,I11813,);
not I_12(I11327,I8830);
not I_13(I11310,I1477);
endmodule


