module test_final(IN_1_1_l,IN_2_1_l,IN_3_1_l,G18_7_l,G15_7_l,IN_1_7_l,IN_4_7_l,IN_5_7_l,IN_7_7_l,IN_9_7_l,IN_10_7_l,IN_1_10_l,IN_2_10_l,IN_3_10_l,IN_4_10_l,blif_clk_net_5_r,blif_reset_net_5_r,N6147_2_r,N1372_4_r,N1508_4_r,n_429_or_0_5_r,G78_5_r,n_576_5_r,n_102_5_r,n_547_5_r,n_42_8_r,G199_8_r,N6147_9_r,N6134_9_r,I_BUFF_1_9_r);
input IN_1_1_l,IN_2_1_l,IN_3_1_l,G18_7_l,G15_7_l,IN_1_7_l,IN_4_7_l,IN_5_7_l,IN_7_7_l,IN_9_7_l,IN_10_7_l,IN_1_10_l,IN_2_10_l,IN_3_10_l,IN_4_10_l,blif_clk_net_5_r,blif_reset_net_5_r;
output N6147_2_r,N1372_4_r,N1508_4_r,n_429_or_0_5_r,G78_5_r,n_576_5_r,n_102_5_r,n_547_5_r,n_42_8_r,G199_8_r,N6147_9_r,N6134_9_r,I_BUFF_1_9_r;
wire N1372_1_l,N1508_1_l,n4_1_l,G42_7_l,n_87_7_l,n_572_7_l,n_573_7_l,n_549_7_l,n_569_7_l,n_452_7_l,n4_7_l,n7_7_l,N1372_10_l,N1508_10_l,n5_10_l,n6_10_l,n5_2_r,n6_2_r,N6138_2_r,n7_2_r,n6_4_r,n7_4_r,n8_4_r,n_431_5_r,n2_5_r,n11_5_r,n12_5_r,n13_5_r,n14_5_r,n15_5_r,n16_5_r,N3_8_r,n3_8_r,N6150_9_r,n3_9_r;
not I_0(N1372_1_l,n4_1_l);
nor I_1(N1508_1_l,IN_3_1_l,n4_1_l);
nand I_2(n4_1_l,IN_1_1_l,IN_2_1_l);
DFFARX1 I_3(n4_7_l,blif_clk_net_5_r,n2_5_r,G42_7_l,);
not I_4(n_87_7_l,G15_7_l);
nor I_5(n_572_7_l,G15_7_l,IN_7_7_l);
or I_6(n_573_7_l,IN_5_7_l,IN_9_7_l);
nor I_7(n_549_7_l,IN_10_7_l,n7_7_l);
or I_8(n_569_7_l,IN_9_7_l,IN_10_7_l);
nor I_9(n_452_7_l,G18_7_l,IN_5_7_l);
nor I_10(n4_7_l,G18_7_l,IN_1_7_l);
and I_11(n7_7_l,IN_4_7_l,n_87_7_l);
not I_12(N1372_10_l,n6_10_l);
nor I_13(N1508_10_l,n5_10_l,n6_10_l);
nor I_14(n5_10_l,IN_3_10_l,IN_4_10_l);
nand I_15(n6_10_l,IN_1_10_l,IN_2_10_l);
nor I_16(N6147_2_r,n5_2_r,n6_2_r);
nor I_17(n5_2_r,n7_2_r,n_569_7_l);
not I_18(n6_2_r,N6138_2_r);
nor I_19(N6138_2_r,N1508_10_l,n_573_7_l);
nor I_20(n7_2_r,N1372_10_l,N1508_1_l);
not I_21(N1372_4_r,n7_4_r);
nor I_22(N1508_4_r,n6_4_r,n7_4_r);
nor I_23(n6_4_r,n8_4_r,n_569_7_l);
nand I_24(n7_4_r,n_572_7_l,n_549_7_l);
and I_25(n8_4_r,N1372_1_l,N1372_10_l);
nand I_26(n_429_or_0_5_r,n12_5_r,G42_7_l);
DFFARX1 I_27(n_431_5_r,blif_clk_net_5_r,n2_5_r,G78_5_r,);
nand I_28(n_576_5_r,n11_5_r,N1372_1_l);
not I_29(n_102_5_r,n_573_7_l);
nand I_30(n_547_5_r,n13_5_r,n_572_7_l);
or I_31(n_431_5_r,n14_5_r,N1508_1_l);
not I_32(n2_5_r,blif_reset_net_5_r);
nor I_33(n11_5_r,n12_5_r,n_573_7_l);
not I_34(n12_5_r,n_569_7_l);
nor I_35(n13_5_r,n_573_7_l,n_452_7_l);
and I_36(n14_5_r,n15_5_r,n_549_7_l);
nor I_37(n15_5_r,n16_5_r,n_549_7_l);
not I_38(n16_5_r,G42_7_l);
nor I_39(n_42_8_r,n_572_7_l,n_452_7_l);
DFFARX1 I_40(N3_8_r,blif_clk_net_5_r,n2_5_r,G199_8_r,);
and I_41(N3_8_r,n3_8_r,G42_7_l);
nand I_42(n3_8_r,N1508_1_l,n_452_7_l);
not I_43(N6150_9_r,n_452_7_l);
nor I_44(N6147_9_r,N6150_9_r,n3_9_r);
nor I_45(N6134_9_r,n3_9_r,N1372_1_l);
nor I_46(n3_9_r,G42_7_l,N1508_10_l);
buf I_47(I_BUFF_1_9_r,n_573_7_l);
endmodule


