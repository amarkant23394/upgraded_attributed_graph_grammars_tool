module test_final(IN_1_2_l_0,IN_2_2_l_0,IN_3_2_l_0,IN_4_2_l_0,IN_5_2_l_0,IN_1_4_l_0,IN_2_4_l_0,IN_3_4_l_0,IN_4_4_l_0,IN_5_4_l_0,IN_1_9_l_0,IN_2_9_l_0,IN_3_9_l_0,IN_4_9_l_0,IN_5_9_l_0,blif_clk_net_5_r_11,blif_reset_net_5_r_11,N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1508_10_r_11);
input IN_1_2_l_0,IN_2_2_l_0,IN_3_2_l_0,IN_4_2_l_0,IN_5_2_l_0,IN_1_4_l_0,IN_2_4_l_0,IN_3_4_l_0,IN_4_4_l_0,IN_5_4_l_0,IN_1_9_l_0,IN_2_9_l_0,IN_3_9_l_0,IN_4_9_l_0,IN_5_9_l_0,blif_clk_net_5_r_11,blif_reset_net_5_r_11;
output N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1508_10_r_11;
wire N1371_0_r_0,N1508_0_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_102_5_r_0,n_547_5_r_0,G42_7_r_0,n_572_7_r_0,n_573_7_r_0,n_549_7_r_0,n_569_7_r_0,n_452_7_r_0,n_431_5_r_0,n4_7_r_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0,n37_0,n38_0,n39_0,n40_0,n41_0,n42_0,n43_0,n44_0,n45_0,n_102_5_r_11,N1372_10_r_11,n_431_5_r_11,n9_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11,n43_11,n44_11,n45_11,n46_11,n47_11,n48_11,n49_11,n50_11,n51_11,n52_11,n53_11,n54_11,n55_11,n56_11,n57_11,n58_11,n59_11,n60_11,n61_11,n62_11,n63_11;
nor I_0(N1371_0_r_0,n_102_5_r_0,n29_0);
nor I_1(N1508_0_r_0,n_102_5_r_0,n_452_7_r_0);
or I_2(n_429_or_0_5_r_0,IN_1_9_l_0,n38_0);
DFFARX1 I_3(n_431_5_r_0,blif_clk_net_5_r_11,n9_11,G78_5_r_0,);
nand I_4(n_576_5_r_0,IN_1_9_l_0,n26_0);
not I_5(n_102_5_r_0,n27_0);
nand I_6(n_547_5_r_0,n30_0,n34_0);
DFFARX1 I_7(n4_7_r_0,blif_clk_net_5_r_11,n9_11,G42_7_r_0,);
nor I_8(n_572_7_r_0,IN_1_9_l_0,n31_0);
or I_9(n_573_7_r_0,n29_0,n30_0);
nor I_10(n_549_7_r_0,n29_0,n33_0);
nand I_11(n_569_7_r_0,n28_0,n32_0);
nor I_12(n_452_7_r_0,n30_0,n31_0);
nand I_13(n_431_5_r_0,n_102_5_r_0,n35_0);
nor I_14(n4_7_r_0,n31_0,n37_0);
nor I_15(n26_0,n27_0,n28_0);
nor I_16(n27_0,n28_0,n44_0);
nand I_17(n28_0,IN_1_4_l_0,IN_2_4_l_0);
not I_18(n29_0,n32_0);
nor I_19(n30_0,IN_5_9_l_0,n39_0);
not I_20(n31_0,n38_0);
nand I_21(n32_0,n41_0,n42_0);
nor I_22(n33_0,IN_1_9_l_0,n_102_5_r_0);
nor I_23(n34_0,IN_1_9_l_0,n27_0);
nand I_24(n35_0,n29_0,n36_0);
nor I_25(n36_0,n37_0,n38_0);
not I_26(n37_0,n28_0);
nand I_27(n38_0,IN_2_9_l_0,n40_0);
nor I_28(n39_0,IN_3_9_l_0,IN_4_9_l_0);
or I_29(n40_0,IN_3_9_l_0,IN_4_9_l_0);
nor I_30(n41_0,IN_1_2_l_0,IN_2_2_l_0);
or I_31(n42_0,IN_5_2_l_0,n43_0);
nor I_32(n43_0,IN_3_2_l_0,IN_4_2_l_0);
nor I_33(n44_0,IN_5_4_l_0,n45_0);
and I_34(n45_0,IN_3_4_l_0,IN_4_4_l_0);
not I_35(N1372_1_r_11,n53_11);
nor I_36(N1508_1_r_11,n39_11,n53_11);
nor I_37(N6147_2_r_11,n48_11,n49_11);
nor I_38(N6147_3_r_11,n44_11,n45_11);
nand I_39(n_429_or_0_5_r_11,n42_11,n43_11);
DFFARX1 I_40(n_431_5_r_11,blif_clk_net_5_r_11,n9_11,G78_5_r_11,);
nand I_41(n_576_5_r_11,n_102_5_r_11,N1372_10_r_11);
not I_42(n_102_5_r_11,n39_11);
nand I_43(n_547_5_r_11,n36_11,n37_11);
nor I_44(N1507_6_r_11,n52_11,n57_11);
nor I_45(N1508_6_r_11,n46_11,n51_11);
nor I_46(N1372_10_r_11,n43_11,n47_11);
nor I_47(N1508_10_r_11,n55_11,n56_11);
nand I_48(n_431_5_r_11,n40_11,n41_11);
not I_49(n9_11,blif_reset_net_5_r_11);
nor I_50(n36_11,n38_11,n39_11);
not I_51(n37_11,n40_11);
nor I_52(n38_11,n60_11,G42_7_r_0);
nor I_53(n39_11,n54_11,n_547_5_r_0);
nand I_54(n40_11,N1371_0_r_0,N1508_0_r_0);
nand I_55(n41_11,n_102_5_r_11,n42_11);
and I_56(n42_11,n58_11,G78_5_r_0);
not I_57(n43_11,n44_11);
nor I_58(n44_11,n40_11,n_572_7_r_0);
nand I_59(n45_11,n46_11,n47_11);
not I_60(n46_11,n38_11);
nand I_61(n47_11,n59_11,n62_11);
and I_62(n48_11,n37_11,n47_11);
or I_63(n49_11,n44_11,n50_11);
nor I_64(n50_11,n60_11,n61_11);
or I_65(n51_11,n_102_5_r_11,n52_11);
nor I_66(n52_11,n42_11,n57_11);
nand I_67(n53_11,n37_11,n50_11);
or I_68(n54_11,n_429_or_0_5_r_0,n_573_7_r_0);
nor I_69(n55_11,n38_11,n42_11);
not I_70(n56_11,N1372_10_r_11);
and I_71(n57_11,n38_11,n50_11);
and I_72(n58_11,n59_11,n_429_or_0_5_r_0);
or I_73(n59_11,n63_11,n_576_5_r_0);
not I_74(n60_11,N1371_0_r_0);
nor I_75(n61_11,n_569_7_r_0,G78_5_r_0);
nand I_76(n62_11,N1508_0_r_0,n_549_7_r_0);
and I_77(n63_11,N1508_0_r_0,n_549_7_r_0);
endmodule


