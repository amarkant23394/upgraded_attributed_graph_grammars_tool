module test_final(IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_6_2_l_6,IN_1_3_l_6,IN_2_3_l_6,IN_4_3_l_6,IN_1_4_l_6,IN_2_4_l_6,IN_3_4_l_6,IN_6_4_l_6,blif_clk_net_1_r_9,blif_reset_net_1_r_9,G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9);
input IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_6_2_l_6,IN_1_3_l_6,IN_2_3_l_6,IN_4_3_l_6,IN_1_4_l_6,IN_2_4_l_6,IN_3_4_l_6,IN_6_4_l_6,blif_clk_net_1_r_9,blif_reset_net_1_r_9;
output G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9;
wire G42_1_r_6,n_572_1_r_6,n_573_1_r_6,n_549_1_r_6,n_569_1_r_6,n_452_1_r_6,G199_4_r_6,G214_4_r_6,ACVQN1_5_r_6,P6_5_r_6,N3_2_l_6,n27_6,n17_6,n28_6,n26_6,N1_4_l_6,n29_6,n18_6,G214_4_l_6,n12_6,n4_1_r_6,N1_4_r_6,n_42_2_l_6,P6_5_r_internal_6,n19_6,n20_6,n21_6,n22_6,n23_6,n24_6,n25_6,n_452_1_r_9,N3_2_l_9,n5_9,n27_9,n16_9,n26_9,n15_9,n29_internal_9,n29_9,N1_4_l_9,n25_9,n28_internal_9,n28_9,n4_1_r_9,N3_2_r_9,N1_4_r_9,n_42_2_l_9,n17_9,n18_9,n19_9,n20_9,n21_9,n22_9,n23_9,n24_9;
DFFARX1 I_0(n4_1_r_6,blif_clk_net_1_r_9,n5_9,G42_1_r_6,);
nor I_1(n_572_1_r_6,n27_6,n28_6);
nand I_2(n_573_1_r_6,n18_6,n19_6);
nor I_3(n_549_1_r_6,n_42_2_l_6,n21_6);
nand I_4(n_569_1_r_6,n19_6,n20_6);
nor I_5(n_452_1_r_6,n28_6,n29_6);
DFFARX1 I_6(N1_4_r_6,blif_clk_net_1_r_9,n5_9,G199_4_r_6,);
DFFARX1 I_7(n_42_2_l_6,blif_clk_net_1_r_9,n5_9,G214_4_r_6,);
DFFARX1 I_8(n_42_2_l_6,blif_clk_net_1_r_9,n5_9,ACVQN1_5_r_6,);
not I_9(P6_5_r_6,P6_5_r_internal_6);
and I_10(N3_2_l_6,IN_6_2_l_6,n23_6);
DFFARX1 I_11(N3_2_l_6,blif_clk_net_1_r_9,n5_9,n27_6,);
not I_12(n17_6,n27_6);
DFFARX1 I_13(IN_1_3_l_6,blif_clk_net_1_r_9,n5_9,n28_6,);
DFFARX1 I_14(IN_2_3_l_6,blif_clk_net_1_r_9,n5_9,n26_6,);
and I_15(N1_4_l_6,IN_6_4_l_6,n25_6);
DFFARX1 I_16(N1_4_l_6,blif_clk_net_1_r_9,n5_9,n29_6,);
not I_17(n18_6,n29_6);
DFFARX1 I_18(IN_3_4_l_6,blif_clk_net_1_r_9,n5_9,G214_4_l_6,);
not I_19(n12_6,G214_4_l_6);
nor I_20(n4_1_r_6,n28_6,n22_6);
nor I_21(N1_4_r_6,n12_6,n24_6);
nor I_22(n_42_2_l_6,IN_1_2_l_6,IN_3_2_l_6);
DFFARX1 I_23(G214_4_l_6,blif_clk_net_1_r_9,n5_9,P6_5_r_internal_6,);
nand I_24(n19_6,IN_4_3_l_6,n26_6);
not I_25(n20_6,n_42_2_l_6);
nor I_26(n21_6,n17_6,n28_6);
and I_27(n22_6,IN_4_3_l_6,n26_6);
nand I_28(n23_6,IN_2_2_l_6,IN_3_2_l_6);
nor I_29(n24_6,n17_6,n18_6);
nand I_30(n25_6,IN_1_4_l_6,IN_2_4_l_6);
DFFARX1 I_31(n4_1_r_9,blif_clk_net_1_r_9,n5_9,G42_1_r_9,);
nor I_32(n_572_1_r_9,n27_9,n_42_2_l_9);
or I_33(n_573_1_r_9,n25_9,n_42_2_l_9);
nand I_34(n_549_1_r_9,n17_9,n18_9);
or I_35(n_569_1_r_9,n26_9,n_42_2_l_9);
nor I_36(n_452_1_r_9,n26_9,n25_9);
nor I_37(n_42_2_r_9,n25_9,n19_9);
DFFARX1 I_38(N3_2_r_9,blif_clk_net_1_r_9,n5_9,G199_2_r_9,);
DFFARX1 I_39(N1_4_r_9,blif_clk_net_1_r_9,n5_9,G199_4_r_9,);
DFFARX1 I_40(n_42_2_l_9,blif_clk_net_1_r_9,n5_9,G214_4_r_9,);
and I_41(N3_2_l_9,n22_9,ACVQN1_5_r_6);
not I_42(n5_9,blif_reset_net_1_r_9);
DFFARX1 I_43(N3_2_l_9,blif_clk_net_1_r_9,n5_9,n27_9,);
not I_44(n16_9,n27_9);
DFFARX1 I_45(G42_1_r_6,blif_clk_net_1_r_9,n5_9,n26_9,);
not I_46(n15_9,n26_9);
DFFARX1 I_47(n_573_1_r_6,blif_clk_net_1_r_9,n5_9,n29_internal_9,);
not I_48(n29_9,n29_internal_9);
and I_49(N1_4_l_9,n24_9,n_549_1_r_6);
DFFARX1 I_50(N1_4_l_9,blif_clk_net_1_r_9,n5_9,n25_9,);
DFFARX1 I_51(G214_4_r_6,blif_clk_net_1_r_9,n5_9,n28_internal_9,);
not I_52(n28_9,n28_internal_9);
nor I_53(n4_1_r_9,n27_9,n26_9);
nor I_54(N3_2_r_9,n15_9,n21_9);
nor I_55(N1_4_r_9,n16_9,n21_9);
nor I_56(n_42_2_l_9,n_572_1_r_6,P6_5_r_6);
not I_57(n17_9,n_452_1_r_9);
nand I_58(n18_9,n27_9,n15_9);
nor I_59(n19_9,n29_9,n20_9);
not I_60(n20_9,n_569_1_r_6);
and I_61(n21_9,n23_9,n_569_1_r_6);
nand I_62(n22_9,n_572_1_r_6,n_452_1_r_6);
nor I_63(n23_9,n29_9,n28_9);
nand I_64(n24_9,G199_4_r_6,G42_1_r_6);
endmodule


