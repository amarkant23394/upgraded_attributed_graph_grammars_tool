module test_I13040(I9477,I9465,I1477,I1470,I13040);
input I9477,I9465,I1477,I1470;
output I13040;
wire I12619,I10715,I13023,I10647,I10766,I9468,I12735,I10636,I10630,I11009,I10732;
nand I_0(I13040,I13023,I12735);
not I_1(I12619,I1477);
nor I_2(I10715,I9477);
DFFARX1 I_3(I10636,I1470,I12619,,,I13023,);
not I_4(I10647,I1477);
not I_5(I10766,I9477);
DFFARX1 I_6(I1470,,,I9468,);
DFFARX1 I_7(I10630,I1470,I12619,,,I12735,);
nor I_8(I10636,I10732,I10766);
not I_9(I10630,I11009);
DFFARX1 I_10(I9468,I1470,I10647,,,I11009,);
nand I_11(I10732,I10715,I9465);
endmodule


