module test_I14933(I12718,I1477,I1470,I15194,I12964,I14933);
input I12718,I1477,I1470,I15194,I12964;
output I14933;
wire I14982,I12596,I15276,I15293,I12599,I15310,I15211,I14965;
DFFARX1 I_0(I15310,I1470,I14965,,,I14933,);
not I_1(I14982,I12596);
DFFARX1 I_2(I1470,,,I12596,);
nand I_3(I15276,I14982,I12599);
nand I_4(I15293,I15276,I15211);
nand I_5(I12599,I12718,I12964);
and I_6(I15310,I15276,I15293);
DFFARX1 I_7(I15194,I1470,I14965,,,I15211,);
not I_8(I14965,I1477);
endmodule


