module Benchmark_testing100(I1579,I1587,I1595,I1603,I1611,I1619,I1627,I1635,I1643,I1651,I1659,I1667,I1675,I1683,I1691,I1698,I1705,I3799,I3814,I3802,I3817,I3808,I3829,I3805,I3826,I3820,I3811,I3823);
input I1579,I1587,I1595,I1603,I1611,I1619,I1627,I1635,I1643,I1651,I1659,I1667,I1675,I1683,I1691,I1698,I1705;
output I3799,I3814,I3802,I3817,I3808,I3829,I3805,I3826,I3820,I3811,I3823;
wire I1579,I1587,I1595,I1603,I1611,I1619,I1627,I1635,I1643,I1651,I1659,I1667,I1675,I1683,I1691,I1698,I1705,I1743,I1760,I1777,I1794,I1811,I1828,I1845,I1723,I1876,I1708,I1732,I1921,I1938,I1955,I1972,I1989,I1711,I2020,I1729,I2051,I2068,I2085,I1735,I2116,I2133,I2150,I2167,I2184,I2201,I2218,I1717,I2249,I1720,I2280,I1726,I2311,I1714,I2369,I2386,I3037,I3034,I2403,I3040,I2429,I2437,I2454,I3046,I2471,I2488,I2505,I3043,I2522,I2539,I2349,I2570,I2587,I3064,I2604,I3052,I2621,I2638,I2655,I3055,I2672,I3049,I2689,I2706,I2340,I2737,I2754,I2771,I3058,I3061,I2337,I2802,I2819,I2361,I2850,I2867,I2884,I2343,I2915,I2352,I2946,I2358,I2355,I2991,I3008,I2346,I3072,I3089,I3106,I3123,I3140,I3157,I3174,I3191,I3222,I3239,I3256,I3273,I3290,I3307,I3324,I3355,I3372,I3417,I3434,I3451,I3468,I3485,I3502,I3533,I3550,I3567,I3584,I3601,I3632,I3663,I3708,I3725,I3756,I3773,I3837,I3854,I3871,I3888,I3905,I3922,I3939,I3956,I3987,I4004,I4021,I4038,I4055,I4072,I4089,I4120,I4137,I4182,I4199,I4216,I4233,I4250,I4267,I4298,I4315,I4332,I4349,I4366,I4397,I4428,I4473,I4490,I4521,I4538;
not I_0 (I1743,I1705);
nor I_1 (I1760,I1603,I1627);
nor I_2 (I1777,I1760,I1579);
not I_3 (I1794,I1777);
not I_4 (I1811,I1595);
nor I_5 (I1828,I1811,I1760);
not I_6 (I1845,I1828);
nand I_7 (I1723,I1794,I1845);
nand I_8 (I1876,I1777,I1611);
not I_9 (I1708,I1876);
nor I_10 (I1732,I1828,I1611);
not I_11 (I1921,I1691);
nand I_12 (I1938,I1635,I1643);
nand I_13 (I1955,I1938,I1921);
nand I_14 (I1972,I1938,I1691);
not I_15 (I1989,I1972);
nor I_16 (I1711,I1989,I1876);
nor I_17 (I2020,I1989,I1611);
nand I_18 (I1729,I1794,I1972);
and I_19 (I2051,I1955,I1667);
nand I_20 (I2068,I2051,I1587);
not I_21 (I2085,I2068);
nor I_22 (I1735,I2085,I2020);
nor I_23 (I2116,I1675,I1651);
or I_24 (I2133,I2116,I1619);
nor I_25 (I2150,I1683,I1659);
nand I_26 (I2167,I2150,I2133);
not I_27 (I2184,I2167);
nor I_28 (I2201,I2184,I1828);
or I_29 (I2218,I2201,I2068);
nor I_30 (I1717,I1794,I2218);
nor I_31 (I2249,I2184,I1611);
DFFARX1 I_32 (I2249,I1698,I1743,I1720,);
nor I_33 (I2280,I2184,I2068);
nor I_34 (I1726,I1989,I2280);
nor I_35 (I2311,I2068,I2167);
nor I_36 (I1714,I1845,I2311);
not I_37 (I2369,I1705);
nand I_38 (I2386,I3037,I3034);
and I_39 (I2403,I2386,I3040);
DFFARX1 I_40 (I2403,I1698,I2369,I2429,);
not I_41 (I2437,I2429);
nor I_42 (I2454,I3046,I3034);
not I_43 (I2471,I2454);
not I_44 (I2488,I3037);
nand I_45 (I2505,I3034,I3043);
nand I_46 (I2522,I2505,I3037);
not I_47 (I2539,I2522);
nor I_48 (I2349,I2539,I2429);
nand I_49 (I2570,I2505,I2488);
and I_50 (I2587,I2570,I3064);
nand I_51 (I2604,I2587,I3052);
and I_52 (I2621,I2604,I2522);
nor I_53 (I2638,I2604,I2522);
or I_54 (I2655,I3043,I3055);
nor I_55 (I2672,I2655,I3049);
not I_56 (I2689,I2672);
nor I_57 (I2706,I2471,I2689);
and I_58 (I2340,I2706,I2437);
nor I_59 (I2737,I2522,I2689);
nand I_60 (I2754,I2539,I2672);
nand I_61 (I2771,I3058,I3061);
nor I_62 (I2337,I2771,I2672);
nor I_63 (I2802,I2771,I2689);
not I_64 (I2819,I2802);
nor I_65 (I2361,I2621,I2819);
or I_66 (I2850,I2771,I3040);
nand I_67 (I2867,I2850,I2754);
not I_68 (I2884,I2867);
nor I_69 (I2343,I2884,I2737);
nor I_70 (I2915,I2850,I2638);
DFFARX1 I_71 (I2915,I1698,I2369,I2352,);
and I_72 (I2946,I2604,I2850);
nor I_73 (I2358,I2946,I2454);
nor I_74 (I2355,I2437,I2946);
not I_75 (I2991,I2771);
nand I_76 (I3008,I2991,I2867);
nor I_77 (I2346,I2471,I3008);
not I_78 (I3072,I1705);
or I_79 (I3089,I1720,I1732);
nor I_80 (I3106,I1720,I1732);
nor I_81 (I3123,I3106,I1729);
not I_82 (I3140,I3123);
nand I_83 (I3157,I3089,I1723);
not I_84 (I3174,I3157);
not I_85 (I3191,I1717);
nor I_86 (I3034,I3191,I3174);
nor I_87 (I3222,I3191,I3157);
nor I_88 (I3239,I3123,I1717);
not I_89 (I3256,I1726);
nand I_90 (I3273,I1714,I1711);
nand I_91 (I3290,I3273,I1726);
nor I_92 (I3307,I3157,I3290);
not I_93 (I3324,I3307);
nor I_94 (I3049,I3290,I3222);
not I_95 (I3355,I3290);
nor I_96 (I3372,I3355,I3123);
nor I_97 (I3037,I3191,I3372);
nor I_98 (I3052,I3290,I3140);
nand I_99 (I3417,I3273,I3256);
and I_100 (I3434,I3417,I1720);
nand I_101 (I3451,I3434,I1708);
not I_102 (I3468,I3451);
nor I_103 (I3485,I3468,I1717);
nand I_104 (I3502,I3239,I3451);
not I_105 (I3043,I3502);
nor I_106 (I3533,I1714,I1711);
or I_107 (I3550,I3533,I1717);
nor I_108 (I3567,I1708,I1735);
nand I_109 (I3584,I3567,I3550);
not I_110 (I3601,I3584);
nor I_111 (I3064,I3601,I3157);
nand I_112 (I3632,I3601,I3485);
nand I_113 (I3040,I3502,I3632);
nor I_114 (I3663,I3601,I3174);
nor I_115 (I3061,I3663,I3191);
nor I_116 (I3055,I3601,I3355);
nor I_117 (I3708,I3584,I3140);
nor I_118 (I3725,I3468,I3708);
nor I_119 (I3046,I3725,I3324);
nor I_120 (I3756,I3157,I3584);
nor I_121 (I3773,I3451,I3756);
DFFARX1 I_122 (I3773,I1698,I3072,I3058,);
not I_123 (I3837,I1705);
or I_124 (I3854,I2337,I2337);
nor I_125 (I3871,I2337,I2337);
nor I_126 (I3888,I3871,I2352);
not I_127 (I3905,I3888);
nand I_128 (I3922,I3854,I2349);
not I_129 (I3939,I3922);
not I_130 (I3956,I2361);
nor I_131 (I3799,I3956,I3939);
nor I_132 (I3987,I3956,I3922);
nor I_133 (I4004,I3888,I2361);
not I_134 (I4021,I2340);
nand I_135 (I4038,I2352,I2343);
nand I_136 (I4055,I4038,I2340);
nor I_137 (I4072,I3922,I4055);
not I_138 (I4089,I4072);
nor I_139 (I3814,I4055,I3987);
not I_140 (I4120,I4055);
nor I_141 (I4137,I4120,I3888);
nor I_142 (I3802,I3956,I4137);
nor I_143 (I3817,I4055,I3905);
nand I_144 (I4182,I4038,I4021);
and I_145 (I4199,I4182,I2349);
nand I_146 (I4216,I4199,I2343);
not I_147 (I4233,I4216);
nor I_148 (I4250,I4233,I2361);
nand I_149 (I4267,I4004,I4216);
not I_150 (I3808,I4267);
nor I_151 (I4298,I2346,I2346);
or I_152 (I4315,I4298,I2340);
nor I_153 (I4332,I2355,I2358);
nand I_154 (I4349,I4332,I4315);
not I_155 (I4366,I4349);
nor I_156 (I3829,I4366,I3922);
nand I_157 (I4397,I4366,I4250);
nand I_158 (I3805,I4267,I4397);
nor I_159 (I4428,I4366,I3939);
nor I_160 (I3826,I4428,I3956);
nor I_161 (I3820,I4366,I4120);
nor I_162 (I4473,I4349,I3905);
nor I_163 (I4490,I4233,I4473);
nor I_164 (I3811,I4490,I4089);
nor I_165 (I4521,I3922,I4349);
nor I_166 (I4538,I4216,I4521);
DFFARX1 I_167 (I4538,I1698,I3837,I3823,);
endmodule


