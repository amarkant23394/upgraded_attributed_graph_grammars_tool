module test_final(IN_1_1_l_5,IN_2_1_l_5,IN_3_1_l_5,IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_4_2_l_5,IN_5_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_3_3_l_5,IN_1_10_l_5,IN_2_10_l_5,IN_3_10_l_5,IN_4_10_l_5,blif_clk_net_7_r_12,blif_reset_net_7_r_12,N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_549_7_r_12,n_569_7_r_12,N6147_9_r_12);
input IN_1_1_l_5,IN_2_1_l_5,IN_3_1_l_5,IN_1_2_l_5,IN_2_2_l_5,IN_3_2_l_5,IN_4_2_l_5,IN_5_2_l_5,IN_1_3_l_5,IN_2_3_l_5,IN_3_3_l_5,IN_1_10_l_5,IN_2_10_l_5,IN_3_10_l_5,IN_4_10_l_5,blif_clk_net_7_r_12,blif_reset_net_7_r_12;
output N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_549_7_r_12,n_569_7_r_12,N6147_9_r_12;
wire N1371_0_r_5,N1508_0_r_5,N1372_1_r_5,N1508_1_r_5,N6147_2_r_5,N1507_6_r_5,N1508_6_r_5,G42_7_r_5,n_572_7_r_5,n_573_7_r_5,n_549_7_r_5,n_569_7_r_5,n_452_7_r_5,n4_7_r_5,n26_5,n27_5,n28_5,n29_5,n30_5,n31_5,n32_5,n33_5,n34_5,n35_5,n36_5,n37_5,n38_5,n39_5,n40_5,n41_5,n42_5,n43_5,n44_5,n45_5,n46_5,n47_5,n_573_7_r_12,n_452_7_r_12,N6134_9_r_12,I_BUFF_1_9_r_12,n1_12,n8_12,n23_12,n24_12,n25_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12,n41_12,n42_12;
nor I_0(N1371_0_r_5,n28_5,n46_5);
nand I_1(N1508_0_r_5,n26_5,n43_5);
not I_2(N1372_1_r_5,n43_5);
nor I_3(N1508_1_r_5,n30_5,n43_5);
nor I_4(N6147_2_r_5,n29_5,n32_5);
nor I_5(N1507_6_r_5,n26_5,n44_5);
nor I_6(N1508_6_r_5,n27_5,n37_5);
DFFARX1 I_7(n4_7_r_5,blif_clk_net_7_r_12,n8_12,G42_7_r_5,);
and I_8(n_572_7_r_5,n27_5,n28_5);
nand I_9(n_573_7_r_5,n26_5,n27_5);
nand I_10(n_549_7_r_5,IN_1_10_l_5,IN_2_10_l_5);
nand I_11(n_569_7_r_5,n_549_7_r_5,n26_5);
not I_12(n_452_7_r_5,n29_5);
nor I_13(n4_7_r_5,n30_5,n31_5);
not I_14(n26_5,n35_5);
nand I_15(n27_5,n40_5,n41_5);
nand I_16(n28_5,IN_1_1_l_5,IN_2_1_l_5);
nand I_17(n29_5,n27_5,n33_5);
nor I_18(n30_5,IN_1_3_l_5,n45_5);
not I_19(n31_5,n_549_7_r_5);
nor I_20(n32_5,n34_5,n35_5);
not I_21(n33_5,n30_5);
nor I_22(n34_5,n31_5,n36_5);
nor I_23(n35_5,IN_3_1_l_5,n28_5);
not I_24(n36_5,n28_5);
nand I_25(n37_5,n36_5,n38_5);
nand I_26(n38_5,n26_5,n39_5);
nand I_27(n39_5,n30_5,n31_5);
nor I_28(n40_5,IN_1_2_l_5,IN_2_2_l_5);
or I_29(n41_5,IN_5_2_l_5,n42_5);
nor I_30(n42_5,IN_3_2_l_5,IN_4_2_l_5);
nand I_31(n43_5,n36_5,n46_5);
nor I_32(n44_5,n_549_7_r_5,n33_5);
or I_33(n45_5,IN_2_3_l_5,IN_3_3_l_5);
and I_34(n46_5,n31_5,n47_5);
or I_35(n47_5,IN_3_10_l_5,IN_4_10_l_5);
nor I_36(N1371_0_r_12,I_BUFF_1_9_r_12,n36_12);
nand I_37(N1508_0_r_12,n30_12,n37_12);
nor I_38(N1507_6_r_12,n25_12,n39_12);
nor I_39(N1508_6_r_12,n25_12,n29_12);
DFFARX1 I_40(n1_12,blif_clk_net_7_r_12,n8_12,G42_7_r_12,);
nor I_41(n_572_7_r_12,n23_12,n24_12);
nand I_42(n_573_7_r_12,n_452_7_r_12,n25_12);
nand I_43(n_549_7_r_12,n27_12,n28_12);
nand I_44(n_569_7_r_12,n25_12,n26_12);
nand I_45(n_452_7_r_12,N1508_1_r_5,N1372_1_r_5);
nand I_46(N6147_9_r_12,n30_12,n31_12);
nor I_47(N6134_9_r_12,n35_12,n36_12);
not I_48(I_BUFF_1_9_r_12,n_452_7_r_12);
not I_49(n1_12,n_573_7_r_12);
not I_50(n8_12,blif_reset_net_7_r_12);
not I_51(n23_12,n36_12);
nor I_52(n24_12,n_452_7_r_12,N6147_2_r_5);
nand I_53(n25_12,n23_12,n40_12);
not I_54(n26_12,n35_12);
not I_55(n27_12,N6134_9_r_12);
nand I_56(n28_12,n26_12,n29_12);
not I_57(n29_12,n24_12);
nand I_58(n30_12,n33_12,n41_12);
nand I_59(n31_12,n32_12,n33_12);
nor I_60(n32_12,n26_12,n34_12);
nor I_61(n33_12,N1508_0_r_5,N1372_1_r_5);
nor I_62(n34_12,n42_12,n_573_7_r_5);
nor I_63(n35_12,n38_12,N1508_0_r_5);
nand I_64(n36_12,n_569_7_r_5,n_452_7_r_5);
nand I_65(n37_12,n23_12,n35_12);
or I_66(n38_12,N1508_6_r_5,G42_7_r_5);
not I_67(n39_12,n30_12);
or I_68(n40_12,n_572_7_r_5,N1371_0_r_5);
nor I_69(n41_12,n34_12,n36_12);
nor I_70(n42_12,N1371_0_r_5,N1507_6_r_5);
endmodule


