module test_final(G18_1_l_0,G15_1_l_0,IN_1_1_l_0,IN_4_1_l_0,IN_5_1_l_0,IN_7_1_l_0,IN_9_1_l_0,IN_10_1_l_0,IN_1_3_l_0,IN_2_3_l_0,IN_4_3_l_0,blif_clk_net_1_r_9,blif_reset_net_1_r_9,G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9);
input G18_1_l_0,G15_1_l_0,IN_1_1_l_0,IN_4_1_l_0,IN_5_1_l_0,IN_7_1_l_0,IN_9_1_l_0,IN_10_1_l_0,IN_1_3_l_0,IN_2_3_l_0,IN_4_3_l_0,blif_clk_net_1_r_9,blif_reset_net_1_r_9;
output G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9;
wire G42_1_r_0,n_572_1_r_0,n_573_1_r_0,n_549_1_r_0,n_569_1_r_0,n_42_2_r_0,G199_2_r_0,G199_4_r_0,G214_4_r_0,n4_1_l_0,n37_0,n38_0,n20_0,ACVQN1_3_l_0,n4_1_r_0,N3_2_r_0,N1_4_r_0,n2_0,n21_0,n22_0,n23_0,n24_0,n25_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0,n_452_1_r_9,N3_2_l_9,n5_9,n27_9,n16_9,n26_9,n15_9,n29_internal_9,n29_9,N1_4_l_9,n25_9,n28_internal_9,n28_9,n4_1_r_9,N3_2_r_9,N1_4_r_9,n_42_2_l_9,n17_9,n18_9,n19_9,n20_9,n21_9,n22_9,n23_9,n24_9;
DFFARX1 I_0(n4_1_r_0,blif_clk_net_1_r_9,n5_9,G42_1_r_0,);
nor I_1(n_572_1_r_0,IN_5_1_l_0,n23_0);
nand I_2(n_573_1_r_0,n21_0,n22_0);
nand I_3(n_549_1_r_0,n_569_1_r_0,n24_0);
nand I_4(n_569_1_r_0,n21_0,n26_0);
nor I_5(n_42_2_r_0,n27_0,n28_0);
DFFARX1 I_6(N3_2_r_0,blif_clk_net_1_r_9,n5_9,G199_2_r_0,);
DFFARX1 I_7(N1_4_r_0,blif_clk_net_1_r_9,n5_9,G199_4_r_0,);
DFFARX1 I_8(n2_0,blif_clk_net_1_r_9,n5_9,G214_4_r_0,);
nor I_9(n4_1_l_0,G18_1_l_0,IN_1_1_l_0);
DFFARX1 I_10(n4_1_l_0,blif_clk_net_1_r_9,n5_9,n37_0,);
DFFARX1 I_11(IN_1_3_l_0,blif_clk_net_1_r_9,n5_9,n38_0,);
not I_12(n20_0,n38_0);
DFFARX1 I_13(IN_2_3_l_0,blif_clk_net_1_r_9,n5_9,ACVQN1_3_l_0,);
nor I_14(n4_1_r_0,IN_10_1_l_0,n23_0);
nor I_15(N3_2_r_0,n31_0,n32_0);
nor I_16(N1_4_r_0,n29_0,n32_0);
not I_17(n2_0,n31_0);
nor I_18(n21_0,IN_9_1_l_0,n37_0);
not I_19(n22_0,IN_5_1_l_0);
nand I_20(n23_0,n20_0,n30_0);
nand I_21(n24_0,n38_0,n25_0);
nor I_22(n25_0,IN_9_1_l_0,IN_10_1_l_0);
not I_23(n26_0,IN_10_1_l_0);
not I_24(n27_0,n29_0);
nor I_25(n28_0,G15_1_l_0,IN_7_1_l_0);
nand I_26(n29_0,n26_0,n33_0);
not I_27(n30_0,IN_9_1_l_0);
nand I_28(n31_0,IN_4_3_l_0,ACVQN1_3_l_0);
and I_29(n32_0,n35_0,n36_0);
nand I_30(n33_0,IN_4_1_l_0,n34_0);
not I_31(n34_0,G15_1_l_0);
nor I_32(n35_0,G18_1_l_0,G15_1_l_0);
nor I_33(n36_0,IN_5_1_l_0,IN_7_1_l_0);
DFFARX1 I_34(n4_1_r_9,blif_clk_net_1_r_9,n5_9,G42_1_r_9,);
nor I_35(n_572_1_r_9,n27_9,n_42_2_l_9);
or I_36(n_573_1_r_9,n25_9,n_42_2_l_9);
nand I_37(n_549_1_r_9,n17_9,n18_9);
or I_38(n_569_1_r_9,n26_9,n_42_2_l_9);
nor I_39(n_452_1_r_9,n26_9,n25_9);
nor I_40(n_42_2_r_9,n25_9,n19_9);
DFFARX1 I_41(N3_2_r_9,blif_clk_net_1_r_9,n5_9,G199_2_r_9,);
DFFARX1 I_42(N1_4_r_9,blif_clk_net_1_r_9,n5_9,G199_4_r_9,);
DFFARX1 I_43(n_42_2_l_9,blif_clk_net_1_r_9,n5_9,G214_4_r_9,);
and I_44(N3_2_l_9,n22_9,n_42_2_r_0);
not I_45(n5_9,blif_reset_net_1_r_9);
DFFARX1 I_46(N3_2_l_9,blif_clk_net_1_r_9,n5_9,n27_9,);
not I_47(n16_9,n27_9);
DFFARX1 I_48(G199_2_r_0,blif_clk_net_1_r_9,n5_9,n26_9,);
not I_49(n15_9,n26_9);
DFFARX1 I_50(n_572_1_r_0,blif_clk_net_1_r_9,n5_9,n29_internal_9,);
not I_51(n29_9,n29_internal_9);
and I_52(N1_4_l_9,n24_9,G42_1_r_0);
DFFARX1 I_53(N1_4_l_9,blif_clk_net_1_r_9,n5_9,n25_9,);
DFFARX1 I_54(n_573_1_r_0,blif_clk_net_1_r_9,n5_9,n28_internal_9,);
not I_55(n28_9,n28_internal_9);
nor I_56(n4_1_r_9,n27_9,n26_9);
nor I_57(N3_2_r_9,n15_9,n21_9);
nor I_58(N1_4_r_9,n16_9,n21_9);
nor I_59(n_42_2_l_9,n_572_1_r_0,n_573_1_r_0);
not I_60(n17_9,n_452_1_r_9);
nand I_61(n18_9,n27_9,n15_9);
nor I_62(n19_9,n29_9,n20_9);
not I_63(n20_9,G42_1_r_0);
and I_64(n21_9,n23_9,G42_1_r_0);
nand I_65(n22_9,n_572_1_r_0,G199_4_r_0);
nor I_66(n23_9,n29_9,n28_9);
nand I_67(n24_9,n_549_1_r_0,G214_4_r_0);
endmodule


