module test_I3481(I3120,I2897,I2557,I3413,I1294,I1301,I3481);
input I3120,I2897,I2557,I3413,I1294,I1301;
output I3481;
wire I3464,I3137,I2551,I2575,I2583,I3430,I3246,I3447;
or I_0(I3464,I3447,I2575);
and I_1(I3137,I2897,I3120);
DFFARX1 I_2(I3464,I1294,I3246,,,I3481,);
DFFARX1 I_3(I2897,I1294,I2583,,,I2551,);
DFFARX1 I_4(I3137,I1294,I2583,,,I2575,);
not I_5(I2583,I1301);
nor I_6(I3430,I3413,I2557);
not I_7(I3246,I1301);
and I_8(I3447,I3430,I2551);
endmodule


