module test_I10583(I1477,I7604,I7731,I1470,I6315,I10583);
input I1477,I7604,I7731,I1470,I6315;
output I10583;
wire I7556,I7621,I7816,I7850,I10490,I10052;
nand I_0(I7556,I7621,I7850);
nand I_1(I7621,I7604,I6315);
DFFARX1 I_2(I1470,,,I7816,);
DFFARX1 I_3(I10490,I1470,I10052,,,I10583,);
nor I_4(I7850,I7816,I7731);
DFFARX1 I_5(I7556,I1470,I10052,,,I10490,);
not I_6(I10052,I1477);
endmodule


