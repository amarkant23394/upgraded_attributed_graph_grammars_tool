module test_final(IN_1_2_l_9,IN_2_2_l_9,IN_3_2_l_9,IN_6_2_l_9,IN_1_3_l_9,IN_2_3_l_9,IN_4_3_l_9,IN_1_4_l_9,IN_2_4_l_9,IN_3_4_l_9,IN_6_4_l_9,blif_clk_net_1_r_4,blif_reset_net_1_r_4,G42_1_r_4,n_572_1_r_4,n_573_1_r_4,n_549_1_r_4,n_569_1_r_4,ACVQN2_3_r_4,n_266_and_0_3_r_4,ACVQN1_5_r_4,P6_5_r_4);
input IN_1_2_l_9,IN_2_2_l_9,IN_3_2_l_9,IN_6_2_l_9,IN_1_3_l_9,IN_2_3_l_9,IN_4_3_l_9,IN_1_4_l_9,IN_2_4_l_9,IN_3_4_l_9,IN_6_4_l_9,blif_clk_net_1_r_4,blif_reset_net_1_r_4;
output G42_1_r_4,n_572_1_r_4,n_573_1_r_4,n_549_1_r_4,n_569_1_r_4,ACVQN2_3_r_4,n_266_and_0_3_r_4,ACVQN1_5_r_4,P6_5_r_4;
wire G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_452_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9,N3_2_l_9,n27_9,n16_9,n26_9,n15_9,n29_internal_9,n29_9,N1_4_l_9,n25_9,n28_internal_9,n28_9,n4_1_r_9,N3_2_r_9,N1_4_r_9,n_42_2_l_9,n17_9,n18_9,n19_9,n20_9,n21_9,n22_9,n23_9,n24_9,n_431_0_l_4,n6_4,G78_0_l_4,ACVQN1_5_l_4,n16_4,n17_internal_4,n17_4,n4_1_r_4,n19_4,n15_internal_4,n15_4,P6_5_r_internal_4,n20_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4;
DFFARX1 I_0(n4_1_r_9,blif_clk_net_1_r_4,n6_4,G42_1_r_9,);
nor I_1(n_572_1_r_9,n27_9,n_42_2_l_9);
or I_2(n_573_1_r_9,n25_9,n_42_2_l_9);
nand I_3(n_549_1_r_9,n17_9,n18_9);
or I_4(n_569_1_r_9,n26_9,n_42_2_l_9);
nor I_5(n_452_1_r_9,n26_9,n25_9);
nor I_6(n_42_2_r_9,n25_9,n19_9);
DFFARX1 I_7(N3_2_r_9,blif_clk_net_1_r_4,n6_4,G199_2_r_9,);
DFFARX1 I_8(N1_4_r_9,blif_clk_net_1_r_4,n6_4,G199_4_r_9,);
DFFARX1 I_9(n_42_2_l_9,blif_clk_net_1_r_4,n6_4,G214_4_r_9,);
and I_10(N3_2_l_9,IN_6_2_l_9,n22_9);
DFFARX1 I_11(N3_2_l_9,blif_clk_net_1_r_4,n6_4,n27_9,);
not I_12(n16_9,n27_9);
DFFARX1 I_13(IN_1_3_l_9,blif_clk_net_1_r_4,n6_4,n26_9,);
not I_14(n15_9,n26_9);
DFFARX1 I_15(IN_2_3_l_9,blif_clk_net_1_r_4,n6_4,n29_internal_9,);
not I_16(n29_9,n29_internal_9);
and I_17(N1_4_l_9,IN_6_4_l_9,n24_9);
DFFARX1 I_18(N1_4_l_9,blif_clk_net_1_r_4,n6_4,n25_9,);
DFFARX1 I_19(IN_3_4_l_9,blif_clk_net_1_r_4,n6_4,n28_internal_9,);
not I_20(n28_9,n28_internal_9);
nor I_21(n4_1_r_9,n27_9,n26_9);
nor I_22(N3_2_r_9,n15_9,n21_9);
nor I_23(N1_4_r_9,n16_9,n21_9);
nor I_24(n_42_2_l_9,IN_1_2_l_9,IN_3_2_l_9);
not I_25(n17_9,n_452_1_r_9);
nand I_26(n18_9,n27_9,n15_9);
nor I_27(n19_9,n29_9,n20_9);
not I_28(n20_9,IN_4_3_l_9);
and I_29(n21_9,IN_4_3_l_9,n23_9);
nand I_30(n22_9,IN_2_2_l_9,IN_3_2_l_9);
nor I_31(n23_9,n29_9,n28_9);
nand I_32(n24_9,IN_1_4_l_9,IN_2_4_l_9);
DFFARX1 I_33(n4_1_r_4,blif_clk_net_1_r_4,n6_4,G42_1_r_4,);
nor I_34(n_572_1_r_4,G78_0_l_4,n17_4);
nand I_35(n_573_1_r_4,n16_4,G214_4_r_9);
nor I_36(n_549_1_r_4,n22_4,n23_4);
nand I_37(n_569_1_r_4,n20_4,n21_4);
DFFARX1 I_38(n19_4,blif_clk_net_1_r_4,n6_4,ACVQN2_3_r_4,);
nor I_39(n_266_and_0_3_r_4,n15_4,n29_4);
DFFARX1 I_40(n19_4,blif_clk_net_1_r_4,n6_4,ACVQN1_5_r_4,);
not I_41(P6_5_r_4,P6_5_r_internal_4);
or I_42(n_431_0_l_4,n26_4,n_572_1_r_9);
not I_43(n6_4,blif_reset_net_1_r_4);
DFFARX1 I_44(n_431_0_l_4,blif_clk_net_1_r_4,n6_4,G78_0_l_4,);
DFFARX1 I_45(n_569_1_r_9,blif_clk_net_1_r_4,n6_4,ACVQN1_5_l_4,);
not I_46(n16_4,ACVQN1_5_l_4);
DFFARX1 I_47(n_549_1_r_9,blif_clk_net_1_r_4,n6_4,n17_internal_4,);
not I_48(n17_4,n17_internal_4);
nor I_49(n4_1_r_4,n30_4,n31_4);
nand I_50(n19_4,n33_4,G42_1_r_9);
DFFARX1 I_51(G78_0_l_4,blif_clk_net_1_r_4,n6_4,n15_internal_4,);
not I_52(n15_4,n15_internal_4);
DFFARX1 I_53(ACVQN1_5_l_4,blif_clk_net_1_r_4,n6_4,P6_5_r_internal_4,);
and I_54(n20_4,n16_4,n_42_2_r_9);
nor I_55(n21_4,G42_1_r_9,G214_4_r_9);
nand I_56(n22_4,G78_0_l_4,n25_4);
nand I_57(n23_4,n24_4,n_42_2_r_9);
not I_58(n24_4,G214_4_r_9);
not I_59(n25_4,G42_1_r_9);
and I_60(n26_4,n27_4,G199_2_r_9);
nor I_61(n27_4,n28_4,n_573_1_r_9);
not I_62(n28_4,G42_1_r_9);
not I_63(n29_4,n30_4);
nand I_64(n30_4,n32_4,G199_4_r_9);
nand I_65(n31_4,n25_4,n_42_2_r_9);
nor I_66(n32_4,n33_4,G214_4_r_9);
not I_67(n33_4,n_572_1_r_9);
endmodule


