module test_I1873(I1215,I1294,I1301,I1873);
input I1215,I1294,I1301;
output I1873;
wire I1342,I1780;
DFFARX1 I_0(I1780,I1294,I1342,,,I1873,);
not I_1(I1342,I1301);
DFFARX1 I_2(I1215,I1294,I1342,,,I1780,);
endmodule


