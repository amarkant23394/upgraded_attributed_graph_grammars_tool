module Benchmark_testing5000(I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1803,I1810,I4472,I4463,I4460,I4466,I4454,I4448,I4469,I4457,I4451,I26116,I26095,I26089,I26104,I26092,I26107,I26098,I26101,I26113,I26110,I37616,I37613,I37604,I37607,I37601,I37610,I37598,I37622,I37619,I41081,I41084,I41066,I41075,I41087,I41078,I41069,I41072,I41090,I74665,I74644,I74647,I74662,I74659,I74656,I74653,I74641,I74650);
input I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1803,I1810;
output I4472,I4463,I4460,I4466,I4454,I4448,I4469,I4457,I4451,I26116,I26095,I26089,I26104,I26092,I26107,I26098,I26101,I26113,I26110,I37616,I37613,I37604,I37607,I37601,I37610,I37598,I37622,I37619,I41081,I41084,I41066,I41075,I41087,I41078,I41069,I41072,I41090,I74665,I74644,I74647,I74662,I74659,I74656,I74653,I74641,I74650;
wire I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1803,I1810,I1845,I82206,I1871,I1888,I1896,I1913,I82209,I82215,I1930,I82224,I1956,I1837,I1828,I82227,I2001,I2009,I82218,I2026,I1825,I2066,I2074,I1831,I1819,I2119,I82233,I82212,I2136,I82221,I2162,I2170,I1813,I2201,I2218,I82230,I2235,I2252,I2269,I1834,I2300,I1822,I1816,I2372,I39338,I2398,I2415,I2423,I2440,I39353,I39356,I2457,I39335,I2483,I2364,I2355,I39341,I2528,I2536,I39347,I2553,I2352,I2593,I2601,I2358,I2346,I2646,I39350,I39332,I2663,I39344,I2689,I2697,I2340,I2728,I2745,I2762,I2779,I2796,I2361,I2827,I2349,I2343,I2899,I79826,I2925,I2942,I2950,I2967,I79829,I79835,I2984,I79844,I3010,I2891,I2882,I79847,I3055,I3063,I79838,I3080,I2879,I3120,I3128,I2885,I2873,I3173,I79853,I79832,I3190,I79841,I3216,I3224,I2867,I3255,I3272,I79850,I3289,I3306,I3323,I2888,I3354,I2876,I2870,I3426,I6559,I3452,I3469,I3477,I3494,I6574,I3511,I6577,I3537,I3418,I3409,I6571,I3582,I3590,I6580,I3607,I3406,I6556,I3647,I3655,I3412,I3400,I3700,I6562,I3717,I6565,I3743,I3751,I3394,I3782,I3799,I6568,I3816,I3833,I3850,I3415,I3881,I3403,I3397,I3953,I3979,I3996,I4004,I4021,I4038,I4064,I3945,I3936,I4109,I4117,I4134,I3933,I4174,I4182,I3939,I3927,I4227,I4244,I4270,I4278,I3921,I4309,I4326,I4343,I4360,I4377,I3942,I4408,I3930,I3924,I4480,I40494,I4506,I4523,I4531,I4548,I40509,I40512,I4565,I40491,I4591,I40497,I4636,I4644,I40503,I4661,I4701,I4709,I4754,I40506,I40488,I4771,I40500,I4797,I4805,I4836,I4853,I4870,I4887,I4904,I4935,I5007,I18653,I5033,I5041,I5058,I18635,I18650,I5075,I18626,I5101,I18629,I5118,I5126,I18644,I5143,I4975,I5174,I5191,I4987,I18647,I5231,I4996,I5253,I18638,I5270,I18632,I5296,I5313,I4999,I5335,I4984,I5366,I18641,I5383,I5400,I5417,I4993,I5448,I4981,I4990,I4978,I5534,I26651,I5560,I5568,I5585,I26645,I26636,I5602,I26657,I5628,I26639,I5645,I5653,I26633,I5670,I5502,I5701,I5718,I5514,I5758,I5523,I5780,I26660,I26642,I5797,I26648,I5823,I5840,I5526,I5862,I5511,I5893,I26654,I5910,I5927,I5944,I5520,I5975,I5508,I5517,I5505,I6061,I60398,I6087,I6095,I6112,I60395,I60401,I6129,I6155,I6172,I6180,I6197,I6029,I6228,I6245,I6041,I60404,I6285,I6050,I6307,I60407,I60416,I6324,I60410,I6350,I6367,I6053,I6389,I6038,I6420,I60413,I6437,I6454,I6471,I6047,I6502,I6035,I6044,I6032,I6588,I46855,I6614,I6622,I6639,I46852,I46867,I6656,I46849,I6682,I46846,I6699,I6707,I6724,I6755,I6772,I6812,I6834,I46861,I6851,I46864,I6877,I6894,I6916,I6947,I46858,I6964,I6981,I6998,I7029,I7115,I15491,I7141,I7149,I7166,I15473,I15488,I7183,I15464,I7209,I15467,I7226,I7234,I15482,I7251,I7083,I7282,I7299,I7095,I15485,I7339,I7104,I7361,I15476,I7378,I15470,I7404,I7421,I7107,I7443,I7092,I7474,I15479,I7491,I7508,I7525,I7101,I7556,I7089,I7098,I7086,I7642,I54590,I7668,I7676,I7693,I54608,I54602,I7710,I54581,I7736,I54599,I7753,I7761,I54584,I7778,I7610,I7809,I7826,I7622,I54596,I7866,I7631,I7888,I54605,I54593,I7905,I54587,I7931,I7948,I7634,I7970,I7619,I8001,I8018,I8035,I8052,I7628,I8083,I7616,I7625,I7613,I8169,I35873,I8195,I8203,I8220,I35885,I35870,I8237,I35864,I8263,I35879,I8280,I8288,I35867,I8305,I8137,I8336,I8353,I8149,I35876,I8393,I8158,I8415,I35882,I35888,I8432,I8458,I8475,I8161,I8497,I8146,I8528,I8545,I8562,I8579,I8155,I8610,I8143,I8152,I8140,I8696,I50017,I8722,I8730,I8747,I50014,I50029,I8764,I50011,I8790,I50008,I8807,I8815,I8832,I8664,I8863,I8880,I8676,I8920,I8685,I8942,I50023,I8959,I50026,I8985,I9002,I8688,I9024,I8673,I9055,I50020,I9072,I9089,I9106,I8682,I9137,I8670,I8679,I8667,I9223,I79243,I9249,I9257,I9274,I79237,I79258,I9291,I79234,I9317,I79255,I9334,I9342,I79252,I9359,I9191,I9390,I9407,I9203,I79240,I9447,I9212,I9469,I79249,I79246,I9486,I79231,I9512,I9529,I9215,I9551,I9200,I9582,I9599,I9616,I9633,I9209,I9664,I9197,I9206,I9194,I9750,I58466,I9776,I9784,I9801,I58484,I58478,I9818,I58457,I9844,I58475,I9861,I9869,I58460,I9886,I9718,I9917,I9934,I9730,I58472,I9974,I9739,I9996,I58481,I58469,I10013,I58463,I10039,I10056,I9742,I10078,I9727,I10109,I10126,I10143,I10160,I9736,I10191,I9724,I9733,I9721,I10277,I66657,I10303,I10311,I10328,I66672,I66651,I10345,I66654,I10371,I66675,I10388,I10396,I10413,I10245,I10444,I10461,I10257,I10501,I10266,I10523,I66663,I66660,I10540,I66666,I10566,I10583,I10269,I10605,I10254,I10636,I66669,I10653,I10670,I10687,I10263,I10718,I10251,I10260,I10248,I10804,I41656,I10830,I10838,I10855,I41647,I41665,I10872,I41644,I10898,I10915,I10923,I41650,I10940,I10772,I10971,I10988,I10784,I11028,I10793,I11050,I41662,I41653,I11067,I41668,I11093,I11110,I10796,I11132,I10781,I11163,I41659,I11180,I11197,I11214,I10790,I11245,I10778,I10787,I10775,I11331,I70119,I11357,I11374,I11323,I11396,I11422,I11430,I11447,I70122,I11464,I70134,I11481,I11498,I70140,I11515,I70131,I11532,I70137,I11549,I11299,I11580,I11597,I11614,I11631,I11311,I11305,I11676,I70128,I11320,I11314,I11721,I11738,I70125,I11755,I70143,I11772,I11798,I11806,I11308,I11302,I11860,I11868,I11317,I11926,I19680,I11952,I11969,I11918,I11991,I19695,I12017,I12025,I12042,I19692,I12059,I12076,I12093,I19689,I12110,I19704,I12127,I19701,I12144,I11894,I12175,I12192,I12209,I12226,I11906,I11900,I12271,I19698,I11915,I11909,I12316,I12333,I19686,I12350,I19707,I12367,I19683,I12393,I12401,I11903,I11897,I12455,I12463,I11912,I12521,I55242,I12547,I12564,I12513,I12586,I55251,I12612,I12620,I12637,I55239,I12654,I55230,I12671,I12688,I55236,I12705,I55254,I12722,I55227,I12739,I12489,I12770,I12787,I12804,I12821,I12501,I12495,I12866,I55233,I12510,I12504,I12911,I12928,I55245,I12945,I12962,I55248,I12988,I12996,I12498,I12492,I13050,I13058,I12507,I13116,I51595,I13142,I13159,I13108,I13181,I51589,I13207,I13215,I13232,I51607,I13249,I13266,I13283,I13300,I51601,I13317,I51592,I13334,I13084,I13365,I13382,I13399,I13416,I13096,I13090,I13461,I51604,I13105,I13099,I13506,I13523,I51610,I13540,I13557,I51598,I13583,I13591,I13093,I13087,I13645,I13653,I13102,I13711,I32989,I13737,I13754,I13703,I13776,I32980,I13802,I13810,I13827,I32998,I13844,I32995,I13861,I13878,I32974,I13895,I32977,I13912,I32986,I13929,I13679,I13960,I13977,I13994,I14011,I13691,I13685,I14056,I32992,I13700,I13694,I14101,I14118,I14135,I32983,I14152,I14178,I14186,I13688,I13682,I14240,I14248,I13697,I14306,I70697,I14332,I14349,I14298,I14371,I14397,I14405,I14422,I70700,I14439,I70712,I14456,I14473,I70718,I14490,I70709,I14507,I70715,I14524,I14274,I14555,I14572,I14589,I14606,I14286,I14280,I14651,I70706,I14295,I14289,I14696,I14713,I70703,I14730,I70721,I14747,I14773,I14781,I14283,I14277,I14835,I14843,I14292,I14901,I28821,I14927,I14944,I14893,I14966,I28815,I14992,I15000,I15017,I28830,I15034,I28827,I15051,I15068,I28818,I15085,I28809,I15102,I28812,I15119,I14869,I15150,I15167,I15184,I15201,I14881,I14875,I15246,I28833,I14890,I14884,I15291,I15308,I28824,I15325,I15342,I15368,I15376,I14878,I14872,I15430,I15438,I14887,I15499,I15525,I15533,I15550,I15576,I15598,I15624,I15632,I15649,I15675,I15697,I15737,I15754,I15762,I15779,I15810,I15827,I15853,I15861,I15906,I15923,I16026,I16052,I16060,I16077,I16103,I15994,I16125,I16151,I16159,I16176,I16202,I16018,I16224,I16000,I16264,I16281,I16289,I16306,I16003,I16337,I16354,I16380,I16388,I15991,I16009,I16433,I16450,I16012,I15997,I16006,I16015,I16553,I16579,I16587,I16604,I16630,I16521,I16652,I16678,I16686,I16703,I16729,I16545,I16751,I16527,I16791,I16808,I16816,I16833,I16530,I16864,I16881,I16907,I16915,I16518,I16536,I16960,I16977,I16539,I16524,I16533,I16542,I17080,I30002,I17106,I17114,I30014,I17131,I29999,I17157,I17048,I17179,I30023,I17205,I17213,I30020,I17230,I17256,I17072,I17278,I17054,I30011,I17318,I17335,I17343,I17360,I17057,I17391,I30008,I17408,I30017,I17434,I17442,I17045,I17063,I17487,I30005,I17504,I17066,I17051,I17060,I17069,I17607,I34145,I17633,I17641,I34130,I34133,I17658,I34148,I17684,I17575,I17706,I34142,I17732,I17740,I17757,I17783,I17599,I17805,I17581,I34139,I17845,I17862,I17870,I17887,I17584,I17918,I34154,I17935,I34151,I17961,I17969,I17572,I17590,I18014,I34136,I18031,I17593,I17578,I17587,I17596,I18134,I81037,I18160,I18168,I81016,I18185,I81043,I18211,I18102,I18233,I81031,I18259,I18267,I81034,I18284,I18310,I18126,I18332,I18108,I81025,I18372,I18389,I18397,I18414,I18111,I18445,I81022,I81019,I18462,I81040,I18488,I18496,I18099,I18117,I18541,I81028,I18558,I18120,I18105,I18114,I18123,I18661,I68963,I18687,I18695,I68978,I18712,I68981,I18738,I18760,I68987,I18786,I18794,I68969,I18811,I18837,I18859,I68966,I18899,I18916,I18924,I18941,I18972,I68972,I18989,I68984,I19015,I19023,I19068,I68975,I19085,I19188,I19214,I19222,I19239,I19265,I19156,I19287,I19313,I19321,I19338,I19364,I19180,I19386,I19162,I19426,I19443,I19451,I19468,I19165,I19499,I19516,I19542,I19550,I19153,I19171,I19595,I19612,I19174,I19159,I19168,I19177,I19715,I59106,I19741,I19749,I59103,I59121,I19766,I59112,I19792,I19814,I59127,I19840,I19848,I59109,I19865,I19891,I19913,I59115,I19953,I19970,I19978,I19995,I20026,I59130,I20043,I59118,I20069,I20077,I20122,I59124,I20139,I20242,I30597,I20268,I20276,I30609,I20293,I30594,I20319,I20210,I20341,I30618,I20367,I20375,I30615,I20392,I20418,I20234,I20440,I20216,I30606,I20480,I20497,I20505,I20522,I20219,I20553,I30603,I20570,I30612,I20596,I20604,I20207,I20225,I20649,I30600,I20666,I20228,I20213,I20222,I20231,I20769,I75778,I20795,I20803,I75775,I75766,I20820,I75763,I20846,I20737,I20868,I75772,I20894,I20902,I75781,I20919,I20945,I20761,I20967,I20743,I75784,I21007,I21024,I21032,I21049,I20746,I21080,I75769,I21097,I75787,I21123,I21131,I20734,I20752,I21176,I21193,I20755,I20740,I20749,I20758,I21296,I62081,I21322,I21330,I62078,I21347,I62090,I21373,I21264,I21395,I21421,I21429,I62096,I21446,I21472,I21288,I21494,I21270,I62084,I21534,I21551,I21559,I21576,I21273,I21607,I62093,I62099,I21624,I21650,I21658,I21261,I21279,I21703,I62087,I21720,I21282,I21267,I21276,I21285,I21823,I55876,I21849,I21857,I55873,I55891,I21874,I55882,I21900,I21791,I21922,I55897,I21948,I21956,I55879,I21973,I21999,I21815,I22021,I21797,I55885,I22061,I22078,I22086,I22103,I21800,I22134,I55900,I22151,I55888,I22177,I22185,I21788,I21806,I22230,I55894,I22247,I21809,I21794,I21803,I21812,I22350,I82822,I22376,I22384,I82801,I22401,I82828,I22427,I22318,I22449,I82816,I22475,I22483,I82819,I22500,I22526,I22342,I22548,I22324,I82810,I22588,I22605,I22613,I22630,I22327,I22661,I82807,I82804,I22678,I82825,I22704,I22712,I22315,I22333,I22757,I82813,I22774,I22336,I22321,I22330,I22339,I22877,I22903,I22911,I22928,I22954,I22845,I22976,I23002,I23010,I23027,I23053,I22869,I23075,I22851,I23115,I23132,I23140,I23157,I22854,I23188,I23205,I23231,I23239,I22842,I22860,I23284,I23301,I22863,I22848,I22857,I22866,I23404,I68388,I23430,I23447,I23396,I23469,I23486,I68400,I23503,I68391,I23529,I23537,I68409,I23563,I23571,I68385,I23588,I23375,I68403,I23628,I23636,I23369,I23384,I23681,I68397,I68394,I23698,I68406,I23724,I23372,I23746,I23763,I23780,I23387,I23811,I23828,I23378,I23859,I23381,I23393,I23390,I23948,I69544,I23974,I23991,I23940,I24013,I24030,I69556,I24047,I69547,I24073,I24081,I69565,I24107,I24115,I69541,I24132,I23919,I69559,I24172,I24180,I23913,I23928,I24225,I69553,I69550,I24242,I69562,I24268,I23916,I24290,I24307,I24324,I23931,I24355,I24372,I23922,I24403,I23925,I23937,I23934,I24492,I52649,I24518,I24535,I24484,I24557,I24574,I52664,I52652,I24591,I52643,I24617,I24625,I52655,I24651,I24659,I52646,I24676,I24463,I52661,I24716,I24724,I24457,I24472,I24769,I52670,I52658,I24786,I52667,I24812,I24460,I24834,I24851,I24868,I24475,I24899,I24916,I24466,I24947,I24469,I24481,I24478,I25036,I48966,I25062,I25079,I25028,I25101,I25118,I48960,I48957,I25135,I48972,I25161,I25169,I25195,I25203,I48954,I25220,I25007,I25260,I25268,I25001,I25016,I25313,I48969,I48963,I25330,I25356,I25004,I25378,I25395,I25412,I25019,I25443,I25460,I48975,I25010,I25491,I25013,I25025,I25022,I25580,I25606,I25623,I25572,I25645,I25662,I25679,I25705,I25713,I25739,I25747,I25764,I25551,I25804,I25812,I25545,I25560,I25857,I25874,I25900,I25548,I25922,I25939,I25956,I25563,I25987,I26004,I25554,I26035,I25557,I25569,I25566,I26124,I26150,I26167,I26189,I26206,I26223,I26249,I26257,I26283,I26291,I26308,I26348,I26356,I26401,I26418,I26444,I26466,I26483,I26500,I26531,I26548,I26579,I26668,I47912,I26694,I26711,I26733,I26750,I47906,I47903,I26767,I47918,I26793,I26801,I26827,I26835,I47900,I26852,I26892,I26900,I26945,I47915,I47909,I26962,I26988,I27010,I27027,I27044,I27075,I27092,I47921,I27123,I27212,I76934,I27238,I27255,I27204,I27277,I27294,I76940,I76943,I27311,I76919,I27337,I27345,I76946,I27371,I27379,I76928,I27396,I27183,I76925,I27436,I27444,I27177,I27192,I27489,I76922,I76931,I27506,I76937,I27532,I27180,I27554,I27571,I27588,I27195,I27619,I27636,I27186,I27667,I27189,I27201,I27198,I27756,I27782,I27799,I27748,I27821,I27838,I27855,I27881,I27889,I27915,I27923,I27940,I27727,I27980,I27988,I27721,I27736,I28033,I28050,I28076,I27724,I28098,I28115,I28132,I27739,I28163,I28180,I27730,I28211,I27733,I27745,I27742,I28300,I28326,I28343,I28292,I28365,I28382,I28399,I28425,I28433,I28459,I28467,I28484,I28271,I28524,I28532,I28265,I28280,I28577,I28594,I28620,I28268,I28642,I28659,I28676,I28283,I28707,I28724,I28274,I28755,I28277,I28289,I28286,I28841,I28867,I28884,I28915,I28923,I28940,I28957,I28974,I28991,I29008,I29025,I29056,I29073,I29090,I29135,I29152,I29183,I29200,I29231,I29248,I29265,I29291,I29299,I29330,I29347,I29378,I29436,I29462,I29479,I29428,I29510,I29518,I29535,I29552,I29569,I29586,I29603,I29620,I29425,I29651,I29668,I29685,I29410,I29422,I29730,I29747,I29416,I29778,I29795,I29404,I29826,I29843,I29860,I29886,I29894,I29413,I29925,I29942,I29419,I29973,I29407,I30031,I56534,I30057,I30074,I56522,I30105,I30113,I56519,I30130,I30147,I56531,I30164,I56528,I30181,I30198,I30215,I30246,I56537,I30263,I56540,I30280,I30325,I30342,I30373,I56543,I30390,I30421,I56546,I30438,I56525,I30455,I30481,I30489,I30520,I30537,I30568,I30626,I71871,I30652,I30669,I71853,I30700,I30708,I71859,I30725,I30742,I71874,I30759,I71865,I30776,I30793,I30810,I30841,I71877,I30858,I71856,I30875,I30920,I30937,I30968,I71862,I30985,I31016,I71868,I31033,I31050,I31076,I31084,I31115,I31132,I31163,I31221,I31247,I31264,I31213,I31295,I31303,I31320,I31337,I31354,I31371,I31388,I31405,I31210,I31436,I31453,I31470,I31195,I31207,I31515,I31532,I31201,I31563,I31580,I31189,I31611,I31628,I31645,I31671,I31679,I31198,I31710,I31727,I31204,I31758,I31192,I31816,I31842,I31859,I31808,I31890,I31898,I31915,I31932,I31949,I31966,I31983,I32000,I31805,I32031,I32048,I32065,I31790,I31802,I32110,I32127,I31796,I32158,I32175,I31784,I32206,I32223,I32240,I32266,I32274,I31793,I32305,I32322,I31799,I32353,I31787,I32411,I53950,I32437,I32454,I32403,I53938,I32485,I32493,I53935,I32510,I32527,I53947,I32544,I53944,I32561,I32578,I32595,I32400,I32626,I53953,I32643,I53956,I32660,I32385,I32397,I32705,I32722,I32391,I32753,I53959,I32770,I32379,I32801,I53962,I32818,I53941,I32835,I32861,I32869,I32388,I32900,I32917,I32394,I32948,I32382,I33006,I33032,I33040,I33066,I33074,I33091,I33108,I33125,I33142,I33173,I33190,I33207,I33224,I33269,I33314,I33331,I33348,I33379,I33396,I33413,I33439,I33447,I33492,I33509,I33526,I33584,I33610,I33618,I33644,I33652,I33669,I33686,I33703,I33720,I33570,I33751,I33768,I33785,I33802,I33567,I33558,I33847,I33561,I33555,I33892,I33909,I33926,I33564,I33957,I33974,I33991,I34017,I34025,I33552,I33576,I34070,I34087,I34104,I33573,I34162,I34188,I34196,I34222,I34230,I34247,I34264,I34281,I34298,I34329,I34346,I34363,I34380,I34425,I34470,I34487,I34504,I34535,I34552,I34569,I34595,I34603,I34648,I34665,I34682,I34740,I34766,I34774,I34800,I34808,I34825,I34842,I34859,I34876,I34726,I34907,I34924,I34941,I34958,I34723,I34714,I35003,I34717,I34711,I35048,I35065,I35082,I34720,I35113,I35130,I35147,I35173,I35181,I34708,I34732,I35226,I35243,I35260,I34729,I35318,I71275,I35344,I35352,I71281,I35378,I35386,I35403,I71278,I35420,I35437,I71296,I35454,I35304,I35485,I35502,I35519,I71299,I35536,I35301,I35292,I35581,I35295,I35289,I35626,I71284,I35643,I35660,I35298,I35691,I71290,I35708,I71287,I35725,I71293,I35751,I35759,I35286,I35310,I35804,I35821,I35838,I35307,I35896,I74115,I35922,I35930,I74109,I35956,I35964,I74118,I35981,I74097,I35998,I36015,I74106,I36032,I36063,I36080,I36097,I74121,I36114,I74100,I36159,I36204,I74103,I36221,I36238,I36269,I74112,I36286,I36303,I36329,I36337,I36382,I36399,I36416,I36474,I43378,I36500,I36508,I43390,I36534,I36542,I43381,I36559,I43384,I36576,I36593,I43387,I36610,I36460,I36641,I36658,I36675,I36692,I43393,I36457,I36448,I36737,I36451,I36445,I36782,I43399,I36799,I36816,I36454,I36847,I36864,I43396,I36881,I43402,I36907,I36915,I36442,I36466,I36960,I36977,I36994,I36463,I37052,I43956,I37078,I37086,I43968,I37112,I37120,I43959,I37137,I43962,I37154,I37171,I43965,I37188,I37038,I37219,I37236,I37253,I37270,I43971,I37035,I37026,I37315,I37029,I37023,I37360,I43977,I37377,I37394,I37032,I37425,I37442,I43974,I37459,I43980,I37485,I37493,I37020,I37044,I37538,I37555,I37572,I37041,I37630,I37656,I37664,I37690,I37698,I37715,I37732,I37749,I37766,I37797,I37814,I37831,I37848,I37893,I37938,I37955,I37972,I38003,I38020,I38037,I38063,I38071,I38116,I38133,I38150,I38208,I47388,I38234,I38242,I38259,I47376,I47394,I38276,I47391,I38302,I38310,I47382,I47379,I38336,I38344,I38361,I38378,I38395,I38191,I47373,I38435,I38443,I38460,I38477,I38494,I38194,I38525,I38542,I38568,I38576,I38176,I38607,I38185,I38638,I38655,I38197,I38686,I47385,I38188,I38179,I38182,I38200,I38786,I63779,I38812,I38820,I38837,I63761,I63773,I38854,I63776,I38880,I38888,I63770,I63767,I38914,I38922,I38939,I38956,I38973,I38769,I63785,I39013,I39021,I39038,I39055,I39072,I38772,I39103,I63764,I39120,I39146,I39154,I38754,I39185,I38763,I39216,I39233,I38775,I39264,I63782,I38766,I38757,I38760,I38778,I39364,I76341,I39390,I39398,I39415,I76365,I76347,I39432,I76353,I39458,I39466,I76359,I76344,I39492,I39500,I39517,I39534,I39551,I76356,I39591,I39599,I39616,I39633,I39650,I39681,I76362,I76350,I39698,I39724,I39732,I39763,I39794,I39811,I39842,I39942,I39968,I39976,I39993,I40010,I40036,I40044,I40070,I40078,I40095,I40112,I40129,I39925,I40169,I40177,I40194,I40211,I40228,I39928,I40259,I40276,I40302,I40310,I39910,I40341,I39919,I40372,I40389,I39931,I40420,I39922,I39913,I39916,I39934,I40520,I65513,I40546,I40554,I40571,I65495,I65507,I40588,I65510,I40614,I40622,I65504,I65501,I40648,I40656,I40673,I40690,I40707,I65519,I40747,I40755,I40772,I40789,I40806,I40837,I65498,I40854,I40880,I40888,I40919,I40950,I40967,I40998,I65516,I41098,I41124,I41132,I41149,I41166,I41192,I41200,I41226,I41234,I41251,I41268,I41285,I41325,I41333,I41350,I41367,I41384,I41415,I41432,I41458,I41466,I41497,I41528,I41545,I41576,I41676,I41702,I41710,I41727,I41744,I41770,I41778,I41804,I41812,I41829,I41846,I41863,I41903,I41911,I41928,I41945,I41962,I41993,I42010,I42036,I42044,I42075,I42106,I42123,I42154,I42254,I42280,I42288,I42305,I42322,I42348,I42356,I42382,I42390,I42407,I42424,I42441,I42237,I42481,I42489,I42506,I42523,I42540,I42240,I42571,I42588,I42614,I42622,I42222,I42653,I42231,I42684,I42701,I42243,I42732,I42234,I42225,I42228,I42246,I42832,I53313,I42858,I42866,I42883,I53289,I53304,I42900,I53316,I42926,I42934,I53301,I53292,I42960,I42968,I42985,I43002,I43019,I42815,I43059,I43067,I43084,I43101,I43118,I42818,I43149,I53307,I53298,I43166,I53310,I43192,I43200,I42800,I43231,I42809,I43262,I43279,I42821,I43310,I53295,I42812,I42803,I42806,I42824,I43410,I67247,I43436,I43444,I43461,I67229,I67241,I43478,I67244,I43504,I43512,I67238,I67235,I43538,I43546,I43563,I43580,I43597,I67253,I43637,I43645,I43662,I43679,I43696,I43727,I67232,I43744,I43770,I43778,I43809,I43840,I43857,I43888,I67250,I43988,I44014,I44022,I44039,I44056,I44082,I44090,I44116,I44124,I44141,I44158,I44175,I44215,I44223,I44240,I44257,I44274,I44305,I44322,I44348,I44356,I44387,I44418,I44435,I44466,I44566,I44592,I44600,I44617,I44634,I44660,I44668,I44694,I44702,I44719,I44736,I44753,I44549,I44793,I44801,I44818,I44835,I44852,I44552,I44883,I44900,I44926,I44934,I44534,I44965,I44543,I44996,I45013,I44555,I45044,I44546,I44537,I44540,I44558,I45144,I75185,I45170,I45178,I45195,I75209,I75191,I45212,I75197,I45238,I45246,I75203,I75188,I45272,I45280,I45297,I45314,I45331,I45127,I75200,I45371,I45379,I45396,I45413,I45430,I45130,I45461,I75206,I75194,I45478,I45504,I45512,I45112,I45543,I45121,I45574,I45591,I45133,I45622,I45124,I45115,I45118,I45136,I45722,I64935,I45748,I45756,I45773,I64917,I64929,I45790,I64932,I45816,I45824,I64926,I64923,I45850,I45858,I45875,I45892,I45909,I45705,I64941,I45949,I45957,I45974,I45991,I46008,I45708,I46039,I64920,I46056,I46082,I46090,I45690,I46121,I45699,I46152,I46169,I45711,I46200,I64938,I45702,I45693,I45696,I45714,I46300,I46326,I46334,I46351,I46368,I46394,I46402,I46428,I46436,I46453,I46470,I46487,I46283,I46527,I46535,I46552,I46569,I46586,I46286,I46617,I46634,I46660,I46668,I46268,I46699,I46277,I46730,I46747,I46289,I46778,I46280,I46271,I46274,I46292,I46875,I64357,I46901,I46909,I46926,I64339,I46943,I64345,I46969,I64342,I47000,I47008,I64351,I47025,I47051,I47059,I64363,I47099,I47135,I64354,I64348,I47152,I47178,I47186,I47203,I47234,I64360,I47251,I47268,I47299,I47330,I47347,I47402,I47428,I47436,I47453,I47470,I47496,I47527,I47535,I47552,I47578,I47586,I47626,I47662,I47679,I47705,I47713,I47730,I47761,I47778,I47795,I47826,I47857,I47874,I47929,I47955,I47963,I47980,I47997,I48023,I48054,I48062,I48079,I48105,I48113,I48153,I48189,I48206,I48232,I48240,I48257,I48288,I48305,I48322,I48353,I48384,I48401,I48456,I48482,I48490,I48507,I48524,I48550,I48445,I48581,I48589,I48606,I48632,I48640,I48448,I48680,I48439,I48430,I48716,I48733,I48759,I48767,I48784,I48433,I48815,I48832,I48849,I48442,I48880,I48427,I48911,I48928,I48436,I48983,I49009,I49017,I49034,I49051,I49077,I49108,I49116,I49133,I49159,I49167,I49207,I49243,I49260,I49286,I49294,I49311,I49342,I49359,I49376,I49407,I49438,I49455,I49510,I57814,I49536,I49544,I49561,I57829,I57811,I49578,I49604,I49499,I57820,I49635,I49643,I57838,I49660,I49686,I49694,I49502,I57835,I49734,I49493,I49484,I49770,I57832,I57823,I49787,I57817,I49813,I49821,I49838,I49487,I49869,I57826,I49886,I49903,I49496,I49934,I49481,I49965,I49982,I49490,I50037,I50063,I50071,I50088,I50105,I50131,I50162,I50170,I50187,I50213,I50221,I50261,I50297,I50314,I50340,I50348,I50365,I50396,I50413,I50430,I50461,I50492,I50509,I50564,I50590,I50598,I50615,I50632,I50658,I50553,I50689,I50697,I50714,I50740,I50748,I50556,I50788,I50547,I50538,I50824,I50841,I50867,I50875,I50892,I50541,I50923,I50940,I50957,I50550,I50988,I50535,I51019,I51036,I50544,I51091,I51117,I51125,I51142,I51159,I51185,I51080,I51216,I51224,I51241,I51267,I51275,I51083,I51315,I51074,I51065,I51351,I51368,I51394,I51402,I51419,I51068,I51450,I51467,I51484,I51077,I51515,I51062,I51546,I51563,I51071,I51618,I72449,I51644,I51652,I51669,I72431,I51686,I72437,I51712,I72434,I51743,I51751,I72443,I51768,I51794,I51802,I72455,I51842,I51878,I72446,I72440,I51895,I51921,I51929,I51946,I51977,I72452,I51994,I52011,I52042,I52073,I52090,I52145,I52171,I52179,I52196,I52213,I52239,I52134,I52270,I52278,I52295,I52321,I52329,I52137,I52369,I52128,I52119,I52405,I52422,I52448,I52456,I52473,I52122,I52504,I52521,I52538,I52131,I52569,I52116,I52600,I52617,I52125,I52678,I52704,I52721,I52729,I52746,I52763,I52780,I52797,I52814,I52845,I52862,I52893,I52910,I52927,I52958,I52998,I53006,I53023,I53040,I53057,I53088,I53105,I53122,I53148,I53170,I53187,I53218,I53263,I53324,I81611,I53350,I81635,I53367,I53375,I53392,I81617,I53409,I81626,I53426,I53443,I81632,I53460,I53491,I53508,I53539,I53556,I81629,I53573,I53604,I53644,I53652,I53669,I53686,I81623,I53703,I53734,I81614,I53751,I81638,I53768,I81620,I53794,I53816,I53833,I53864,I53909,I53970,I53996,I54013,I54021,I54038,I54055,I54072,I54089,I54106,I54137,I54154,I54185,I54202,I54219,I54250,I54290,I54298,I54315,I54332,I54349,I54380,I54397,I54414,I54440,I54462,I54479,I54510,I54555,I54616,I78041,I54642,I78065,I54659,I54667,I54684,I78047,I54701,I78056,I54718,I54735,I78062,I54752,I54783,I54800,I54831,I54848,I78059,I54865,I54896,I54936,I54944,I54961,I54978,I78053,I54995,I55026,I78044,I55043,I78068,I55060,I78050,I55086,I55108,I55125,I55156,I55201,I55262,I66091,I55288,I66073,I55305,I55313,I55330,I66082,I55347,I66094,I55364,I66076,I55381,I66085,I55398,I55429,I55446,I55477,I55494,I66097,I55511,I55542,I55582,I55590,I55607,I55624,I55641,I55672,I66079,I55689,I66088,I55706,I55732,I55754,I55771,I55802,I55847,I55908,I80421,I55934,I80445,I55951,I55959,I55976,I80427,I55993,I80436,I56010,I56027,I80442,I56044,I56075,I56092,I56123,I56140,I80439,I56157,I56188,I56228,I56236,I56253,I56270,I80433,I56287,I56318,I80424,I56335,I80448,I56352,I80430,I56378,I56400,I56417,I56448,I56493,I56554,I56580,I56597,I56605,I56622,I56639,I56656,I56673,I56690,I56721,I56738,I56769,I56786,I56803,I56834,I56874,I56882,I56899,I56916,I56933,I56964,I56981,I56998,I57024,I57046,I57063,I57094,I57139,I57200,I57226,I57243,I57251,I57268,I57285,I57302,I57319,I57336,I57186,I57367,I57384,I57189,I57415,I57432,I57449,I57165,I57480,I57177,I57520,I57528,I57545,I57562,I57579,I57192,I57610,I57627,I57644,I57670,I57180,I57692,I57709,I57174,I57740,I57168,I57171,I57785,I57183,I57846,I57872,I57889,I57897,I57914,I57931,I57948,I57965,I57982,I58013,I58030,I58061,I58078,I58095,I58126,I58166,I58174,I58191,I58208,I58225,I58256,I58273,I58290,I58316,I58338,I58355,I58386,I58431,I58492,I58518,I58535,I58543,I58560,I58577,I58594,I58611,I58628,I58659,I58676,I58707,I58724,I58741,I58772,I58812,I58820,I58837,I58854,I58871,I58902,I58919,I58936,I58962,I58984,I59001,I59032,I59077,I59138,I59164,I59181,I59189,I59206,I59223,I59240,I59257,I59274,I59305,I59322,I59353,I59370,I59387,I59418,I59458,I59466,I59483,I59500,I59517,I59548,I59565,I59582,I59608,I59630,I59647,I59678,I59723,I59784,I59810,I59827,I59835,I59852,I59869,I59886,I59903,I59920,I59770,I59951,I59968,I59773,I59999,I60016,I60033,I59749,I60064,I59761,I60104,I60112,I60129,I60146,I60163,I59776,I60194,I60211,I60228,I60254,I59764,I60276,I60293,I59758,I60324,I59752,I59755,I60369,I59767,I60424,I60450,I60467,I60489,I60515,I60523,I60540,I60557,I60574,I60591,I60608,I60625,I60656,I60687,I60704,I60721,I60738,I60769,I60814,I60831,I60848,I60874,I60882,I60913,I60930,I60985,I67822,I61011,I61028,I60977,I61050,I67813,I61076,I61084,I67810,I61101,I61118,I67819,I61135,I67828,I61152,I61169,I67807,I61186,I60959,I61217,I60962,I61248,I67816,I61265,I61282,I61299,I60971,I61330,I60974,I60968,I61375,I67831,I61392,I61409,I67825,I61435,I61443,I60956,I61474,I61491,I60965,I61546,I61572,I61589,I61538,I61611,I61637,I61645,I61662,I61679,I61696,I61713,I61730,I61747,I61520,I61778,I61523,I61809,I61826,I61843,I61860,I61532,I61891,I61535,I61529,I61936,I61953,I61970,I61996,I62004,I61517,I62035,I62052,I61526,I62107,I62133,I62150,I62172,I62198,I62206,I62223,I62240,I62257,I62274,I62291,I62308,I62339,I62370,I62387,I62404,I62421,I62452,I62497,I62514,I62531,I62557,I62565,I62596,I62613,I62668,I73559,I62694,I62711,I62660,I62733,I73565,I62759,I62767,I73574,I62784,I62801,I73553,I62818,I73556,I62835,I62852,I73568,I62869,I62642,I62900,I62645,I62931,I73562,I62948,I62965,I62982,I62654,I63013,I62657,I62651,I63058,I73577,I63075,I63092,I73571,I63118,I63126,I62639,I63157,I63174,I62648,I63229,I63255,I63272,I63221,I63294,I63320,I63328,I63345,I63362,I63379,I63396,I63413,I63430,I63203,I63461,I63206,I63492,I63509,I63526,I63543,I63215,I63574,I63218,I63212,I63619,I63636,I63653,I63679,I63687,I63200,I63718,I63735,I63209,I63793,I63819,I63827,I63867,I63875,I63892,I63909,I63949,I63971,I63988,I64014,I64022,I64039,I64056,I64073,I64090,I64135,I64166,I64183,I64209,I64217,I64248,I64265,I64282,I64299,I64371,I64397,I64405,I64445,I64453,I64470,I64487,I64527,I64549,I64566,I64592,I64600,I64617,I64634,I64651,I64668,I64713,I64744,I64761,I64787,I64795,I64826,I64843,I64860,I64877,I64949,I64975,I64983,I65023,I65031,I65048,I65065,I65105,I65127,I65144,I65170,I65178,I65195,I65212,I65229,I65246,I65291,I65322,I65339,I65365,I65373,I65404,I65421,I65438,I65455,I65527,I65553,I65561,I65601,I65609,I65626,I65643,I65683,I65705,I65722,I65748,I65756,I65773,I65790,I65807,I65824,I65869,I65900,I65917,I65943,I65951,I65982,I65999,I66016,I66033,I66105,I66131,I66139,I66179,I66187,I66204,I66221,I66261,I66283,I66300,I66326,I66334,I66351,I66368,I66385,I66402,I66447,I66478,I66495,I66521,I66529,I66560,I66577,I66594,I66611,I66683,I66709,I66717,I66757,I66765,I66782,I66799,I66839,I66861,I66878,I66904,I66912,I66929,I66946,I66963,I66980,I67025,I67056,I67073,I67099,I67107,I67138,I67155,I67172,I67189,I67261,I67287,I67295,I67335,I67343,I67360,I67377,I67417,I67439,I67456,I67482,I67490,I67507,I67524,I67541,I67558,I67603,I67634,I67651,I67677,I67685,I67716,I67733,I67750,I67767,I67839,I67865,I67873,I67913,I67921,I67938,I67955,I67995,I68017,I68034,I68060,I68068,I68085,I68102,I68119,I68136,I68181,I68212,I68229,I68255,I68263,I68294,I68311,I68328,I68345,I68417,I83423,I68443,I68451,I83405,I83396,I68491,I68499,I83411,I68516,I83399,I68533,I68573,I68595,I83408,I68612,I68638,I68646,I68663,I83417,I68680,I68697,I68714,I68759,I83420,I68790,I68807,I83414,I83402,I68833,I68841,I68872,I68889,I68906,I68923,I68995,I78663,I69021,I69029,I78645,I78636,I69069,I69077,I78651,I69094,I78639,I69111,I69151,I69173,I78648,I69190,I69216,I69224,I69241,I78657,I69258,I69275,I69292,I69337,I78660,I69368,I69385,I78654,I78642,I69411,I69419,I69450,I69467,I69484,I69501,I69573,I69599,I69607,I69647,I69655,I69672,I69689,I69729,I69751,I69768,I69794,I69802,I69819,I69836,I69853,I69870,I69915,I69946,I69963,I69989,I69997,I70028,I70045,I70062,I70079,I70151,I70177,I70185,I70225,I70233,I70250,I70267,I70307,I70329,I70346,I70372,I70380,I70397,I70414,I70431,I70448,I70493,I70524,I70541,I70567,I70575,I70606,I70623,I70640,I70657,I70729,I70755,I70763,I70803,I70811,I70828,I70845,I70885,I70907,I70924,I70950,I70958,I70975,I70992,I71009,I71026,I71071,I71102,I71119,I71145,I71153,I71184,I71201,I71218,I71235,I71307,I71333,I71341,I71381,I71389,I71406,I71423,I71463,I71485,I71502,I71528,I71536,I71553,I71570,I71587,I71604,I71649,I71680,I71697,I71723,I71731,I71762,I71779,I71796,I71813,I71885,I71911,I71919,I71959,I71967,I71984,I72001,I72041,I72063,I72080,I72106,I72114,I72131,I72148,I72165,I72182,I72227,I72258,I72275,I72301,I72309,I72340,I72357,I72374,I72391,I72463,I72489,I72497,I72537,I72545,I72562,I72579,I72619,I72641,I72658,I72684,I72692,I72709,I72726,I72743,I72760,I72805,I72836,I72853,I72879,I72887,I72918,I72935,I72952,I72969,I73041,I73067,I73075,I73101,I73118,I73033,I73140,I73157,I73174,I73191,I73208,I73012,I73239,I73256,I73273,I73290,I73015,I73030,I73335,I73352,I73369,I73027,I73024,I73021,I73428,I73454,I73462,I73479,I73496,I73009,I73527,I73018,I73585,I73611,I73619,I73645,I73662,I73684,I73701,I73718,I73735,I73752,I73783,I73800,I73817,I73834,I73879,I73896,I73913,I73972,I73998,I74006,I74023,I74040,I74071,I74129,I74155,I74163,I74189,I74206,I74228,I74245,I74262,I74279,I74296,I74327,I74344,I74361,I74378,I74423,I74440,I74457,I74516,I74542,I74550,I74567,I74584,I74615,I74673,I74699,I74707,I74733,I74750,I74772,I74789,I74806,I74823,I74840,I74871,I74888,I74905,I74922,I74967,I74984,I75001,I75060,I75086,I75094,I75111,I75128,I75159,I75217,I77498,I75243,I75251,I77492,I75268,I77507,I75294,I75302,I75319,I77483,I75336,I77480,I75353,I75370,I77486,I75401,I75418,I77495,I75435,I75466,I77489,I75483,I75523,I75531,I75562,I77504,I75579,I75596,I75613,I75644,I75675,I77501,I75701,I75723,I75795,I75821,I75829,I75846,I75872,I75880,I75897,I75914,I75931,I75948,I75979,I75996,I76013,I76044,I76061,I76101,I76109,I76140,I76157,I76174,I76191,I76222,I76253,I76279,I76301,I76373,I76399,I76407,I76424,I76450,I76458,I76475,I76492,I76509,I76526,I76557,I76574,I76591,I76622,I76639,I76679,I76687,I76718,I76735,I76752,I76769,I76800,I76831,I76857,I76879,I76954,I76980,I76988,I77005,I77031,I77039,I77056,I77073,I77104,I77135,I77152,I77169,I77186,I77203,I77234,I77293,I77310,I77336,I77358,I77384,I77392,I77409,I77440,I77515,I77541,I77549,I77566,I77592,I77600,I77617,I77634,I77665,I77696,I77713,I77730,I77747,I77764,I77795,I77854,I77871,I77897,I77919,I77945,I77953,I77970,I78001,I78076,I78102,I78119,I78127,I78172,I78189,I78206,I78223,I78240,I78257,I78274,I78305,I78322,I78367,I78384,I78401,I78432,I78458,I78466,I78497,I78514,I78531,I78557,I78565,I78582,I78671,I78697,I78714,I78722,I78767,I78784,I78801,I78818,I78835,I78852,I78869,I78900,I78917,I78962,I78979,I78996,I79027,I79053,I79061,I79092,I79109,I79126,I79152,I79160,I79177,I79266,I79292,I79309,I79317,I79362,I79379,I79396,I79413,I79430,I79447,I79464,I79495,I79512,I79557,I79574,I79591,I79622,I79648,I79656,I79687,I79704,I79721,I79747,I79755,I79772,I79861,I79887,I79904,I79912,I79957,I79974,I79991,I80008,I80025,I80042,I80059,I80090,I80107,I80152,I80169,I80186,I80217,I80243,I80251,I80282,I80299,I80316,I80342,I80350,I80367,I80456,I80482,I80499,I80507,I80552,I80569,I80586,I80603,I80620,I80637,I80654,I80685,I80702,I80747,I80764,I80781,I80812,I80838,I80846,I80877,I80894,I80911,I80937,I80945,I80962,I81051,I81077,I81094,I81102,I81147,I81164,I81181,I81198,I81215,I81232,I81249,I81280,I81297,I81342,I81359,I81376,I81407,I81433,I81441,I81472,I81489,I81506,I81532,I81540,I81557,I81646,I81672,I81689,I81697,I81742,I81759,I81776,I81793,I81810,I81827,I81844,I81875,I81892,I81937,I81954,I81971,I82002,I82028,I82036,I82067,I82084,I82101,I82127,I82135,I82152,I82241,I82267,I82284,I82292,I82337,I82354,I82371,I82388,I82405,I82422,I82439,I82470,I82487,I82532,I82549,I82566,I82597,I82623,I82631,I82662,I82679,I82696,I82722,I82730,I82747,I82836,I82862,I82879,I82887,I82932,I82949,I82966,I82983,I83000,I83017,I83034,I83065,I83082,I83127,I83144,I83161,I83192,I83218,I83226,I83257,I83274,I83291,I83317,I83325,I83342,I83431,I83457,I83474,I83482,I83527,I83544,I83561,I83578,I83595,I83612,I83629,I83660,I83677,I83722,I83739,I83756,I83787,I83813,I83821,I83852,I83869,I83886,I83912,I83920,I83937;
not I_0 (I1845,I1810);
DFFARX1 I_1 (I82206,I1803,I1845,I1871,);
DFFARX1 I_2 (I1871,I1803,I1845,I1888,);
not I_3 (I1896,I1888);
nand I_4 (I1913,I82209,I82215);
and I_5 (I1930,I1913,I82224);
DFFARX1 I_6 (I1930,I1803,I1845,I1956,);
DFFARX1 I_7 (I1956,I1803,I1845,I1837,);
DFFARX1 I_8 (I1956,I1803,I1845,I1828,);
DFFARX1 I_9 (I82227,I1803,I1845,I2001,);
nand I_10 (I2009,I2001,I82218);
not I_11 (I2026,I2009);
nor I_12 (I1825,I1871,I2026);
DFFARX1 I_13 (I82206,I1803,I1845,I2066,);
not I_14 (I2074,I2066);
nor I_15 (I1831,I2074,I1896);
nand I_16 (I1819,I2074,I2009);
nand I_17 (I2119,I82233,I82212);
and I_18 (I2136,I2119,I82221);
DFFARX1 I_19 (I2136,I1803,I1845,I2162,);
nor I_20 (I2170,I2162,I1871);
DFFARX1 I_21 (I2170,I1803,I1845,I1813,);
not I_22 (I2201,I2162);
nor I_23 (I2218,I82230,I82212);
not I_24 (I2235,I2218);
nor I_25 (I2252,I2009,I2235);
nor I_26 (I2269,I2201,I2252);
DFFARX1 I_27 (I2269,I1803,I1845,I1834,);
nor I_28 (I2300,I2162,I2235);
nor I_29 (I1822,I2026,I2300);
nor I_30 (I1816,I2162,I2218);
not I_31 (I2372,I1810);
DFFARX1 I_32 (I39338,I1803,I2372,I2398,);
DFFARX1 I_33 (I2398,I1803,I2372,I2415,);
not I_34 (I2423,I2415);
nand I_35 (I2440,I39353,I39356);
and I_36 (I2457,I2440,I39335);
DFFARX1 I_37 (I2457,I1803,I2372,I2483,);
DFFARX1 I_38 (I2483,I1803,I2372,I2364,);
DFFARX1 I_39 (I2483,I1803,I2372,I2355,);
DFFARX1 I_40 (I39341,I1803,I2372,I2528,);
nand I_41 (I2536,I2528,I39347);
not I_42 (I2553,I2536);
nor I_43 (I2352,I2398,I2553);
DFFARX1 I_44 (I39335,I1803,I2372,I2593,);
not I_45 (I2601,I2593);
nor I_46 (I2358,I2601,I2423);
nand I_47 (I2346,I2601,I2536);
nand I_48 (I2646,I39350,I39332);
and I_49 (I2663,I2646,I39344);
DFFARX1 I_50 (I2663,I1803,I2372,I2689,);
nor I_51 (I2697,I2689,I2398);
DFFARX1 I_52 (I2697,I1803,I2372,I2340,);
not I_53 (I2728,I2689);
nor I_54 (I2745,I39332,I39332);
not I_55 (I2762,I2745);
nor I_56 (I2779,I2536,I2762);
nor I_57 (I2796,I2728,I2779);
DFFARX1 I_58 (I2796,I1803,I2372,I2361,);
nor I_59 (I2827,I2689,I2762);
nor I_60 (I2349,I2553,I2827);
nor I_61 (I2343,I2689,I2745);
not I_62 (I2899,I1810);
DFFARX1 I_63 (I79826,I1803,I2899,I2925,);
DFFARX1 I_64 (I2925,I1803,I2899,I2942,);
not I_65 (I2950,I2942);
nand I_66 (I2967,I79829,I79835);
and I_67 (I2984,I2967,I79844);
DFFARX1 I_68 (I2984,I1803,I2899,I3010,);
DFFARX1 I_69 (I3010,I1803,I2899,I2891,);
DFFARX1 I_70 (I3010,I1803,I2899,I2882,);
DFFARX1 I_71 (I79847,I1803,I2899,I3055,);
nand I_72 (I3063,I3055,I79838);
not I_73 (I3080,I3063);
nor I_74 (I2879,I2925,I3080);
DFFARX1 I_75 (I79826,I1803,I2899,I3120,);
not I_76 (I3128,I3120);
nor I_77 (I2885,I3128,I2950);
nand I_78 (I2873,I3128,I3063);
nand I_79 (I3173,I79853,I79832);
and I_80 (I3190,I3173,I79841);
DFFARX1 I_81 (I3190,I1803,I2899,I3216,);
nor I_82 (I3224,I3216,I2925);
DFFARX1 I_83 (I3224,I1803,I2899,I2867,);
not I_84 (I3255,I3216);
nor I_85 (I3272,I79850,I79832);
not I_86 (I3289,I3272);
nor I_87 (I3306,I3063,I3289);
nor I_88 (I3323,I3255,I3306);
DFFARX1 I_89 (I3323,I1803,I2899,I2888,);
nor I_90 (I3354,I3216,I3289);
nor I_91 (I2876,I3080,I3354);
nor I_92 (I2870,I3216,I3272);
not I_93 (I3426,I1810);
DFFARX1 I_94 (I6559,I1803,I3426,I3452,);
DFFARX1 I_95 (I3452,I1803,I3426,I3469,);
not I_96 (I3477,I3469);
nand I_97 (I3494,I6559,I6574);
and I_98 (I3511,I3494,I6577);
DFFARX1 I_99 (I3511,I1803,I3426,I3537,);
DFFARX1 I_100 (I3537,I1803,I3426,I3418,);
DFFARX1 I_101 (I3537,I1803,I3426,I3409,);
DFFARX1 I_102 (I6571,I1803,I3426,I3582,);
nand I_103 (I3590,I3582,I6580);
not I_104 (I3607,I3590);
nor I_105 (I3406,I3452,I3607);
DFFARX1 I_106 (I6556,I1803,I3426,I3647,);
not I_107 (I3655,I3647);
nor I_108 (I3412,I3655,I3477);
nand I_109 (I3400,I3655,I3590);
nand I_110 (I3700,I6556,I6562);
and I_111 (I3717,I3700,I6565);
DFFARX1 I_112 (I3717,I1803,I3426,I3743,);
nor I_113 (I3751,I3743,I3452);
DFFARX1 I_114 (I3751,I1803,I3426,I3394,);
not I_115 (I3782,I3743);
nor I_116 (I3799,I6568,I6562);
not I_117 (I3816,I3799);
nor I_118 (I3833,I3590,I3816);
nor I_119 (I3850,I3782,I3833);
DFFARX1 I_120 (I3850,I1803,I3426,I3415,);
nor I_121 (I3881,I3743,I3816);
nor I_122 (I3403,I3607,I3881);
nor I_123 (I3397,I3743,I3799);
not I_124 (I3953,I1810);
DFFARX1 I_125 (I1684,I1803,I3953,I3979,);
DFFARX1 I_126 (I3979,I1803,I3953,I3996,);
not I_127 (I4004,I3996);
nand I_128 (I4021,I1764,I1756);
and I_129 (I4038,I4021,I1404);
DFFARX1 I_130 (I4038,I1803,I3953,I4064,);
DFFARX1 I_131 (I4064,I1803,I3953,I3945,);
DFFARX1 I_132 (I4064,I1803,I3953,I3936,);
DFFARX1 I_133 (I1588,I1803,I3953,I4109,);
nand I_134 (I4117,I4109,I1524);
not I_135 (I4134,I4117);
nor I_136 (I3933,I3979,I4134);
DFFARX1 I_137 (I1372,I1803,I3953,I4174,);
not I_138 (I4182,I4174);
nor I_139 (I3939,I4182,I4004);
nand I_140 (I3927,I4182,I4117);
nand I_141 (I4227,I1644,I1636);
and I_142 (I4244,I4227,I1652);
DFFARX1 I_143 (I4244,I1803,I3953,I4270,);
nor I_144 (I4278,I4270,I3979);
DFFARX1 I_145 (I4278,I1803,I3953,I3921,);
not I_146 (I4309,I4270);
nor I_147 (I4326,I1444,I1636);
not I_148 (I4343,I4326);
nor I_149 (I4360,I4117,I4343);
nor I_150 (I4377,I4309,I4360);
DFFARX1 I_151 (I4377,I1803,I3953,I3942,);
nor I_152 (I4408,I4270,I4343);
nor I_153 (I3930,I4134,I4408);
nor I_154 (I3924,I4270,I4326);
not I_155 (I4480,I1810);
DFFARX1 I_156 (I40494,I1803,I4480,I4506,);
DFFARX1 I_157 (I4506,I1803,I4480,I4523,);
not I_158 (I4531,I4523);
nand I_159 (I4548,I40509,I40512);
and I_160 (I4565,I4548,I40491);
DFFARX1 I_161 (I4565,I1803,I4480,I4591,);
DFFARX1 I_162 (I4591,I1803,I4480,I4472,);
DFFARX1 I_163 (I4591,I1803,I4480,I4463,);
DFFARX1 I_164 (I40497,I1803,I4480,I4636,);
nand I_165 (I4644,I4636,I40503);
not I_166 (I4661,I4644);
nor I_167 (I4460,I4506,I4661);
DFFARX1 I_168 (I40491,I1803,I4480,I4701,);
not I_169 (I4709,I4701);
nor I_170 (I4466,I4709,I4531);
nand I_171 (I4454,I4709,I4644);
nand I_172 (I4754,I40506,I40488);
and I_173 (I4771,I4754,I40500);
DFFARX1 I_174 (I4771,I1803,I4480,I4797,);
nor I_175 (I4805,I4797,I4506);
DFFARX1 I_176 (I4805,I1803,I4480,I4448,);
not I_177 (I4836,I4797);
nor I_178 (I4853,I40488,I40488);
not I_179 (I4870,I4853);
nor I_180 (I4887,I4644,I4870);
nor I_181 (I4904,I4836,I4887);
DFFARX1 I_182 (I4904,I1803,I4480,I4469,);
nor I_183 (I4935,I4797,I4870);
nor I_184 (I4457,I4661,I4935);
nor I_185 (I4451,I4797,I4853);
not I_186 (I5007,I1810);
DFFARX1 I_187 (I18653,I1803,I5007,I5033,);
not I_188 (I5041,I5033);
nand I_189 (I5058,I18635,I18650);
and I_190 (I5075,I5058,I18626);
DFFARX1 I_191 (I5075,I1803,I5007,I5101,);
DFFARX1 I_192 (I18629,I1803,I5007,I5118,);
and I_193 (I5126,I5118,I18644);
nor I_194 (I5143,I5101,I5126);
DFFARX1 I_195 (I5143,I1803,I5007,I4975,);
nand I_196 (I5174,I5118,I18644);
nand I_197 (I5191,I5041,I5174);
not I_198 (I4987,I5191);
DFFARX1 I_199 (I18647,I1803,I5007,I5231,);
DFFARX1 I_200 (I5231,I1803,I5007,I4996,);
nand I_201 (I5253,I18626,I18638);
and I_202 (I5270,I5253,I18632);
DFFARX1 I_203 (I5270,I1803,I5007,I5296,);
DFFARX1 I_204 (I5296,I1803,I5007,I5313,);
not I_205 (I4999,I5313);
not I_206 (I5335,I5296);
nand I_207 (I4984,I5335,I5174);
nor I_208 (I5366,I18641,I18638);
not I_209 (I5383,I5366);
nor I_210 (I5400,I5335,I5383);
nor I_211 (I5417,I5041,I5400);
DFFARX1 I_212 (I5417,I1803,I5007,I4993,);
nor I_213 (I5448,I5101,I5383);
nor I_214 (I4981,I5296,I5448);
nor I_215 (I4990,I5231,I5366);
nor I_216 (I4978,I5101,I5366);
not I_217 (I5534,I1810);
DFFARX1 I_218 (I26651,I1803,I5534,I5560,);
not I_219 (I5568,I5560);
nand I_220 (I5585,I26645,I26636);
and I_221 (I5602,I5585,I26657);
DFFARX1 I_222 (I5602,I1803,I5534,I5628,);
DFFARX1 I_223 (I26639,I1803,I5534,I5645,);
and I_224 (I5653,I5645,I26633);
nor I_225 (I5670,I5628,I5653);
DFFARX1 I_226 (I5670,I1803,I5534,I5502,);
nand I_227 (I5701,I5645,I26633);
nand I_228 (I5718,I5568,I5701);
not I_229 (I5514,I5718);
DFFARX1 I_230 (I26633,I1803,I5534,I5758,);
DFFARX1 I_231 (I5758,I1803,I5534,I5523,);
nand I_232 (I5780,I26660,I26642);
and I_233 (I5797,I5780,I26648);
DFFARX1 I_234 (I5797,I1803,I5534,I5823,);
DFFARX1 I_235 (I5823,I1803,I5534,I5840,);
not I_236 (I5526,I5840);
not I_237 (I5862,I5823);
nand I_238 (I5511,I5862,I5701);
nor I_239 (I5893,I26654,I26642);
not I_240 (I5910,I5893);
nor I_241 (I5927,I5862,I5910);
nor I_242 (I5944,I5568,I5927);
DFFARX1 I_243 (I5944,I1803,I5534,I5520,);
nor I_244 (I5975,I5628,I5910);
nor I_245 (I5508,I5823,I5975);
nor I_246 (I5517,I5758,I5893);
nor I_247 (I5505,I5628,I5893);
not I_248 (I6061,I1810);
DFFARX1 I_249 (I60398,I1803,I6061,I6087,);
not I_250 (I6095,I6087);
nand I_251 (I6112,I60395,I60401);
and I_252 (I6129,I6112,I60398);
DFFARX1 I_253 (I6129,I1803,I6061,I6155,);
DFFARX1 I_254 (I60401,I1803,I6061,I6172,);
and I_255 (I6180,I6172,I60395);
nor I_256 (I6197,I6155,I6180);
DFFARX1 I_257 (I6197,I1803,I6061,I6029,);
nand I_258 (I6228,I6172,I60395);
nand I_259 (I6245,I6095,I6228);
not I_260 (I6041,I6245);
DFFARX1 I_261 (I60404,I1803,I6061,I6285,);
DFFARX1 I_262 (I6285,I1803,I6061,I6050,);
nand I_263 (I6307,I60407,I60416);
and I_264 (I6324,I6307,I60410);
DFFARX1 I_265 (I6324,I1803,I6061,I6350,);
DFFARX1 I_266 (I6350,I1803,I6061,I6367,);
not I_267 (I6053,I6367);
not I_268 (I6389,I6350);
nand I_269 (I6038,I6389,I6228);
nor I_270 (I6420,I60413,I60416);
not I_271 (I6437,I6420);
nor I_272 (I6454,I6389,I6437);
nor I_273 (I6471,I6095,I6454);
DFFARX1 I_274 (I6471,I1803,I6061,I6047,);
nor I_275 (I6502,I6155,I6437);
nor I_276 (I6035,I6350,I6502);
nor I_277 (I6044,I6285,I6420);
nor I_278 (I6032,I6155,I6420);
not I_279 (I6588,I1810);
DFFARX1 I_280 (I46855,I1803,I6588,I6614,);
not I_281 (I6622,I6614);
nand I_282 (I6639,I46852,I46867);
and I_283 (I6656,I6639,I46849);
DFFARX1 I_284 (I6656,I1803,I6588,I6682,);
DFFARX1 I_285 (I46846,I1803,I6588,I6699,);
and I_286 (I6707,I6699,I46846);
nor I_287 (I6724,I6682,I6707);
DFFARX1 I_288 (I6724,I1803,I6588,I6556,);
nand I_289 (I6755,I6699,I46846);
nand I_290 (I6772,I6622,I6755);
not I_291 (I6568,I6772);
DFFARX1 I_292 (I46849,I1803,I6588,I6812,);
DFFARX1 I_293 (I6812,I1803,I6588,I6577,);
nand I_294 (I6834,I46861,I46852);
and I_295 (I6851,I6834,I46864);
DFFARX1 I_296 (I6851,I1803,I6588,I6877,);
DFFARX1 I_297 (I6877,I1803,I6588,I6894,);
not I_298 (I6580,I6894);
not I_299 (I6916,I6877);
nand I_300 (I6565,I6916,I6755);
nor I_301 (I6947,I46858,I46852);
not I_302 (I6964,I6947);
nor I_303 (I6981,I6916,I6964);
nor I_304 (I6998,I6622,I6981);
DFFARX1 I_305 (I6998,I1803,I6588,I6574,);
nor I_306 (I7029,I6682,I6964);
nor I_307 (I6562,I6877,I7029);
nor I_308 (I6571,I6812,I6947);
nor I_309 (I6559,I6682,I6947);
not I_310 (I7115,I1810);
DFFARX1 I_311 (I15491,I1803,I7115,I7141,);
not I_312 (I7149,I7141);
nand I_313 (I7166,I15473,I15488);
and I_314 (I7183,I7166,I15464);
DFFARX1 I_315 (I7183,I1803,I7115,I7209,);
DFFARX1 I_316 (I15467,I1803,I7115,I7226,);
and I_317 (I7234,I7226,I15482);
nor I_318 (I7251,I7209,I7234);
DFFARX1 I_319 (I7251,I1803,I7115,I7083,);
nand I_320 (I7282,I7226,I15482);
nand I_321 (I7299,I7149,I7282);
not I_322 (I7095,I7299);
DFFARX1 I_323 (I15485,I1803,I7115,I7339,);
DFFARX1 I_324 (I7339,I1803,I7115,I7104,);
nand I_325 (I7361,I15464,I15476);
and I_326 (I7378,I7361,I15470);
DFFARX1 I_327 (I7378,I1803,I7115,I7404,);
DFFARX1 I_328 (I7404,I1803,I7115,I7421,);
not I_329 (I7107,I7421);
not I_330 (I7443,I7404);
nand I_331 (I7092,I7443,I7282);
nor I_332 (I7474,I15479,I15476);
not I_333 (I7491,I7474);
nor I_334 (I7508,I7443,I7491);
nor I_335 (I7525,I7149,I7508);
DFFARX1 I_336 (I7525,I1803,I7115,I7101,);
nor I_337 (I7556,I7209,I7491);
nor I_338 (I7089,I7404,I7556);
nor I_339 (I7098,I7339,I7474);
nor I_340 (I7086,I7209,I7474);
not I_341 (I7642,I1810);
DFFARX1 I_342 (I54590,I1803,I7642,I7668,);
not I_343 (I7676,I7668);
nand I_344 (I7693,I54608,I54602);
and I_345 (I7710,I7693,I54581);
DFFARX1 I_346 (I7710,I1803,I7642,I7736,);
DFFARX1 I_347 (I54599,I1803,I7642,I7753,);
and I_348 (I7761,I7753,I54584);
nor I_349 (I7778,I7736,I7761);
DFFARX1 I_350 (I7778,I1803,I7642,I7610,);
nand I_351 (I7809,I7753,I54584);
nand I_352 (I7826,I7676,I7809);
not I_353 (I7622,I7826);
DFFARX1 I_354 (I54596,I1803,I7642,I7866,);
DFFARX1 I_355 (I7866,I1803,I7642,I7631,);
nand I_356 (I7888,I54605,I54593);
and I_357 (I7905,I7888,I54587);
DFFARX1 I_358 (I7905,I1803,I7642,I7931,);
DFFARX1 I_359 (I7931,I1803,I7642,I7948,);
not I_360 (I7634,I7948);
not I_361 (I7970,I7931);
nand I_362 (I7619,I7970,I7809);
nor I_363 (I8001,I54581,I54593);
not I_364 (I8018,I8001);
nor I_365 (I8035,I7970,I8018);
nor I_366 (I8052,I7676,I8035);
DFFARX1 I_367 (I8052,I1803,I7642,I7628,);
nor I_368 (I8083,I7736,I8018);
nor I_369 (I7616,I7931,I8083);
nor I_370 (I7625,I7866,I8001);
nor I_371 (I7613,I7736,I8001);
not I_372 (I8169,I1810);
DFFARX1 I_373 (I35873,I1803,I8169,I8195,);
not I_374 (I8203,I8195);
nand I_375 (I8220,I35885,I35870);
and I_376 (I8237,I8220,I35864);
DFFARX1 I_377 (I8237,I1803,I8169,I8263,);
DFFARX1 I_378 (I35879,I1803,I8169,I8280,);
and I_379 (I8288,I8280,I35867);
nor I_380 (I8305,I8263,I8288);
DFFARX1 I_381 (I8305,I1803,I8169,I8137,);
nand I_382 (I8336,I8280,I35867);
nand I_383 (I8353,I8203,I8336);
not I_384 (I8149,I8353);
DFFARX1 I_385 (I35876,I1803,I8169,I8393,);
DFFARX1 I_386 (I8393,I1803,I8169,I8158,);
nand I_387 (I8415,I35882,I35888);
and I_388 (I8432,I8415,I35864);
DFFARX1 I_389 (I8432,I1803,I8169,I8458,);
DFFARX1 I_390 (I8458,I1803,I8169,I8475,);
not I_391 (I8161,I8475);
not I_392 (I8497,I8458);
nand I_393 (I8146,I8497,I8336);
nor I_394 (I8528,I35867,I35888);
not I_395 (I8545,I8528);
nor I_396 (I8562,I8497,I8545);
nor I_397 (I8579,I8203,I8562);
DFFARX1 I_398 (I8579,I1803,I8169,I8155,);
nor I_399 (I8610,I8263,I8545);
nor I_400 (I8143,I8458,I8610);
nor I_401 (I8152,I8393,I8528);
nor I_402 (I8140,I8263,I8528);
not I_403 (I8696,I1810);
DFFARX1 I_404 (I50017,I1803,I8696,I8722,);
not I_405 (I8730,I8722);
nand I_406 (I8747,I50014,I50029);
and I_407 (I8764,I8747,I50011);
DFFARX1 I_408 (I8764,I1803,I8696,I8790,);
DFFARX1 I_409 (I50008,I1803,I8696,I8807,);
and I_410 (I8815,I8807,I50008);
nor I_411 (I8832,I8790,I8815);
DFFARX1 I_412 (I8832,I1803,I8696,I8664,);
nand I_413 (I8863,I8807,I50008);
nand I_414 (I8880,I8730,I8863);
not I_415 (I8676,I8880);
DFFARX1 I_416 (I50011,I1803,I8696,I8920,);
DFFARX1 I_417 (I8920,I1803,I8696,I8685,);
nand I_418 (I8942,I50023,I50014);
and I_419 (I8959,I8942,I50026);
DFFARX1 I_420 (I8959,I1803,I8696,I8985,);
DFFARX1 I_421 (I8985,I1803,I8696,I9002,);
not I_422 (I8688,I9002);
not I_423 (I9024,I8985);
nand I_424 (I8673,I9024,I8863);
nor I_425 (I9055,I50020,I50014);
not I_426 (I9072,I9055);
nor I_427 (I9089,I9024,I9072);
nor I_428 (I9106,I8730,I9089);
DFFARX1 I_429 (I9106,I1803,I8696,I8682,);
nor I_430 (I9137,I8790,I9072);
nor I_431 (I8670,I8985,I9137);
nor I_432 (I8679,I8920,I9055);
nor I_433 (I8667,I8790,I9055);
not I_434 (I9223,I1810);
DFFARX1 I_435 (I79243,I1803,I9223,I9249,);
not I_436 (I9257,I9249);
nand I_437 (I9274,I79237,I79258);
and I_438 (I9291,I9274,I79234);
DFFARX1 I_439 (I9291,I1803,I9223,I9317,);
DFFARX1 I_440 (I79255,I1803,I9223,I9334,);
and I_441 (I9342,I9334,I79252);
nor I_442 (I9359,I9317,I9342);
DFFARX1 I_443 (I9359,I1803,I9223,I9191,);
nand I_444 (I9390,I9334,I79252);
nand I_445 (I9407,I9257,I9390);
not I_446 (I9203,I9407);
DFFARX1 I_447 (I79240,I1803,I9223,I9447,);
DFFARX1 I_448 (I9447,I1803,I9223,I9212,);
nand I_449 (I9469,I79249,I79246);
and I_450 (I9486,I9469,I79231);
DFFARX1 I_451 (I9486,I1803,I9223,I9512,);
DFFARX1 I_452 (I9512,I1803,I9223,I9529,);
not I_453 (I9215,I9529);
not I_454 (I9551,I9512);
nand I_455 (I9200,I9551,I9390);
nor I_456 (I9582,I79231,I79246);
not I_457 (I9599,I9582);
nor I_458 (I9616,I9551,I9599);
nor I_459 (I9633,I9257,I9616);
DFFARX1 I_460 (I9633,I1803,I9223,I9209,);
nor I_461 (I9664,I9317,I9599);
nor I_462 (I9197,I9512,I9664);
nor I_463 (I9206,I9447,I9582);
nor I_464 (I9194,I9317,I9582);
not I_465 (I9750,I1810);
DFFARX1 I_466 (I58466,I1803,I9750,I9776,);
not I_467 (I9784,I9776);
nand I_468 (I9801,I58484,I58478);
and I_469 (I9818,I9801,I58457);
DFFARX1 I_470 (I9818,I1803,I9750,I9844,);
DFFARX1 I_471 (I58475,I1803,I9750,I9861,);
and I_472 (I9869,I9861,I58460);
nor I_473 (I9886,I9844,I9869);
DFFARX1 I_474 (I9886,I1803,I9750,I9718,);
nand I_475 (I9917,I9861,I58460);
nand I_476 (I9934,I9784,I9917);
not I_477 (I9730,I9934);
DFFARX1 I_478 (I58472,I1803,I9750,I9974,);
DFFARX1 I_479 (I9974,I1803,I9750,I9739,);
nand I_480 (I9996,I58481,I58469);
and I_481 (I10013,I9996,I58463);
DFFARX1 I_482 (I10013,I1803,I9750,I10039,);
DFFARX1 I_483 (I10039,I1803,I9750,I10056,);
not I_484 (I9742,I10056);
not I_485 (I10078,I10039);
nand I_486 (I9727,I10078,I9917);
nor I_487 (I10109,I58457,I58469);
not I_488 (I10126,I10109);
nor I_489 (I10143,I10078,I10126);
nor I_490 (I10160,I9784,I10143);
DFFARX1 I_491 (I10160,I1803,I9750,I9736,);
nor I_492 (I10191,I9844,I10126);
nor I_493 (I9724,I10039,I10191);
nor I_494 (I9733,I9974,I10109);
nor I_495 (I9721,I9844,I10109);
not I_496 (I10277,I1810);
DFFARX1 I_497 (I66657,I1803,I10277,I10303,);
not I_498 (I10311,I10303);
nand I_499 (I10328,I66672,I66651);
and I_500 (I10345,I10328,I66654);
DFFARX1 I_501 (I10345,I1803,I10277,I10371,);
DFFARX1 I_502 (I66675,I1803,I10277,I10388,);
and I_503 (I10396,I10388,I66654);
nor I_504 (I10413,I10371,I10396);
DFFARX1 I_505 (I10413,I1803,I10277,I10245,);
nand I_506 (I10444,I10388,I66654);
nand I_507 (I10461,I10311,I10444);
not I_508 (I10257,I10461);
DFFARX1 I_509 (I66651,I1803,I10277,I10501,);
DFFARX1 I_510 (I10501,I1803,I10277,I10266,);
nand I_511 (I10523,I66663,I66660);
and I_512 (I10540,I10523,I66666);
DFFARX1 I_513 (I10540,I1803,I10277,I10566,);
DFFARX1 I_514 (I10566,I1803,I10277,I10583,);
not I_515 (I10269,I10583);
not I_516 (I10605,I10566);
nand I_517 (I10254,I10605,I10444);
nor I_518 (I10636,I66669,I66660);
not I_519 (I10653,I10636);
nor I_520 (I10670,I10605,I10653);
nor I_521 (I10687,I10311,I10670);
DFFARX1 I_522 (I10687,I1803,I10277,I10263,);
nor I_523 (I10718,I10371,I10653);
nor I_524 (I10251,I10566,I10718);
nor I_525 (I10260,I10501,I10636);
nor I_526 (I10248,I10371,I10636);
not I_527 (I10804,I1810);
DFFARX1 I_528 (I41656,I1803,I10804,I10830,);
not I_529 (I10838,I10830);
nand I_530 (I10855,I41647,I41665);
and I_531 (I10872,I10855,I41644);
DFFARX1 I_532 (I10872,I1803,I10804,I10898,);
DFFARX1 I_533 (I41647,I1803,I10804,I10915,);
and I_534 (I10923,I10915,I41650);
nor I_535 (I10940,I10898,I10923);
DFFARX1 I_536 (I10940,I1803,I10804,I10772,);
nand I_537 (I10971,I10915,I41650);
nand I_538 (I10988,I10838,I10971);
not I_539 (I10784,I10988);
DFFARX1 I_540 (I41644,I1803,I10804,I11028,);
DFFARX1 I_541 (I11028,I1803,I10804,I10793,);
nand I_542 (I11050,I41662,I41653);
and I_543 (I11067,I11050,I41668);
DFFARX1 I_544 (I11067,I1803,I10804,I11093,);
DFFARX1 I_545 (I11093,I1803,I10804,I11110,);
not I_546 (I10796,I11110);
not I_547 (I11132,I11093);
nand I_548 (I10781,I11132,I10971);
nor I_549 (I11163,I41659,I41653);
not I_550 (I11180,I11163);
nor I_551 (I11197,I11132,I11180);
nor I_552 (I11214,I10838,I11197);
DFFARX1 I_553 (I11214,I1803,I10804,I10790,);
nor I_554 (I11245,I10898,I11180);
nor I_555 (I10778,I11093,I11245);
nor I_556 (I10787,I11028,I11163);
nor I_557 (I10775,I10898,I11163);
not I_558 (I11331,I1810);
DFFARX1 I_559 (I70119,I1803,I11331,I11357,);
DFFARX1 I_560 (I11357,I1803,I11331,I11374,);
not I_561 (I11323,I11374);
not I_562 (I11396,I11357);
DFFARX1 I_563 (I70119,I1803,I11331,I11422,);
not I_564 (I11430,I11422);
and I_565 (I11447,I11396,I70122);
not I_566 (I11464,I70134);
nand I_567 (I11481,I11464,I70122);
not I_568 (I11498,I70140);
nor I_569 (I11515,I11498,I70131);
nand I_570 (I11532,I11515,I70137);
nor I_571 (I11549,I11532,I11481);
DFFARX1 I_572 (I11549,I1803,I11331,I11299,);
not I_573 (I11580,I11532);
not I_574 (I11597,I70131);
nand I_575 (I11614,I11597,I70122);
nor I_576 (I11631,I70131,I70134);
nand I_577 (I11311,I11447,I11631);
nand I_578 (I11305,I11396,I70131);
nand I_579 (I11676,I11498,I70128);
DFFARX1 I_580 (I11676,I1803,I11331,I11320,);
DFFARX1 I_581 (I11676,I1803,I11331,I11314,);
not I_582 (I11721,I70128);
nor I_583 (I11738,I11721,I70125);
and I_584 (I11755,I11738,I70143);
or I_585 (I11772,I11755,I70122);
DFFARX1 I_586 (I11772,I1803,I11331,I11798,);
nand I_587 (I11806,I11798,I11464);
nor I_588 (I11308,I11806,I11614);
nor I_589 (I11302,I11798,I11430);
DFFARX1 I_590 (I11798,I1803,I11331,I11860,);
not I_591 (I11868,I11860);
nor I_592 (I11317,I11868,I11580);
not I_593 (I11926,I1810);
DFFARX1 I_594 (I19680,I1803,I11926,I11952,);
DFFARX1 I_595 (I11952,I1803,I11926,I11969,);
not I_596 (I11918,I11969);
not I_597 (I11991,I11952);
DFFARX1 I_598 (I19695,I1803,I11926,I12017,);
not I_599 (I12025,I12017);
and I_600 (I12042,I11991,I19692);
not I_601 (I12059,I19680);
nand I_602 (I12076,I12059,I19692);
not I_603 (I12093,I19689);
nor I_604 (I12110,I12093,I19704);
nand I_605 (I12127,I12110,I19701);
nor I_606 (I12144,I12127,I12076);
DFFARX1 I_607 (I12144,I1803,I11926,I11894,);
not I_608 (I12175,I12127);
not I_609 (I12192,I19704);
nand I_610 (I12209,I12192,I19692);
nor I_611 (I12226,I19704,I19680);
nand I_612 (I11906,I12042,I12226);
nand I_613 (I11900,I11991,I19704);
nand I_614 (I12271,I12093,I19698);
DFFARX1 I_615 (I12271,I1803,I11926,I11915,);
DFFARX1 I_616 (I12271,I1803,I11926,I11909,);
not I_617 (I12316,I19698);
nor I_618 (I12333,I12316,I19686);
and I_619 (I12350,I12333,I19707);
or I_620 (I12367,I12350,I19683);
DFFARX1 I_621 (I12367,I1803,I11926,I12393,);
nand I_622 (I12401,I12393,I12059);
nor I_623 (I11903,I12401,I12209);
nor I_624 (I11897,I12393,I12025);
DFFARX1 I_625 (I12393,I1803,I11926,I12455,);
not I_626 (I12463,I12455);
nor I_627 (I11912,I12463,I12175);
not I_628 (I12521,I1810);
DFFARX1 I_629 (I55242,I1803,I12521,I12547,);
DFFARX1 I_630 (I12547,I1803,I12521,I12564,);
not I_631 (I12513,I12564);
not I_632 (I12586,I12547);
DFFARX1 I_633 (I55251,I1803,I12521,I12612,);
not I_634 (I12620,I12612);
and I_635 (I12637,I12586,I55239);
not I_636 (I12654,I55230);
nand I_637 (I12671,I12654,I55239);
not I_638 (I12688,I55236);
nor I_639 (I12705,I12688,I55254);
nand I_640 (I12722,I12705,I55227);
nor I_641 (I12739,I12722,I12671);
DFFARX1 I_642 (I12739,I1803,I12521,I12489,);
not I_643 (I12770,I12722);
not I_644 (I12787,I55254);
nand I_645 (I12804,I12787,I55239);
nor I_646 (I12821,I55254,I55230);
nand I_647 (I12501,I12637,I12821);
nand I_648 (I12495,I12586,I55254);
nand I_649 (I12866,I12688,I55233);
DFFARX1 I_650 (I12866,I1803,I12521,I12510,);
DFFARX1 I_651 (I12866,I1803,I12521,I12504,);
not I_652 (I12911,I55233);
nor I_653 (I12928,I12911,I55245);
and I_654 (I12945,I12928,I55227);
or I_655 (I12962,I12945,I55248);
DFFARX1 I_656 (I12962,I1803,I12521,I12988,);
nand I_657 (I12996,I12988,I12654);
nor I_658 (I12498,I12996,I12804);
nor I_659 (I12492,I12988,I12620);
DFFARX1 I_660 (I12988,I1803,I12521,I13050,);
not I_661 (I13058,I13050);
nor I_662 (I12507,I13058,I12770);
not I_663 (I13116,I1810);
DFFARX1 I_664 (I51595,I1803,I13116,I13142,);
DFFARX1 I_665 (I13142,I1803,I13116,I13159,);
not I_666 (I13108,I13159);
not I_667 (I13181,I13142);
DFFARX1 I_668 (I51589,I1803,I13116,I13207,);
not I_669 (I13215,I13207);
and I_670 (I13232,I13181,I51607);
not I_671 (I13249,I51595);
nand I_672 (I13266,I13249,I51607);
not I_673 (I13283,I51589);
nor I_674 (I13300,I13283,I51601);
nand I_675 (I13317,I13300,I51592);
nor I_676 (I13334,I13317,I13266);
DFFARX1 I_677 (I13334,I1803,I13116,I13084,);
not I_678 (I13365,I13317);
not I_679 (I13382,I51601);
nand I_680 (I13399,I13382,I51607);
nor I_681 (I13416,I51601,I51595);
nand I_682 (I13096,I13232,I13416);
nand I_683 (I13090,I13181,I51601);
nand I_684 (I13461,I13283,I51604);
DFFARX1 I_685 (I13461,I1803,I13116,I13105,);
DFFARX1 I_686 (I13461,I1803,I13116,I13099,);
not I_687 (I13506,I51604);
nor I_688 (I13523,I13506,I51610);
and I_689 (I13540,I13523,I51592);
or I_690 (I13557,I13540,I51598);
DFFARX1 I_691 (I13557,I1803,I13116,I13583,);
nand I_692 (I13591,I13583,I13249);
nor I_693 (I13093,I13591,I13399);
nor I_694 (I13087,I13583,I13215);
DFFARX1 I_695 (I13583,I1803,I13116,I13645,);
not I_696 (I13653,I13645);
nor I_697 (I13102,I13653,I13365);
not I_698 (I13711,I1810);
DFFARX1 I_699 (I32989,I1803,I13711,I13737,);
DFFARX1 I_700 (I13737,I1803,I13711,I13754,);
not I_701 (I13703,I13754);
not I_702 (I13776,I13737);
DFFARX1 I_703 (I32980,I1803,I13711,I13802,);
not I_704 (I13810,I13802);
and I_705 (I13827,I13776,I32998);
not I_706 (I13844,I32995);
nand I_707 (I13861,I13844,I32998);
not I_708 (I13878,I32974);
nor I_709 (I13895,I13878,I32977);
nand I_710 (I13912,I13895,I32986);
nor I_711 (I13929,I13912,I13861);
DFFARX1 I_712 (I13929,I1803,I13711,I13679,);
not I_713 (I13960,I13912);
not I_714 (I13977,I32977);
nand I_715 (I13994,I13977,I32998);
nor I_716 (I14011,I32977,I32995);
nand I_717 (I13691,I13827,I14011);
nand I_718 (I13685,I13776,I32977);
nand I_719 (I14056,I13878,I32992);
DFFARX1 I_720 (I14056,I1803,I13711,I13700,);
DFFARX1 I_721 (I14056,I1803,I13711,I13694,);
not I_722 (I14101,I32992);
nor I_723 (I14118,I14101,I32974);
and I_724 (I14135,I14118,I32983);
or I_725 (I14152,I14135,I32977);
DFFARX1 I_726 (I14152,I1803,I13711,I14178,);
nand I_727 (I14186,I14178,I13844);
nor I_728 (I13688,I14186,I13994);
nor I_729 (I13682,I14178,I13810);
DFFARX1 I_730 (I14178,I1803,I13711,I14240,);
not I_731 (I14248,I14240);
nor I_732 (I13697,I14248,I13960);
not I_733 (I14306,I1810);
DFFARX1 I_734 (I70697,I1803,I14306,I14332,);
DFFARX1 I_735 (I14332,I1803,I14306,I14349,);
not I_736 (I14298,I14349);
not I_737 (I14371,I14332);
DFFARX1 I_738 (I70697,I1803,I14306,I14397,);
not I_739 (I14405,I14397);
and I_740 (I14422,I14371,I70700);
not I_741 (I14439,I70712);
nand I_742 (I14456,I14439,I70700);
not I_743 (I14473,I70718);
nor I_744 (I14490,I14473,I70709);
nand I_745 (I14507,I14490,I70715);
nor I_746 (I14524,I14507,I14456);
DFFARX1 I_747 (I14524,I1803,I14306,I14274,);
not I_748 (I14555,I14507);
not I_749 (I14572,I70709);
nand I_750 (I14589,I14572,I70700);
nor I_751 (I14606,I70709,I70712);
nand I_752 (I14286,I14422,I14606);
nand I_753 (I14280,I14371,I70709);
nand I_754 (I14651,I14473,I70706);
DFFARX1 I_755 (I14651,I1803,I14306,I14295,);
DFFARX1 I_756 (I14651,I1803,I14306,I14289,);
not I_757 (I14696,I70706);
nor I_758 (I14713,I14696,I70703);
and I_759 (I14730,I14713,I70721);
or I_760 (I14747,I14730,I70700);
DFFARX1 I_761 (I14747,I1803,I14306,I14773,);
nand I_762 (I14781,I14773,I14439);
nor I_763 (I14283,I14781,I14589);
nor I_764 (I14277,I14773,I14405);
DFFARX1 I_765 (I14773,I1803,I14306,I14835,);
not I_766 (I14843,I14835);
nor I_767 (I14292,I14843,I14555);
not I_768 (I14901,I1810);
DFFARX1 I_769 (I28821,I1803,I14901,I14927,);
DFFARX1 I_770 (I14927,I1803,I14901,I14944,);
not I_771 (I14893,I14944);
not I_772 (I14966,I14927);
DFFARX1 I_773 (I28815,I1803,I14901,I14992,);
not I_774 (I15000,I14992);
and I_775 (I15017,I14966,I28830);
not I_776 (I15034,I28827);
nand I_777 (I15051,I15034,I28830);
not I_778 (I15068,I28818);
nor I_779 (I15085,I15068,I28809);
nand I_780 (I15102,I15085,I28812);
nor I_781 (I15119,I15102,I15051);
DFFARX1 I_782 (I15119,I1803,I14901,I14869,);
not I_783 (I15150,I15102);
not I_784 (I15167,I28809);
nand I_785 (I15184,I15167,I28830);
nor I_786 (I15201,I28809,I28827);
nand I_787 (I14881,I15017,I15201);
nand I_788 (I14875,I14966,I28809);
nand I_789 (I15246,I15068,I28833);
DFFARX1 I_790 (I15246,I1803,I14901,I14890,);
DFFARX1 I_791 (I15246,I1803,I14901,I14884,);
not I_792 (I15291,I28833);
nor I_793 (I15308,I15291,I28824);
and I_794 (I15325,I15308,I28809);
or I_795 (I15342,I15325,I28812);
DFFARX1 I_796 (I15342,I1803,I14901,I15368,);
nand I_797 (I15376,I15368,I15034);
nor I_798 (I14878,I15376,I15184);
nor I_799 (I14872,I15368,I15000);
DFFARX1 I_800 (I15368,I1803,I14901,I15430,);
not I_801 (I15438,I15430);
nor I_802 (I14887,I15438,I15150);
not I_803 (I15499,I1810);
DFFARX1 I_804 (I4978,I1803,I15499,I15525,);
nand I_805 (I15533,I4990,I4999);
and I_806 (I15550,I15533,I4978);
DFFARX1 I_807 (I15550,I1803,I15499,I15576,);
nor I_808 (I15467,I15576,I15525);
not I_809 (I15598,I15576);
DFFARX1 I_810 (I4993,I1803,I15499,I15624,);
nand I_811 (I15632,I15624,I4981);
not I_812 (I15649,I15632);
DFFARX1 I_813 (I15649,I1803,I15499,I15675,);
not I_814 (I15491,I15675);
nor I_815 (I15697,I15525,I15632);
nor I_816 (I15473,I15576,I15697);
DFFARX1 I_817 (I4984,I1803,I15499,I15737,);
DFFARX1 I_818 (I15737,I1803,I15499,I15754,);
not I_819 (I15762,I15754);
not I_820 (I15779,I15737);
nand I_821 (I15476,I15779,I15598);
nand I_822 (I15810,I4975,I4975);
and I_823 (I15827,I15810,I4987);
DFFARX1 I_824 (I15827,I1803,I15499,I15853,);
nor I_825 (I15861,I15853,I15525);
DFFARX1 I_826 (I15861,I1803,I15499,I15464,);
DFFARX1 I_827 (I15853,I1803,I15499,I15482,);
nor I_828 (I15906,I4996,I4975);
not I_829 (I15923,I15906);
nor I_830 (I15485,I15762,I15923);
nand I_831 (I15470,I15779,I15923);
nor I_832 (I15479,I15525,I15906);
DFFARX1 I_833 (I15906,I1803,I15499,I15488,);
not I_834 (I16026,I1810);
DFFARX1 I_835 (I14274,I1803,I16026,I16052,);
nand I_836 (I16060,I14274,I14280);
and I_837 (I16077,I16060,I14298);
DFFARX1 I_838 (I16077,I1803,I16026,I16103,);
nor I_839 (I15994,I16103,I16052);
not I_840 (I16125,I16103);
DFFARX1 I_841 (I14286,I1803,I16026,I16151,);
nand I_842 (I16159,I16151,I14283);
not I_843 (I16176,I16159);
DFFARX1 I_844 (I16176,I1803,I16026,I16202,);
not I_845 (I16018,I16202);
nor I_846 (I16224,I16052,I16159);
nor I_847 (I16000,I16103,I16224);
DFFARX1 I_848 (I14292,I1803,I16026,I16264,);
DFFARX1 I_849 (I16264,I1803,I16026,I16281,);
not I_850 (I16289,I16281);
not I_851 (I16306,I16264);
nand I_852 (I16003,I16306,I16125);
nand I_853 (I16337,I14277,I14277);
and I_854 (I16354,I16337,I14289);
DFFARX1 I_855 (I16354,I1803,I16026,I16380,);
nor I_856 (I16388,I16380,I16052);
DFFARX1 I_857 (I16388,I1803,I16026,I15991,);
DFFARX1 I_858 (I16380,I1803,I16026,I16009,);
nor I_859 (I16433,I14295,I14277);
not I_860 (I16450,I16433);
nor I_861 (I16012,I16289,I16450);
nand I_862 (I15997,I16306,I16450);
nor I_863 (I16006,I16052,I16433);
DFFARX1 I_864 (I16433,I1803,I16026,I16015,);
not I_865 (I16553,I1810);
DFFARX1 I_866 (I8667,I1803,I16553,I16579,);
nand I_867 (I16587,I8679,I8688);
and I_868 (I16604,I16587,I8667);
DFFARX1 I_869 (I16604,I1803,I16553,I16630,);
nor I_870 (I16521,I16630,I16579);
not I_871 (I16652,I16630);
DFFARX1 I_872 (I8682,I1803,I16553,I16678,);
nand I_873 (I16686,I16678,I8670);
not I_874 (I16703,I16686);
DFFARX1 I_875 (I16703,I1803,I16553,I16729,);
not I_876 (I16545,I16729);
nor I_877 (I16751,I16579,I16686);
nor I_878 (I16527,I16630,I16751);
DFFARX1 I_879 (I8673,I1803,I16553,I16791,);
DFFARX1 I_880 (I16791,I1803,I16553,I16808,);
not I_881 (I16816,I16808);
not I_882 (I16833,I16791);
nand I_883 (I16530,I16833,I16652);
nand I_884 (I16864,I8664,I8664);
and I_885 (I16881,I16864,I8676);
DFFARX1 I_886 (I16881,I1803,I16553,I16907,);
nor I_887 (I16915,I16907,I16579);
DFFARX1 I_888 (I16915,I1803,I16553,I16518,);
DFFARX1 I_889 (I16907,I1803,I16553,I16536,);
nor I_890 (I16960,I8685,I8664);
not I_891 (I16977,I16960);
nor I_892 (I16539,I16816,I16977);
nand I_893 (I16524,I16833,I16977);
nor I_894 (I16533,I16579,I16960);
DFFARX1 I_895 (I16960,I1803,I16553,I16542,);
not I_896 (I17080,I1810);
DFFARX1 I_897 (I30002,I1803,I17080,I17106,);
nand I_898 (I17114,I30002,I30014);
and I_899 (I17131,I17114,I29999);
DFFARX1 I_900 (I17131,I1803,I17080,I17157,);
nor I_901 (I17048,I17157,I17106);
not I_902 (I17179,I17157);
DFFARX1 I_903 (I30023,I1803,I17080,I17205,);
nand I_904 (I17213,I17205,I30020);
not I_905 (I17230,I17213);
DFFARX1 I_906 (I17230,I1803,I17080,I17256,);
not I_907 (I17072,I17256);
nor I_908 (I17278,I17106,I17213);
nor I_909 (I17054,I17157,I17278);
DFFARX1 I_910 (I30011,I1803,I17080,I17318,);
DFFARX1 I_911 (I17318,I1803,I17080,I17335,);
not I_912 (I17343,I17335);
not I_913 (I17360,I17318);
nand I_914 (I17057,I17360,I17179);
nand I_915 (I17391,I29999,I30008);
and I_916 (I17408,I17391,I30017);
DFFARX1 I_917 (I17408,I1803,I17080,I17434,);
nor I_918 (I17442,I17434,I17106);
DFFARX1 I_919 (I17442,I1803,I17080,I17045,);
DFFARX1 I_920 (I17434,I1803,I17080,I17063,);
nor I_921 (I17487,I30005,I30008);
not I_922 (I17504,I17487);
nor I_923 (I17066,I17343,I17504);
nand I_924 (I17051,I17360,I17504);
nor I_925 (I17060,I17106,I17487);
DFFARX1 I_926 (I17487,I1803,I17080,I17069,);
not I_927 (I17607,I1810);
DFFARX1 I_928 (I34145,I1803,I17607,I17633,);
nand I_929 (I17641,I34130,I34133);
and I_930 (I17658,I17641,I34148);
DFFARX1 I_931 (I17658,I1803,I17607,I17684,);
nor I_932 (I17575,I17684,I17633);
not I_933 (I17706,I17684);
DFFARX1 I_934 (I34142,I1803,I17607,I17732,);
nand I_935 (I17740,I17732,I34133);
not I_936 (I17757,I17740);
DFFARX1 I_937 (I17757,I1803,I17607,I17783,);
not I_938 (I17599,I17783);
nor I_939 (I17805,I17633,I17740);
nor I_940 (I17581,I17684,I17805);
DFFARX1 I_941 (I34139,I1803,I17607,I17845,);
DFFARX1 I_942 (I17845,I1803,I17607,I17862,);
not I_943 (I17870,I17862);
not I_944 (I17887,I17845);
nand I_945 (I17584,I17887,I17706);
nand I_946 (I17918,I34154,I34130);
and I_947 (I17935,I17918,I34151);
DFFARX1 I_948 (I17935,I1803,I17607,I17961,);
nor I_949 (I17969,I17961,I17633);
DFFARX1 I_950 (I17969,I1803,I17607,I17572,);
DFFARX1 I_951 (I17961,I1803,I17607,I17590,);
nor I_952 (I18014,I34136,I34130);
not I_953 (I18031,I18014);
nor I_954 (I17593,I17870,I18031);
nand I_955 (I17578,I17887,I18031);
nor I_956 (I17587,I17633,I18014);
DFFARX1 I_957 (I18014,I1803,I17607,I17596,);
not I_958 (I18134,I1810);
DFFARX1 I_959 (I81037,I1803,I18134,I18160,);
nand I_960 (I18168,I81016,I81016);
and I_961 (I18185,I18168,I81043);
DFFARX1 I_962 (I18185,I1803,I18134,I18211,);
nor I_963 (I18102,I18211,I18160);
not I_964 (I18233,I18211);
DFFARX1 I_965 (I81031,I1803,I18134,I18259,);
nand I_966 (I18267,I18259,I81034);
not I_967 (I18284,I18267);
DFFARX1 I_968 (I18284,I1803,I18134,I18310,);
not I_969 (I18126,I18310);
nor I_970 (I18332,I18160,I18267);
nor I_971 (I18108,I18211,I18332);
DFFARX1 I_972 (I81025,I1803,I18134,I18372,);
DFFARX1 I_973 (I18372,I1803,I18134,I18389,);
not I_974 (I18397,I18389);
not I_975 (I18414,I18372);
nand I_976 (I18111,I18414,I18233);
nand I_977 (I18445,I81022,I81019);
and I_978 (I18462,I18445,I81040);
DFFARX1 I_979 (I18462,I1803,I18134,I18488,);
nor I_980 (I18496,I18488,I18160);
DFFARX1 I_981 (I18496,I1803,I18134,I18099,);
DFFARX1 I_982 (I18488,I1803,I18134,I18117,);
nor I_983 (I18541,I81028,I81019);
not I_984 (I18558,I18541);
nor I_985 (I18120,I18397,I18558);
nand I_986 (I18105,I18414,I18558);
nor I_987 (I18114,I18160,I18541);
DFFARX1 I_988 (I18541,I1803,I18134,I18123,);
not I_989 (I18661,I1810);
DFFARX1 I_990 (I68963,I1803,I18661,I18687,);
nand I_991 (I18695,I68978,I68963);
and I_992 (I18712,I18695,I68981);
DFFARX1 I_993 (I18712,I1803,I18661,I18738,);
nor I_994 (I18629,I18738,I18687);
not I_995 (I18760,I18738);
DFFARX1 I_996 (I68987,I1803,I18661,I18786,);
nand I_997 (I18794,I18786,I68969);
not I_998 (I18811,I18794);
DFFARX1 I_999 (I18811,I1803,I18661,I18837,);
not I_1000 (I18653,I18837);
nor I_1001 (I18859,I18687,I18794);
nor I_1002 (I18635,I18738,I18859);
DFFARX1 I_1003 (I68966,I1803,I18661,I18899,);
DFFARX1 I_1004 (I18899,I1803,I18661,I18916,);
not I_1005 (I18924,I18916);
not I_1006 (I18941,I18899);
nand I_1007 (I18638,I18941,I18760);
nand I_1008 (I18972,I68966,I68972);
and I_1009 (I18989,I18972,I68984);
DFFARX1 I_1010 (I18989,I1803,I18661,I19015,);
nor I_1011 (I19023,I19015,I18687);
DFFARX1 I_1012 (I19023,I1803,I18661,I18626,);
DFFARX1 I_1013 (I19015,I1803,I18661,I18644,);
nor I_1014 (I19068,I68975,I68972);
not I_1015 (I19085,I19068);
nor I_1016 (I18647,I18924,I19085);
nand I_1017 (I18632,I18941,I19085);
nor I_1018 (I18641,I18687,I19068);
DFFARX1 I_1019 (I19068,I1803,I18661,I18650,);
not I_1020 (I19188,I1810);
DFFARX1 I_1021 (I13679,I1803,I19188,I19214,);
nand I_1022 (I19222,I13679,I13685);
and I_1023 (I19239,I19222,I13703);
DFFARX1 I_1024 (I19239,I1803,I19188,I19265,);
nor I_1025 (I19156,I19265,I19214);
not I_1026 (I19287,I19265);
DFFARX1 I_1027 (I13691,I1803,I19188,I19313,);
nand I_1028 (I19321,I19313,I13688);
not I_1029 (I19338,I19321);
DFFARX1 I_1030 (I19338,I1803,I19188,I19364,);
not I_1031 (I19180,I19364);
nor I_1032 (I19386,I19214,I19321);
nor I_1033 (I19162,I19265,I19386);
DFFARX1 I_1034 (I13697,I1803,I19188,I19426,);
DFFARX1 I_1035 (I19426,I1803,I19188,I19443,);
not I_1036 (I19451,I19443);
not I_1037 (I19468,I19426);
nand I_1038 (I19165,I19468,I19287);
nand I_1039 (I19499,I13682,I13682);
and I_1040 (I19516,I19499,I13694);
DFFARX1 I_1041 (I19516,I1803,I19188,I19542,);
nor I_1042 (I19550,I19542,I19214);
DFFARX1 I_1043 (I19550,I1803,I19188,I19153,);
DFFARX1 I_1044 (I19542,I1803,I19188,I19171,);
nor I_1045 (I19595,I13700,I13682);
not I_1046 (I19612,I19595);
nor I_1047 (I19174,I19451,I19612);
nand I_1048 (I19159,I19468,I19612);
nor I_1049 (I19168,I19214,I19595);
DFFARX1 I_1050 (I19595,I1803,I19188,I19177,);
not I_1051 (I19715,I1810);
DFFARX1 I_1052 (I59106,I1803,I19715,I19741,);
nand I_1053 (I19749,I59103,I59121);
and I_1054 (I19766,I19749,I59112);
DFFARX1 I_1055 (I19766,I1803,I19715,I19792,);
nor I_1056 (I19683,I19792,I19741);
not I_1057 (I19814,I19792);
DFFARX1 I_1058 (I59127,I1803,I19715,I19840,);
nand I_1059 (I19848,I19840,I59109);
not I_1060 (I19865,I19848);
DFFARX1 I_1061 (I19865,I1803,I19715,I19891,);
not I_1062 (I19707,I19891);
nor I_1063 (I19913,I19741,I19848);
nor I_1064 (I19689,I19792,I19913);
DFFARX1 I_1065 (I59115,I1803,I19715,I19953,);
DFFARX1 I_1066 (I19953,I1803,I19715,I19970,);
not I_1067 (I19978,I19970);
not I_1068 (I19995,I19953);
nand I_1069 (I19692,I19995,I19814);
nand I_1070 (I20026,I59103,I59130);
and I_1071 (I20043,I20026,I59118);
DFFARX1 I_1072 (I20043,I1803,I19715,I20069,);
nor I_1073 (I20077,I20069,I19741);
DFFARX1 I_1074 (I20077,I1803,I19715,I19680,);
DFFARX1 I_1075 (I20069,I1803,I19715,I19698,);
nor I_1076 (I20122,I59124,I59130);
not I_1077 (I20139,I20122);
nor I_1078 (I19701,I19978,I20139);
nand I_1079 (I19686,I19995,I20139);
nor I_1080 (I19695,I19741,I20122);
DFFARX1 I_1081 (I20122,I1803,I19715,I19704,);
not I_1082 (I20242,I1810);
DFFARX1 I_1083 (I30597,I1803,I20242,I20268,);
nand I_1084 (I20276,I30597,I30609);
and I_1085 (I20293,I20276,I30594);
DFFARX1 I_1086 (I20293,I1803,I20242,I20319,);
nor I_1087 (I20210,I20319,I20268);
not I_1088 (I20341,I20319);
DFFARX1 I_1089 (I30618,I1803,I20242,I20367,);
nand I_1090 (I20375,I20367,I30615);
not I_1091 (I20392,I20375);
DFFARX1 I_1092 (I20392,I1803,I20242,I20418,);
not I_1093 (I20234,I20418);
nor I_1094 (I20440,I20268,I20375);
nor I_1095 (I20216,I20319,I20440);
DFFARX1 I_1096 (I30606,I1803,I20242,I20480,);
DFFARX1 I_1097 (I20480,I1803,I20242,I20497,);
not I_1098 (I20505,I20497);
not I_1099 (I20522,I20480);
nand I_1100 (I20219,I20522,I20341);
nand I_1101 (I20553,I30594,I30603);
and I_1102 (I20570,I20553,I30612);
DFFARX1 I_1103 (I20570,I1803,I20242,I20596,);
nor I_1104 (I20604,I20596,I20268);
DFFARX1 I_1105 (I20604,I1803,I20242,I20207,);
DFFARX1 I_1106 (I20596,I1803,I20242,I20225,);
nor I_1107 (I20649,I30600,I30603);
not I_1108 (I20666,I20649);
nor I_1109 (I20228,I20505,I20666);
nand I_1110 (I20213,I20522,I20666);
nor I_1111 (I20222,I20268,I20649);
DFFARX1 I_1112 (I20649,I1803,I20242,I20231,);
not I_1113 (I20769,I1810);
DFFARX1 I_1114 (I75778,I1803,I20769,I20795,);
nand I_1115 (I20803,I75775,I75766);
and I_1116 (I20820,I20803,I75763);
DFFARX1 I_1117 (I20820,I1803,I20769,I20846,);
nor I_1118 (I20737,I20846,I20795);
not I_1119 (I20868,I20846);
DFFARX1 I_1120 (I75772,I1803,I20769,I20894,);
nand I_1121 (I20902,I20894,I75781);
not I_1122 (I20919,I20902);
DFFARX1 I_1123 (I20919,I1803,I20769,I20945,);
not I_1124 (I20761,I20945);
nor I_1125 (I20967,I20795,I20902);
nor I_1126 (I20743,I20846,I20967);
DFFARX1 I_1127 (I75784,I1803,I20769,I21007,);
DFFARX1 I_1128 (I21007,I1803,I20769,I21024,);
not I_1129 (I21032,I21024);
not I_1130 (I21049,I21007);
nand I_1131 (I20746,I21049,I20868);
nand I_1132 (I21080,I75763,I75769);
and I_1133 (I21097,I21080,I75787);
DFFARX1 I_1134 (I21097,I1803,I20769,I21123,);
nor I_1135 (I21131,I21123,I20795);
DFFARX1 I_1136 (I21131,I1803,I20769,I20734,);
DFFARX1 I_1137 (I21123,I1803,I20769,I20752,);
nor I_1138 (I21176,I75766,I75769);
not I_1139 (I21193,I21176);
nor I_1140 (I20755,I21032,I21193);
nand I_1141 (I20740,I21049,I21193);
nor I_1142 (I20749,I20795,I21176);
DFFARX1 I_1143 (I21176,I1803,I20769,I20758,);
not I_1144 (I21296,I1810);
DFFARX1 I_1145 (I62081,I1803,I21296,I21322,);
nand I_1146 (I21330,I62078,I62081);
and I_1147 (I21347,I21330,I62090);
DFFARX1 I_1148 (I21347,I1803,I21296,I21373,);
nor I_1149 (I21264,I21373,I21322);
not I_1150 (I21395,I21373);
DFFARX1 I_1151 (I62078,I1803,I21296,I21421,);
nand I_1152 (I21429,I21421,I62096);
not I_1153 (I21446,I21429);
DFFARX1 I_1154 (I21446,I1803,I21296,I21472,);
not I_1155 (I21288,I21472);
nor I_1156 (I21494,I21322,I21429);
nor I_1157 (I21270,I21373,I21494);
DFFARX1 I_1158 (I62084,I1803,I21296,I21534,);
DFFARX1 I_1159 (I21534,I1803,I21296,I21551,);
not I_1160 (I21559,I21551);
not I_1161 (I21576,I21534);
nand I_1162 (I21273,I21576,I21395);
nand I_1163 (I21607,I62093,I62099);
and I_1164 (I21624,I21607,I62084);
DFFARX1 I_1165 (I21624,I1803,I21296,I21650,);
nor I_1166 (I21658,I21650,I21322);
DFFARX1 I_1167 (I21658,I1803,I21296,I21261,);
DFFARX1 I_1168 (I21650,I1803,I21296,I21279,);
nor I_1169 (I21703,I62087,I62099);
not I_1170 (I21720,I21703);
nor I_1171 (I21282,I21559,I21720);
nand I_1172 (I21267,I21576,I21720);
nor I_1173 (I21276,I21322,I21703);
DFFARX1 I_1174 (I21703,I1803,I21296,I21285,);
not I_1175 (I21823,I1810);
DFFARX1 I_1176 (I55876,I1803,I21823,I21849,);
nand I_1177 (I21857,I55873,I55891);
and I_1178 (I21874,I21857,I55882);
DFFARX1 I_1179 (I21874,I1803,I21823,I21900,);
nor I_1180 (I21791,I21900,I21849);
not I_1181 (I21922,I21900);
DFFARX1 I_1182 (I55897,I1803,I21823,I21948,);
nand I_1183 (I21956,I21948,I55879);
not I_1184 (I21973,I21956);
DFFARX1 I_1185 (I21973,I1803,I21823,I21999,);
not I_1186 (I21815,I21999);
nor I_1187 (I22021,I21849,I21956);
nor I_1188 (I21797,I21900,I22021);
DFFARX1 I_1189 (I55885,I1803,I21823,I22061,);
DFFARX1 I_1190 (I22061,I1803,I21823,I22078,);
not I_1191 (I22086,I22078);
not I_1192 (I22103,I22061);
nand I_1193 (I21800,I22103,I21922);
nand I_1194 (I22134,I55873,I55900);
and I_1195 (I22151,I22134,I55888);
DFFARX1 I_1196 (I22151,I1803,I21823,I22177,);
nor I_1197 (I22185,I22177,I21849);
DFFARX1 I_1198 (I22185,I1803,I21823,I21788,);
DFFARX1 I_1199 (I22177,I1803,I21823,I21806,);
nor I_1200 (I22230,I55894,I55900);
not I_1201 (I22247,I22230);
nor I_1202 (I21809,I22086,I22247);
nand I_1203 (I21794,I22103,I22247);
nor I_1204 (I21803,I21849,I22230);
DFFARX1 I_1205 (I22230,I1803,I21823,I21812,);
not I_1206 (I22350,I1810);
DFFARX1 I_1207 (I82822,I1803,I22350,I22376,);
nand I_1208 (I22384,I82801,I82801);
and I_1209 (I22401,I22384,I82828);
DFFARX1 I_1210 (I22401,I1803,I22350,I22427,);
nor I_1211 (I22318,I22427,I22376);
not I_1212 (I22449,I22427);
DFFARX1 I_1213 (I82816,I1803,I22350,I22475,);
nand I_1214 (I22483,I22475,I82819);
not I_1215 (I22500,I22483);
DFFARX1 I_1216 (I22500,I1803,I22350,I22526,);
not I_1217 (I22342,I22526);
nor I_1218 (I22548,I22376,I22483);
nor I_1219 (I22324,I22427,I22548);
DFFARX1 I_1220 (I82810,I1803,I22350,I22588,);
DFFARX1 I_1221 (I22588,I1803,I22350,I22605,);
not I_1222 (I22613,I22605);
not I_1223 (I22630,I22588);
nand I_1224 (I22327,I22630,I22449);
nand I_1225 (I22661,I82807,I82804);
and I_1226 (I22678,I22661,I82825);
DFFARX1 I_1227 (I22678,I1803,I22350,I22704,);
nor I_1228 (I22712,I22704,I22376);
DFFARX1 I_1229 (I22712,I1803,I22350,I22315,);
DFFARX1 I_1230 (I22704,I1803,I22350,I22333,);
nor I_1231 (I22757,I82813,I82804);
not I_1232 (I22774,I22757);
nor I_1233 (I22336,I22613,I22774);
nand I_1234 (I22321,I22630,I22774);
nor I_1235 (I22330,I22376,I22757);
DFFARX1 I_1236 (I22757,I1803,I22350,I22339,);
not I_1237 (I22877,I1810);
DFFARX1 I_1238 (I1596,I1803,I22877,I22903,);
nand I_1239 (I22911,I1540,I1748);
and I_1240 (I22928,I22911,I1508);
DFFARX1 I_1241 (I22928,I1803,I22877,I22954,);
nor I_1242 (I22845,I22954,I22903);
not I_1243 (I22976,I22954);
DFFARX1 I_1244 (I1700,I1803,I22877,I23002,);
nand I_1245 (I23010,I23002,I1460);
not I_1246 (I23027,I23010);
DFFARX1 I_1247 (I23027,I1803,I22877,I23053,);
not I_1248 (I22869,I23053);
nor I_1249 (I23075,I22903,I23010);
nor I_1250 (I22851,I22954,I23075);
DFFARX1 I_1251 (I1468,I1803,I22877,I23115,);
DFFARX1 I_1252 (I23115,I1803,I22877,I23132,);
not I_1253 (I23140,I23132);
not I_1254 (I23157,I23115);
nand I_1255 (I22854,I23157,I22976);
nand I_1256 (I23188,I1364,I1796);
and I_1257 (I23205,I23188,I1548);
DFFARX1 I_1258 (I23205,I1803,I22877,I23231,);
nor I_1259 (I23239,I23231,I22903);
DFFARX1 I_1260 (I23239,I1803,I22877,I22842,);
DFFARX1 I_1261 (I23231,I1803,I22877,I22860,);
nor I_1262 (I23284,I1412,I1796);
not I_1263 (I23301,I23284);
nor I_1264 (I22863,I23140,I23301);
nand I_1265 (I22848,I23157,I23301);
nor I_1266 (I22857,I22903,I23284);
DFFARX1 I_1267 (I23284,I1803,I22877,I22866,);
not I_1268 (I23404,I1810);
DFFARX1 I_1269 (I68388,I1803,I23404,I23430,);
DFFARX1 I_1270 (I23430,I1803,I23404,I23447,);
not I_1271 (I23396,I23447);
not I_1272 (I23469,I23430);
nand I_1273 (I23486,I68400,I68388);
and I_1274 (I23503,I23486,I68391);
DFFARX1 I_1275 (I23503,I1803,I23404,I23529,);
not I_1276 (I23537,I23529);
DFFARX1 I_1277 (I68409,I1803,I23404,I23563,);
and I_1278 (I23571,I23563,I68385);
nand I_1279 (I23588,I23563,I68385);
nand I_1280 (I23375,I23537,I23588);
DFFARX1 I_1281 (I68403,I1803,I23404,I23628,);
nor I_1282 (I23636,I23628,I23571);
DFFARX1 I_1283 (I23636,I1803,I23404,I23369,);
nor I_1284 (I23384,I23628,I23529);
nand I_1285 (I23681,I68397,I68394);
and I_1286 (I23698,I23681,I68406);
DFFARX1 I_1287 (I23698,I1803,I23404,I23724,);
nor I_1288 (I23372,I23724,I23628);
not I_1289 (I23746,I23724);
nor I_1290 (I23763,I23746,I23537);
nor I_1291 (I23780,I23469,I23763);
DFFARX1 I_1292 (I23780,I1803,I23404,I23387,);
nor I_1293 (I23811,I23746,I23628);
nor I_1294 (I23828,I68385,I68394);
nor I_1295 (I23378,I23828,I23811);
not I_1296 (I23859,I23828);
nand I_1297 (I23381,I23588,I23859);
DFFARX1 I_1298 (I23828,I1803,I23404,I23393,);
DFFARX1 I_1299 (I23828,I1803,I23404,I23390,);
not I_1300 (I23948,I1810);
DFFARX1 I_1301 (I69544,I1803,I23948,I23974,);
DFFARX1 I_1302 (I23974,I1803,I23948,I23991,);
not I_1303 (I23940,I23991);
not I_1304 (I24013,I23974);
nand I_1305 (I24030,I69556,I69544);
and I_1306 (I24047,I24030,I69547);
DFFARX1 I_1307 (I24047,I1803,I23948,I24073,);
not I_1308 (I24081,I24073);
DFFARX1 I_1309 (I69565,I1803,I23948,I24107,);
and I_1310 (I24115,I24107,I69541);
nand I_1311 (I24132,I24107,I69541);
nand I_1312 (I23919,I24081,I24132);
DFFARX1 I_1313 (I69559,I1803,I23948,I24172,);
nor I_1314 (I24180,I24172,I24115);
DFFARX1 I_1315 (I24180,I1803,I23948,I23913,);
nor I_1316 (I23928,I24172,I24073);
nand I_1317 (I24225,I69553,I69550);
and I_1318 (I24242,I24225,I69562);
DFFARX1 I_1319 (I24242,I1803,I23948,I24268,);
nor I_1320 (I23916,I24268,I24172);
not I_1321 (I24290,I24268);
nor I_1322 (I24307,I24290,I24081);
nor I_1323 (I24324,I24013,I24307);
DFFARX1 I_1324 (I24324,I1803,I23948,I23931,);
nor I_1325 (I24355,I24290,I24172);
nor I_1326 (I24372,I69541,I69550);
nor I_1327 (I23922,I24372,I24355);
not I_1328 (I24403,I24372);
nand I_1329 (I23925,I24132,I24403);
DFFARX1 I_1330 (I24372,I1803,I23948,I23937,);
DFFARX1 I_1331 (I24372,I1803,I23948,I23934,);
not I_1332 (I24492,I1810);
DFFARX1 I_1333 (I52649,I1803,I24492,I24518,);
DFFARX1 I_1334 (I24518,I1803,I24492,I24535,);
not I_1335 (I24484,I24535);
not I_1336 (I24557,I24518);
nand I_1337 (I24574,I52664,I52652);
and I_1338 (I24591,I24574,I52643);
DFFARX1 I_1339 (I24591,I1803,I24492,I24617,);
not I_1340 (I24625,I24617);
DFFARX1 I_1341 (I52655,I1803,I24492,I24651,);
and I_1342 (I24659,I24651,I52646);
nand I_1343 (I24676,I24651,I52646);
nand I_1344 (I24463,I24625,I24676);
DFFARX1 I_1345 (I52661,I1803,I24492,I24716,);
nor I_1346 (I24724,I24716,I24659);
DFFARX1 I_1347 (I24724,I1803,I24492,I24457,);
nor I_1348 (I24472,I24716,I24617);
nand I_1349 (I24769,I52670,I52658);
and I_1350 (I24786,I24769,I52667);
DFFARX1 I_1351 (I24786,I1803,I24492,I24812,);
nor I_1352 (I24460,I24812,I24716);
not I_1353 (I24834,I24812);
nor I_1354 (I24851,I24834,I24625);
nor I_1355 (I24868,I24557,I24851);
DFFARX1 I_1356 (I24868,I1803,I24492,I24475,);
nor I_1357 (I24899,I24834,I24716);
nor I_1358 (I24916,I52643,I52658);
nor I_1359 (I24466,I24916,I24899);
not I_1360 (I24947,I24916);
nand I_1361 (I24469,I24676,I24947);
DFFARX1 I_1362 (I24916,I1803,I24492,I24481,);
DFFARX1 I_1363 (I24916,I1803,I24492,I24478,);
not I_1364 (I25036,I1810);
DFFARX1 I_1365 (I48966,I1803,I25036,I25062,);
DFFARX1 I_1366 (I25062,I1803,I25036,I25079,);
not I_1367 (I25028,I25079);
not I_1368 (I25101,I25062);
nand I_1369 (I25118,I48960,I48957);
and I_1370 (I25135,I25118,I48972);
DFFARX1 I_1371 (I25135,I1803,I25036,I25161,);
not I_1372 (I25169,I25161);
DFFARX1 I_1373 (I48960,I1803,I25036,I25195,);
and I_1374 (I25203,I25195,I48954);
nand I_1375 (I25220,I25195,I48954);
nand I_1376 (I25007,I25169,I25220);
DFFARX1 I_1377 (I48954,I1803,I25036,I25260,);
nor I_1378 (I25268,I25260,I25203);
DFFARX1 I_1379 (I25268,I1803,I25036,I25001,);
nor I_1380 (I25016,I25260,I25161);
nand I_1381 (I25313,I48969,I48963);
and I_1382 (I25330,I25313,I48957);
DFFARX1 I_1383 (I25330,I1803,I25036,I25356,);
nor I_1384 (I25004,I25356,I25260);
not I_1385 (I25378,I25356);
nor I_1386 (I25395,I25378,I25169);
nor I_1387 (I25412,I25101,I25395);
DFFARX1 I_1388 (I25412,I1803,I25036,I25019,);
nor I_1389 (I25443,I25378,I25260);
nor I_1390 (I25460,I48975,I48963);
nor I_1391 (I25010,I25460,I25443);
not I_1392 (I25491,I25460);
nand I_1393 (I25013,I25220,I25491);
DFFARX1 I_1394 (I25460,I1803,I25036,I25025,);
DFFARX1 I_1395 (I25460,I1803,I25036,I25022,);
not I_1396 (I25580,I1810);
DFFARX1 I_1397 (I16539,I1803,I25580,I25606,);
DFFARX1 I_1398 (I25606,I1803,I25580,I25623,);
not I_1399 (I25572,I25623);
not I_1400 (I25645,I25606);
nand I_1401 (I25662,I16518,I16542);
and I_1402 (I25679,I25662,I16545);
DFFARX1 I_1403 (I25679,I1803,I25580,I25705,);
not I_1404 (I25713,I25705);
DFFARX1 I_1405 (I16527,I1803,I25580,I25739,);
and I_1406 (I25747,I25739,I16533);
nand I_1407 (I25764,I25739,I16533);
nand I_1408 (I25551,I25713,I25764);
DFFARX1 I_1409 (I16521,I1803,I25580,I25804,);
nor I_1410 (I25812,I25804,I25747);
DFFARX1 I_1411 (I25812,I1803,I25580,I25545,);
nor I_1412 (I25560,I25804,I25705);
nand I_1413 (I25857,I16530,I16518);
and I_1414 (I25874,I25857,I16524);
DFFARX1 I_1415 (I25874,I1803,I25580,I25900,);
nor I_1416 (I25548,I25900,I25804);
not I_1417 (I25922,I25900);
nor I_1418 (I25939,I25922,I25713);
nor I_1419 (I25956,I25645,I25939);
DFFARX1 I_1420 (I25956,I1803,I25580,I25563,);
nor I_1421 (I25987,I25922,I25804);
nor I_1422 (I26004,I16536,I16518);
nor I_1423 (I25554,I26004,I25987);
not I_1424 (I26035,I26004);
nand I_1425 (I25557,I25764,I26035);
DFFARX1 I_1426 (I26004,I1803,I25580,I25569,);
DFFARX1 I_1427 (I26004,I1803,I25580,I25566,);
not I_1428 (I26124,I1810);
DFFARX1 I_1429 (I11903,I1803,I26124,I26150,);
DFFARX1 I_1430 (I26150,I1803,I26124,I26167,);
not I_1431 (I26116,I26167);
not I_1432 (I26189,I26150);
nand I_1433 (I26206,I11915,I11894);
and I_1434 (I26223,I26206,I11897);
DFFARX1 I_1435 (I26223,I1803,I26124,I26249,);
not I_1436 (I26257,I26249);
DFFARX1 I_1437 (I11906,I1803,I26124,I26283,);
and I_1438 (I26291,I26283,I11918);
nand I_1439 (I26308,I26283,I11918);
nand I_1440 (I26095,I26257,I26308);
DFFARX1 I_1441 (I11912,I1803,I26124,I26348,);
nor I_1442 (I26356,I26348,I26291);
DFFARX1 I_1443 (I26356,I1803,I26124,I26089,);
nor I_1444 (I26104,I26348,I26249);
nand I_1445 (I26401,I11900,I11897);
and I_1446 (I26418,I26401,I11909);
DFFARX1 I_1447 (I26418,I1803,I26124,I26444,);
nor I_1448 (I26092,I26444,I26348);
not I_1449 (I26466,I26444);
nor I_1450 (I26483,I26466,I26257);
nor I_1451 (I26500,I26189,I26483);
DFFARX1 I_1452 (I26500,I1803,I26124,I26107,);
nor I_1453 (I26531,I26466,I26348);
nor I_1454 (I26548,I11894,I11897);
nor I_1455 (I26098,I26548,I26531);
not I_1456 (I26579,I26548);
nand I_1457 (I26101,I26308,I26579);
DFFARX1 I_1458 (I26548,I1803,I26124,I26113,);
DFFARX1 I_1459 (I26548,I1803,I26124,I26110,);
not I_1460 (I26668,I1810);
DFFARX1 I_1461 (I47912,I1803,I26668,I26694,);
DFFARX1 I_1462 (I26694,I1803,I26668,I26711,);
not I_1463 (I26660,I26711);
not I_1464 (I26733,I26694);
nand I_1465 (I26750,I47906,I47903);
and I_1466 (I26767,I26750,I47918);
DFFARX1 I_1467 (I26767,I1803,I26668,I26793,);
not I_1468 (I26801,I26793);
DFFARX1 I_1469 (I47906,I1803,I26668,I26827,);
and I_1470 (I26835,I26827,I47900);
nand I_1471 (I26852,I26827,I47900);
nand I_1472 (I26639,I26801,I26852);
DFFARX1 I_1473 (I47900,I1803,I26668,I26892,);
nor I_1474 (I26900,I26892,I26835);
DFFARX1 I_1475 (I26900,I1803,I26668,I26633,);
nor I_1476 (I26648,I26892,I26793);
nand I_1477 (I26945,I47915,I47909);
and I_1478 (I26962,I26945,I47903);
DFFARX1 I_1479 (I26962,I1803,I26668,I26988,);
nor I_1480 (I26636,I26988,I26892);
not I_1481 (I27010,I26988);
nor I_1482 (I27027,I27010,I26801);
nor I_1483 (I27044,I26733,I27027);
DFFARX1 I_1484 (I27044,I1803,I26668,I26651,);
nor I_1485 (I27075,I27010,I26892);
nor I_1486 (I27092,I47921,I47909);
nor I_1487 (I26642,I27092,I27075);
not I_1488 (I27123,I27092);
nand I_1489 (I26645,I26852,I27123);
DFFARX1 I_1490 (I27092,I1803,I26668,I26657,);
DFFARX1 I_1491 (I27092,I1803,I26668,I26654,);
not I_1492 (I27212,I1810);
DFFARX1 I_1493 (I76934,I1803,I27212,I27238,);
DFFARX1 I_1494 (I27238,I1803,I27212,I27255,);
not I_1495 (I27204,I27255);
not I_1496 (I27277,I27238);
nand I_1497 (I27294,I76940,I76943);
and I_1498 (I27311,I27294,I76919);
DFFARX1 I_1499 (I27311,I1803,I27212,I27337,);
not I_1500 (I27345,I27337);
DFFARX1 I_1501 (I76946,I1803,I27212,I27371,);
and I_1502 (I27379,I27371,I76928);
nand I_1503 (I27396,I27371,I76928);
nand I_1504 (I27183,I27345,I27396);
DFFARX1 I_1505 (I76925,I1803,I27212,I27436,);
nor I_1506 (I27444,I27436,I27379);
DFFARX1 I_1507 (I27444,I1803,I27212,I27177,);
nor I_1508 (I27192,I27436,I27337);
nand I_1509 (I27489,I76922,I76931);
and I_1510 (I27506,I27489,I76937);
DFFARX1 I_1511 (I27506,I1803,I27212,I27532,);
nor I_1512 (I27180,I27532,I27436);
not I_1513 (I27554,I27532);
nor I_1514 (I27571,I27554,I27345);
nor I_1515 (I27588,I27277,I27571);
DFFARX1 I_1516 (I27588,I1803,I27212,I27195,);
nor I_1517 (I27619,I27554,I27436);
nor I_1518 (I27636,I76919,I76931);
nor I_1519 (I27186,I27636,I27619);
not I_1520 (I27667,I27636);
nand I_1521 (I27189,I27396,I27667);
DFFARX1 I_1522 (I27636,I1803,I27212,I27201,);
DFFARX1 I_1523 (I27636,I1803,I27212,I27198,);
not I_1524 (I27756,I1810);
DFFARX1 I_1525 (I9197,I1803,I27756,I27782,);
DFFARX1 I_1526 (I27782,I1803,I27756,I27799,);
not I_1527 (I27748,I27799);
not I_1528 (I27821,I27782);
nand I_1529 (I27838,I9212,I9191);
and I_1530 (I27855,I27838,I9194);
DFFARX1 I_1531 (I27855,I1803,I27756,I27881,);
not I_1532 (I27889,I27881);
DFFARX1 I_1533 (I9200,I1803,I27756,I27915,);
and I_1534 (I27923,I27915,I9194);
nand I_1535 (I27940,I27915,I9194);
nand I_1536 (I27727,I27889,I27940);
DFFARX1 I_1537 (I9209,I1803,I27756,I27980,);
nor I_1538 (I27988,I27980,I27923);
DFFARX1 I_1539 (I27988,I1803,I27756,I27721,);
nor I_1540 (I27736,I27980,I27881);
nand I_1541 (I28033,I9191,I9206);
and I_1542 (I28050,I28033,I9203);
DFFARX1 I_1543 (I28050,I1803,I27756,I28076,);
nor I_1544 (I27724,I28076,I27980);
not I_1545 (I28098,I28076);
nor I_1546 (I28115,I28098,I27889);
nor I_1547 (I28132,I27821,I28115);
DFFARX1 I_1548 (I28132,I1803,I27756,I27739,);
nor I_1549 (I28163,I28098,I27980);
nor I_1550 (I28180,I9215,I9206);
nor I_1551 (I27730,I28180,I28163);
not I_1552 (I28211,I28180);
nand I_1553 (I27733,I27940,I28211);
DFFARX1 I_1554 (I28180,I1803,I27756,I27745,);
DFFARX1 I_1555 (I28180,I1803,I27756,I27742,);
not I_1556 (I28300,I1810);
DFFARX1 I_1557 (I6035,I1803,I28300,I28326,);
DFFARX1 I_1558 (I28326,I1803,I28300,I28343,);
not I_1559 (I28292,I28343);
not I_1560 (I28365,I28326);
nand I_1561 (I28382,I6050,I6029);
and I_1562 (I28399,I28382,I6032);
DFFARX1 I_1563 (I28399,I1803,I28300,I28425,);
not I_1564 (I28433,I28425);
DFFARX1 I_1565 (I6038,I1803,I28300,I28459,);
and I_1566 (I28467,I28459,I6032);
nand I_1567 (I28484,I28459,I6032);
nand I_1568 (I28271,I28433,I28484);
DFFARX1 I_1569 (I6047,I1803,I28300,I28524,);
nor I_1570 (I28532,I28524,I28467);
DFFARX1 I_1571 (I28532,I1803,I28300,I28265,);
nor I_1572 (I28280,I28524,I28425);
nand I_1573 (I28577,I6029,I6044);
and I_1574 (I28594,I28577,I6041);
DFFARX1 I_1575 (I28594,I1803,I28300,I28620,);
nor I_1576 (I28268,I28620,I28524);
not I_1577 (I28642,I28620);
nor I_1578 (I28659,I28642,I28433);
nor I_1579 (I28676,I28365,I28659);
DFFARX1 I_1580 (I28676,I1803,I28300,I28283,);
nor I_1581 (I28707,I28642,I28524);
nor I_1582 (I28724,I6053,I6044);
nor I_1583 (I28274,I28724,I28707);
not I_1584 (I28755,I28724);
nand I_1585 (I28277,I28484,I28755);
DFFARX1 I_1586 (I28724,I1803,I28300,I28289,);
DFFARX1 I_1587 (I28724,I1803,I28300,I28286,);
not I_1588 (I28841,I1810);
DFFARX1 I_1589 (I21276,I1803,I28841,I28867,);
DFFARX1 I_1590 (I28867,I1803,I28841,I28884,);
not I_1591 (I28833,I28884);
DFFARX1 I_1592 (I21264,I1803,I28841,I28915,);
not I_1593 (I28923,I21267);
nor I_1594 (I28940,I28867,I28923);
not I_1595 (I28957,I21270);
not I_1596 (I28974,I21282);
nand I_1597 (I28991,I28974,I21270);
nor I_1598 (I29008,I28923,I28991);
nor I_1599 (I29025,I28915,I29008);
DFFARX1 I_1600 (I28974,I1803,I28841,I28830,);
nor I_1601 (I29056,I21282,I21273);
nand I_1602 (I29073,I29056,I21261);
nor I_1603 (I29090,I29073,I28957);
nand I_1604 (I28815,I29090,I21267);
DFFARX1 I_1605 (I29073,I1803,I28841,I28827,);
nand I_1606 (I29135,I28957,I21282);
nor I_1607 (I29152,I28957,I21282);
nand I_1608 (I28821,I28940,I29152);
not I_1609 (I29183,I21279);
nor I_1610 (I29200,I29183,I29135);
DFFARX1 I_1611 (I29200,I1803,I28841,I28809,);
nor I_1612 (I29231,I29183,I21285);
and I_1613 (I29248,I29231,I21288);
or I_1614 (I29265,I29248,I21261);
DFFARX1 I_1615 (I29265,I1803,I28841,I29291,);
nor I_1616 (I29299,I29291,I28915);
nor I_1617 (I28818,I28867,I29299);
not I_1618 (I29330,I29291);
nor I_1619 (I29347,I29330,I29025);
DFFARX1 I_1620 (I29347,I1803,I28841,I28824,);
nand I_1621 (I29378,I29330,I28957);
nor I_1622 (I28812,I29183,I29378);
not I_1623 (I29436,I1810);
DFFARX1 I_1624 (I23369,I1803,I29436,I29462,);
DFFARX1 I_1625 (I29462,I1803,I29436,I29479,);
not I_1626 (I29428,I29479);
DFFARX1 I_1627 (I23393,I1803,I29436,I29510,);
not I_1628 (I29518,I23372);
nor I_1629 (I29535,I29462,I29518);
not I_1630 (I29552,I23378);
not I_1631 (I29569,I23384);
nand I_1632 (I29586,I29569,I23378);
nor I_1633 (I29603,I29518,I29586);
nor I_1634 (I29620,I29510,I29603);
DFFARX1 I_1635 (I29569,I1803,I29436,I29425,);
nor I_1636 (I29651,I23384,I23396);
nand I_1637 (I29668,I29651,I23390);
nor I_1638 (I29685,I29668,I29552);
nand I_1639 (I29410,I29685,I23372);
DFFARX1 I_1640 (I29668,I1803,I29436,I29422,);
nand I_1641 (I29730,I29552,I23384);
nor I_1642 (I29747,I29552,I23384);
nand I_1643 (I29416,I29535,I29747);
not I_1644 (I29778,I23375);
nor I_1645 (I29795,I29778,I29730);
DFFARX1 I_1646 (I29795,I1803,I29436,I29404,);
nor I_1647 (I29826,I29778,I23369);
and I_1648 (I29843,I29826,I23387);
or I_1649 (I29860,I29843,I23381);
DFFARX1 I_1650 (I29860,I1803,I29436,I29886,);
nor I_1651 (I29894,I29886,I29510);
nor I_1652 (I29413,I29462,I29894);
not I_1653 (I29925,I29886);
nor I_1654 (I29942,I29925,I29620);
DFFARX1 I_1655 (I29942,I1803,I29436,I29419,);
nand I_1656 (I29973,I29925,I29552);
nor I_1657 (I29407,I29778,I29973);
not I_1658 (I30031,I1810);
DFFARX1 I_1659 (I56534,I1803,I30031,I30057,);
DFFARX1 I_1660 (I30057,I1803,I30031,I30074,);
not I_1661 (I30023,I30074);
DFFARX1 I_1662 (I56522,I1803,I30031,I30105,);
not I_1663 (I30113,I56519);
nor I_1664 (I30130,I30057,I30113);
not I_1665 (I30147,I56531);
not I_1666 (I30164,I56528);
nand I_1667 (I30181,I30164,I56531);
nor I_1668 (I30198,I30113,I30181);
nor I_1669 (I30215,I30105,I30198);
DFFARX1 I_1670 (I30164,I1803,I30031,I30020,);
nor I_1671 (I30246,I56528,I56537);
nand I_1672 (I30263,I30246,I56540);
nor I_1673 (I30280,I30263,I30147);
nand I_1674 (I30005,I30280,I56519);
DFFARX1 I_1675 (I30263,I1803,I30031,I30017,);
nand I_1676 (I30325,I30147,I56528);
nor I_1677 (I30342,I30147,I56528);
nand I_1678 (I30011,I30130,I30342);
not I_1679 (I30373,I56543);
nor I_1680 (I30390,I30373,I30325);
DFFARX1 I_1681 (I30390,I1803,I30031,I29999,);
nor I_1682 (I30421,I30373,I56546);
and I_1683 (I30438,I30421,I56525);
or I_1684 (I30455,I30438,I56519);
DFFARX1 I_1685 (I30455,I1803,I30031,I30481,);
nor I_1686 (I30489,I30481,I30105);
nor I_1687 (I30008,I30057,I30489);
not I_1688 (I30520,I30481);
nor I_1689 (I30537,I30520,I30215);
DFFARX1 I_1690 (I30537,I1803,I30031,I30014,);
nand I_1691 (I30568,I30520,I30147);
nor I_1692 (I30002,I30373,I30568);
not I_1693 (I30626,I1810);
DFFARX1 I_1694 (I71871,I1803,I30626,I30652,);
DFFARX1 I_1695 (I30652,I1803,I30626,I30669,);
not I_1696 (I30618,I30669);
DFFARX1 I_1697 (I71853,I1803,I30626,I30700,);
not I_1698 (I30708,I71859);
nor I_1699 (I30725,I30652,I30708);
not I_1700 (I30742,I71874);
not I_1701 (I30759,I71865);
nand I_1702 (I30776,I30759,I71874);
nor I_1703 (I30793,I30708,I30776);
nor I_1704 (I30810,I30700,I30793);
DFFARX1 I_1705 (I30759,I1803,I30626,I30615,);
nor I_1706 (I30841,I71865,I71877);
nand I_1707 (I30858,I30841,I71856);
nor I_1708 (I30875,I30858,I30742);
nand I_1709 (I30600,I30875,I71859);
DFFARX1 I_1710 (I30858,I1803,I30626,I30612,);
nand I_1711 (I30920,I30742,I71865);
nor I_1712 (I30937,I30742,I71865);
nand I_1713 (I30606,I30725,I30937);
not I_1714 (I30968,I71862);
nor I_1715 (I30985,I30968,I30920);
DFFARX1 I_1716 (I30985,I1803,I30626,I30594,);
nor I_1717 (I31016,I30968,I71868);
and I_1718 (I31033,I31016,I71853);
or I_1719 (I31050,I31033,I71856);
DFFARX1 I_1720 (I31050,I1803,I30626,I31076,);
nor I_1721 (I31084,I31076,I30700);
nor I_1722 (I30603,I30652,I31084);
not I_1723 (I31115,I31076);
nor I_1724 (I31132,I31115,I30810);
DFFARX1 I_1725 (I31132,I1803,I30626,I30609,);
nand I_1726 (I31163,I31115,I30742);
nor I_1727 (I30597,I30968,I31163);
not I_1728 (I31221,I1810);
DFFARX1 I_1729 (I22330,I1803,I31221,I31247,);
DFFARX1 I_1730 (I31247,I1803,I31221,I31264,);
not I_1731 (I31213,I31264);
DFFARX1 I_1732 (I22318,I1803,I31221,I31295,);
not I_1733 (I31303,I22321);
nor I_1734 (I31320,I31247,I31303);
not I_1735 (I31337,I22324);
not I_1736 (I31354,I22336);
nand I_1737 (I31371,I31354,I22324);
nor I_1738 (I31388,I31303,I31371);
nor I_1739 (I31405,I31295,I31388);
DFFARX1 I_1740 (I31354,I1803,I31221,I31210,);
nor I_1741 (I31436,I22336,I22327);
nand I_1742 (I31453,I31436,I22315);
nor I_1743 (I31470,I31453,I31337);
nand I_1744 (I31195,I31470,I22321);
DFFARX1 I_1745 (I31453,I1803,I31221,I31207,);
nand I_1746 (I31515,I31337,I22336);
nor I_1747 (I31532,I31337,I22336);
nand I_1748 (I31201,I31320,I31532);
not I_1749 (I31563,I22333);
nor I_1750 (I31580,I31563,I31515);
DFFARX1 I_1751 (I31580,I1803,I31221,I31189,);
nor I_1752 (I31611,I31563,I22339);
and I_1753 (I31628,I31611,I22342);
or I_1754 (I31645,I31628,I22315);
DFFARX1 I_1755 (I31645,I1803,I31221,I31671,);
nor I_1756 (I31679,I31671,I31295);
nor I_1757 (I31198,I31247,I31679);
not I_1758 (I31710,I31671);
nor I_1759 (I31727,I31710,I31405);
DFFARX1 I_1760 (I31727,I1803,I31221,I31204,);
nand I_1761 (I31758,I31710,I31337);
nor I_1762 (I31192,I31563,I31758);
not I_1763 (I31816,I1810);
DFFARX1 I_1764 (I19168,I1803,I31816,I31842,);
DFFARX1 I_1765 (I31842,I1803,I31816,I31859,);
not I_1766 (I31808,I31859);
DFFARX1 I_1767 (I19156,I1803,I31816,I31890,);
not I_1768 (I31898,I19159);
nor I_1769 (I31915,I31842,I31898);
not I_1770 (I31932,I19162);
not I_1771 (I31949,I19174);
nand I_1772 (I31966,I31949,I19162);
nor I_1773 (I31983,I31898,I31966);
nor I_1774 (I32000,I31890,I31983);
DFFARX1 I_1775 (I31949,I1803,I31816,I31805,);
nor I_1776 (I32031,I19174,I19165);
nand I_1777 (I32048,I32031,I19153);
nor I_1778 (I32065,I32048,I31932);
nand I_1779 (I31790,I32065,I19159);
DFFARX1 I_1780 (I32048,I1803,I31816,I31802,);
nand I_1781 (I32110,I31932,I19174);
nor I_1782 (I32127,I31932,I19174);
nand I_1783 (I31796,I31915,I32127);
not I_1784 (I32158,I19171);
nor I_1785 (I32175,I32158,I32110);
DFFARX1 I_1786 (I32175,I1803,I31816,I31784,);
nor I_1787 (I32206,I32158,I19177);
and I_1788 (I32223,I32206,I19180);
or I_1789 (I32240,I32223,I19153);
DFFARX1 I_1790 (I32240,I1803,I31816,I32266,);
nor I_1791 (I32274,I32266,I31890);
nor I_1792 (I31793,I31842,I32274);
not I_1793 (I32305,I32266);
nor I_1794 (I32322,I32305,I32000);
DFFARX1 I_1795 (I32322,I1803,I31816,I31799,);
nand I_1796 (I32353,I32305,I31932);
nor I_1797 (I31787,I32158,I32353);
not I_1798 (I32411,I1810);
DFFARX1 I_1799 (I53950,I1803,I32411,I32437,);
DFFARX1 I_1800 (I32437,I1803,I32411,I32454,);
not I_1801 (I32403,I32454);
DFFARX1 I_1802 (I53938,I1803,I32411,I32485,);
not I_1803 (I32493,I53935);
nor I_1804 (I32510,I32437,I32493);
not I_1805 (I32527,I53947);
not I_1806 (I32544,I53944);
nand I_1807 (I32561,I32544,I53947);
nor I_1808 (I32578,I32493,I32561);
nor I_1809 (I32595,I32485,I32578);
DFFARX1 I_1810 (I32544,I1803,I32411,I32400,);
nor I_1811 (I32626,I53944,I53953);
nand I_1812 (I32643,I32626,I53956);
nor I_1813 (I32660,I32643,I32527);
nand I_1814 (I32385,I32660,I53935);
DFFARX1 I_1815 (I32643,I1803,I32411,I32397,);
nand I_1816 (I32705,I32527,I53944);
nor I_1817 (I32722,I32527,I53944);
nand I_1818 (I32391,I32510,I32722);
not I_1819 (I32753,I53959);
nor I_1820 (I32770,I32753,I32705);
DFFARX1 I_1821 (I32770,I1803,I32411,I32379,);
nor I_1822 (I32801,I32753,I53962);
and I_1823 (I32818,I32801,I53941);
or I_1824 (I32835,I32818,I53935);
DFFARX1 I_1825 (I32835,I1803,I32411,I32861,);
nor I_1826 (I32869,I32861,I32485);
nor I_1827 (I32388,I32437,I32869);
not I_1828 (I32900,I32861);
nor I_1829 (I32917,I32900,I32595);
DFFARX1 I_1830 (I32917,I1803,I32411,I32394,);
nand I_1831 (I32948,I32900,I32527);
nor I_1832 (I32382,I32753,I32948);
not I_1833 (I33006,I1810);
DFFARX1 I_1834 (I10269,I1803,I33006,I33032,);
not I_1835 (I33040,I33032);
DFFARX1 I_1836 (I10248,I1803,I33006,I33066,);
not I_1837 (I33074,I10245);
nand I_1838 (I33091,I33074,I10260);
not I_1839 (I33108,I33091);
nor I_1840 (I33125,I33108,I10248);
nor I_1841 (I33142,I33040,I33125);
DFFARX1 I_1842 (I33142,I1803,I33006,I32992,);
not I_1843 (I33173,I10248);
nand I_1844 (I33190,I33173,I33108);
and I_1845 (I33207,I33173,I10251);
nand I_1846 (I33224,I33207,I10266);
nor I_1847 (I32989,I33224,I33173);
and I_1848 (I32980,I33066,I33224);
not I_1849 (I33269,I33224);
nand I_1850 (I32983,I33066,I33269);
nor I_1851 (I32977,I33032,I33224);
not I_1852 (I33314,I10257);
nor I_1853 (I33331,I33314,I10251);
nand I_1854 (I33348,I33331,I33173);
nor I_1855 (I32986,I33091,I33348);
nor I_1856 (I33379,I33314,I10245);
and I_1857 (I33396,I33379,I10254);
or I_1858 (I33413,I33396,I10263);
DFFARX1 I_1859 (I33413,I1803,I33006,I33439,);
nor I_1860 (I33447,I33439,I33190);
DFFARX1 I_1861 (I33447,I1803,I33006,I32974,);
DFFARX1 I_1862 (I33439,I1803,I33006,I32998,);
not I_1863 (I33492,I33439);
nor I_1864 (I33509,I33492,I33066);
nor I_1865 (I33526,I33331,I33509);
DFFARX1 I_1866 (I33526,I1803,I33006,I32995,);
not I_1867 (I33584,I1810);
DFFARX1 I_1868 (I1772,I1803,I33584,I33610,);
not I_1869 (I33618,I33610);
DFFARX1 I_1870 (I1692,I1803,I33584,I33644,);
not I_1871 (I33652,I1452);
nand I_1872 (I33669,I33652,I1628);
not I_1873 (I33686,I33669);
nor I_1874 (I33703,I33686,I1492);
nor I_1875 (I33720,I33618,I33703);
DFFARX1 I_1876 (I33720,I1803,I33584,I33570,);
not I_1877 (I33751,I1492);
nand I_1878 (I33768,I33751,I33686);
and I_1879 (I33785,I33751,I1396);
nand I_1880 (I33802,I33785,I1668);
nor I_1881 (I33567,I33802,I33751);
and I_1882 (I33558,I33644,I33802);
not I_1883 (I33847,I33802);
nand I_1884 (I33561,I33644,I33847);
nor I_1885 (I33555,I33610,I33802);
not I_1886 (I33892,I1484);
nor I_1887 (I33909,I33892,I1396);
nand I_1888 (I33926,I33909,I33751);
nor I_1889 (I33564,I33669,I33926);
nor I_1890 (I33957,I33892,I1716);
and I_1891 (I33974,I33957,I1620);
or I_1892 (I33991,I33974,I1564);
DFFARX1 I_1893 (I33991,I1803,I33584,I34017,);
nor I_1894 (I34025,I34017,I33768);
DFFARX1 I_1895 (I34025,I1803,I33584,I33552,);
DFFARX1 I_1896 (I34017,I1803,I33584,I33576,);
not I_1897 (I34070,I34017);
nor I_1898 (I34087,I34070,I33644);
nor I_1899 (I34104,I33909,I34087);
DFFARX1 I_1900 (I34104,I1803,I33584,I33573,);
not I_1901 (I34162,I1810);
DFFARX1 I_1902 (I11314,I1803,I34162,I34188,);
not I_1903 (I34196,I34188);
DFFARX1 I_1904 (I11299,I1803,I34162,I34222,);
not I_1905 (I34230,I11317);
nand I_1906 (I34247,I34230,I11302);
not I_1907 (I34264,I34247);
nor I_1908 (I34281,I34264,I11299);
nor I_1909 (I34298,I34196,I34281);
DFFARX1 I_1910 (I34298,I1803,I34162,I34148,);
not I_1911 (I34329,I11299);
nand I_1912 (I34346,I34329,I34264);
and I_1913 (I34363,I34329,I11302);
nand I_1914 (I34380,I34363,I11323);
nor I_1915 (I34145,I34380,I34329);
and I_1916 (I34136,I34222,I34380);
not I_1917 (I34425,I34380);
nand I_1918 (I34139,I34222,I34425);
nor I_1919 (I34133,I34188,I34380);
not I_1920 (I34470,I11311);
nor I_1921 (I34487,I34470,I11302);
nand I_1922 (I34504,I34487,I34329);
nor I_1923 (I34142,I34247,I34504);
nor I_1924 (I34535,I34470,I11305);
and I_1925 (I34552,I34535,I11320);
or I_1926 (I34569,I34552,I11308);
DFFARX1 I_1927 (I34569,I1803,I34162,I34595,);
nor I_1928 (I34603,I34595,I34346);
DFFARX1 I_1929 (I34603,I1803,I34162,I34130,);
DFFARX1 I_1930 (I34595,I1803,I34162,I34154,);
not I_1931 (I34648,I34595);
nor I_1932 (I34665,I34648,I34222);
nor I_1933 (I34682,I34487,I34665);
DFFARX1 I_1934 (I34682,I1803,I34162,I34151,);
not I_1935 (I34740,I1810);
DFFARX1 I_1936 (I18105,I1803,I34740,I34766,);
not I_1937 (I34774,I34766);
DFFARX1 I_1938 (I18120,I1803,I34740,I34800,);
not I_1939 (I34808,I18123);
nand I_1940 (I34825,I34808,I18102);
not I_1941 (I34842,I34825);
nor I_1942 (I34859,I34842,I18126);
nor I_1943 (I34876,I34774,I34859);
DFFARX1 I_1944 (I34876,I1803,I34740,I34726,);
not I_1945 (I34907,I18126);
nand I_1946 (I34924,I34907,I34842);
and I_1947 (I34941,I34907,I18108);
nand I_1948 (I34958,I34941,I18099);
nor I_1949 (I34723,I34958,I34907);
and I_1950 (I34714,I34800,I34958);
not I_1951 (I35003,I34958);
nand I_1952 (I34717,I34800,I35003);
nor I_1953 (I34711,I34766,I34958);
not I_1954 (I35048,I18099);
nor I_1955 (I35065,I35048,I18108);
nand I_1956 (I35082,I35065,I34907);
nor I_1957 (I34720,I34825,I35082);
nor I_1958 (I35113,I35048,I18114);
and I_1959 (I35130,I35113,I18117);
or I_1960 (I35147,I35130,I18111);
DFFARX1 I_1961 (I35147,I1803,I34740,I35173,);
nor I_1962 (I35181,I35173,I34924);
DFFARX1 I_1963 (I35181,I1803,I34740,I34708,);
DFFARX1 I_1964 (I35173,I1803,I34740,I34732,);
not I_1965 (I35226,I35173);
nor I_1966 (I35243,I35226,I34800);
nor I_1967 (I35260,I35065,I35243);
DFFARX1 I_1968 (I35260,I1803,I34740,I34729,);
not I_1969 (I35318,I1810);
DFFARX1 I_1970 (I71275,I1803,I35318,I35344,);
not I_1971 (I35352,I35344);
DFFARX1 I_1972 (I71281,I1803,I35318,I35378,);
not I_1973 (I35386,I71275);
nand I_1974 (I35403,I35386,I71278);
not I_1975 (I35420,I35403);
nor I_1976 (I35437,I35420,I71296);
nor I_1977 (I35454,I35352,I35437);
DFFARX1 I_1978 (I35454,I1803,I35318,I35304,);
not I_1979 (I35485,I71296);
nand I_1980 (I35502,I35485,I35420);
and I_1981 (I35519,I35485,I71299);
nand I_1982 (I35536,I35519,I71278);
nor I_1983 (I35301,I35536,I35485);
and I_1984 (I35292,I35378,I35536);
not I_1985 (I35581,I35536);
nand I_1986 (I35295,I35378,I35581);
nor I_1987 (I35289,I35344,I35536);
not I_1988 (I35626,I71284);
nor I_1989 (I35643,I35626,I71299);
nand I_1990 (I35660,I35643,I35485);
nor I_1991 (I35298,I35403,I35660);
nor I_1992 (I35691,I35626,I71290);
and I_1993 (I35708,I35691,I71287);
or I_1994 (I35725,I35708,I71293);
DFFARX1 I_1995 (I35725,I1803,I35318,I35751,);
nor I_1996 (I35759,I35751,I35502);
DFFARX1 I_1997 (I35759,I1803,I35318,I35286,);
DFFARX1 I_1998 (I35751,I1803,I35318,I35310,);
not I_1999 (I35804,I35751);
nor I_2000 (I35821,I35804,I35378);
nor I_2001 (I35838,I35643,I35821);
DFFARX1 I_2002 (I35838,I1803,I35318,I35307,);
not I_2003 (I35896,I1810);
DFFARX1 I_2004 (I74115,I1803,I35896,I35922,);
not I_2005 (I35930,I35922);
DFFARX1 I_2006 (I74109,I1803,I35896,I35956,);
not I_2007 (I35964,I74118);
nand I_2008 (I35981,I35964,I74097);
not I_2009 (I35998,I35981);
nor I_2010 (I36015,I35998,I74106);
nor I_2011 (I36032,I35930,I36015);
DFFARX1 I_2012 (I36032,I1803,I35896,I35882,);
not I_2013 (I36063,I74106);
nand I_2014 (I36080,I36063,I35998);
and I_2015 (I36097,I36063,I74121);
nand I_2016 (I36114,I36097,I74100);
nor I_2017 (I35879,I36114,I36063);
and I_2018 (I35870,I35956,I36114);
not I_2019 (I36159,I36114);
nand I_2020 (I35873,I35956,I36159);
nor I_2021 (I35867,I35922,I36114);
not I_2022 (I36204,I74103);
nor I_2023 (I36221,I36204,I74121);
nand I_2024 (I36238,I36221,I36063);
nor I_2025 (I35876,I35981,I36238);
nor I_2026 (I36269,I36204,I74112);
and I_2027 (I36286,I36269,I74100);
or I_2028 (I36303,I36286,I74097);
DFFARX1 I_2029 (I36303,I1803,I35896,I36329,);
nor I_2030 (I36337,I36329,I36080);
DFFARX1 I_2031 (I36337,I1803,I35896,I35864,);
DFFARX1 I_2032 (I36329,I1803,I35896,I35888,);
not I_2033 (I36382,I36329);
nor I_2034 (I36399,I36382,I35956);
nor I_2035 (I36416,I36221,I36399);
DFFARX1 I_2036 (I36416,I1803,I35896,I35885,);
not I_2037 (I36474,I1810);
DFFARX1 I_2038 (I43378,I1803,I36474,I36500,);
not I_2039 (I36508,I36500);
DFFARX1 I_2040 (I43390,I1803,I36474,I36534,);
not I_2041 (I36542,I43381);
nand I_2042 (I36559,I36542,I43384);
not I_2043 (I36576,I36559);
nor I_2044 (I36593,I36576,I43387);
nor I_2045 (I36610,I36508,I36593);
DFFARX1 I_2046 (I36610,I1803,I36474,I36460,);
not I_2047 (I36641,I43387);
nand I_2048 (I36658,I36641,I36576);
and I_2049 (I36675,I36641,I43381);
nand I_2050 (I36692,I36675,I43393);
nor I_2051 (I36457,I36692,I36641);
and I_2052 (I36448,I36534,I36692);
not I_2053 (I36737,I36692);
nand I_2054 (I36451,I36534,I36737);
nor I_2055 (I36445,I36500,I36692);
not I_2056 (I36782,I43399);
nor I_2057 (I36799,I36782,I43381);
nand I_2058 (I36816,I36799,I36641);
nor I_2059 (I36454,I36559,I36816);
nor I_2060 (I36847,I36782,I43378);
and I_2061 (I36864,I36847,I43396);
or I_2062 (I36881,I36864,I43402);
DFFARX1 I_2063 (I36881,I1803,I36474,I36907,);
nor I_2064 (I36915,I36907,I36658);
DFFARX1 I_2065 (I36915,I1803,I36474,I36442,);
DFFARX1 I_2066 (I36907,I1803,I36474,I36466,);
not I_2067 (I36960,I36907);
nor I_2068 (I36977,I36960,I36534);
nor I_2069 (I36994,I36799,I36977);
DFFARX1 I_2070 (I36994,I1803,I36474,I36463,);
not I_2071 (I37052,I1810);
DFFARX1 I_2072 (I43956,I1803,I37052,I37078,);
not I_2073 (I37086,I37078);
DFFARX1 I_2074 (I43968,I1803,I37052,I37112,);
not I_2075 (I37120,I43959);
nand I_2076 (I37137,I37120,I43962);
not I_2077 (I37154,I37137);
nor I_2078 (I37171,I37154,I43965);
nor I_2079 (I37188,I37086,I37171);
DFFARX1 I_2080 (I37188,I1803,I37052,I37038,);
not I_2081 (I37219,I43965);
nand I_2082 (I37236,I37219,I37154);
and I_2083 (I37253,I37219,I43959);
nand I_2084 (I37270,I37253,I43971);
nor I_2085 (I37035,I37270,I37219);
and I_2086 (I37026,I37112,I37270);
not I_2087 (I37315,I37270);
nand I_2088 (I37029,I37112,I37315);
nor I_2089 (I37023,I37078,I37270);
not I_2090 (I37360,I43977);
nor I_2091 (I37377,I37360,I43959);
nand I_2092 (I37394,I37377,I37219);
nor I_2093 (I37032,I37137,I37394);
nor I_2094 (I37425,I37360,I43956);
and I_2095 (I37442,I37425,I43974);
or I_2096 (I37459,I37442,I43980);
DFFARX1 I_2097 (I37459,I1803,I37052,I37485,);
nor I_2098 (I37493,I37485,I37236);
DFFARX1 I_2099 (I37493,I1803,I37052,I37020,);
DFFARX1 I_2100 (I37485,I1803,I37052,I37044,);
not I_2101 (I37538,I37485);
nor I_2102 (I37555,I37538,I37112);
nor I_2103 (I37572,I37377,I37555);
DFFARX1 I_2104 (I37572,I1803,I37052,I37041,);
not I_2105 (I37630,I1810);
DFFARX1 I_2106 (I7107,I1803,I37630,I37656,);
not I_2107 (I37664,I37656);
DFFARX1 I_2108 (I7086,I1803,I37630,I37690,);
not I_2109 (I37698,I7083);
nand I_2110 (I37715,I37698,I7098);
not I_2111 (I37732,I37715);
nor I_2112 (I37749,I37732,I7086);
nor I_2113 (I37766,I37664,I37749);
DFFARX1 I_2114 (I37766,I1803,I37630,I37616,);
not I_2115 (I37797,I7086);
nand I_2116 (I37814,I37797,I37732);
and I_2117 (I37831,I37797,I7089);
nand I_2118 (I37848,I37831,I7104);
nor I_2119 (I37613,I37848,I37797);
and I_2120 (I37604,I37690,I37848);
not I_2121 (I37893,I37848);
nand I_2122 (I37607,I37690,I37893);
nor I_2123 (I37601,I37656,I37848);
not I_2124 (I37938,I7095);
nor I_2125 (I37955,I37938,I7089);
nand I_2126 (I37972,I37955,I37797);
nor I_2127 (I37610,I37715,I37972);
nor I_2128 (I38003,I37938,I7083);
and I_2129 (I38020,I38003,I7092);
or I_2130 (I38037,I38020,I7101);
DFFARX1 I_2131 (I38037,I1803,I37630,I38063,);
nor I_2132 (I38071,I38063,I37814);
DFFARX1 I_2133 (I38071,I1803,I37630,I37598,);
DFFARX1 I_2134 (I38063,I1803,I37630,I37622,);
not I_2135 (I38116,I38063);
nor I_2136 (I38133,I38116,I37690);
nor I_2137 (I38150,I37955,I38133);
DFFARX1 I_2138 (I38150,I1803,I37630,I37619,);
not I_2139 (I38208,I1810);
DFFARX1 I_2140 (I47388,I1803,I38208,I38234,);
not I_2141 (I38242,I38234);
nand I_2142 (I38259,I47376,I47394);
and I_2143 (I38276,I38259,I47391);
DFFARX1 I_2144 (I38276,I1803,I38208,I38302,);
not I_2145 (I38310,I47382);
DFFARX1 I_2146 (I47379,I1803,I38208,I38336,);
not I_2147 (I38344,I38336);
nor I_2148 (I38361,I38344,I38242);
and I_2149 (I38378,I38361,I47382);
nor I_2150 (I38395,I38344,I38310);
nor I_2151 (I38191,I38302,I38395);
DFFARX1 I_2152 (I47373,I1803,I38208,I38435,);
nor I_2153 (I38443,I38435,I38302);
not I_2154 (I38460,I38443);
not I_2155 (I38477,I38435);
nor I_2156 (I38494,I38477,I38378);
DFFARX1 I_2157 (I38494,I1803,I38208,I38194,);
nand I_2158 (I38525,I47373,I47376);
and I_2159 (I38542,I38525,I47379);
DFFARX1 I_2160 (I38542,I1803,I38208,I38568,);
nor I_2161 (I38576,I38568,I38435);
DFFARX1 I_2162 (I38576,I1803,I38208,I38176,);
nand I_2163 (I38607,I38568,I38477);
nand I_2164 (I38185,I38460,I38607);
not I_2165 (I38638,I38568);
nor I_2166 (I38655,I38638,I38378);
DFFARX1 I_2167 (I38655,I1803,I38208,I38197,);
nor I_2168 (I38686,I47385,I47376);
or I_2169 (I38188,I38435,I38686);
nor I_2170 (I38179,I38568,I38686);
or I_2171 (I38182,I38302,I38686);
DFFARX1 I_2172 (I38686,I1803,I38208,I38200,);
not I_2173 (I38786,I1810);
DFFARX1 I_2174 (I63779,I1803,I38786,I38812,);
not I_2175 (I38820,I38812);
nand I_2176 (I38837,I63761,I63773);
and I_2177 (I38854,I38837,I63776);
DFFARX1 I_2178 (I38854,I1803,I38786,I38880,);
not I_2179 (I38888,I63770);
DFFARX1 I_2180 (I63767,I1803,I38786,I38914,);
not I_2181 (I38922,I38914);
nor I_2182 (I38939,I38922,I38820);
and I_2183 (I38956,I38939,I63770);
nor I_2184 (I38973,I38922,I38888);
nor I_2185 (I38769,I38880,I38973);
DFFARX1 I_2186 (I63785,I1803,I38786,I39013,);
nor I_2187 (I39021,I39013,I38880);
not I_2188 (I39038,I39021);
not I_2189 (I39055,I39013);
nor I_2190 (I39072,I39055,I38956);
DFFARX1 I_2191 (I39072,I1803,I38786,I38772,);
nand I_2192 (I39103,I63764,I63764);
and I_2193 (I39120,I39103,I63761);
DFFARX1 I_2194 (I39120,I1803,I38786,I39146,);
nor I_2195 (I39154,I39146,I39013);
DFFARX1 I_2196 (I39154,I1803,I38786,I38754,);
nand I_2197 (I39185,I39146,I39055);
nand I_2198 (I38763,I39038,I39185);
not I_2199 (I39216,I39146);
nor I_2200 (I39233,I39216,I38956);
DFFARX1 I_2201 (I39233,I1803,I38786,I38775,);
nor I_2202 (I39264,I63782,I63764);
or I_2203 (I38766,I39013,I39264);
nor I_2204 (I38757,I39146,I39264);
or I_2205 (I38760,I38880,I39264);
DFFARX1 I_2206 (I39264,I1803,I38786,I38778,);
not I_2207 (I39364,I1810);
DFFARX1 I_2208 (I76341,I1803,I39364,I39390,);
not I_2209 (I39398,I39390);
nand I_2210 (I39415,I76365,I76347);
and I_2211 (I39432,I39415,I76353);
DFFARX1 I_2212 (I39432,I1803,I39364,I39458,);
not I_2213 (I39466,I76359);
DFFARX1 I_2214 (I76344,I1803,I39364,I39492,);
not I_2215 (I39500,I39492);
nor I_2216 (I39517,I39500,I39398);
and I_2217 (I39534,I39517,I76359);
nor I_2218 (I39551,I39500,I39466);
nor I_2219 (I39347,I39458,I39551);
DFFARX1 I_2220 (I76356,I1803,I39364,I39591,);
nor I_2221 (I39599,I39591,I39458);
not I_2222 (I39616,I39599);
not I_2223 (I39633,I39591);
nor I_2224 (I39650,I39633,I39534);
DFFARX1 I_2225 (I39650,I1803,I39364,I39350,);
nand I_2226 (I39681,I76362,I76350);
and I_2227 (I39698,I39681,I76344);
DFFARX1 I_2228 (I39698,I1803,I39364,I39724,);
nor I_2229 (I39732,I39724,I39591);
DFFARX1 I_2230 (I39732,I1803,I39364,I39332,);
nand I_2231 (I39763,I39724,I39633);
nand I_2232 (I39341,I39616,I39763);
not I_2233 (I39794,I39724);
nor I_2234 (I39811,I39794,I39534);
DFFARX1 I_2235 (I39811,I1803,I39364,I39353,);
nor I_2236 (I39842,I76341,I76350);
or I_2237 (I39344,I39591,I39842);
nor I_2238 (I39335,I39724,I39842);
or I_2239 (I39338,I39458,I39842);
DFFARX1 I_2240 (I39842,I1803,I39364,I39356,);
not I_2241 (I39942,I1810);
DFFARX1 I_2242 (I28274,I1803,I39942,I39968,);
not I_2243 (I39976,I39968);
nand I_2244 (I39993,I28265,I28283);
and I_2245 (I40010,I39993,I28286);
DFFARX1 I_2246 (I40010,I1803,I39942,I40036,);
not I_2247 (I40044,I28280);
DFFARX1 I_2248 (I28268,I1803,I39942,I40070,);
not I_2249 (I40078,I40070);
nor I_2250 (I40095,I40078,I39976);
and I_2251 (I40112,I40095,I28280);
nor I_2252 (I40129,I40078,I40044);
nor I_2253 (I39925,I40036,I40129);
DFFARX1 I_2254 (I28277,I1803,I39942,I40169,);
nor I_2255 (I40177,I40169,I40036);
not I_2256 (I40194,I40177);
not I_2257 (I40211,I40169);
nor I_2258 (I40228,I40211,I40112);
DFFARX1 I_2259 (I40228,I1803,I39942,I39928,);
nand I_2260 (I40259,I28292,I28289);
and I_2261 (I40276,I40259,I28271);
DFFARX1 I_2262 (I40276,I1803,I39942,I40302,);
nor I_2263 (I40310,I40302,I40169);
DFFARX1 I_2264 (I40310,I1803,I39942,I39910,);
nand I_2265 (I40341,I40302,I40211);
nand I_2266 (I39919,I40194,I40341);
not I_2267 (I40372,I40302);
nor I_2268 (I40389,I40372,I40112);
DFFARX1 I_2269 (I40389,I1803,I39942,I39931,);
nor I_2270 (I40420,I28265,I28289);
or I_2271 (I39922,I40169,I40420);
nor I_2272 (I39913,I40302,I40420);
or I_2273 (I39916,I40036,I40420);
DFFARX1 I_2274 (I40420,I1803,I39942,I39934,);
not I_2275 (I40520,I1810);
DFFARX1 I_2276 (I65513,I1803,I40520,I40546,);
not I_2277 (I40554,I40546);
nand I_2278 (I40571,I65495,I65507);
and I_2279 (I40588,I40571,I65510);
DFFARX1 I_2280 (I40588,I1803,I40520,I40614,);
not I_2281 (I40622,I65504);
DFFARX1 I_2282 (I65501,I1803,I40520,I40648,);
not I_2283 (I40656,I40648);
nor I_2284 (I40673,I40656,I40554);
and I_2285 (I40690,I40673,I65504);
nor I_2286 (I40707,I40656,I40622);
nor I_2287 (I40503,I40614,I40707);
DFFARX1 I_2288 (I65519,I1803,I40520,I40747,);
nor I_2289 (I40755,I40747,I40614);
not I_2290 (I40772,I40755);
not I_2291 (I40789,I40747);
nor I_2292 (I40806,I40789,I40690);
DFFARX1 I_2293 (I40806,I1803,I40520,I40506,);
nand I_2294 (I40837,I65498,I65498);
and I_2295 (I40854,I40837,I65495);
DFFARX1 I_2296 (I40854,I1803,I40520,I40880,);
nor I_2297 (I40888,I40880,I40747);
DFFARX1 I_2298 (I40888,I1803,I40520,I40488,);
nand I_2299 (I40919,I40880,I40789);
nand I_2300 (I40497,I40772,I40919);
not I_2301 (I40950,I40880);
nor I_2302 (I40967,I40950,I40690);
DFFARX1 I_2303 (I40967,I1803,I40520,I40509,);
nor I_2304 (I40998,I65516,I65498);
or I_2305 (I40500,I40747,I40998);
nor I_2306 (I40491,I40880,I40998);
or I_2307 (I40494,I40614,I40998);
DFFARX1 I_2308 (I40998,I1803,I40520,I40512,);
not I_2309 (I41098,I1810);
DFFARX1 I_2310 (I23922,I1803,I41098,I41124,);
not I_2311 (I41132,I41124);
nand I_2312 (I41149,I23913,I23931);
and I_2313 (I41166,I41149,I23934);
DFFARX1 I_2314 (I41166,I1803,I41098,I41192,);
not I_2315 (I41200,I23928);
DFFARX1 I_2316 (I23916,I1803,I41098,I41226,);
not I_2317 (I41234,I41226);
nor I_2318 (I41251,I41234,I41132);
and I_2319 (I41268,I41251,I23928);
nor I_2320 (I41285,I41234,I41200);
nor I_2321 (I41081,I41192,I41285);
DFFARX1 I_2322 (I23925,I1803,I41098,I41325,);
nor I_2323 (I41333,I41325,I41192);
not I_2324 (I41350,I41333);
not I_2325 (I41367,I41325);
nor I_2326 (I41384,I41367,I41268);
DFFARX1 I_2327 (I41384,I1803,I41098,I41084,);
nand I_2328 (I41415,I23940,I23937);
and I_2329 (I41432,I41415,I23919);
DFFARX1 I_2330 (I41432,I1803,I41098,I41458,);
nor I_2331 (I41466,I41458,I41325);
DFFARX1 I_2332 (I41466,I1803,I41098,I41066,);
nand I_2333 (I41497,I41458,I41367);
nand I_2334 (I41075,I41350,I41497);
not I_2335 (I41528,I41458);
nor I_2336 (I41545,I41528,I41268);
DFFARX1 I_2337 (I41545,I1803,I41098,I41087,);
nor I_2338 (I41576,I23913,I23937);
or I_2339 (I41078,I41325,I41576);
nor I_2340 (I41069,I41458,I41576);
or I_2341 (I41072,I41192,I41576);
DFFARX1 I_2342 (I41576,I1803,I41098,I41090,);
not I_2343 (I41676,I1810);
DFFARX1 I_2344 (I1825,I1803,I41676,I41702,);
not I_2345 (I41710,I41702);
nand I_2346 (I41727,I1822,I1813);
and I_2347 (I41744,I41727,I1813);
DFFARX1 I_2348 (I41744,I1803,I41676,I41770,);
not I_2349 (I41778,I1816);
DFFARX1 I_2350 (I1831,I1803,I41676,I41804,);
not I_2351 (I41812,I41804);
nor I_2352 (I41829,I41812,I41710);
and I_2353 (I41846,I41829,I1816);
nor I_2354 (I41863,I41812,I41778);
nor I_2355 (I41659,I41770,I41863);
DFFARX1 I_2356 (I1816,I1803,I41676,I41903,);
nor I_2357 (I41911,I41903,I41770);
not I_2358 (I41928,I41911);
not I_2359 (I41945,I41903);
nor I_2360 (I41962,I41945,I41846);
DFFARX1 I_2361 (I41962,I1803,I41676,I41662,);
nand I_2362 (I41993,I1834,I1819);
and I_2363 (I42010,I41993,I1837);
DFFARX1 I_2364 (I42010,I1803,I41676,I42036,);
nor I_2365 (I42044,I42036,I41903);
DFFARX1 I_2366 (I42044,I1803,I41676,I41644,);
nand I_2367 (I42075,I42036,I41945);
nand I_2368 (I41653,I41928,I42075);
not I_2369 (I42106,I42036);
nor I_2370 (I42123,I42106,I41846);
DFFARX1 I_2371 (I42123,I1803,I41676,I41665,);
nor I_2372 (I42154,I1828,I1819);
or I_2373 (I41656,I41903,I42154);
nor I_2374 (I41647,I42036,I42154);
or I_2375 (I41650,I41770,I42154);
DFFARX1 I_2376 (I42154,I1803,I41676,I41668,);
not I_2377 (I42254,I1810);
DFFARX1 I_2378 (I10775,I1803,I42254,I42280,);
not I_2379 (I42288,I42280);
nand I_2380 (I42305,I10784,I10793);
and I_2381 (I42322,I42305,I10772);
DFFARX1 I_2382 (I42322,I1803,I42254,I42348,);
not I_2383 (I42356,I10775);
DFFARX1 I_2384 (I10790,I1803,I42254,I42382,);
not I_2385 (I42390,I42382);
nor I_2386 (I42407,I42390,I42288);
and I_2387 (I42424,I42407,I10775);
nor I_2388 (I42441,I42390,I42356);
nor I_2389 (I42237,I42348,I42441);
DFFARX1 I_2390 (I10781,I1803,I42254,I42481,);
nor I_2391 (I42489,I42481,I42348);
not I_2392 (I42506,I42489);
not I_2393 (I42523,I42481);
nor I_2394 (I42540,I42523,I42424);
DFFARX1 I_2395 (I42540,I1803,I42254,I42240,);
nand I_2396 (I42571,I10796,I10772);
and I_2397 (I42588,I42571,I10778);
DFFARX1 I_2398 (I42588,I1803,I42254,I42614,);
nor I_2399 (I42622,I42614,I42481);
DFFARX1 I_2400 (I42622,I1803,I42254,I42222,);
nand I_2401 (I42653,I42614,I42523);
nand I_2402 (I42231,I42506,I42653);
not I_2403 (I42684,I42614);
nor I_2404 (I42701,I42684,I42424);
DFFARX1 I_2405 (I42701,I1803,I42254,I42243,);
nor I_2406 (I42732,I10787,I10772);
or I_2407 (I42234,I42481,I42732);
nor I_2408 (I42225,I42614,I42732);
or I_2409 (I42228,I42348,I42732);
DFFARX1 I_2410 (I42732,I1803,I42254,I42246,);
not I_2411 (I42832,I1810);
DFFARX1 I_2412 (I53313,I1803,I42832,I42858,);
not I_2413 (I42866,I42858);
nand I_2414 (I42883,I53289,I53304);
and I_2415 (I42900,I42883,I53316);
DFFARX1 I_2416 (I42900,I1803,I42832,I42926,);
not I_2417 (I42934,I53301);
DFFARX1 I_2418 (I53292,I1803,I42832,I42960,);
not I_2419 (I42968,I42960);
nor I_2420 (I42985,I42968,I42866);
and I_2421 (I43002,I42985,I53301);
nor I_2422 (I43019,I42968,I42934);
nor I_2423 (I42815,I42926,I43019);
DFFARX1 I_2424 (I53289,I1803,I42832,I43059,);
nor I_2425 (I43067,I43059,I42926);
not I_2426 (I43084,I43067);
not I_2427 (I43101,I43059);
nor I_2428 (I43118,I43101,I43002);
DFFARX1 I_2429 (I43118,I1803,I42832,I42818,);
nand I_2430 (I43149,I53307,I53298);
and I_2431 (I43166,I43149,I53310);
DFFARX1 I_2432 (I43166,I1803,I42832,I43192,);
nor I_2433 (I43200,I43192,I43059);
DFFARX1 I_2434 (I43200,I1803,I42832,I42800,);
nand I_2435 (I43231,I43192,I43101);
nand I_2436 (I42809,I43084,I43231);
not I_2437 (I43262,I43192);
nor I_2438 (I43279,I43262,I43002);
DFFARX1 I_2439 (I43279,I1803,I42832,I42821,);
nor I_2440 (I43310,I53295,I53298);
or I_2441 (I42812,I43059,I43310);
nor I_2442 (I42803,I43192,I43310);
or I_2443 (I42806,I42926,I43310);
DFFARX1 I_2444 (I43310,I1803,I42832,I42824,);
not I_2445 (I43410,I1810);
DFFARX1 I_2446 (I67247,I1803,I43410,I43436,);
not I_2447 (I43444,I43436);
nand I_2448 (I43461,I67229,I67241);
and I_2449 (I43478,I43461,I67244);
DFFARX1 I_2450 (I43478,I1803,I43410,I43504,);
not I_2451 (I43512,I67238);
DFFARX1 I_2452 (I67235,I1803,I43410,I43538,);
not I_2453 (I43546,I43538);
nor I_2454 (I43563,I43546,I43444);
and I_2455 (I43580,I43563,I67238);
nor I_2456 (I43597,I43546,I43512);
nor I_2457 (I43393,I43504,I43597);
DFFARX1 I_2458 (I67253,I1803,I43410,I43637,);
nor I_2459 (I43645,I43637,I43504);
not I_2460 (I43662,I43645);
not I_2461 (I43679,I43637);
nor I_2462 (I43696,I43679,I43580);
DFFARX1 I_2463 (I43696,I1803,I43410,I43396,);
nand I_2464 (I43727,I67232,I67232);
and I_2465 (I43744,I43727,I67229);
DFFARX1 I_2466 (I43744,I1803,I43410,I43770,);
nor I_2467 (I43778,I43770,I43637);
DFFARX1 I_2468 (I43778,I1803,I43410,I43378,);
nand I_2469 (I43809,I43770,I43679);
nand I_2470 (I43387,I43662,I43809);
not I_2471 (I43840,I43770);
nor I_2472 (I43857,I43840,I43580);
DFFARX1 I_2473 (I43857,I1803,I43410,I43399,);
nor I_2474 (I43888,I67250,I67232);
or I_2475 (I43390,I43637,I43888);
nor I_2476 (I43381,I43770,I43888);
or I_2477 (I43384,I43504,I43888);
DFFARX1 I_2478 (I43888,I1803,I43410,I43402,);
not I_2479 (I43988,I1810);
DFFARX1 I_2480 (I12489,I1803,I43988,I44014,);
not I_2481 (I44022,I44014);
nand I_2482 (I44039,I12492,I12513);
and I_2483 (I44056,I44039,I12501);
DFFARX1 I_2484 (I44056,I1803,I43988,I44082,);
not I_2485 (I44090,I12498);
DFFARX1 I_2486 (I12489,I1803,I43988,I44116,);
not I_2487 (I44124,I44116);
nor I_2488 (I44141,I44124,I44022);
and I_2489 (I44158,I44141,I12498);
nor I_2490 (I44175,I44124,I44090);
nor I_2491 (I43971,I44082,I44175);
DFFARX1 I_2492 (I12507,I1803,I43988,I44215,);
nor I_2493 (I44223,I44215,I44082);
not I_2494 (I44240,I44223);
not I_2495 (I44257,I44215);
nor I_2496 (I44274,I44257,I44158);
DFFARX1 I_2497 (I44274,I1803,I43988,I43974,);
nand I_2498 (I44305,I12492,I12495);
and I_2499 (I44322,I44305,I12504);
DFFARX1 I_2500 (I44322,I1803,I43988,I44348,);
nor I_2501 (I44356,I44348,I44215);
DFFARX1 I_2502 (I44356,I1803,I43988,I43956,);
nand I_2503 (I44387,I44348,I44257);
nand I_2504 (I43965,I44240,I44387);
not I_2505 (I44418,I44348);
nor I_2506 (I44435,I44418,I44158);
DFFARX1 I_2507 (I44435,I1803,I43988,I43977,);
nor I_2508 (I44466,I12510,I12495);
or I_2509 (I43968,I44215,I44466);
nor I_2510 (I43959,I44348,I44466);
or I_2511 (I43962,I44082,I44466);
DFFARX1 I_2512 (I44466,I1803,I43988,I43980,);
not I_2513 (I44566,I1810);
DFFARX1 I_2514 (I24466,I1803,I44566,I44592,);
not I_2515 (I44600,I44592);
nand I_2516 (I44617,I24457,I24475);
and I_2517 (I44634,I44617,I24478);
DFFARX1 I_2518 (I44634,I1803,I44566,I44660,);
not I_2519 (I44668,I24472);
DFFARX1 I_2520 (I24460,I1803,I44566,I44694,);
not I_2521 (I44702,I44694);
nor I_2522 (I44719,I44702,I44600);
and I_2523 (I44736,I44719,I24472);
nor I_2524 (I44753,I44702,I44668);
nor I_2525 (I44549,I44660,I44753);
DFFARX1 I_2526 (I24469,I1803,I44566,I44793,);
nor I_2527 (I44801,I44793,I44660);
not I_2528 (I44818,I44801);
not I_2529 (I44835,I44793);
nor I_2530 (I44852,I44835,I44736);
DFFARX1 I_2531 (I44852,I1803,I44566,I44552,);
nand I_2532 (I44883,I24484,I24481);
and I_2533 (I44900,I44883,I24463);
DFFARX1 I_2534 (I44900,I1803,I44566,I44926,);
nor I_2535 (I44934,I44926,I44793);
DFFARX1 I_2536 (I44934,I1803,I44566,I44534,);
nand I_2537 (I44965,I44926,I44835);
nand I_2538 (I44543,I44818,I44965);
not I_2539 (I44996,I44926);
nor I_2540 (I45013,I44996,I44736);
DFFARX1 I_2541 (I45013,I1803,I44566,I44555,);
nor I_2542 (I45044,I24457,I24481);
or I_2543 (I44546,I44793,I45044);
nor I_2544 (I44537,I44926,I45044);
or I_2545 (I44540,I44660,I45044);
DFFARX1 I_2546 (I45044,I1803,I44566,I44558,);
not I_2547 (I45144,I1810);
DFFARX1 I_2548 (I75185,I1803,I45144,I45170,);
not I_2549 (I45178,I45170);
nand I_2550 (I45195,I75209,I75191);
and I_2551 (I45212,I45195,I75197);
DFFARX1 I_2552 (I45212,I1803,I45144,I45238,);
not I_2553 (I45246,I75203);
DFFARX1 I_2554 (I75188,I1803,I45144,I45272,);
not I_2555 (I45280,I45272);
nor I_2556 (I45297,I45280,I45178);
and I_2557 (I45314,I45297,I75203);
nor I_2558 (I45331,I45280,I45246);
nor I_2559 (I45127,I45238,I45331);
DFFARX1 I_2560 (I75200,I1803,I45144,I45371,);
nor I_2561 (I45379,I45371,I45238);
not I_2562 (I45396,I45379);
not I_2563 (I45413,I45371);
nor I_2564 (I45430,I45413,I45314);
DFFARX1 I_2565 (I45430,I1803,I45144,I45130,);
nand I_2566 (I45461,I75206,I75194);
and I_2567 (I45478,I45461,I75188);
DFFARX1 I_2568 (I45478,I1803,I45144,I45504,);
nor I_2569 (I45512,I45504,I45371);
DFFARX1 I_2570 (I45512,I1803,I45144,I45112,);
nand I_2571 (I45543,I45504,I45413);
nand I_2572 (I45121,I45396,I45543);
not I_2573 (I45574,I45504);
nor I_2574 (I45591,I45574,I45314);
DFFARX1 I_2575 (I45591,I1803,I45144,I45133,);
nor I_2576 (I45622,I75185,I75194);
or I_2577 (I45124,I45371,I45622);
nor I_2578 (I45115,I45504,I45622);
or I_2579 (I45118,I45238,I45622);
DFFARX1 I_2580 (I45622,I1803,I45144,I45136,);
not I_2581 (I45722,I1810);
DFFARX1 I_2582 (I64935,I1803,I45722,I45748,);
not I_2583 (I45756,I45748);
nand I_2584 (I45773,I64917,I64929);
and I_2585 (I45790,I45773,I64932);
DFFARX1 I_2586 (I45790,I1803,I45722,I45816,);
not I_2587 (I45824,I64926);
DFFARX1 I_2588 (I64923,I1803,I45722,I45850,);
not I_2589 (I45858,I45850);
nor I_2590 (I45875,I45858,I45756);
and I_2591 (I45892,I45875,I64926);
nor I_2592 (I45909,I45858,I45824);
nor I_2593 (I45705,I45816,I45909);
DFFARX1 I_2594 (I64941,I1803,I45722,I45949,);
nor I_2595 (I45957,I45949,I45816);
not I_2596 (I45974,I45957);
not I_2597 (I45991,I45949);
nor I_2598 (I46008,I45991,I45892);
DFFARX1 I_2599 (I46008,I1803,I45722,I45708,);
nand I_2600 (I46039,I64920,I64920);
and I_2601 (I46056,I46039,I64917);
DFFARX1 I_2602 (I46056,I1803,I45722,I46082,);
nor I_2603 (I46090,I46082,I45949);
DFFARX1 I_2604 (I46090,I1803,I45722,I45690,);
nand I_2605 (I46121,I46082,I45991);
nand I_2606 (I45699,I45974,I46121);
not I_2607 (I46152,I46082);
nor I_2608 (I46169,I46152,I45892);
DFFARX1 I_2609 (I46169,I1803,I45722,I45711,);
nor I_2610 (I46200,I64938,I64920);
or I_2611 (I45702,I45949,I46200);
nor I_2612 (I45693,I46082,I46200);
or I_2613 (I45696,I45816,I46200);
DFFARX1 I_2614 (I46200,I1803,I45722,I45714,);
not I_2615 (I46300,I1810);
DFFARX1 I_2616 (I9721,I1803,I46300,I46326,);
not I_2617 (I46334,I46326);
nand I_2618 (I46351,I9730,I9739);
and I_2619 (I46368,I46351,I9718);
DFFARX1 I_2620 (I46368,I1803,I46300,I46394,);
not I_2621 (I46402,I9721);
DFFARX1 I_2622 (I9736,I1803,I46300,I46428,);
not I_2623 (I46436,I46428);
nor I_2624 (I46453,I46436,I46334);
and I_2625 (I46470,I46453,I9721);
nor I_2626 (I46487,I46436,I46402);
nor I_2627 (I46283,I46394,I46487);
DFFARX1 I_2628 (I9727,I1803,I46300,I46527,);
nor I_2629 (I46535,I46527,I46394);
not I_2630 (I46552,I46535);
not I_2631 (I46569,I46527);
nor I_2632 (I46586,I46569,I46470);
DFFARX1 I_2633 (I46586,I1803,I46300,I46286,);
nand I_2634 (I46617,I9742,I9718);
and I_2635 (I46634,I46617,I9724);
DFFARX1 I_2636 (I46634,I1803,I46300,I46660,);
nor I_2637 (I46668,I46660,I46527);
DFFARX1 I_2638 (I46668,I1803,I46300,I46268,);
nand I_2639 (I46699,I46660,I46569);
nand I_2640 (I46277,I46552,I46699);
not I_2641 (I46730,I46660);
nor I_2642 (I46747,I46730,I46470);
DFFARX1 I_2643 (I46747,I1803,I46300,I46289,);
nor I_2644 (I46778,I9733,I9718);
or I_2645 (I46280,I46527,I46778);
nor I_2646 (I46271,I46660,I46778);
or I_2647 (I46274,I46394,I46778);
DFFARX1 I_2648 (I46778,I1803,I46300,I46292,);
not I_2649 (I46875,I1810);
DFFARX1 I_2650 (I64357,I1803,I46875,I46901,);
not I_2651 (I46909,I46901);
nand I_2652 (I46926,I64339,I64339);
and I_2653 (I46943,I46926,I64345);
DFFARX1 I_2654 (I46943,I1803,I46875,I46969,);
DFFARX1 I_2655 (I46969,I1803,I46875,I46864,);
DFFARX1 I_2656 (I64342,I1803,I46875,I47000,);
nand I_2657 (I47008,I47000,I64351);
not I_2658 (I47025,I47008);
DFFARX1 I_2659 (I47025,I1803,I46875,I47051,);
not I_2660 (I47059,I47051);
nor I_2661 (I46867,I46909,I47059);
DFFARX1 I_2662 (I64363,I1803,I46875,I47099,);
nor I_2663 (I46858,I47099,I46969);
nor I_2664 (I46849,I47099,I47025);
nand I_2665 (I47135,I64354,I64348);
and I_2666 (I47152,I47135,I64342);
DFFARX1 I_2667 (I47152,I1803,I46875,I47178,);
not I_2668 (I47186,I47178);
nand I_2669 (I47203,I47186,I47099);
nand I_2670 (I46852,I47186,I47008);
nor I_2671 (I47234,I64360,I64348);
and I_2672 (I47251,I47099,I47234);
nor I_2673 (I47268,I47186,I47251);
DFFARX1 I_2674 (I47268,I1803,I46875,I46861,);
nor I_2675 (I47299,I46901,I47234);
DFFARX1 I_2676 (I47299,I1803,I46875,I46846,);
nor I_2677 (I47330,I47178,I47234);
not I_2678 (I47347,I47330);
nand I_2679 (I46855,I47347,I47203);
not I_2680 (I47402,I1810);
DFFARX1 I_2681 (I25551,I1803,I47402,I47428,);
not I_2682 (I47436,I47428);
nand I_2683 (I47453,I25548,I25557);
and I_2684 (I47470,I47453,I25566);
DFFARX1 I_2685 (I47470,I1803,I47402,I47496,);
DFFARX1 I_2686 (I47496,I1803,I47402,I47391,);
DFFARX1 I_2687 (I25569,I1803,I47402,I47527,);
nand I_2688 (I47535,I47527,I25572);
not I_2689 (I47552,I47535);
DFFARX1 I_2690 (I47552,I1803,I47402,I47578,);
not I_2691 (I47586,I47578);
nor I_2692 (I47394,I47436,I47586);
DFFARX1 I_2693 (I25545,I1803,I47402,I47626,);
nor I_2694 (I47385,I47626,I47496);
nor I_2695 (I47376,I47626,I47552);
nand I_2696 (I47662,I25560,I25563);
and I_2697 (I47679,I47662,I25554);
DFFARX1 I_2698 (I47679,I1803,I47402,I47705,);
not I_2699 (I47713,I47705);
nand I_2700 (I47730,I47713,I47626);
nand I_2701 (I47379,I47713,I47535);
nor I_2702 (I47761,I25545,I25563);
and I_2703 (I47778,I47626,I47761);
nor I_2704 (I47795,I47713,I47778);
DFFARX1 I_2705 (I47795,I1803,I47402,I47388,);
nor I_2706 (I47826,I47428,I47761);
DFFARX1 I_2707 (I47826,I1803,I47402,I47373,);
nor I_2708 (I47857,I47705,I47761);
not I_2709 (I47874,I47857);
nand I_2710 (I47382,I47874,I47730);
not I_2711 (I47929,I1810);
DFFARX1 I_2712 (I38176,I1803,I47929,I47955,);
not I_2713 (I47963,I47955);
nand I_2714 (I47980,I38179,I38176);
and I_2715 (I47997,I47980,I38188);
DFFARX1 I_2716 (I47997,I1803,I47929,I48023,);
DFFARX1 I_2717 (I48023,I1803,I47929,I47918,);
DFFARX1 I_2718 (I38185,I1803,I47929,I48054,);
nand I_2719 (I48062,I48054,I38191);
not I_2720 (I48079,I48062);
DFFARX1 I_2721 (I48079,I1803,I47929,I48105,);
not I_2722 (I48113,I48105);
nor I_2723 (I47921,I47963,I48113);
DFFARX1 I_2724 (I38200,I1803,I47929,I48153,);
nor I_2725 (I47912,I48153,I48023);
nor I_2726 (I47903,I48153,I48079);
nand I_2727 (I48189,I38194,I38182);
and I_2728 (I48206,I48189,I38179);
DFFARX1 I_2729 (I48206,I1803,I47929,I48232,);
not I_2730 (I48240,I48232);
nand I_2731 (I48257,I48240,I48153);
nand I_2732 (I47906,I48240,I48062);
nor I_2733 (I48288,I38197,I38182);
and I_2734 (I48305,I48153,I48288);
nor I_2735 (I48322,I48240,I48305);
DFFARX1 I_2736 (I48322,I1803,I47929,I47915,);
nor I_2737 (I48353,I47955,I48288);
DFFARX1 I_2738 (I48353,I1803,I47929,I47900,);
nor I_2739 (I48384,I48232,I48288);
not I_2740 (I48401,I48384);
nand I_2741 (I47909,I48401,I48257);
not I_2742 (I48456,I1810);
DFFARX1 I_2743 (I39910,I1803,I48456,I48482,);
not I_2744 (I48490,I48482);
nand I_2745 (I48507,I39913,I39910);
and I_2746 (I48524,I48507,I39922);
DFFARX1 I_2747 (I48524,I1803,I48456,I48550,);
DFFARX1 I_2748 (I48550,I1803,I48456,I48445,);
DFFARX1 I_2749 (I39919,I1803,I48456,I48581,);
nand I_2750 (I48589,I48581,I39925);
not I_2751 (I48606,I48589);
DFFARX1 I_2752 (I48606,I1803,I48456,I48632,);
not I_2753 (I48640,I48632);
nor I_2754 (I48448,I48490,I48640);
DFFARX1 I_2755 (I39934,I1803,I48456,I48680,);
nor I_2756 (I48439,I48680,I48550);
nor I_2757 (I48430,I48680,I48606);
nand I_2758 (I48716,I39928,I39916);
and I_2759 (I48733,I48716,I39913);
DFFARX1 I_2760 (I48733,I1803,I48456,I48759,);
not I_2761 (I48767,I48759);
nand I_2762 (I48784,I48767,I48680);
nand I_2763 (I48433,I48767,I48589);
nor I_2764 (I48815,I39931,I39916);
and I_2765 (I48832,I48680,I48815);
nor I_2766 (I48849,I48767,I48832);
DFFARX1 I_2767 (I48849,I1803,I48456,I48442,);
nor I_2768 (I48880,I48482,I48815);
DFFARX1 I_2769 (I48880,I1803,I48456,I48427,);
nor I_2770 (I48911,I48759,I48815);
not I_2771 (I48928,I48911);
nand I_2772 (I48436,I48928,I48784);
not I_2773 (I48983,I1810);
DFFARX1 I_2774 (I33567,I1803,I48983,I49009,);
not I_2775 (I49017,I49009);
nand I_2776 (I49034,I33552,I33573);
and I_2777 (I49051,I49034,I33561);
DFFARX1 I_2778 (I49051,I1803,I48983,I49077,);
DFFARX1 I_2779 (I49077,I1803,I48983,I48972,);
DFFARX1 I_2780 (I33555,I1803,I48983,I49108,);
nand I_2781 (I49116,I49108,I33564);
not I_2782 (I49133,I49116);
DFFARX1 I_2783 (I49133,I1803,I48983,I49159,);
not I_2784 (I49167,I49159);
nor I_2785 (I48975,I49017,I49167);
DFFARX1 I_2786 (I33570,I1803,I48983,I49207,);
nor I_2787 (I48966,I49207,I49077);
nor I_2788 (I48957,I49207,I49133);
nand I_2789 (I49243,I33552,I33555);
and I_2790 (I49260,I49243,I33576);
DFFARX1 I_2791 (I49260,I1803,I48983,I49286,);
not I_2792 (I49294,I49286);
nand I_2793 (I49311,I49294,I49207);
nand I_2794 (I48960,I49294,I49116);
nor I_2795 (I49342,I33558,I33555);
and I_2796 (I49359,I49207,I49342);
nor I_2797 (I49376,I49294,I49359);
DFFARX1 I_2798 (I49376,I1803,I48983,I48969,);
nor I_2799 (I49407,I49009,I49342);
DFFARX1 I_2800 (I49407,I1803,I48983,I48954,);
nor I_2801 (I49438,I49286,I49342);
not I_2802 (I49455,I49438);
nand I_2803 (I48963,I49455,I49311);
not I_2804 (I49510,I1810);
DFFARX1 I_2805 (I57814,I1803,I49510,I49536,);
not I_2806 (I49544,I49536);
nand I_2807 (I49561,I57829,I57811);
and I_2808 (I49578,I49561,I57811);
DFFARX1 I_2809 (I49578,I1803,I49510,I49604,);
DFFARX1 I_2810 (I49604,I1803,I49510,I49499,);
DFFARX1 I_2811 (I57820,I1803,I49510,I49635,);
nand I_2812 (I49643,I49635,I57838);
not I_2813 (I49660,I49643);
DFFARX1 I_2814 (I49660,I1803,I49510,I49686,);
not I_2815 (I49694,I49686);
nor I_2816 (I49502,I49544,I49694);
DFFARX1 I_2817 (I57835,I1803,I49510,I49734,);
nor I_2818 (I49493,I49734,I49604);
nor I_2819 (I49484,I49734,I49660);
nand I_2820 (I49770,I57832,I57823);
and I_2821 (I49787,I49770,I57817);
DFFARX1 I_2822 (I49787,I1803,I49510,I49813,);
not I_2823 (I49821,I49813);
nand I_2824 (I49838,I49821,I49734);
nand I_2825 (I49487,I49821,I49643);
nor I_2826 (I49869,I57826,I57823);
and I_2827 (I49886,I49734,I49869);
nor I_2828 (I49903,I49821,I49886);
DFFARX1 I_2829 (I49903,I1803,I49510,I49496,);
nor I_2830 (I49934,I49536,I49869);
DFFARX1 I_2831 (I49934,I1803,I49510,I49481,);
nor I_2832 (I49965,I49813,I49869);
not I_2833 (I49982,I49965);
nand I_2834 (I49490,I49982,I49838);
not I_2835 (I50037,I1810);
DFFARX1 I_2836 (I25007,I1803,I50037,I50063,);
not I_2837 (I50071,I50063);
nand I_2838 (I50088,I25004,I25013);
and I_2839 (I50105,I50088,I25022);
DFFARX1 I_2840 (I50105,I1803,I50037,I50131,);
DFFARX1 I_2841 (I50131,I1803,I50037,I50026,);
DFFARX1 I_2842 (I25025,I1803,I50037,I50162,);
nand I_2843 (I50170,I50162,I25028);
not I_2844 (I50187,I50170);
DFFARX1 I_2845 (I50187,I1803,I50037,I50213,);
not I_2846 (I50221,I50213);
nor I_2847 (I50029,I50071,I50221);
DFFARX1 I_2848 (I25001,I1803,I50037,I50261,);
nor I_2849 (I50020,I50261,I50131);
nor I_2850 (I50011,I50261,I50187);
nand I_2851 (I50297,I25016,I25019);
and I_2852 (I50314,I50297,I25010);
DFFARX1 I_2853 (I50314,I1803,I50037,I50340,);
not I_2854 (I50348,I50340);
nand I_2855 (I50365,I50348,I50261);
nand I_2856 (I50014,I50348,I50170);
nor I_2857 (I50396,I25001,I25019);
and I_2858 (I50413,I50261,I50396);
nor I_2859 (I50430,I50348,I50413);
DFFARX1 I_2860 (I50430,I1803,I50037,I50023,);
nor I_2861 (I50461,I50063,I50396);
DFFARX1 I_2862 (I50461,I1803,I50037,I50008,);
nor I_2863 (I50492,I50340,I50396);
not I_2864 (I50509,I50492);
nand I_2865 (I50017,I50509,I50365);
not I_2866 (I50564,I1810);
DFFARX1 I_2867 (I29410,I1803,I50564,I50590,);
not I_2868 (I50598,I50590);
nand I_2869 (I50615,I29428,I29419);
and I_2870 (I50632,I50615,I29422);
DFFARX1 I_2871 (I50632,I1803,I50564,I50658,);
DFFARX1 I_2872 (I50658,I1803,I50564,I50553,);
DFFARX1 I_2873 (I29416,I1803,I50564,I50689,);
nand I_2874 (I50697,I50689,I29407);
not I_2875 (I50714,I50697);
DFFARX1 I_2876 (I50714,I1803,I50564,I50740,);
not I_2877 (I50748,I50740);
nor I_2878 (I50556,I50598,I50748);
DFFARX1 I_2879 (I29413,I1803,I50564,I50788,);
nor I_2880 (I50547,I50788,I50658);
nor I_2881 (I50538,I50788,I50714);
nand I_2882 (I50824,I29407,I29404);
and I_2883 (I50841,I50824,I29425);
DFFARX1 I_2884 (I50841,I1803,I50564,I50867,);
not I_2885 (I50875,I50867);
nand I_2886 (I50892,I50875,I50788);
nand I_2887 (I50541,I50875,I50697);
nor I_2888 (I50923,I29404,I29404);
and I_2889 (I50940,I50788,I50923);
nor I_2890 (I50957,I50875,I50940);
DFFARX1 I_2891 (I50957,I1803,I50564,I50550,);
nor I_2892 (I50988,I50590,I50923);
DFFARX1 I_2893 (I50988,I1803,I50564,I50535,);
nor I_2894 (I51019,I50867,I50923);
not I_2895 (I51036,I51019);
nand I_2896 (I50544,I51036,I50892);
not I_2897 (I51091,I1810);
DFFARX1 I_2898 (I31790,I1803,I51091,I51117,);
not I_2899 (I51125,I51117);
nand I_2900 (I51142,I31808,I31799);
and I_2901 (I51159,I51142,I31802);
DFFARX1 I_2902 (I51159,I1803,I51091,I51185,);
DFFARX1 I_2903 (I51185,I1803,I51091,I51080,);
DFFARX1 I_2904 (I31796,I1803,I51091,I51216,);
nand I_2905 (I51224,I51216,I31787);
not I_2906 (I51241,I51224);
DFFARX1 I_2907 (I51241,I1803,I51091,I51267,);
not I_2908 (I51275,I51267);
nor I_2909 (I51083,I51125,I51275);
DFFARX1 I_2910 (I31793,I1803,I51091,I51315,);
nor I_2911 (I51074,I51315,I51185);
nor I_2912 (I51065,I51315,I51241);
nand I_2913 (I51351,I31787,I31784);
and I_2914 (I51368,I51351,I31805);
DFFARX1 I_2915 (I51368,I1803,I51091,I51394,);
not I_2916 (I51402,I51394);
nand I_2917 (I51419,I51402,I51315);
nand I_2918 (I51068,I51402,I51224);
nor I_2919 (I51450,I31784,I31784);
and I_2920 (I51467,I51315,I51450);
nor I_2921 (I51484,I51402,I51467);
DFFARX1 I_2922 (I51484,I1803,I51091,I51077,);
nor I_2923 (I51515,I51117,I51450);
DFFARX1 I_2924 (I51515,I1803,I51091,I51062,);
nor I_2925 (I51546,I51394,I51450);
not I_2926 (I51563,I51546);
nand I_2927 (I51071,I51563,I51419);
not I_2928 (I51618,I1810);
DFFARX1 I_2929 (I72449,I1803,I51618,I51644,);
not I_2930 (I51652,I51644);
nand I_2931 (I51669,I72431,I72431);
and I_2932 (I51686,I51669,I72437);
DFFARX1 I_2933 (I51686,I1803,I51618,I51712,);
DFFARX1 I_2934 (I51712,I1803,I51618,I51607,);
DFFARX1 I_2935 (I72434,I1803,I51618,I51743,);
nand I_2936 (I51751,I51743,I72443);
not I_2937 (I51768,I51751);
DFFARX1 I_2938 (I51768,I1803,I51618,I51794,);
not I_2939 (I51802,I51794);
nor I_2940 (I51610,I51652,I51802);
DFFARX1 I_2941 (I72455,I1803,I51618,I51842,);
nor I_2942 (I51601,I51842,I51712);
nor I_2943 (I51592,I51842,I51768);
nand I_2944 (I51878,I72446,I72440);
and I_2945 (I51895,I51878,I72434);
DFFARX1 I_2946 (I51895,I1803,I51618,I51921,);
not I_2947 (I51929,I51921);
nand I_2948 (I51946,I51929,I51842);
nand I_2949 (I51595,I51929,I51751);
nor I_2950 (I51977,I72452,I72440);
and I_2951 (I51994,I51842,I51977);
nor I_2952 (I52011,I51929,I51994);
DFFARX1 I_2953 (I52011,I1803,I51618,I51604,);
nor I_2954 (I52042,I51644,I51977);
DFFARX1 I_2955 (I52042,I1803,I51618,I51589,);
nor I_2956 (I52073,I51921,I51977);
not I_2957 (I52090,I52073);
nand I_2958 (I51598,I52090,I51946);
not I_2959 (I52145,I1810);
DFFARX1 I_2960 (I45112,I1803,I52145,I52171,);
not I_2961 (I52179,I52171);
nand I_2962 (I52196,I45115,I45112);
and I_2963 (I52213,I52196,I45124);
DFFARX1 I_2964 (I52213,I1803,I52145,I52239,);
DFFARX1 I_2965 (I52239,I1803,I52145,I52134,);
DFFARX1 I_2966 (I45121,I1803,I52145,I52270,);
nand I_2967 (I52278,I52270,I45127);
not I_2968 (I52295,I52278);
DFFARX1 I_2969 (I52295,I1803,I52145,I52321,);
not I_2970 (I52329,I52321);
nor I_2971 (I52137,I52179,I52329);
DFFARX1 I_2972 (I45136,I1803,I52145,I52369,);
nor I_2973 (I52128,I52369,I52239);
nor I_2974 (I52119,I52369,I52295);
nand I_2975 (I52405,I45130,I45118);
and I_2976 (I52422,I52405,I45115);
DFFARX1 I_2977 (I52422,I1803,I52145,I52448,);
not I_2978 (I52456,I52448);
nand I_2979 (I52473,I52456,I52369);
nand I_2980 (I52122,I52456,I52278);
nor I_2981 (I52504,I45133,I45118);
and I_2982 (I52521,I52369,I52504);
nor I_2983 (I52538,I52456,I52521);
DFFARX1 I_2984 (I52538,I1803,I52145,I52131,);
nor I_2985 (I52569,I52171,I52504);
DFFARX1 I_2986 (I52569,I1803,I52145,I52116,);
nor I_2987 (I52600,I52448,I52504);
not I_2988 (I52617,I52600);
nand I_2989 (I52125,I52617,I52473);
not I_2990 (I52678,I1810);
DFFARX1 I_2991 (I50541,I1803,I52678,I52704,);
DFFARX1 I_2992 (I50538,I1803,I52678,I52721,);
not I_2993 (I52729,I52721);
not I_2994 (I52746,I50538);
nor I_2995 (I52763,I52746,I50541);
not I_2996 (I52780,I50553);
nor I_2997 (I52797,I52763,I50547);
nor I_2998 (I52814,I52721,I52797);
DFFARX1 I_2999 (I52814,I1803,I52678,I52664,);
nor I_3000 (I52845,I50547,I50541);
nand I_3001 (I52862,I52845,I50538);
DFFARX1 I_3002 (I52862,I1803,I52678,I52667,);
nor I_3003 (I52893,I52780,I50547);
nand I_3004 (I52910,I52893,I50535);
nor I_3005 (I52927,I52704,I52910);
DFFARX1 I_3006 (I52927,I1803,I52678,I52643,);
not I_3007 (I52958,I52910);
nand I_3008 (I52655,I52721,I52958);
DFFARX1 I_3009 (I52910,I1803,I52678,I52998,);
not I_3010 (I53006,I52998);
not I_3011 (I53023,I50547);
not I_3012 (I53040,I50544);
nor I_3013 (I53057,I53040,I50553);
nor I_3014 (I52670,I53006,I53057);
nor I_3015 (I53088,I53040,I50550);
and I_3016 (I53105,I53088,I50556);
or I_3017 (I53122,I53105,I50535);
DFFARX1 I_3018 (I53122,I1803,I52678,I53148,);
nor I_3019 (I52658,I53148,I52704);
not I_3020 (I53170,I53148);
and I_3021 (I53187,I53170,I52704);
nor I_3022 (I52652,I52729,I53187);
nand I_3023 (I53218,I53170,I52780);
nor I_3024 (I52646,I53040,I53218);
nand I_3025 (I52649,I53170,I52958);
nand I_3026 (I53263,I52780,I50544);
nor I_3027 (I52661,I53023,I53263);
not I_3028 (I53324,I1810);
DFFARX1 I_3029 (I81611,I1803,I53324,I53350,);
DFFARX1 I_3030 (I81635,I1803,I53324,I53367,);
not I_3031 (I53375,I53367);
not I_3032 (I53392,I81617);
nor I_3033 (I53409,I53392,I81626);
not I_3034 (I53426,I81611);
nor I_3035 (I53443,I53409,I81632);
nor I_3036 (I53460,I53367,I53443);
DFFARX1 I_3037 (I53460,I1803,I53324,I53310,);
nor I_3038 (I53491,I81632,I81626);
nand I_3039 (I53508,I53491,I81617);
DFFARX1 I_3040 (I53508,I1803,I53324,I53313,);
nor I_3041 (I53539,I53426,I81632);
nand I_3042 (I53556,I53539,I81629);
nor I_3043 (I53573,I53350,I53556);
DFFARX1 I_3044 (I53573,I1803,I53324,I53289,);
not I_3045 (I53604,I53556);
nand I_3046 (I53301,I53367,I53604);
DFFARX1 I_3047 (I53556,I1803,I53324,I53644,);
not I_3048 (I53652,I53644);
not I_3049 (I53669,I81632);
not I_3050 (I53686,I81623);
nor I_3051 (I53703,I53686,I81611);
nor I_3052 (I53316,I53652,I53703);
nor I_3053 (I53734,I53686,I81614);
and I_3054 (I53751,I53734,I81638);
or I_3055 (I53768,I53751,I81620);
DFFARX1 I_3056 (I53768,I1803,I53324,I53794,);
nor I_3057 (I53304,I53794,I53350);
not I_3058 (I53816,I53794);
and I_3059 (I53833,I53816,I53350);
nor I_3060 (I53298,I53375,I53833);
nand I_3061 (I53864,I53816,I53426);
nor I_3062 (I53292,I53686,I53864);
nand I_3063 (I53295,I53816,I53604);
nand I_3064 (I53909,I53426,I81623);
nor I_3065 (I53307,I53669,I53909);
not I_3066 (I53970,I1810);
DFFARX1 I_3067 (I15991,I1803,I53970,I53996,);
DFFARX1 I_3068 (I15997,I1803,I53970,I54013,);
not I_3069 (I54021,I54013);
not I_3070 (I54038,I16018);
nor I_3071 (I54055,I54038,I16006);
not I_3072 (I54072,I16015);
nor I_3073 (I54089,I54055,I16000);
nor I_3074 (I54106,I54013,I54089);
DFFARX1 I_3075 (I54106,I1803,I53970,I53956,);
nor I_3076 (I54137,I16000,I16006);
nand I_3077 (I54154,I54137,I16018);
DFFARX1 I_3078 (I54154,I1803,I53970,I53959,);
nor I_3079 (I54185,I54072,I16000);
nand I_3080 (I54202,I54185,I15991);
nor I_3081 (I54219,I53996,I54202);
DFFARX1 I_3082 (I54219,I1803,I53970,I53935,);
not I_3083 (I54250,I54202);
nand I_3084 (I53947,I54013,I54250);
DFFARX1 I_3085 (I54202,I1803,I53970,I54290,);
not I_3086 (I54298,I54290);
not I_3087 (I54315,I16000);
not I_3088 (I54332,I16003);
nor I_3089 (I54349,I54332,I16015);
nor I_3090 (I53962,I54298,I54349);
nor I_3091 (I54380,I54332,I16012);
and I_3092 (I54397,I54380,I15994);
or I_3093 (I54414,I54397,I16009);
DFFARX1 I_3094 (I54414,I1803,I53970,I54440,);
nor I_3095 (I53950,I54440,I53996);
not I_3096 (I54462,I54440);
and I_3097 (I54479,I54462,I53996);
nor I_3098 (I53944,I54021,I54479);
nand I_3099 (I54510,I54462,I54072);
nor I_3100 (I53938,I54332,I54510);
nand I_3101 (I53941,I54462,I54250);
nand I_3102 (I54555,I54072,I16003);
nor I_3103 (I53953,I54315,I54555);
not I_3104 (I54616,I1810);
DFFARX1 I_3105 (I78041,I1803,I54616,I54642,);
DFFARX1 I_3106 (I78065,I1803,I54616,I54659,);
not I_3107 (I54667,I54659);
not I_3108 (I54684,I78047);
nor I_3109 (I54701,I54684,I78056);
not I_3110 (I54718,I78041);
nor I_3111 (I54735,I54701,I78062);
nor I_3112 (I54752,I54659,I54735);
DFFARX1 I_3113 (I54752,I1803,I54616,I54602,);
nor I_3114 (I54783,I78062,I78056);
nand I_3115 (I54800,I54783,I78047);
DFFARX1 I_3116 (I54800,I1803,I54616,I54605,);
nor I_3117 (I54831,I54718,I78062);
nand I_3118 (I54848,I54831,I78059);
nor I_3119 (I54865,I54642,I54848);
DFFARX1 I_3120 (I54865,I1803,I54616,I54581,);
not I_3121 (I54896,I54848);
nand I_3122 (I54593,I54659,I54896);
DFFARX1 I_3123 (I54848,I1803,I54616,I54936,);
not I_3124 (I54944,I54936);
not I_3125 (I54961,I78062);
not I_3126 (I54978,I78053);
nor I_3127 (I54995,I54978,I78041);
nor I_3128 (I54608,I54944,I54995);
nor I_3129 (I55026,I54978,I78044);
and I_3130 (I55043,I55026,I78068);
or I_3131 (I55060,I55043,I78050);
DFFARX1 I_3132 (I55060,I1803,I54616,I55086,);
nor I_3133 (I54596,I55086,I54642);
not I_3134 (I55108,I55086);
and I_3135 (I55125,I55108,I54642);
nor I_3136 (I54590,I54667,I55125);
nand I_3137 (I55156,I55108,I54718);
nor I_3138 (I54584,I54978,I55156);
nand I_3139 (I54587,I55108,I54896);
nand I_3140 (I55201,I54718,I78053);
nor I_3141 (I54599,I54961,I55201);
not I_3142 (I55262,I1810);
DFFARX1 I_3143 (I66091,I1803,I55262,I55288,);
DFFARX1 I_3144 (I66073,I1803,I55262,I55305,);
not I_3145 (I55313,I55305);
not I_3146 (I55330,I66082);
nor I_3147 (I55347,I55330,I66094);
not I_3148 (I55364,I66076);
nor I_3149 (I55381,I55347,I66085);
nor I_3150 (I55398,I55305,I55381);
DFFARX1 I_3151 (I55398,I1803,I55262,I55248,);
nor I_3152 (I55429,I66085,I66094);
nand I_3153 (I55446,I55429,I66082);
DFFARX1 I_3154 (I55446,I1803,I55262,I55251,);
nor I_3155 (I55477,I55364,I66085);
nand I_3156 (I55494,I55477,I66097);
nor I_3157 (I55511,I55288,I55494);
DFFARX1 I_3158 (I55511,I1803,I55262,I55227,);
not I_3159 (I55542,I55494);
nand I_3160 (I55239,I55305,I55542);
DFFARX1 I_3161 (I55494,I1803,I55262,I55582,);
not I_3162 (I55590,I55582);
not I_3163 (I55607,I66085);
not I_3164 (I55624,I66073);
nor I_3165 (I55641,I55624,I66076);
nor I_3166 (I55254,I55590,I55641);
nor I_3167 (I55672,I55624,I66079);
and I_3168 (I55689,I55672,I66088);
or I_3169 (I55706,I55689,I66076);
DFFARX1 I_3170 (I55706,I1803,I55262,I55732,);
nor I_3171 (I55242,I55732,I55288);
not I_3172 (I55754,I55732);
and I_3173 (I55771,I55754,I55288);
nor I_3174 (I55236,I55313,I55771);
nand I_3175 (I55802,I55754,I55364);
nor I_3176 (I55230,I55624,I55802);
nand I_3177 (I55233,I55754,I55542);
nand I_3178 (I55847,I55364,I66073);
nor I_3179 (I55245,I55607,I55847);
not I_3180 (I55908,I1810);
DFFARX1 I_3181 (I80421,I1803,I55908,I55934,);
DFFARX1 I_3182 (I80445,I1803,I55908,I55951,);
not I_3183 (I55959,I55951);
not I_3184 (I55976,I80427);
nor I_3185 (I55993,I55976,I80436);
not I_3186 (I56010,I80421);
nor I_3187 (I56027,I55993,I80442);
nor I_3188 (I56044,I55951,I56027);
DFFARX1 I_3189 (I56044,I1803,I55908,I55894,);
nor I_3190 (I56075,I80442,I80436);
nand I_3191 (I56092,I56075,I80427);
DFFARX1 I_3192 (I56092,I1803,I55908,I55897,);
nor I_3193 (I56123,I56010,I80442);
nand I_3194 (I56140,I56123,I80439);
nor I_3195 (I56157,I55934,I56140);
DFFARX1 I_3196 (I56157,I1803,I55908,I55873,);
not I_3197 (I56188,I56140);
nand I_3198 (I55885,I55951,I56188);
DFFARX1 I_3199 (I56140,I1803,I55908,I56228,);
not I_3200 (I56236,I56228);
not I_3201 (I56253,I80442);
not I_3202 (I56270,I80433);
nor I_3203 (I56287,I56270,I80421);
nor I_3204 (I55900,I56236,I56287);
nor I_3205 (I56318,I56270,I80424);
and I_3206 (I56335,I56318,I80448);
or I_3207 (I56352,I56335,I80430);
DFFARX1 I_3208 (I56352,I1803,I55908,I56378,);
nor I_3209 (I55888,I56378,I55934);
not I_3210 (I56400,I56378);
and I_3211 (I56417,I56400,I55934);
nor I_3212 (I55882,I55959,I56417);
nand I_3213 (I56448,I56400,I56010);
nor I_3214 (I55876,I56270,I56448);
nand I_3215 (I55879,I56400,I56188);
nand I_3216 (I56493,I56010,I80433);
nor I_3217 (I55891,I56253,I56493);
not I_3218 (I56554,I1810);
DFFARX1 I_3219 (I13090,I1803,I56554,I56580,);
DFFARX1 I_3220 (I13102,I1803,I56554,I56597,);
not I_3221 (I56605,I56597);
not I_3222 (I56622,I13108);
nor I_3223 (I56639,I56622,I13093);
not I_3224 (I56656,I13084);
nor I_3225 (I56673,I56639,I13105);
nor I_3226 (I56690,I56597,I56673);
DFFARX1 I_3227 (I56690,I1803,I56554,I56540,);
nor I_3228 (I56721,I13105,I13093);
nand I_3229 (I56738,I56721,I13108);
DFFARX1 I_3230 (I56738,I1803,I56554,I56543,);
nor I_3231 (I56769,I56656,I13105);
nand I_3232 (I56786,I56769,I13087);
nor I_3233 (I56803,I56580,I56786);
DFFARX1 I_3234 (I56803,I1803,I56554,I56519,);
not I_3235 (I56834,I56786);
nand I_3236 (I56531,I56597,I56834);
DFFARX1 I_3237 (I56786,I1803,I56554,I56874,);
not I_3238 (I56882,I56874);
not I_3239 (I56899,I13105);
not I_3240 (I56916,I13096);
nor I_3241 (I56933,I56916,I13084);
nor I_3242 (I56546,I56882,I56933);
nor I_3243 (I56964,I56916,I13099);
and I_3244 (I56981,I56964,I13087);
or I_3245 (I56998,I56981,I13084);
DFFARX1 I_3246 (I56998,I1803,I56554,I57024,);
nor I_3247 (I56534,I57024,I56580);
not I_3248 (I57046,I57024);
and I_3249 (I57063,I57046,I56580);
nor I_3250 (I56528,I56605,I57063);
nand I_3251 (I57094,I57046,I56656);
nor I_3252 (I56522,I56916,I57094);
nand I_3253 (I56525,I57046,I56834);
nand I_3254 (I57139,I56656,I13096);
nor I_3255 (I56537,I56899,I57139);
not I_3256 (I57200,I1810);
DFFARX1 I_3257 (I3921,I1803,I57200,I57226,);
DFFARX1 I_3258 (I3927,I1803,I57200,I57243,);
not I_3259 (I57251,I57243);
not I_3260 (I57268,I3921);
nor I_3261 (I57285,I57268,I3933);
not I_3262 (I57302,I3945);
nor I_3263 (I57319,I57285,I3939);
nor I_3264 (I57336,I57243,I57319);
DFFARX1 I_3265 (I57336,I1803,I57200,I57186,);
nor I_3266 (I57367,I3939,I3933);
nand I_3267 (I57384,I57367,I3921);
DFFARX1 I_3268 (I57384,I1803,I57200,I57189,);
nor I_3269 (I57415,I57302,I3939);
nand I_3270 (I57432,I57415,I3924);
nor I_3271 (I57449,I57226,I57432);
DFFARX1 I_3272 (I57449,I1803,I57200,I57165,);
not I_3273 (I57480,I57432);
nand I_3274 (I57177,I57243,I57480);
DFFARX1 I_3275 (I57432,I1803,I57200,I57520,);
not I_3276 (I57528,I57520);
not I_3277 (I57545,I3939);
not I_3278 (I57562,I3924);
nor I_3279 (I57579,I57562,I3945);
nor I_3280 (I57192,I57528,I57579);
nor I_3281 (I57610,I57562,I3942);
and I_3282 (I57627,I57610,I3936);
or I_3283 (I57644,I57627,I3930);
DFFARX1 I_3284 (I57644,I1803,I57200,I57670,);
nor I_3285 (I57180,I57670,I57226);
not I_3286 (I57692,I57670);
and I_3287 (I57709,I57692,I57226);
nor I_3288 (I57174,I57251,I57709);
nand I_3289 (I57740,I57692,I57302);
nor I_3290 (I57168,I57562,I57740);
nand I_3291 (I57171,I57692,I57480);
nand I_3292 (I57785,I57302,I3924);
nor I_3293 (I57183,I57545,I57785);
not I_3294 (I57846,I1810);
DFFARX1 I_3295 (I45696,I1803,I57846,I57872,);
DFFARX1 I_3296 (I45690,I1803,I57846,I57889,);
not I_3297 (I57897,I57889);
not I_3298 (I57914,I45705);
nor I_3299 (I57931,I57914,I45690);
not I_3300 (I57948,I45699);
nor I_3301 (I57965,I57931,I45708);
nor I_3302 (I57982,I57889,I57965);
DFFARX1 I_3303 (I57982,I1803,I57846,I57832,);
nor I_3304 (I58013,I45708,I45690);
nand I_3305 (I58030,I58013,I45705);
DFFARX1 I_3306 (I58030,I1803,I57846,I57835,);
nor I_3307 (I58061,I57948,I45708);
nand I_3308 (I58078,I58061,I45693);
nor I_3309 (I58095,I57872,I58078);
DFFARX1 I_3310 (I58095,I1803,I57846,I57811,);
not I_3311 (I58126,I58078);
nand I_3312 (I57823,I57889,I58126);
DFFARX1 I_3313 (I58078,I1803,I57846,I58166,);
not I_3314 (I58174,I58166);
not I_3315 (I58191,I45708);
not I_3316 (I58208,I45702);
nor I_3317 (I58225,I58208,I45699);
nor I_3318 (I57838,I58174,I58225);
nor I_3319 (I58256,I58208,I45711);
and I_3320 (I58273,I58256,I45714);
or I_3321 (I58290,I58273,I45693);
DFFARX1 I_3322 (I58290,I1803,I57846,I58316,);
nor I_3323 (I57826,I58316,I57872);
not I_3324 (I58338,I58316);
and I_3325 (I58355,I58338,I57872);
nor I_3326 (I57820,I57897,I58355);
nand I_3327 (I58386,I58338,I57948);
nor I_3328 (I57814,I58208,I58386);
nand I_3329 (I57817,I58338,I58126);
nand I_3330 (I58431,I57948,I45702);
nor I_3331 (I57829,I58191,I58431);
not I_3332 (I58492,I1810);
DFFARX1 I_3333 (I7610,I1803,I58492,I58518,);
DFFARX1 I_3334 (I7616,I1803,I58492,I58535,);
not I_3335 (I58543,I58535);
not I_3336 (I58560,I7634);
nor I_3337 (I58577,I58560,I7613);
not I_3338 (I58594,I7619);
nor I_3339 (I58611,I58577,I7625);
nor I_3340 (I58628,I58535,I58611);
DFFARX1 I_3341 (I58628,I1803,I58492,I58478,);
nor I_3342 (I58659,I7625,I7613);
nand I_3343 (I58676,I58659,I7634);
DFFARX1 I_3344 (I58676,I1803,I58492,I58481,);
nor I_3345 (I58707,I58594,I7625);
nand I_3346 (I58724,I58707,I7631);
nor I_3347 (I58741,I58518,I58724);
DFFARX1 I_3348 (I58741,I1803,I58492,I58457,);
not I_3349 (I58772,I58724);
nand I_3350 (I58469,I58535,I58772);
DFFARX1 I_3351 (I58724,I1803,I58492,I58812,);
not I_3352 (I58820,I58812);
not I_3353 (I58837,I7625);
not I_3354 (I58854,I7613);
nor I_3355 (I58871,I58854,I7619);
nor I_3356 (I58484,I58820,I58871);
nor I_3357 (I58902,I58854,I7622);
and I_3358 (I58919,I58902,I7610);
or I_3359 (I58936,I58919,I7628);
DFFARX1 I_3360 (I58936,I1803,I58492,I58962,);
nor I_3361 (I58472,I58962,I58518);
not I_3362 (I58984,I58962);
and I_3363 (I59001,I58984,I58518);
nor I_3364 (I58466,I58543,I59001);
nand I_3365 (I59032,I58984,I58594);
nor I_3366 (I58460,I58854,I59032);
nand I_3367 (I58463,I58984,I58772);
nand I_3368 (I59077,I58594,I7613);
nor I_3369 (I58475,I58837,I59077);
not I_3370 (I59138,I1810);
DFFARX1 I_3371 (I8137,I1803,I59138,I59164,);
DFFARX1 I_3372 (I8143,I1803,I59138,I59181,);
not I_3373 (I59189,I59181);
not I_3374 (I59206,I8161);
nor I_3375 (I59223,I59206,I8140);
not I_3376 (I59240,I8146);
nor I_3377 (I59257,I59223,I8152);
nor I_3378 (I59274,I59181,I59257);
DFFARX1 I_3379 (I59274,I1803,I59138,I59124,);
nor I_3380 (I59305,I8152,I8140);
nand I_3381 (I59322,I59305,I8161);
DFFARX1 I_3382 (I59322,I1803,I59138,I59127,);
nor I_3383 (I59353,I59240,I8152);
nand I_3384 (I59370,I59353,I8158);
nor I_3385 (I59387,I59164,I59370);
DFFARX1 I_3386 (I59387,I1803,I59138,I59103,);
not I_3387 (I59418,I59370);
nand I_3388 (I59115,I59181,I59418);
DFFARX1 I_3389 (I59370,I1803,I59138,I59458,);
not I_3390 (I59466,I59458);
not I_3391 (I59483,I8152);
not I_3392 (I59500,I8140);
nor I_3393 (I59517,I59500,I8146);
nor I_3394 (I59130,I59466,I59517);
nor I_3395 (I59548,I59500,I8149);
and I_3396 (I59565,I59548,I8137);
or I_3397 (I59582,I59565,I8155);
DFFARX1 I_3398 (I59582,I1803,I59138,I59608,);
nor I_3399 (I59118,I59608,I59164);
not I_3400 (I59630,I59608);
and I_3401 (I59647,I59630,I59164);
nor I_3402 (I59112,I59189,I59647);
nand I_3403 (I59678,I59630,I59240);
nor I_3404 (I59106,I59500,I59678);
nand I_3405 (I59109,I59630,I59418);
nand I_3406 (I59723,I59240,I8140);
nor I_3407 (I59121,I59483,I59723);
not I_3408 (I59784,I1810);
DFFARX1 I_3409 (I49487,I1803,I59784,I59810,);
DFFARX1 I_3410 (I49484,I1803,I59784,I59827,);
not I_3411 (I59835,I59827);
not I_3412 (I59852,I49484);
nor I_3413 (I59869,I59852,I49487);
not I_3414 (I59886,I49499);
nor I_3415 (I59903,I59869,I49493);
nor I_3416 (I59920,I59827,I59903);
DFFARX1 I_3417 (I59920,I1803,I59784,I59770,);
nor I_3418 (I59951,I49493,I49487);
nand I_3419 (I59968,I59951,I49484);
DFFARX1 I_3420 (I59968,I1803,I59784,I59773,);
nor I_3421 (I59999,I59886,I49493);
nand I_3422 (I60016,I59999,I49481);
nor I_3423 (I60033,I59810,I60016);
DFFARX1 I_3424 (I60033,I1803,I59784,I59749,);
not I_3425 (I60064,I60016);
nand I_3426 (I59761,I59827,I60064);
DFFARX1 I_3427 (I60016,I1803,I59784,I60104,);
not I_3428 (I60112,I60104);
not I_3429 (I60129,I49493);
not I_3430 (I60146,I49490);
nor I_3431 (I60163,I60146,I49499);
nor I_3432 (I59776,I60112,I60163);
nor I_3433 (I60194,I60146,I49496);
and I_3434 (I60211,I60194,I49502);
or I_3435 (I60228,I60211,I49481);
DFFARX1 I_3436 (I60228,I1803,I59784,I60254,);
nor I_3437 (I59764,I60254,I59810);
not I_3438 (I60276,I60254);
and I_3439 (I60293,I60276,I59810);
nor I_3440 (I59758,I59835,I60293);
nand I_3441 (I60324,I60276,I59886);
nor I_3442 (I59752,I60146,I60324);
nand I_3443 (I59755,I60276,I60064);
nand I_3444 (I60369,I59886,I49490);
nor I_3445 (I59767,I60129,I60369);
not I_3446 (I60424,I1810);
DFFARX1 I_3447 (I42803,I1803,I60424,I60450,);
DFFARX1 I_3448 (I60450,I1803,I60424,I60467,);
not I_3449 (I60416,I60467);
not I_3450 (I60489,I60450);
DFFARX1 I_3451 (I42815,I1803,I60424,I60515,);
nand I_3452 (I60523,I60515,I42824);
not I_3453 (I60540,I42824);
not I_3454 (I60557,I42806);
nand I_3455 (I60574,I42809,I42800);
and I_3456 (I60591,I42809,I42800);
not I_3457 (I60608,I42818);
nand I_3458 (I60625,I60608,I60557);
nor I_3459 (I60398,I60625,I60523);
nor I_3460 (I60656,I60540,I60625);
nand I_3461 (I60401,I60591,I60656);
not I_3462 (I60687,I42821);
nor I_3463 (I60704,I60687,I42809);
nor I_3464 (I60721,I60704,I42818);
nor I_3465 (I60738,I60489,I60721);
DFFARX1 I_3466 (I60738,I1803,I60424,I60410,);
not I_3467 (I60769,I60704);
DFFARX1 I_3468 (I60769,I1803,I60424,I60413,);
and I_3469 (I60407,I60515,I60704);
nor I_3470 (I60814,I60687,I42800);
and I_3471 (I60831,I60814,I42812);
or I_3472 (I60848,I60831,I42803);
DFFARX1 I_3473 (I60848,I1803,I60424,I60874,);
nor I_3474 (I60882,I60874,I60608);
DFFARX1 I_3475 (I60882,I1803,I60424,I60395,);
nand I_3476 (I60913,I60874,I60515);
nand I_3477 (I60930,I60608,I60913);
nor I_3478 (I60404,I60930,I60574);
not I_3479 (I60985,I1810);
DFFARX1 I_3480 (I67822,I1803,I60985,I61011,);
DFFARX1 I_3481 (I61011,I1803,I60985,I61028,);
not I_3482 (I60977,I61028);
not I_3483 (I61050,I61011);
DFFARX1 I_3484 (I67813,I1803,I60985,I61076,);
nand I_3485 (I61084,I61076,I67810);
not I_3486 (I61101,I67810);
not I_3487 (I61118,I67819);
nand I_3488 (I61135,I67828,I67810);
and I_3489 (I61152,I67828,I67810);
not I_3490 (I61169,I67807);
nand I_3491 (I61186,I61169,I61118);
nor I_3492 (I60959,I61186,I61084);
nor I_3493 (I61217,I61101,I61186);
nand I_3494 (I60962,I61152,I61217);
not I_3495 (I61248,I67816);
nor I_3496 (I61265,I61248,I67828);
nor I_3497 (I61282,I61265,I67807);
nor I_3498 (I61299,I61050,I61282);
DFFARX1 I_3499 (I61299,I1803,I60985,I60971,);
not I_3500 (I61330,I61265);
DFFARX1 I_3501 (I61330,I1803,I60985,I60974,);
and I_3502 (I60968,I61076,I61265);
nor I_3503 (I61375,I61248,I67831);
and I_3504 (I61392,I61375,I67807);
or I_3505 (I61409,I61392,I67825);
DFFARX1 I_3506 (I61409,I1803,I60985,I61435,);
nor I_3507 (I61443,I61435,I61169);
DFFARX1 I_3508 (I61443,I1803,I60985,I60956,);
nand I_3509 (I61474,I61435,I61076);
nand I_3510 (I61491,I61169,I61474);
nor I_3511 (I60965,I61491,I61135);
not I_3512 (I61546,I1810);
DFFARX1 I_3513 (I37020,I1803,I61546,I61572,);
DFFARX1 I_3514 (I61572,I1803,I61546,I61589,);
not I_3515 (I61538,I61589);
not I_3516 (I61611,I61572);
DFFARX1 I_3517 (I37035,I1803,I61546,I61637,);
nand I_3518 (I61645,I61637,I37026);
not I_3519 (I61662,I37026);
not I_3520 (I61679,I37032);
nand I_3521 (I61696,I37029,I37038);
and I_3522 (I61713,I37029,I37038);
not I_3523 (I61730,I37023);
nand I_3524 (I61747,I61730,I61679);
nor I_3525 (I61520,I61747,I61645);
nor I_3526 (I61778,I61662,I61747);
nand I_3527 (I61523,I61713,I61778);
not I_3528 (I61809,I37020);
nor I_3529 (I61826,I61809,I37029);
nor I_3530 (I61843,I61826,I37023);
nor I_3531 (I61860,I61611,I61843);
DFFARX1 I_3532 (I61860,I1803,I61546,I61532,);
not I_3533 (I61891,I61826);
DFFARX1 I_3534 (I61891,I1803,I61546,I61535,);
and I_3535 (I61529,I61637,I61826);
nor I_3536 (I61936,I61809,I37044);
and I_3537 (I61953,I61936,I37023);
or I_3538 (I61970,I61953,I37041);
DFFARX1 I_3539 (I61970,I1803,I61546,I61996,);
nor I_3540 (I62004,I61996,I61730);
DFFARX1 I_3541 (I62004,I1803,I61546,I61517,);
nand I_3542 (I62035,I61996,I61637);
nand I_3543 (I62052,I61730,I62035);
nor I_3544 (I61526,I62052,I61696);
not I_3545 (I62107,I1810);
DFFARX1 I_3546 (I35286,I1803,I62107,I62133,);
DFFARX1 I_3547 (I62133,I1803,I62107,I62150,);
not I_3548 (I62099,I62150);
not I_3549 (I62172,I62133);
DFFARX1 I_3550 (I35301,I1803,I62107,I62198,);
nand I_3551 (I62206,I62198,I35292);
not I_3552 (I62223,I35292);
not I_3553 (I62240,I35298);
nand I_3554 (I62257,I35295,I35304);
and I_3555 (I62274,I35295,I35304);
not I_3556 (I62291,I35289);
nand I_3557 (I62308,I62291,I62240);
nor I_3558 (I62081,I62308,I62206);
nor I_3559 (I62339,I62223,I62308);
nand I_3560 (I62084,I62274,I62339);
not I_3561 (I62370,I35286);
nor I_3562 (I62387,I62370,I35295);
nor I_3563 (I62404,I62387,I35289);
nor I_3564 (I62421,I62172,I62404);
DFFARX1 I_3565 (I62421,I1803,I62107,I62093,);
not I_3566 (I62452,I62387);
DFFARX1 I_3567 (I62452,I1803,I62107,I62096,);
and I_3568 (I62090,I62198,I62387);
nor I_3569 (I62497,I62370,I35310);
and I_3570 (I62514,I62497,I35289);
or I_3571 (I62531,I62514,I35307);
DFFARX1 I_3572 (I62531,I1803,I62107,I62557,);
nor I_3573 (I62565,I62557,I62291);
DFFARX1 I_3574 (I62565,I1803,I62107,I62078,);
nand I_3575 (I62596,I62557,I62198);
nand I_3576 (I62613,I62291,I62596);
nor I_3577 (I62087,I62613,I62257);
not I_3578 (I62668,I1810);
DFFARX1 I_3579 (I73559,I1803,I62668,I62694,);
DFFARX1 I_3580 (I62694,I1803,I62668,I62711,);
not I_3581 (I62660,I62711);
not I_3582 (I62733,I62694);
DFFARX1 I_3583 (I73565,I1803,I62668,I62759,);
nand I_3584 (I62767,I62759,I73574);
not I_3585 (I62784,I73574);
not I_3586 (I62801,I73553);
nand I_3587 (I62818,I73556,I73556);
and I_3588 (I62835,I73556,I73556);
not I_3589 (I62852,I73568);
nand I_3590 (I62869,I62852,I62801);
nor I_3591 (I62642,I62869,I62767);
nor I_3592 (I62900,I62784,I62869);
nand I_3593 (I62645,I62835,I62900);
not I_3594 (I62931,I73562);
nor I_3595 (I62948,I62931,I73556);
nor I_3596 (I62965,I62948,I73568);
nor I_3597 (I62982,I62733,I62965);
DFFARX1 I_3598 (I62982,I1803,I62668,I62654,);
not I_3599 (I63013,I62948);
DFFARX1 I_3600 (I63013,I1803,I62668,I62657,);
and I_3601 (I62651,I62759,I62948);
nor I_3602 (I63058,I62931,I73577);
and I_3603 (I63075,I63058,I73553);
or I_3604 (I63092,I63075,I73571);
DFFARX1 I_3605 (I63092,I1803,I62668,I63118,);
nor I_3606 (I63126,I63118,I62852);
DFFARX1 I_3607 (I63126,I1803,I62668,I62639,);
nand I_3608 (I63157,I63118,I62759);
nand I_3609 (I63174,I62852,I63157);
nor I_3610 (I62648,I63174,I62818);
not I_3611 (I63229,I1810);
DFFARX1 I_3612 (I51071,I1803,I63229,I63255,);
DFFARX1 I_3613 (I63255,I1803,I63229,I63272,);
not I_3614 (I63221,I63272);
not I_3615 (I63294,I63255);
DFFARX1 I_3616 (I51068,I1803,I63229,I63320,);
nand I_3617 (I63328,I63320,I51083);
not I_3618 (I63345,I51083);
not I_3619 (I63362,I51080);
nand I_3620 (I63379,I51077,I51065);
and I_3621 (I63396,I51077,I51065);
not I_3622 (I63413,I51062);
nand I_3623 (I63430,I63413,I63362);
nor I_3624 (I63203,I63430,I63328);
nor I_3625 (I63461,I63345,I63430);
nand I_3626 (I63206,I63396,I63461);
not I_3627 (I63492,I51068);
nor I_3628 (I63509,I63492,I51077);
nor I_3629 (I63526,I63509,I51062);
nor I_3630 (I63543,I63294,I63526);
DFFARX1 I_3631 (I63543,I1803,I63229,I63215,);
not I_3632 (I63574,I63509);
DFFARX1 I_3633 (I63574,I1803,I63229,I63218,);
and I_3634 (I63212,I63320,I63509);
nor I_3635 (I63619,I63492,I51074);
and I_3636 (I63636,I63619,I51062);
or I_3637 (I63653,I63636,I51065);
DFFARX1 I_3638 (I63653,I1803,I63229,I63679,);
nor I_3639 (I63687,I63679,I63413);
DFFARX1 I_3640 (I63687,I1803,I63229,I63200,);
nand I_3641 (I63718,I63679,I63320);
nand I_3642 (I63735,I63413,I63718);
nor I_3643 (I63209,I63735,I63379);
not I_3644 (I63793,I1810);
DFFARX1 I_3645 (I27721,I1803,I63793,I63819,);
and I_3646 (I63827,I63819,I27736);
DFFARX1 I_3647 (I63827,I1803,I63793,I63776,);
DFFARX1 I_3648 (I27739,I1803,I63793,I63867,);
not I_3649 (I63875,I27733);
not I_3650 (I63892,I27748);
nand I_3651 (I63909,I63892,I63875);
nor I_3652 (I63764,I63867,I63909);
DFFARX1 I_3653 (I63909,I1803,I63793,I63949,);
not I_3654 (I63785,I63949);
not I_3655 (I63971,I27724);
nand I_3656 (I63988,I63892,I63971);
DFFARX1 I_3657 (I63988,I1803,I63793,I64014,);
not I_3658 (I64022,I64014);
not I_3659 (I64039,I27727);
nand I_3660 (I64056,I64039,I27721);
and I_3661 (I64073,I63875,I64056);
nor I_3662 (I64090,I63988,I64073);
DFFARX1 I_3663 (I64090,I1803,I63793,I63761,);
DFFARX1 I_3664 (I64073,I1803,I63793,I63782,);
nor I_3665 (I64135,I27727,I27730);
nor I_3666 (I63773,I63988,I64135);
or I_3667 (I64166,I27727,I27730);
nor I_3668 (I64183,I27745,I27742);
DFFARX1 I_3669 (I64183,I1803,I63793,I64209,);
not I_3670 (I64217,I64209);
nor I_3671 (I63779,I64217,I64022);
nand I_3672 (I64248,I64217,I63867);
not I_3673 (I64265,I27745);
nand I_3674 (I64282,I64265,I63971);
nand I_3675 (I64299,I64217,I64282);
nand I_3676 (I63770,I64299,I64248);
nand I_3677 (I63767,I64282,I64166);
not I_3678 (I64371,I1810);
DFFARX1 I_3679 (I5526,I1803,I64371,I64397,);
and I_3680 (I64405,I64397,I5502);
DFFARX1 I_3681 (I64405,I1803,I64371,I64354,);
DFFARX1 I_3682 (I5520,I1803,I64371,I64445,);
not I_3683 (I64453,I5508);
not I_3684 (I64470,I5505);
nand I_3685 (I64487,I64470,I64453);
nor I_3686 (I64342,I64445,I64487);
DFFARX1 I_3687 (I64487,I1803,I64371,I64527,);
not I_3688 (I64363,I64527);
not I_3689 (I64549,I5514);
nand I_3690 (I64566,I64470,I64549);
DFFARX1 I_3691 (I64566,I1803,I64371,I64592,);
not I_3692 (I64600,I64592);
not I_3693 (I64617,I5505);
nand I_3694 (I64634,I64617,I5523);
and I_3695 (I64651,I64453,I64634);
nor I_3696 (I64668,I64566,I64651);
DFFARX1 I_3697 (I64668,I1803,I64371,I64339,);
DFFARX1 I_3698 (I64651,I1803,I64371,I64360,);
nor I_3699 (I64713,I5505,I5517);
nor I_3700 (I64351,I64566,I64713);
or I_3701 (I64744,I5505,I5517);
nor I_3702 (I64761,I5511,I5502);
DFFARX1 I_3703 (I64761,I1803,I64371,I64787,);
not I_3704 (I64795,I64787);
nor I_3705 (I64357,I64795,I64600);
nand I_3706 (I64826,I64795,I64445);
not I_3707 (I64843,I5511);
nand I_3708 (I64860,I64843,I64549);
nand I_3709 (I64877,I64795,I64860);
nand I_3710 (I64348,I64877,I64826);
nand I_3711 (I64345,I64860,I64744);
not I_3712 (I64949,I1810);
DFFARX1 I_3713 (I20761,I1803,I64949,I64975,);
and I_3714 (I64983,I64975,I20746);
DFFARX1 I_3715 (I64983,I1803,I64949,I64932,);
DFFARX1 I_3716 (I20752,I1803,I64949,I65023,);
not I_3717 (I65031,I20734);
not I_3718 (I65048,I20755);
nand I_3719 (I65065,I65048,I65031);
nor I_3720 (I64920,I65023,I65065);
DFFARX1 I_3721 (I65065,I1803,I64949,I65105,);
not I_3722 (I64941,I65105);
not I_3723 (I65127,I20758);
nand I_3724 (I65144,I65048,I65127);
DFFARX1 I_3725 (I65144,I1803,I64949,I65170,);
not I_3726 (I65178,I65170);
not I_3727 (I65195,I20749);
nand I_3728 (I65212,I65195,I20737);
and I_3729 (I65229,I65031,I65212);
nor I_3730 (I65246,I65144,I65229);
DFFARX1 I_3731 (I65246,I1803,I64949,I64917,);
DFFARX1 I_3732 (I65229,I1803,I64949,I64938,);
nor I_3733 (I65291,I20749,I20743);
nor I_3734 (I64929,I65144,I65291);
or I_3735 (I65322,I20749,I20743);
nor I_3736 (I65339,I20740,I20734);
DFFARX1 I_3737 (I65339,I1803,I64949,I65365,);
not I_3738 (I65373,I65365);
nor I_3739 (I64935,I65373,I65178);
nand I_3740 (I65404,I65373,I65023);
not I_3741 (I65421,I20740);
nand I_3742 (I65438,I65421,I65127);
nand I_3743 (I65455,I65373,I65438);
nand I_3744 (I64926,I65455,I65404);
nand I_3745 (I64923,I65438,I65322);
not I_3746 (I65527,I1810);
DFFARX1 I_3747 (I2340,I1803,I65527,I65553,);
and I_3748 (I65561,I65553,I2343);
DFFARX1 I_3749 (I65561,I1803,I65527,I65510,);
DFFARX1 I_3750 (I2343,I1803,I65527,I65601,);
not I_3751 (I65609,I2346);
not I_3752 (I65626,I2361);
nand I_3753 (I65643,I65626,I65609);
nor I_3754 (I65498,I65601,I65643);
DFFARX1 I_3755 (I65643,I1803,I65527,I65683,);
not I_3756 (I65519,I65683);
not I_3757 (I65705,I2355);
nand I_3758 (I65722,I65626,I65705);
DFFARX1 I_3759 (I65722,I1803,I65527,I65748,);
not I_3760 (I65756,I65748);
not I_3761 (I65773,I2358);
nand I_3762 (I65790,I65773,I2340);
and I_3763 (I65807,I65609,I65790);
nor I_3764 (I65824,I65722,I65807);
DFFARX1 I_3765 (I65824,I1803,I65527,I65495,);
DFFARX1 I_3766 (I65807,I1803,I65527,I65516,);
nor I_3767 (I65869,I2358,I2352);
nor I_3768 (I65507,I65722,I65869);
or I_3769 (I65900,I2358,I2352);
nor I_3770 (I65917,I2349,I2364);
DFFARX1 I_3771 (I65917,I1803,I65527,I65943,);
not I_3772 (I65951,I65943);
nor I_3773 (I65513,I65951,I65756);
nand I_3774 (I65982,I65951,I65601);
not I_3775 (I65999,I2349);
nand I_3776 (I66016,I65999,I65705);
nand I_3777 (I66033,I65951,I66016);
nand I_3778 (I65504,I66033,I65982);
nand I_3779 (I65501,I66016,I65900);
not I_3780 (I66105,I1810);
DFFARX1 I_3781 (I21815,I1803,I66105,I66131,);
and I_3782 (I66139,I66131,I21800);
DFFARX1 I_3783 (I66139,I1803,I66105,I66088,);
DFFARX1 I_3784 (I21806,I1803,I66105,I66179,);
not I_3785 (I66187,I21788);
not I_3786 (I66204,I21809);
nand I_3787 (I66221,I66204,I66187);
nor I_3788 (I66076,I66179,I66221);
DFFARX1 I_3789 (I66221,I1803,I66105,I66261,);
not I_3790 (I66097,I66261);
not I_3791 (I66283,I21812);
nand I_3792 (I66300,I66204,I66283);
DFFARX1 I_3793 (I66300,I1803,I66105,I66326,);
not I_3794 (I66334,I66326);
not I_3795 (I66351,I21803);
nand I_3796 (I66368,I66351,I21791);
and I_3797 (I66385,I66187,I66368);
nor I_3798 (I66402,I66300,I66385);
DFFARX1 I_3799 (I66402,I1803,I66105,I66073,);
DFFARX1 I_3800 (I66385,I1803,I66105,I66094,);
nor I_3801 (I66447,I21803,I21797);
nor I_3802 (I66085,I66300,I66447);
or I_3803 (I66478,I21803,I21797);
nor I_3804 (I66495,I21794,I21788);
DFFARX1 I_3805 (I66495,I1803,I66105,I66521,);
not I_3806 (I66529,I66521);
nor I_3807 (I66091,I66529,I66334);
nand I_3808 (I66560,I66529,I66179);
not I_3809 (I66577,I21794);
nand I_3810 (I66594,I66577,I66283);
nand I_3811 (I66611,I66529,I66594);
nand I_3812 (I66082,I66611,I66560);
nand I_3813 (I66079,I66594,I66478);
not I_3814 (I66683,I1810);
DFFARX1 I_3815 (I20234,I1803,I66683,I66709,);
and I_3816 (I66717,I66709,I20219);
DFFARX1 I_3817 (I66717,I1803,I66683,I66666,);
DFFARX1 I_3818 (I20225,I1803,I66683,I66757,);
not I_3819 (I66765,I20207);
not I_3820 (I66782,I20228);
nand I_3821 (I66799,I66782,I66765);
nor I_3822 (I66654,I66757,I66799);
DFFARX1 I_3823 (I66799,I1803,I66683,I66839,);
not I_3824 (I66675,I66839);
not I_3825 (I66861,I20231);
nand I_3826 (I66878,I66782,I66861);
DFFARX1 I_3827 (I66878,I1803,I66683,I66904,);
not I_3828 (I66912,I66904);
not I_3829 (I66929,I20222);
nand I_3830 (I66946,I66929,I20210);
and I_3831 (I66963,I66765,I66946);
nor I_3832 (I66980,I66878,I66963);
DFFARX1 I_3833 (I66980,I1803,I66683,I66651,);
DFFARX1 I_3834 (I66963,I1803,I66683,I66672,);
nor I_3835 (I67025,I20222,I20216);
nor I_3836 (I66663,I66878,I67025);
or I_3837 (I67056,I20222,I20216);
nor I_3838 (I67073,I20213,I20207);
DFFARX1 I_3839 (I67073,I1803,I66683,I67099,);
not I_3840 (I67107,I67099);
nor I_3841 (I66669,I67107,I66912);
nand I_3842 (I67138,I67107,I66757);
not I_3843 (I67155,I20213);
nand I_3844 (I67172,I67155,I66861);
nand I_3845 (I67189,I67107,I67172);
nand I_3846 (I66660,I67189,I67138);
nand I_3847 (I66657,I67172,I67056);
not I_3848 (I67261,I1810);
DFFARX1 I_3849 (I62642,I1803,I67261,I67287,);
and I_3850 (I67295,I67287,I62639);
DFFARX1 I_3851 (I67295,I1803,I67261,I67244,);
DFFARX1 I_3852 (I62645,I1803,I67261,I67335,);
not I_3853 (I67343,I62648);
not I_3854 (I67360,I62642);
nand I_3855 (I67377,I67360,I67343);
nor I_3856 (I67232,I67335,I67377);
DFFARX1 I_3857 (I67377,I1803,I67261,I67417,);
not I_3858 (I67253,I67417);
not I_3859 (I67439,I62657);
nand I_3860 (I67456,I67360,I67439);
DFFARX1 I_3861 (I67456,I1803,I67261,I67482,);
not I_3862 (I67490,I67482);
not I_3863 (I67507,I62654);
nand I_3864 (I67524,I67507,I62660);
and I_3865 (I67541,I67343,I67524);
nor I_3866 (I67558,I67456,I67541);
DFFARX1 I_3867 (I67558,I1803,I67261,I67229,);
DFFARX1 I_3868 (I67541,I1803,I67261,I67250,);
nor I_3869 (I67603,I62654,I62639);
nor I_3870 (I67241,I67456,I67603);
or I_3871 (I67634,I62654,I62639);
nor I_3872 (I67651,I62651,I62645);
DFFARX1 I_3873 (I67651,I1803,I67261,I67677,);
not I_3874 (I67685,I67677);
nor I_3875 (I67247,I67685,I67490);
nand I_3876 (I67716,I67685,I67335);
not I_3877 (I67733,I62651);
nand I_3878 (I67750,I67733,I67439);
nand I_3879 (I67767,I67685,I67750);
nand I_3880 (I67238,I67767,I67716);
nand I_3881 (I67235,I67750,I67634);
not I_3882 (I67839,I1810);
DFFARX1 I_3883 (I3394,I1803,I67839,I67865,);
and I_3884 (I67873,I67865,I3397);
DFFARX1 I_3885 (I67873,I1803,I67839,I67822,);
DFFARX1 I_3886 (I3397,I1803,I67839,I67913,);
not I_3887 (I67921,I3400);
not I_3888 (I67938,I3415);
nand I_3889 (I67955,I67938,I67921);
nor I_3890 (I67810,I67913,I67955);
DFFARX1 I_3891 (I67955,I1803,I67839,I67995,);
not I_3892 (I67831,I67995);
not I_3893 (I68017,I3409);
nand I_3894 (I68034,I67938,I68017);
DFFARX1 I_3895 (I68034,I1803,I67839,I68060,);
not I_3896 (I68068,I68060);
not I_3897 (I68085,I3412);
nand I_3898 (I68102,I68085,I3394);
and I_3899 (I68119,I67921,I68102);
nor I_3900 (I68136,I68034,I68119);
DFFARX1 I_3901 (I68136,I1803,I67839,I67807,);
DFFARX1 I_3902 (I68119,I1803,I67839,I67828,);
nor I_3903 (I68181,I3412,I3406);
nor I_3904 (I67819,I68034,I68181);
or I_3905 (I68212,I3412,I3406);
nor I_3906 (I68229,I3403,I3418);
DFFARX1 I_3907 (I68229,I1803,I67839,I68255,);
not I_3908 (I68263,I68255);
nor I_3909 (I67825,I68263,I68068);
nand I_3910 (I68294,I68263,I67913);
not I_3911 (I68311,I3403);
nand I_3912 (I68328,I68311,I68017);
nand I_3913 (I68345,I68263,I68328);
nand I_3914 (I67816,I68345,I68294);
nand I_3915 (I67813,I68328,I68212);
not I_3916 (I68417,I1810);
DFFARX1 I_3917 (I83423,I1803,I68417,I68443,);
and I_3918 (I68451,I68443,I83405);
DFFARX1 I_3919 (I68451,I1803,I68417,I68400,);
DFFARX1 I_3920 (I83396,I1803,I68417,I68491,);
not I_3921 (I68499,I83411);
not I_3922 (I68516,I83399);
nand I_3923 (I68533,I68516,I68499);
nor I_3924 (I68388,I68491,I68533);
DFFARX1 I_3925 (I68533,I1803,I68417,I68573,);
not I_3926 (I68409,I68573);
not I_3927 (I68595,I83408);
nand I_3928 (I68612,I68516,I68595);
DFFARX1 I_3929 (I68612,I1803,I68417,I68638,);
not I_3930 (I68646,I68638);
not I_3931 (I68663,I83417);
nand I_3932 (I68680,I68663,I83396);
and I_3933 (I68697,I68499,I68680);
nor I_3934 (I68714,I68612,I68697);
DFFARX1 I_3935 (I68714,I1803,I68417,I68385,);
DFFARX1 I_3936 (I68697,I1803,I68417,I68406,);
nor I_3937 (I68759,I83417,I83420);
nor I_3938 (I68397,I68612,I68759);
or I_3939 (I68790,I83417,I83420);
nor I_3940 (I68807,I83414,I83402);
DFFARX1 I_3941 (I68807,I1803,I68417,I68833,);
not I_3942 (I68841,I68833);
nor I_3943 (I68403,I68841,I68646);
nand I_3944 (I68872,I68841,I68491);
not I_3945 (I68889,I83414);
nand I_3946 (I68906,I68889,I68595);
nand I_3947 (I68923,I68841,I68906);
nand I_3948 (I68394,I68923,I68872);
nand I_3949 (I68391,I68906,I68790);
not I_3950 (I68995,I1810);
DFFARX1 I_3951 (I78663,I1803,I68995,I69021,);
and I_3952 (I69029,I69021,I78645);
DFFARX1 I_3953 (I69029,I1803,I68995,I68978,);
DFFARX1 I_3954 (I78636,I1803,I68995,I69069,);
not I_3955 (I69077,I78651);
not I_3956 (I69094,I78639);
nand I_3957 (I69111,I69094,I69077);
nor I_3958 (I68966,I69069,I69111);
DFFARX1 I_3959 (I69111,I1803,I68995,I69151,);
not I_3960 (I68987,I69151);
not I_3961 (I69173,I78648);
nand I_3962 (I69190,I69094,I69173);
DFFARX1 I_3963 (I69190,I1803,I68995,I69216,);
not I_3964 (I69224,I69216);
not I_3965 (I69241,I78657);
nand I_3966 (I69258,I69241,I78636);
and I_3967 (I69275,I69077,I69258);
nor I_3968 (I69292,I69190,I69275);
DFFARX1 I_3969 (I69292,I1803,I68995,I68963,);
DFFARX1 I_3970 (I69275,I1803,I68995,I68984,);
nor I_3971 (I69337,I78657,I78660);
nor I_3972 (I68975,I69190,I69337);
or I_3973 (I69368,I78657,I78660);
nor I_3974 (I69385,I78654,I78642);
DFFARX1 I_3975 (I69385,I1803,I68995,I69411,);
not I_3976 (I69419,I69411);
nor I_3977 (I68981,I69419,I69224);
nand I_3978 (I69450,I69419,I69069);
not I_3979 (I69467,I78654);
nand I_3980 (I69484,I69467,I69173);
nand I_3981 (I69501,I69419,I69484);
nand I_3982 (I68972,I69501,I69450);
nand I_3983 (I68969,I69484,I69368);
not I_3984 (I69573,I1810);
DFFARX1 I_3985 (I36457,I1803,I69573,I69599,);
and I_3986 (I69607,I69599,I36445);
DFFARX1 I_3987 (I69607,I1803,I69573,I69556,);
DFFARX1 I_3988 (I36460,I1803,I69573,I69647,);
not I_3989 (I69655,I36451);
not I_3990 (I69672,I36442);
nand I_3991 (I69689,I69672,I69655);
nor I_3992 (I69544,I69647,I69689);
DFFARX1 I_3993 (I69689,I1803,I69573,I69729,);
not I_3994 (I69565,I69729);
not I_3995 (I69751,I36448);
nand I_3996 (I69768,I69672,I69751);
DFFARX1 I_3997 (I69768,I1803,I69573,I69794,);
not I_3998 (I69802,I69794);
not I_3999 (I69819,I36463);
nand I_4000 (I69836,I69819,I36466);
and I_4001 (I69853,I69655,I69836);
nor I_4002 (I69870,I69768,I69853);
DFFARX1 I_4003 (I69870,I1803,I69573,I69541,);
DFFARX1 I_4004 (I69853,I1803,I69573,I69562,);
nor I_4005 (I69915,I36463,I36442);
nor I_4006 (I69553,I69768,I69915);
or I_4007 (I69946,I36463,I36442);
nor I_4008 (I69963,I36454,I36445);
DFFARX1 I_4009 (I69963,I1803,I69573,I69989,);
not I_4010 (I69997,I69989);
nor I_4011 (I69559,I69997,I69802);
nand I_4012 (I70028,I69997,I69647);
not I_4013 (I70045,I36454);
nand I_4014 (I70062,I70045,I69751);
nand I_4015 (I70079,I69997,I70062);
nand I_4016 (I69550,I70079,I70028);
nand I_4017 (I69547,I70062,I69946);
not I_4018 (I70151,I1810);
DFFARX1 I_4019 (I22869,I1803,I70151,I70177,);
and I_4020 (I70185,I70177,I22854);
DFFARX1 I_4021 (I70185,I1803,I70151,I70134,);
DFFARX1 I_4022 (I22860,I1803,I70151,I70225,);
not I_4023 (I70233,I22842);
not I_4024 (I70250,I22863);
nand I_4025 (I70267,I70250,I70233);
nor I_4026 (I70122,I70225,I70267);
DFFARX1 I_4027 (I70267,I1803,I70151,I70307,);
not I_4028 (I70143,I70307);
not I_4029 (I70329,I22866);
nand I_4030 (I70346,I70250,I70329);
DFFARX1 I_4031 (I70346,I1803,I70151,I70372,);
not I_4032 (I70380,I70372);
not I_4033 (I70397,I22857);
nand I_4034 (I70414,I70397,I22845);
and I_4035 (I70431,I70233,I70414);
nor I_4036 (I70448,I70346,I70431);
DFFARX1 I_4037 (I70448,I1803,I70151,I70119,);
DFFARX1 I_4038 (I70431,I1803,I70151,I70140,);
nor I_4039 (I70493,I22857,I22851);
nor I_4040 (I70131,I70346,I70493);
or I_4041 (I70524,I22857,I22851);
nor I_4042 (I70541,I22848,I22842);
DFFARX1 I_4043 (I70541,I1803,I70151,I70567,);
not I_4044 (I70575,I70567);
nor I_4045 (I70137,I70575,I70380);
nand I_4046 (I70606,I70575,I70225);
not I_4047 (I70623,I22848);
nand I_4048 (I70640,I70623,I70329);
nand I_4049 (I70657,I70575,I70640);
nand I_4050 (I70128,I70657,I70606);
nand I_4051 (I70125,I70640,I70524);
not I_4052 (I70729,I1810);
DFFARX1 I_4053 (I17599,I1803,I70729,I70755,);
and I_4054 (I70763,I70755,I17584);
DFFARX1 I_4055 (I70763,I1803,I70729,I70712,);
DFFARX1 I_4056 (I17590,I1803,I70729,I70803,);
not I_4057 (I70811,I17572);
not I_4058 (I70828,I17593);
nand I_4059 (I70845,I70828,I70811);
nor I_4060 (I70700,I70803,I70845);
DFFARX1 I_4061 (I70845,I1803,I70729,I70885,);
not I_4062 (I70721,I70885);
not I_4063 (I70907,I17596);
nand I_4064 (I70924,I70828,I70907);
DFFARX1 I_4065 (I70924,I1803,I70729,I70950,);
not I_4066 (I70958,I70950);
not I_4067 (I70975,I17587);
nand I_4068 (I70992,I70975,I17575);
and I_4069 (I71009,I70811,I70992);
nor I_4070 (I71026,I70924,I71009);
DFFARX1 I_4071 (I71026,I1803,I70729,I70697,);
DFFARX1 I_4072 (I71009,I1803,I70729,I70718,);
nor I_4073 (I71071,I17587,I17581);
nor I_4074 (I70709,I70924,I71071);
or I_4075 (I71102,I17587,I17581);
nor I_4076 (I71119,I17578,I17572);
DFFARX1 I_4077 (I71119,I1803,I70729,I71145,);
not I_4078 (I71153,I71145);
nor I_4079 (I70715,I71153,I70958);
nand I_4080 (I71184,I71153,I70803);
not I_4081 (I71201,I17578);
nand I_4082 (I71218,I71201,I70907);
nand I_4083 (I71235,I71153,I71218);
nand I_4084 (I70706,I71235,I71184);
nand I_4085 (I70703,I71218,I71102);
not I_4086 (I71307,I1810);
DFFARX1 I_4087 (I44549,I1803,I71307,I71333,);
and I_4088 (I71341,I71333,I44537);
DFFARX1 I_4089 (I71341,I1803,I71307,I71290,);
DFFARX1 I_4090 (I44540,I1803,I71307,I71381,);
not I_4091 (I71389,I44534);
not I_4092 (I71406,I44558);
nand I_4093 (I71423,I71406,I71389);
nor I_4094 (I71278,I71381,I71423);
DFFARX1 I_4095 (I71423,I1803,I71307,I71463,);
not I_4096 (I71299,I71463);
not I_4097 (I71485,I44546);
nand I_4098 (I71502,I71406,I71485);
DFFARX1 I_4099 (I71502,I1803,I71307,I71528,);
not I_4100 (I71536,I71528);
not I_4101 (I71553,I44555);
nand I_4102 (I71570,I71553,I44552);
and I_4103 (I71587,I71389,I71570);
nor I_4104 (I71604,I71502,I71587);
DFFARX1 I_4105 (I71604,I1803,I71307,I71275,);
DFFARX1 I_4106 (I71587,I1803,I71307,I71296,);
nor I_4107 (I71649,I44555,I44543);
nor I_4108 (I71287,I71502,I71649);
or I_4109 (I71680,I44555,I44543);
nor I_4110 (I71697,I44534,I44537);
DFFARX1 I_4111 (I71697,I1803,I71307,I71723,);
not I_4112 (I71731,I71723);
nor I_4113 (I71293,I71731,I71536);
nand I_4114 (I71762,I71731,I71381);
not I_4115 (I71779,I44534);
nand I_4116 (I71796,I71779,I71485);
nand I_4117 (I71813,I71731,I71796);
nand I_4118 (I71284,I71813,I71762);
nand I_4119 (I71281,I71796,I71680);
not I_4120 (I71885,I1810);
DFFARX1 I_4121 (I57171,I1803,I71885,I71911,);
and I_4122 (I71919,I71911,I57165);
DFFARX1 I_4123 (I71919,I1803,I71885,I71868,);
DFFARX1 I_4124 (I57183,I1803,I71885,I71959,);
not I_4125 (I71967,I57174);
not I_4126 (I71984,I57186);
nand I_4127 (I72001,I71984,I71967);
nor I_4128 (I71856,I71959,I72001);
DFFARX1 I_4129 (I72001,I1803,I71885,I72041,);
not I_4130 (I71877,I72041);
not I_4131 (I72063,I57192);
nand I_4132 (I72080,I71984,I72063);
DFFARX1 I_4133 (I72080,I1803,I71885,I72106,);
not I_4134 (I72114,I72106);
not I_4135 (I72131,I57168);
nand I_4136 (I72148,I72131,I57189);
and I_4137 (I72165,I71967,I72148);
nor I_4138 (I72182,I72080,I72165);
DFFARX1 I_4139 (I72182,I1803,I71885,I71853,);
DFFARX1 I_4140 (I72165,I1803,I71885,I71874,);
nor I_4141 (I72227,I57168,I57180);
nor I_4142 (I71865,I72080,I72227);
or I_4143 (I72258,I57168,I57180);
nor I_4144 (I72275,I57165,I57177);
DFFARX1 I_4145 (I72275,I1803,I71885,I72301,);
not I_4146 (I72309,I72301);
nor I_4147 (I71871,I72309,I72114);
nand I_4148 (I72340,I72309,I71959);
not I_4149 (I72357,I57165);
nand I_4150 (I72374,I72357,I72063);
nand I_4151 (I72391,I72309,I72374);
nand I_4152 (I71862,I72391,I72340);
nand I_4153 (I71859,I72374,I72258);
not I_4154 (I72463,I1810);
DFFARX1 I_4155 (I63203,I1803,I72463,I72489,);
and I_4156 (I72497,I72489,I63200);
DFFARX1 I_4157 (I72497,I1803,I72463,I72446,);
DFFARX1 I_4158 (I63206,I1803,I72463,I72537,);
not I_4159 (I72545,I63209);
not I_4160 (I72562,I63203);
nand I_4161 (I72579,I72562,I72545);
nor I_4162 (I72434,I72537,I72579);
DFFARX1 I_4163 (I72579,I1803,I72463,I72619,);
not I_4164 (I72455,I72619);
not I_4165 (I72641,I63218);
nand I_4166 (I72658,I72562,I72641);
DFFARX1 I_4167 (I72658,I1803,I72463,I72684,);
not I_4168 (I72692,I72684);
not I_4169 (I72709,I63215);
nand I_4170 (I72726,I72709,I63221);
and I_4171 (I72743,I72545,I72726);
nor I_4172 (I72760,I72658,I72743);
DFFARX1 I_4173 (I72760,I1803,I72463,I72431,);
DFFARX1 I_4174 (I72743,I1803,I72463,I72452,);
nor I_4175 (I72805,I63215,I63200);
nor I_4176 (I72443,I72658,I72805);
or I_4177 (I72836,I63215,I63200);
nor I_4178 (I72853,I63212,I63206);
DFFARX1 I_4179 (I72853,I1803,I72463,I72879,);
not I_4180 (I72887,I72879);
nor I_4181 (I72449,I72887,I72692);
nand I_4182 (I72918,I72887,I72537);
not I_4183 (I72935,I63212);
nand I_4184 (I72952,I72935,I72641);
nand I_4185 (I72969,I72887,I72952);
nand I_4186 (I72440,I72969,I72918);
nand I_4187 (I72437,I72952,I72836);
not I_4188 (I73041,I1810);
DFFARX1 I_4189 (I14878,I1803,I73041,I73067,);
nand I_4190 (I73075,I73067,I14893);
DFFARX1 I_4191 (I14890,I1803,I73041,I73101,);
DFFARX1 I_4192 (I73101,I1803,I73041,I73118,);
not I_4193 (I73033,I73118);
not I_4194 (I73140,I14869);
nor I_4195 (I73157,I14869,I14875);
not I_4196 (I73174,I14881);
nand I_4197 (I73191,I73140,I73174);
nor I_4198 (I73208,I14881,I14869);
and I_4199 (I73012,I73208,I73075);
not I_4200 (I73239,I14887);
nand I_4201 (I73256,I73239,I14869);
nor I_4202 (I73273,I14887,I14872);
not I_4203 (I73290,I73273);
nand I_4204 (I73015,I73157,I73290);
DFFARX1 I_4205 (I73273,I1803,I73041,I73030,);
nor I_4206 (I73335,I14872,I14881);
nor I_4207 (I73352,I73335,I14875);
and I_4208 (I73369,I73352,I73256);
DFFARX1 I_4209 (I73369,I1803,I73041,I73027,);
nor I_4210 (I73024,I73335,I73191);
or I_4211 (I73021,I73273,I73335);
nor I_4212 (I73428,I14872,I14884);
DFFARX1 I_4213 (I73428,I1803,I73041,I73454,);
not I_4214 (I73462,I73454);
nand I_4215 (I73479,I73462,I73140);
nor I_4216 (I73496,I73479,I14875);
DFFARX1 I_4217 (I73496,I1803,I73041,I73009,);
nor I_4218 (I73527,I73462,I73191);
nor I_4219 (I73018,I73335,I73527);
not I_4220 (I73585,I1810);
DFFARX1 I_4221 (I31189,I1803,I73585,I73611,);
nand I_4222 (I73619,I73611,I31213);
DFFARX1 I_4223 (I31192,I1803,I73585,I73645,);
DFFARX1 I_4224 (I73645,I1803,I73585,I73662,);
not I_4225 (I73577,I73662);
not I_4226 (I73684,I31195);
nor I_4227 (I73701,I31195,I31210);
not I_4228 (I73718,I31201);
nand I_4229 (I73735,I73684,I73718);
nor I_4230 (I73752,I31201,I31195);
and I_4231 (I73556,I73752,I73619);
not I_4232 (I73783,I31198);
nand I_4233 (I73800,I73783,I31192);
nor I_4234 (I73817,I31198,I31207);
not I_4235 (I73834,I73817);
nand I_4236 (I73559,I73701,I73834);
DFFARX1 I_4237 (I73817,I1803,I73585,I73574,);
nor I_4238 (I73879,I31204,I31201);
nor I_4239 (I73896,I73879,I31210);
and I_4240 (I73913,I73896,I73800);
DFFARX1 I_4241 (I73913,I1803,I73585,I73571,);
nor I_4242 (I73568,I73879,I73735);
or I_4243 (I73565,I73817,I73879);
nor I_4244 (I73972,I31204,I31189);
DFFARX1 I_4245 (I73972,I1803,I73585,I73998,);
not I_4246 (I74006,I73998);
nand I_4247 (I74023,I74006,I73684);
nor I_4248 (I74040,I74023,I31210);
DFFARX1 I_4249 (I74040,I1803,I73585,I73553,);
nor I_4250 (I74071,I74006,I73735);
nor I_4251 (I73562,I73879,I74071);
not I_4252 (I74129,I1810);
DFFARX1 I_4253 (I59749,I1803,I74129,I74155,);
nand I_4254 (I74163,I74155,I59749);
DFFARX1 I_4255 (I59761,I1803,I74129,I74189,);
DFFARX1 I_4256 (I74189,I1803,I74129,I74206,);
not I_4257 (I74121,I74206);
not I_4258 (I74228,I59755);
nor I_4259 (I74245,I59755,I59776);
not I_4260 (I74262,I59764);
nand I_4261 (I74279,I74228,I74262);
nor I_4262 (I74296,I59764,I59755);
and I_4263 (I74100,I74296,I74163);
not I_4264 (I74327,I59758);
nand I_4265 (I74344,I74327,I59773);
nor I_4266 (I74361,I59758,I59767);
not I_4267 (I74378,I74361);
nand I_4268 (I74103,I74245,I74378);
DFFARX1 I_4269 (I74361,I1803,I74129,I74118,);
nor I_4270 (I74423,I59770,I59764);
nor I_4271 (I74440,I74423,I59776);
and I_4272 (I74457,I74440,I74344);
DFFARX1 I_4273 (I74457,I1803,I74129,I74115,);
nor I_4274 (I74112,I74423,I74279);
or I_4275 (I74109,I74361,I74423);
nor I_4276 (I74516,I59770,I59752);
DFFARX1 I_4277 (I74516,I1803,I74129,I74542,);
not I_4278 (I74550,I74542);
nand I_4279 (I74567,I74550,I74228);
nor I_4280 (I74584,I74567,I59776);
DFFARX1 I_4281 (I74584,I1803,I74129,I74097,);
nor I_4282 (I74615,I74550,I74279);
nor I_4283 (I74106,I74423,I74615);
not I_4284 (I74673,I1810);
DFFARX1 I_4285 (I52122,I1803,I74673,I74699,);
nand I_4286 (I74707,I74699,I52116);
DFFARX1 I_4287 (I52119,I1803,I74673,I74733,);
DFFARX1 I_4288 (I74733,I1803,I74673,I74750,);
not I_4289 (I74665,I74750);
not I_4290 (I74772,I52125);
nor I_4291 (I74789,I52125,I52119);
not I_4292 (I74806,I52128);
nand I_4293 (I74823,I74772,I74806);
nor I_4294 (I74840,I52128,I52125);
and I_4295 (I74644,I74840,I74707);
not I_4296 (I74871,I52137);
nand I_4297 (I74888,I74871,I52131);
nor I_4298 (I74905,I52137,I52134);
not I_4299 (I74922,I74905);
nand I_4300 (I74647,I74789,I74922);
DFFARX1 I_4301 (I74905,I1803,I74673,I74662,);
nor I_4302 (I74967,I52116,I52128);
nor I_4303 (I74984,I74967,I52119);
and I_4304 (I75001,I74984,I74888);
DFFARX1 I_4305 (I75001,I1803,I74673,I74659,);
nor I_4306 (I74656,I74967,I74823);
or I_4307 (I74653,I74905,I74967);
nor I_4308 (I75060,I52116,I52122);
DFFARX1 I_4309 (I75060,I1803,I74673,I75086,);
not I_4310 (I75094,I75086);
nand I_4311 (I75111,I75094,I74772);
nor I_4312 (I75128,I75111,I52119);
DFFARX1 I_4313 (I75128,I1803,I74673,I74641,);
nor I_4314 (I75159,I75094,I74823);
nor I_4315 (I74650,I74967,I75159);
not I_4316 (I75217,I1810);
DFFARX1 I_4317 (I77498,I1803,I75217,I75243,);
nand I_4318 (I75251,I75243,I77492);
not I_4319 (I75268,I75251);
DFFARX1 I_4320 (I77507,I1803,I75217,I75294,);
not I_4321 (I75302,I75294);
not I_4322 (I75319,I77483);
or I_4323 (I75336,I77480,I77483);
nor I_4324 (I75353,I77480,I77483);
or I_4325 (I75370,I77486,I77480);
DFFARX1 I_4326 (I75370,I1803,I75217,I75209,);
not I_4327 (I75401,I77480);
nand I_4328 (I75418,I75401,I77495);
nand I_4329 (I75435,I75319,I75418);
and I_4330 (I75188,I75302,I75435);
nor I_4331 (I75466,I77480,I77489);
and I_4332 (I75483,I75302,I75466);
nor I_4333 (I75194,I75268,I75483);
DFFARX1 I_4334 (I75466,I1803,I75217,I75523,);
not I_4335 (I75531,I75523);
nor I_4336 (I75203,I75302,I75531);
or I_4337 (I75562,I75370,I77504);
nor I_4338 (I75579,I77504,I77486);
nand I_4339 (I75596,I75435,I75579);
nand I_4340 (I75613,I75562,I75596);
DFFARX1 I_4341 (I75613,I1803,I75217,I75206,);
nor I_4342 (I75644,I75579,I75336);
DFFARX1 I_4343 (I75644,I1803,I75217,I75185,);
nor I_4344 (I75675,I77504,I77501);
DFFARX1 I_4345 (I75675,I1803,I75217,I75701,);
DFFARX1 I_4346 (I75701,I1803,I75217,I75200,);
not I_4347 (I75723,I75701);
nand I_4348 (I75197,I75723,I75251);
nand I_4349 (I75191,I75723,I75353);
not I_4350 (I75795,I1810);
DFFARX1 I_4351 (I2873,I1803,I75795,I75821,);
nand I_4352 (I75829,I75821,I2867);
not I_4353 (I75846,I75829);
DFFARX1 I_4354 (I2885,I1803,I75795,I75872,);
not I_4355 (I75880,I75872);
not I_4356 (I75897,I2888);
or I_4357 (I75914,I2891,I2888);
nor I_4358 (I75931,I2891,I2888);
or I_4359 (I75948,I2876,I2891);
DFFARX1 I_4360 (I75948,I1803,I75795,I75787,);
not I_4361 (I75979,I2879);
nand I_4362 (I75996,I75979,I2882);
nand I_4363 (I76013,I75897,I75996);
and I_4364 (I75766,I75880,I76013);
nor I_4365 (I76044,I2879,I2870);
and I_4366 (I76061,I75880,I76044);
nor I_4367 (I75772,I75846,I76061);
DFFARX1 I_4368 (I76044,I1803,I75795,I76101,);
not I_4369 (I76109,I76101);
nor I_4370 (I75781,I75880,I76109);
or I_4371 (I76140,I75948,I2870);
nor I_4372 (I76157,I2870,I2876);
nand I_4373 (I76174,I76013,I76157);
nand I_4374 (I76191,I76140,I76174);
DFFARX1 I_4375 (I76191,I1803,I75795,I75784,);
nor I_4376 (I76222,I76157,I75914);
DFFARX1 I_4377 (I76222,I1803,I75795,I75763,);
nor I_4378 (I76253,I2870,I2867);
DFFARX1 I_4379 (I76253,I1803,I75795,I76279,);
DFFARX1 I_4380 (I76279,I1803,I75795,I75778,);
not I_4381 (I76301,I76279);
nand I_4382 (I75775,I76301,I75829);
nand I_4383 (I75769,I76301,I75931);
not I_4384 (I76373,I1810);
DFFARX1 I_4385 (I46268,I1803,I76373,I76399,);
nand I_4386 (I76407,I76399,I46271);
not I_4387 (I76424,I76407);
DFFARX1 I_4388 (I46283,I1803,I76373,I76450,);
not I_4389 (I76458,I76450);
not I_4390 (I76475,I46268);
or I_4391 (I76492,I46277,I46268);
nor I_4392 (I76509,I46277,I46268);
or I_4393 (I76526,I46286,I46277);
DFFARX1 I_4394 (I76526,I1803,I76373,I76365,);
not I_4395 (I76557,I46289);
nand I_4396 (I76574,I76557,I46271);
nand I_4397 (I76591,I76475,I76574);
and I_4398 (I76344,I76458,I76591);
nor I_4399 (I76622,I46289,I46274);
and I_4400 (I76639,I76458,I76622);
nor I_4401 (I76350,I76424,I76639);
DFFARX1 I_4402 (I76622,I1803,I76373,I76679,);
not I_4403 (I76687,I76679);
nor I_4404 (I76359,I76458,I76687);
or I_4405 (I76718,I76526,I46280);
nor I_4406 (I76735,I46280,I46286);
nand I_4407 (I76752,I76591,I76735);
nand I_4408 (I76769,I76718,I76752);
DFFARX1 I_4409 (I76769,I1803,I76373,I76362,);
nor I_4410 (I76800,I76735,I76492);
DFFARX1 I_4411 (I76800,I1803,I76373,I76341,);
nor I_4412 (I76831,I46280,I46292);
DFFARX1 I_4413 (I76831,I1803,I76373,I76857,);
DFFARX1 I_4414 (I76857,I1803,I76373,I76356,);
not I_4415 (I76879,I76857);
nand I_4416 (I76353,I76879,I76407);
nand I_4417 (I76347,I76879,I76509);
not I_4418 (I76954,I1810);
DFFARX1 I_4419 (I38772,I1803,I76954,I76980,);
nand I_4420 (I76988,I76980,I38757);
not I_4421 (I77005,I76988);
DFFARX1 I_4422 (I38775,I1803,I76954,I77031,);
not I_4423 (I77039,I77031);
nor I_4424 (I77056,I38754,I38769);
not I_4425 (I77073,I77056);
DFFARX1 I_4426 (I77073,I1803,I76954,I76940,);
or I_4427 (I77104,I38766,I38754);
DFFARX1 I_4428 (I77104,I1803,I76954,I76943,);
not I_4429 (I77135,I38754);
nor I_4430 (I77152,I77135,I38763);
nor I_4431 (I77169,I77152,I38769);
nor I_4432 (I77186,I38763,I38757);
nor I_4433 (I77203,I77039,I77186);
nor I_4434 (I76928,I77005,I77203);
not I_4435 (I77234,I77186);
nand I_4436 (I76931,I77234,I76988);
nand I_4437 (I76925,I77234,I77056);
nor I_4438 (I76922,I77186,I77169);
nor I_4439 (I77293,I38760,I38766);
not I_4440 (I77310,I77293);
DFFARX1 I_4441 (I77293,I1803,I76954,I77336,);
not I_4442 (I76946,I77336);
nor I_4443 (I77358,I38760,I38778);
DFFARX1 I_4444 (I77358,I1803,I76954,I77384,);
and I_4445 (I77392,I77384,I38754);
nor I_4446 (I77409,I77392,I77310);
DFFARX1 I_4447 (I77409,I1803,I76954,I76937,);
nor I_4448 (I77440,I77384,I77169);
DFFARX1 I_4449 (I77440,I1803,I76954,I76919,);
nor I_4450 (I76934,I77384,I77073);
not I_4451 (I77515,I1810);
DFFARX1 I_4452 (I42240,I1803,I77515,I77541,);
nand I_4453 (I77549,I77541,I42225);
not I_4454 (I77566,I77549);
DFFARX1 I_4455 (I42243,I1803,I77515,I77592,);
not I_4456 (I77600,I77592);
nor I_4457 (I77617,I42222,I42237);
not I_4458 (I77634,I77617);
DFFARX1 I_4459 (I77634,I1803,I77515,I77501,);
or I_4460 (I77665,I42234,I42222);
DFFARX1 I_4461 (I77665,I1803,I77515,I77504,);
not I_4462 (I77696,I42222);
nor I_4463 (I77713,I77696,I42231);
nor I_4464 (I77730,I77713,I42237);
nor I_4465 (I77747,I42231,I42225);
nor I_4466 (I77764,I77600,I77747);
nor I_4467 (I77489,I77566,I77764);
not I_4468 (I77795,I77747);
nand I_4469 (I77492,I77795,I77549);
nand I_4470 (I77486,I77795,I77617);
nor I_4471 (I77483,I77747,I77730);
nor I_4472 (I77854,I42228,I42234);
not I_4473 (I77871,I77854);
DFFARX1 I_4474 (I77854,I1803,I77515,I77897,);
not I_4475 (I77507,I77897);
nor I_4476 (I77919,I42228,I42246);
DFFARX1 I_4477 (I77919,I1803,I77515,I77945,);
and I_4478 (I77953,I77945,I42222);
nor I_4479 (I77970,I77953,I77871);
DFFARX1 I_4480 (I77970,I1803,I77515,I77498,);
nor I_4481 (I78001,I77945,I77730);
DFFARX1 I_4482 (I78001,I1803,I77515,I77480,);
nor I_4483 (I77495,I77945,I77634);
not I_4484 (I78076,I1810);
DFFARX1 I_4485 (I48436,I1803,I78076,I78102,);
DFFARX1 I_4486 (I48433,I1803,I78076,I78119,);
not I_4487 (I78127,I78119);
nor I_4488 (I78044,I78102,I78127);
DFFARX1 I_4489 (I78127,I1803,I78076,I78059,);
nor I_4490 (I78172,I48448,I48430);
and I_4491 (I78189,I78172,I48427);
nor I_4492 (I78206,I78189,I48448);
not I_4493 (I78223,I48448);
and I_4494 (I78240,I78223,I48433);
nand I_4495 (I78257,I78240,I48445);
nor I_4496 (I78274,I78223,I78257);
DFFARX1 I_4497 (I78274,I1803,I78076,I78041,);
not I_4498 (I78305,I78257);
nand I_4499 (I78322,I78127,I78305);
nand I_4500 (I78053,I78189,I78305);
DFFARX1 I_4501 (I78223,I1803,I78076,I78068,);
not I_4502 (I78367,I48439);
nor I_4503 (I78384,I78367,I48433);
nor I_4504 (I78401,I78384,I78206);
DFFARX1 I_4505 (I78401,I1803,I78076,I78065,);
not I_4506 (I78432,I78384);
DFFARX1 I_4507 (I78432,I1803,I78076,I78458,);
not I_4508 (I78466,I78458);
nor I_4509 (I78062,I78466,I78384);
nor I_4510 (I78497,I78367,I48427);
and I_4511 (I78514,I78497,I48442);
or I_4512 (I78531,I78514,I48430);
DFFARX1 I_4513 (I78531,I1803,I78076,I78557,);
not I_4514 (I78565,I78557);
nand I_4515 (I78582,I78565,I78305);
not I_4516 (I78056,I78582);
nand I_4517 (I78050,I78582,I78322);
nand I_4518 (I78047,I78565,I78189);
not I_4519 (I78671,I1810);
DFFARX1 I_4520 (I73009,I1803,I78671,I78697,);
DFFARX1 I_4521 (I73012,I1803,I78671,I78714,);
not I_4522 (I78722,I78714);
nor I_4523 (I78639,I78697,I78722);
DFFARX1 I_4524 (I78722,I1803,I78671,I78654,);
nor I_4525 (I78767,I73012,I73027);
and I_4526 (I78784,I78767,I73021);
nor I_4527 (I78801,I78784,I73012);
not I_4528 (I78818,I73012);
and I_4529 (I78835,I78818,I73030);
nand I_4530 (I78852,I78835,I73018);
nor I_4531 (I78869,I78818,I78852);
DFFARX1 I_4532 (I78869,I1803,I78671,I78636,);
not I_4533 (I78900,I78852);
nand I_4534 (I78917,I78722,I78900);
nand I_4535 (I78648,I78784,I78900);
DFFARX1 I_4536 (I78818,I1803,I78671,I78663,);
not I_4537 (I78962,I73024);
nor I_4538 (I78979,I78962,I73030);
nor I_4539 (I78996,I78979,I78801);
DFFARX1 I_4540 (I78996,I1803,I78671,I78660,);
not I_4541 (I79027,I78979);
DFFARX1 I_4542 (I79027,I1803,I78671,I79053,);
not I_4543 (I79061,I79053);
nor I_4544 (I78657,I79061,I78979);
nor I_4545 (I79092,I78962,I73009);
and I_4546 (I79109,I79092,I73033);
or I_4547 (I79126,I79109,I73015);
DFFARX1 I_4548 (I79126,I1803,I78671,I79152,);
not I_4549 (I79160,I79152);
nand I_4550 (I79177,I79160,I78900);
not I_4551 (I78651,I79177);
nand I_4552 (I78645,I79177,I78917);
nand I_4553 (I78642,I79160,I78784);
not I_4554 (I79266,I1810);
DFFARX1 I_4555 (I1420,I1803,I79266,I79292,);
DFFARX1 I_4556 (I1724,I1803,I79266,I79309,);
not I_4557 (I79317,I79309);
nor I_4558 (I79234,I79292,I79317);
DFFARX1 I_4559 (I79317,I1803,I79266,I79249,);
nor I_4560 (I79362,I1788,I1604);
and I_4561 (I79379,I79362,I1556);
nor I_4562 (I79396,I79379,I1788);
not I_4563 (I79413,I1788);
and I_4564 (I79430,I79413,I1516);
nand I_4565 (I79447,I79430,I1732);
nor I_4566 (I79464,I79413,I79447);
DFFARX1 I_4567 (I79464,I1803,I79266,I79231,);
not I_4568 (I79495,I79447);
nand I_4569 (I79512,I79317,I79495);
nand I_4570 (I79243,I79379,I79495);
DFFARX1 I_4571 (I79413,I1803,I79266,I79258,);
not I_4572 (I79557,I1500);
nor I_4573 (I79574,I79557,I1516);
nor I_4574 (I79591,I79574,I79396);
DFFARX1 I_4575 (I79591,I1803,I79266,I79255,);
not I_4576 (I79622,I79574);
DFFARX1 I_4577 (I79622,I1803,I79266,I79648,);
not I_4578 (I79656,I79648);
nor I_4579 (I79252,I79656,I79574);
nor I_4580 (I79687,I79557,I1612);
and I_4581 (I79704,I79687,I1388);
or I_4582 (I79721,I79704,I1380);
DFFARX1 I_4583 (I79721,I1803,I79266,I79747,);
not I_4584 (I79755,I79747);
nand I_4585 (I79772,I79755,I79495);
not I_4586 (I79246,I79772);
nand I_4587 (I79240,I79772,I79512);
nand I_4588 (I79237,I79755,I79379);
not I_4589 (I79861,I1810);
DFFARX1 I_4590 (I34729,I1803,I79861,I79887,);
DFFARX1 I_4591 (I34723,I1803,I79861,I79904,);
not I_4592 (I79912,I79904);
nor I_4593 (I79829,I79887,I79912);
DFFARX1 I_4594 (I79912,I1803,I79861,I79844,);
nor I_4595 (I79957,I34720,I34711);
and I_4596 (I79974,I79957,I34708);
nor I_4597 (I79991,I79974,I34720);
not I_4598 (I80008,I34720);
and I_4599 (I80025,I80008,I34714);
nand I_4600 (I80042,I80025,I34726);
nor I_4601 (I80059,I80008,I80042);
DFFARX1 I_4602 (I80059,I1803,I79861,I79826,);
not I_4603 (I80090,I80042);
nand I_4604 (I80107,I79912,I80090);
nand I_4605 (I79838,I79974,I80090);
DFFARX1 I_4606 (I80008,I1803,I79861,I79853,);
not I_4607 (I80152,I34732);
nor I_4608 (I80169,I80152,I34714);
nor I_4609 (I80186,I80169,I79991);
DFFARX1 I_4610 (I80186,I1803,I79861,I79850,);
not I_4611 (I80217,I80169);
DFFARX1 I_4612 (I80217,I1803,I79861,I80243,);
not I_4613 (I80251,I80243);
nor I_4614 (I79847,I80251,I80169);
nor I_4615 (I80282,I80152,I34711);
and I_4616 (I80299,I80282,I34717);
or I_4617 (I80316,I80299,I34708);
DFFARX1 I_4618 (I80316,I1803,I79861,I80342,);
not I_4619 (I80350,I80342);
nand I_4620 (I80367,I80350,I80090);
not I_4621 (I79841,I80367);
nand I_4622 (I79835,I80367,I80107);
nand I_4623 (I79832,I80350,I79974);
not I_4624 (I80456,I1810);
DFFARX1 I_4625 (I1740,I1803,I80456,I80482,);
DFFARX1 I_4626 (I1660,I1803,I80456,I80499,);
not I_4627 (I80507,I80499);
nor I_4628 (I80424,I80482,I80507);
DFFARX1 I_4629 (I80507,I1803,I80456,I80439,);
nor I_4630 (I80552,I1580,I1476);
and I_4631 (I80569,I80552,I1436);
nor I_4632 (I80586,I80569,I1580);
not I_4633 (I80603,I1580);
and I_4634 (I80620,I80603,I1572);
nand I_4635 (I80637,I80620,I1708);
nor I_4636 (I80654,I80603,I80637);
DFFARX1 I_4637 (I80654,I1803,I80456,I80421,);
not I_4638 (I80685,I80637);
nand I_4639 (I80702,I80507,I80685);
nand I_4640 (I80433,I80569,I80685);
DFFARX1 I_4641 (I80603,I1803,I80456,I80448,);
not I_4642 (I80747,I1676);
nor I_4643 (I80764,I80747,I1572);
nor I_4644 (I80781,I80764,I80586);
DFFARX1 I_4645 (I80781,I1803,I80456,I80445,);
not I_4646 (I80812,I80764);
DFFARX1 I_4647 (I80812,I1803,I80456,I80838,);
not I_4648 (I80846,I80838);
nor I_4649 (I80442,I80846,I80764);
nor I_4650 (I80877,I80747,I1780);
and I_4651 (I80894,I80877,I1532);
or I_4652 (I80911,I80894,I1428);
DFFARX1 I_4653 (I80911,I1803,I80456,I80937,);
not I_4654 (I80945,I80937);
nand I_4655 (I80962,I80945,I80685);
not I_4656 (I80436,I80962);
nand I_4657 (I80430,I80962,I80702);
nand I_4658 (I80427,I80945,I80569);
not I_4659 (I81051,I1810);
DFFARX1 I_4660 (I32379,I1803,I81051,I81077,);
DFFARX1 I_4661 (I32382,I1803,I81051,I81094,);
not I_4662 (I81102,I81094);
nor I_4663 (I81019,I81077,I81102);
DFFARX1 I_4664 (I81102,I1803,I81051,I81034,);
nor I_4665 (I81147,I32385,I32403);
and I_4666 (I81164,I81147,I32388);
nor I_4667 (I81181,I81164,I32385);
not I_4668 (I81198,I32385);
and I_4669 (I81215,I81198,I32397);
nand I_4670 (I81232,I81215,I32400);
nor I_4671 (I81249,I81198,I81232);
DFFARX1 I_4672 (I81249,I1803,I81051,I81016,);
not I_4673 (I81280,I81232);
nand I_4674 (I81297,I81102,I81280);
nand I_4675 (I81028,I81164,I81280);
DFFARX1 I_4676 (I81198,I1803,I81051,I81043,);
not I_4677 (I81342,I32391);
nor I_4678 (I81359,I81342,I32397);
nor I_4679 (I81376,I81359,I81181);
DFFARX1 I_4680 (I81376,I1803,I81051,I81040,);
not I_4681 (I81407,I81359);
DFFARX1 I_4682 (I81407,I1803,I81051,I81433,);
not I_4683 (I81441,I81433);
nor I_4684 (I81037,I81441,I81359);
nor I_4685 (I81472,I81342,I32379);
and I_4686 (I81489,I81472,I32394);
or I_4687 (I81506,I81489,I32382);
DFFARX1 I_4688 (I81506,I1803,I81051,I81532,);
not I_4689 (I81540,I81532);
nand I_4690 (I81557,I81540,I81280);
not I_4691 (I81031,I81557);
nand I_4692 (I81025,I81557,I81297);
nand I_4693 (I81022,I81540,I81164);
not I_4694 (I81646,I1810);
DFFARX1 I_4695 (I61529,I1803,I81646,I81672,);
DFFARX1 I_4696 (I61520,I1803,I81646,I81689,);
not I_4697 (I81697,I81689);
nor I_4698 (I81614,I81672,I81697);
DFFARX1 I_4699 (I81697,I1803,I81646,I81629,);
nor I_4700 (I81742,I61526,I61535);
and I_4701 (I81759,I81742,I61538);
nor I_4702 (I81776,I81759,I61526);
not I_4703 (I81793,I61526);
and I_4704 (I81810,I81793,I61517);
nand I_4705 (I81827,I81810,I61523);
nor I_4706 (I81844,I81793,I81827);
DFFARX1 I_4707 (I81844,I1803,I81646,I81611,);
not I_4708 (I81875,I81827);
nand I_4709 (I81892,I81697,I81875);
nand I_4710 (I81623,I81759,I81875);
DFFARX1 I_4711 (I81793,I1803,I81646,I81638,);
not I_4712 (I81937,I61532);
nor I_4713 (I81954,I81937,I61517);
nor I_4714 (I81971,I81954,I81776);
DFFARX1 I_4715 (I81971,I1803,I81646,I81635,);
not I_4716 (I82002,I81954);
DFFARX1 I_4717 (I82002,I1803,I81646,I82028,);
not I_4718 (I82036,I82028);
nor I_4719 (I81632,I82036,I81954);
nor I_4720 (I82067,I81937,I61517);
and I_4721 (I82084,I82067,I61520);
or I_4722 (I82101,I82084,I61523);
DFFARX1 I_4723 (I82101,I1803,I81646,I82127,);
not I_4724 (I82135,I82127);
nand I_4725 (I82152,I82135,I81875);
not I_4726 (I81626,I82152);
nand I_4727 (I81620,I82152,I81892);
nand I_4728 (I81617,I82135,I81759);
not I_4729 (I82241,I1810);
DFFARX1 I_4730 (I17066,I1803,I82241,I82267,);
DFFARX1 I_4731 (I17060,I1803,I82241,I82284,);
not I_4732 (I82292,I82284);
nor I_4733 (I82209,I82267,I82292);
DFFARX1 I_4734 (I82292,I1803,I82241,I82224,);
nor I_4735 (I82337,I17048,I17069);
and I_4736 (I82354,I82337,I17063);
nor I_4737 (I82371,I82354,I17048);
not I_4738 (I82388,I17048);
and I_4739 (I82405,I82388,I17045);
nand I_4740 (I82422,I82405,I17057);
nor I_4741 (I82439,I82388,I82422);
DFFARX1 I_4742 (I82439,I1803,I82241,I82206,);
not I_4743 (I82470,I82422);
nand I_4744 (I82487,I82292,I82470);
nand I_4745 (I82218,I82354,I82470);
DFFARX1 I_4746 (I82388,I1803,I82241,I82233,);
not I_4747 (I82532,I17072);
nor I_4748 (I82549,I82532,I17045);
nor I_4749 (I82566,I82549,I82371);
DFFARX1 I_4750 (I82566,I1803,I82241,I82230,);
not I_4751 (I82597,I82549);
DFFARX1 I_4752 (I82597,I1803,I82241,I82623,);
not I_4753 (I82631,I82623);
nor I_4754 (I82227,I82631,I82549);
nor I_4755 (I82662,I82532,I17054);
and I_4756 (I82679,I82662,I17051);
or I_4757 (I82696,I82679,I17045);
DFFARX1 I_4758 (I82696,I1803,I82241,I82722,);
not I_4759 (I82730,I82722);
nand I_4760 (I82747,I82730,I82470);
not I_4761 (I82221,I82747);
nand I_4762 (I82215,I82747,I82487);
nand I_4763 (I82212,I82730,I82354);
not I_4764 (I82836,I1810);
DFFARX1 I_4765 (I60968,I1803,I82836,I82862,);
DFFARX1 I_4766 (I60959,I1803,I82836,I82879,);
not I_4767 (I82887,I82879);
nor I_4768 (I82804,I82862,I82887);
DFFARX1 I_4769 (I82887,I1803,I82836,I82819,);
nor I_4770 (I82932,I60965,I60974);
and I_4771 (I82949,I82932,I60977);
nor I_4772 (I82966,I82949,I60965);
not I_4773 (I82983,I60965);
and I_4774 (I83000,I82983,I60956);
nand I_4775 (I83017,I83000,I60962);
nor I_4776 (I83034,I82983,I83017);
DFFARX1 I_4777 (I83034,I1803,I82836,I82801,);
not I_4778 (I83065,I83017);
nand I_4779 (I83082,I82887,I83065);
nand I_4780 (I82813,I82949,I83065);
DFFARX1 I_4781 (I82983,I1803,I82836,I82828,);
not I_4782 (I83127,I60971);
nor I_4783 (I83144,I83127,I60956);
nor I_4784 (I83161,I83144,I82966);
DFFARX1 I_4785 (I83161,I1803,I82836,I82825,);
not I_4786 (I83192,I83144);
DFFARX1 I_4787 (I83192,I1803,I82836,I83218,);
not I_4788 (I83226,I83218);
nor I_4789 (I82822,I83226,I83144);
nor I_4790 (I83257,I83127,I60956);
and I_4791 (I83274,I83257,I60959);
or I_4792 (I83291,I83274,I60962);
DFFARX1 I_4793 (I83291,I1803,I82836,I83317,);
not I_4794 (I83325,I83317);
nand I_4795 (I83342,I83325,I83065);
not I_4796 (I82816,I83342);
nand I_4797 (I82810,I83342,I83082);
nand I_4798 (I82807,I83325,I82949);
not I_4799 (I83431,I1810);
DFFARX1 I_4800 (I27177,I1803,I83431,I83457,);
DFFARX1 I_4801 (I27183,I1803,I83431,I83474,);
not I_4802 (I83482,I83474);
nor I_4803 (I83399,I83457,I83482);
DFFARX1 I_4804 (I83482,I1803,I83431,I83414,);
nor I_4805 (I83527,I27192,I27177);
and I_4806 (I83544,I83527,I27204);
nor I_4807 (I83561,I83544,I27192);
not I_4808 (I83578,I27192);
and I_4809 (I83595,I83578,I27180);
nand I_4810 (I83612,I83595,I27201);
nor I_4811 (I83629,I83578,I83612);
DFFARX1 I_4812 (I83629,I1803,I83431,I83396,);
not I_4813 (I83660,I83612);
nand I_4814 (I83677,I83482,I83660);
nand I_4815 (I83408,I83544,I83660);
DFFARX1 I_4816 (I83578,I1803,I83431,I83423,);
not I_4817 (I83722,I27189);
nor I_4818 (I83739,I83722,I27180);
nor I_4819 (I83756,I83739,I83561);
DFFARX1 I_4820 (I83756,I1803,I83431,I83420,);
not I_4821 (I83787,I83739);
DFFARX1 I_4822 (I83787,I1803,I83431,I83813,);
not I_4823 (I83821,I83813);
nor I_4824 (I83417,I83821,I83739);
nor I_4825 (I83852,I83722,I27186);
and I_4826 (I83869,I83852,I27198);
or I_4827 (I83886,I83869,I27195);
DFFARX1 I_4828 (I83886,I1803,I83431,I83912,);
not I_4829 (I83920,I83912);
nand I_4830 (I83937,I83920,I83660);
not I_4831 (I83411,I83937);
nand I_4832 (I83405,I83937,I83677);
nand I_4833 (I83402,I83920,I83544);
endmodule


