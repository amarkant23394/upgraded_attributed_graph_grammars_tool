module test_I10647(I1477,I10647);
input I1477;
output I10647;
wire ;
not I_0(I10647,I1477);
endmodule


