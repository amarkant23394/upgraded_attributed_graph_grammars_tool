module test_I13970(I1477,I1470,I11990,I12174,I12459,I13970);
input I1477,I1470,I11990,I12174,I12459;
output I13970;
wire I11935,I12270,I11950,I12476,I10014,I12208,I10023,I12349,I12493,I11973,I12191;
DFFARX1 I_0(I12208,I1470,I11973,,,I11935,);
nand I_1(I12270,I11990,I10014);
DFFARX1 I_2(I12493,I1470,I11973,,,I11950,);
and I_3(I12476,I12349,I12459);
DFFARX1 I_4(I1470,,,I10014,);
DFFARX1 I_5(I12191,I1470,I11973,,,I12208,);
DFFARX1 I_6(I1470,,,I10023,);
DFFARX1 I_7(I1470,I11973,,,I12349,);
or I_8(I12493,I12270,I12476);
not I_9(I11973,I1477);
nand I_10(I13970,I11935,I11950);
or I_11(I12191,I12174,I10023);
endmodule


