module test_final(IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_4_2_l_6,IN_5_2_l_6,IN_1_6_l_6,IN_2_6_l_6,IN_3_6_l_6,IN_4_6_l_6,IN_5_6_l_6,IN_1_9_l_6,IN_2_9_l_6,IN_3_9_l_6,IN_4_9_l_6,IN_5_9_l_6,blif_clk_net_7_r_3,blif_reset_net_7_r_3,N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6134_9_r_3);
input IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_4_2_l_6,IN_5_2_l_6,IN_1_6_l_6,IN_2_6_l_6,IN_3_6_l_6,IN_4_6_l_6,IN_5_6_l_6,IN_1_9_l_6,IN_2_9_l_6,IN_3_9_l_6,IN_4_9_l_6,IN_5_9_l_6,blif_clk_net_7_r_3,blif_reset_net_7_r_3;
output N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6134_9_r_3;
wire N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,I_BUFF_1_9_r_6,N1372_10_r_6,N1508_10_r_6,N3_8_r_6,n30_6,n31_6,n32_6,n33_6,n34_6,n35_6,n36_6,n37_6,n38_6,n39_6,n40_6,n41_6,n42_6,n43_6,n44_6,n45_6,n46_6,n47_6,n48_6,n49_6,n50_6,n51_6,n52_6,n53_6,n54_6,n_572_7_r_3,N6147_9_r_3,I_BUFF_1_9_r_3,n4_7_r_3,n10_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3,n40_3,n41_3,n42_3,n43_3,n44_3,n45_3,n46_3,n47_3,n48_3,n49_3,n50_3,n51_3;
nor I_0(N1371_0_r_6,n30_6,n33_6);
nor I_1(N1508_0_r_6,n33_6,n44_6);
not I_2(N1372_1_r_6,n41_6);
nor I_3(N1508_1_r_6,n40_6,n41_6);
nor I_4(N1507_6_r_6,n39_6,n45_6);
nor I_5(N1508_6_r_6,n37_6,n38_6);
nor I_6(n_42_8_r_6,n30_6,n31_6);
DFFARX1 I_7(N3_8_r_6,blif_clk_net_7_r_3,n10_3,G199_8_r_6,);
nor I_8(N6147_9_r_6,n32_6,n33_6);
nor I_9(N6134_9_r_6,I_BUFF_1_9_r_6,n35_6);
not I_10(I_BUFF_1_9_r_6,n37_6);
not I_11(N1372_10_r_6,n43_6);
nor I_12(N1508_10_r_6,n42_6,n43_6);
nor I_13(N3_8_r_6,IN_1_9_l_6,n36_6);
nor I_14(n30_6,IN_5_9_l_6,n53_6);
not I_15(n31_6,n36_6);
nor I_16(n32_6,I_BUFF_1_9_r_6,n34_6);
not I_17(n33_6,IN_1_9_l_6);
not I_18(n34_6,n35_6);
nand I_19(n35_6,IN_2_6_l_6,n49_6);
nand I_20(n36_6,IN_5_6_l_6,n51_6);
nand I_21(n37_6,IN_2_9_l_6,n54_6);
or I_22(n38_6,n35_6,n39_6);
nor I_23(n39_6,n40_6,n45_6);
and I_24(n40_6,n46_6,n47_6);
nand I_25(n41_6,n30_6,n31_6);
nor I_26(n42_6,n34_6,n40_6);
nand I_27(n43_6,IN_1_9_l_6,n30_6);
nor I_28(n44_6,n31_6,n40_6);
nor I_29(n45_6,n35_6,n36_6);
nor I_30(n46_6,IN_1_2_l_6,IN_2_2_l_6);
or I_31(n47_6,IN_5_2_l_6,n48_6);
nor I_32(n48_6,IN_3_2_l_6,IN_4_2_l_6);
and I_33(n49_6,IN_1_6_l_6,n50_6);
nand I_34(n50_6,n51_6,n52_6);
nand I_35(n51_6,IN_3_6_l_6,IN_4_6_l_6);
not I_36(n52_6,IN_5_6_l_6);
nor I_37(n53_6,IN_3_9_l_6,IN_4_9_l_6);
or I_38(n54_6,IN_3_9_l_6,IN_4_9_l_6);
not I_39(N1372_1_r_3,n40_3);
nor I_40(N1508_1_r_3,N6147_9_r_3,n40_3);
nor I_41(N1507_6_r_3,n31_3,n42_3);
nor I_42(N1508_6_r_3,n30_3,n38_3);
DFFARX1 I_43(n4_7_r_3,blif_clk_net_7_r_3,n10_3,G42_7_r_3,);
nor I_44(n_572_7_r_3,I_BUFF_1_9_r_3,n35_3);
nand I_45(n_573_7_r_3,n30_3,n31_3);
nor I_46(n_549_7_r_3,N6147_9_r_3,n33_3);
nand I_47(n_569_7_r_3,n30_3,n32_3);
nor I_48(n_452_7_r_3,n35_3,N1372_10_r_6);
not I_49(N6147_9_r_3,n32_3);
nor I_50(N6134_9_r_3,n36_3,n37_3);
not I_51(I_BUFF_1_9_r_3,n45_3);
nor I_52(n4_7_r_3,I_BUFF_1_9_r_3,N1372_10_r_6);
not I_53(n10_3,blif_reset_net_7_r_3);
not I_54(n30_3,n39_3);
not I_55(n31_3,n35_3);
nand I_56(n32_3,n41_3,N1508_0_r_6);
nor I_57(n33_3,I_BUFF_1_9_r_3,n34_3);
nand I_58(n34_3,n46_3,N1371_0_r_6);
nor I_59(n35_3,n43_3,n44_3);
not I_60(n36_3,n34_3);
nor I_61(n37_3,N6147_9_r_3,N1372_10_r_6);
or I_62(n38_3,n_572_7_r_3,n34_3);
nor I_63(n39_3,n44_3,N6134_9_r_6);
nand I_64(n40_3,n39_3,N1372_10_r_6);
nand I_65(n41_3,N1508_0_r_6,N6147_9_r_6);
nor I_66(n42_3,n34_3,n45_3);
not I_67(n43_3,N1372_1_r_6);
nor I_68(n44_3,N1371_0_r_6,G199_8_r_6);
nand I_69(n45_3,n49_3,n50_3);
and I_70(n46_3,n47_3,N1508_10_r_6);
nand I_71(n47_3,n41_3,n48_3);
not I_72(n48_3,N1508_0_r_6);
nor I_73(n49_3,N1372_1_r_6,N1507_6_r_6);
or I_74(n50_3,n51_3,N1508_6_r_6);
nor I_75(n51_3,N1508_1_r_6,n_42_8_r_6);
endmodule


