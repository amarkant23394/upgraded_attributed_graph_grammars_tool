module test_I7946(I1477,I1470,I3972,I7946);
input I1477,I1470,I3972;
output I7946;
wire I6606,I6300,I7881,I7570,I7587,I6329,I6688,I6705,I6291;
DFFARX1 I_0(I1470,I6329,,,I6606,);
DFFARX1 I_1(I6606,I1470,I6329,,,I6300,);
DFFARX1 I_2(I7881,I1470,I7570,,,I7946,);
nand I_3(I7881,I7587,I6291);
not I_4(I7570,I1477);
not I_5(I7587,I6300);
not I_6(I6329,I1477);
DFFARX1 I_7(I1470,I6329,,,I6688,);
and I_8(I6705,I6688,I3972);
DFFARX1 I_9(I6705,I1470,I6329,,,I6291,);
endmodule


