module test_I16795(I1477,I16886,I1470,I14954,I15310,I16795);
input I1477,I16886,I1470,I14954,I15310;
output I16795;
wire I14927,I17321,I14933,I17270,I17304,I17205,I17287,I17092,I16818,I14965,I17109;
DFFARX1 I_0(I1470,I14965,,,I14927,);
or I_1(I17321,I17109,I17304);
DFFARX1 I_2(I15310,I1470,I14965,,,I14933,);
not I_3(I17270,I17205);
and I_4(I17304,I17205,I17287);
DFFARX1 I_5(I14927,I1470,I16818,,,I17205,);
nor I_6(I17287,I16886,I17270);
DFFARX1 I_7(I14954,I1470,I16818,,,I17092,);
not I_8(I16818,I1477);
DFFARX1 I_9(I17321,I1470,I16818,,,I16795,);
not I_10(I14965,I1477);
and I_11(I17109,I17092,I14933);
endmodule


