module test_I9083(I5070,I5368,I7410,I7269,I5642,I6924,I9083);
input I5070,I5368,I7410,I7269,I5642,I6924;
output I9083;
wire I6992,I6975,I7427,I7317,I7026,I7057,I6881,I8879,I6887,I5097;
nand I_0(I6992,I6975,I5097);
nor I_1(I6975,I6924,I5070);
not I_2(I7427,I7410);
nor I_3(I7317,I7269,I7057);
not I_4(I7026,I5070);
not I_5(I7057,I7026);
nand I_6(I6881,I6992,I7057);
not I_7(I8879,I6887);
nand I_8(I6887,I7427,I7317);
nand I_9(I5097,I5642,I5368);
nand I_10(I9083,I8879,I6881);
endmodule


