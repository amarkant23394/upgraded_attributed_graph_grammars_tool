module test_I2793(I1351,I1319,I2793);
input I1351,I1319;
output I2793;
wire ;
nor I_0(I2793,I1351,I1319);
endmodule


