module test_final(G18_1_l_13,G15_1_l_13,IN_1_1_l_13,IN_4_1_l_13,IN_5_1_l_13,IN_7_1_l_13,IN_9_1_l_13,IN_10_1_l_13,IN_1_3_l_13,IN_2_3_l_13,IN_4_3_l_13,blif_clk_net_1_r_4,blif_reset_net_1_r_4,G42_1_r_4,n_572_1_r_4,n_573_1_r_4,n_549_1_r_4,n_569_1_r_4,ACVQN2_3_r_4,n_266_and_0_3_r_4,ACVQN1_5_r_4,P6_5_r_4);
input G18_1_l_13,G15_1_l_13,IN_1_1_l_13,IN_4_1_l_13,IN_5_1_l_13,IN_7_1_l_13,IN_9_1_l_13,IN_10_1_l_13,IN_1_3_l_13,IN_2_3_l_13,IN_4_3_l_13,blif_clk_net_1_r_4,blif_reset_net_1_r_4;
output G42_1_r_4,n_572_1_r_4,n_573_1_r_4,n_549_1_r_4,n_569_1_r_4,ACVQN2_3_r_4,n_266_and_0_3_r_4,ACVQN1_5_r_4,P6_5_r_4;
wire G42_1_r_13,n_572_1_r_13,n_573_1_r_13,n_549_1_r_13,n_569_1_r_13,n_452_1_r_13,ACVQN2_3_r_13,n_266_and_0_3_r_13,ACVQN1_5_r_13,P6_5_r_13,n4_1_l_13,n17_internal_13,n17_13,n28_13,ACVQN1_3_l_13,n4_1_r_13,n_266_and_0_3_l_13,n_573_1_l_13,n14_internal_13,n14_13,n_549_1_l_13,n_569_1_l_13,P6_5_r_internal_13,n18_13,n19_13,n20_13,n21_13,n22_13,n23_13,n24_13,n25_13,n26_13,n27_13,n_431_0_l_4,n6_4,G78_0_l_4,ACVQN1_5_l_4,n16_4,n17_internal_4,n17_4,n4_1_r_4,n19_4,n15_internal_4,n15_4,P6_5_r_internal_4,n20_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4;
DFFARX1 I_0(n4_1_r_13,blif_clk_net_1_r_4,n6_4,G42_1_r_13,);
nor I_1(n_572_1_r_13,n28_13,n_569_1_l_13);
nand I_2(n_573_1_r_13,n18_13,n19_13);
nand I_3(n_549_1_r_13,n_569_1_r_13,n22_13);
nand I_4(n_569_1_r_13,n17_13,n18_13);
nor I_5(n_452_1_r_13,n_573_1_l_13,n25_13);
DFFARX1 I_6(n_266_and_0_3_l_13,blif_clk_net_1_r_4,n6_4,ACVQN2_3_r_13,);
nor I_7(n_266_and_0_3_r_13,n17_13,n14_13);
DFFARX1 I_8(n_549_1_l_13,blif_clk_net_1_r_4,n6_4,ACVQN1_5_r_13,);
not I_9(P6_5_r_13,P6_5_r_internal_13);
nor I_10(n4_1_l_13,G18_1_l_13,IN_1_1_l_13);
DFFARX1 I_11(n4_1_l_13,blif_clk_net_1_r_4,n6_4,n17_internal_13,);
not I_12(n17_13,n17_internal_13);
DFFARX1 I_13(IN_1_3_l_13,blif_clk_net_1_r_4,n6_4,n28_13,);
DFFARX1 I_14(IN_2_3_l_13,blif_clk_net_1_r_4,n6_4,ACVQN1_3_l_13,);
nor I_15(n4_1_r_13,n_573_1_l_13,n_549_1_l_13);
and I_16(n_266_and_0_3_l_13,IN_4_3_l_13,ACVQN1_3_l_13);
nand I_17(n_573_1_l_13,n20_13,n24_13);
DFFARX1 I_18(n_573_1_l_13,blif_clk_net_1_r_4,n6_4,n14_internal_13,);
not I_19(n14_13,n14_internal_13);
and I_20(n_549_1_l_13,n21_13,n26_13);
nand I_21(n_569_1_l_13,n20_13,n21_13);
DFFARX1 I_22(n_569_1_l_13,blif_clk_net_1_r_4,n6_4,P6_5_r_internal_13,);
nand I_23(n18_13,n23_13,n24_13);
or I_24(n19_13,G15_1_l_13,IN_7_1_l_13);
not I_25(n20_13,IN_9_1_l_13);
not I_26(n21_13,IN_10_1_l_13);
nand I_27(n22_13,n17_13,n28_13);
not I_28(n23_13,G18_1_l_13);
not I_29(n24_13,IN_5_1_l_13);
nor I_30(n25_13,G15_1_l_13,IN_7_1_l_13);
nand I_31(n26_13,IN_4_1_l_13,n27_13);
not I_32(n27_13,G15_1_l_13);
DFFARX1 I_33(n4_1_r_4,blif_clk_net_1_r_4,n6_4,G42_1_r_4,);
nor I_34(n_572_1_r_4,G78_0_l_4,n17_4);
nand I_35(n_573_1_r_4,n16_4,n_452_1_r_13);
nor I_36(n_549_1_r_4,n22_4,n23_4);
nand I_37(n_569_1_r_4,n20_4,n21_4);
DFFARX1 I_38(n19_4,blif_clk_net_1_r_4,n6_4,ACVQN2_3_r_4,);
nor I_39(n_266_and_0_3_r_4,n15_4,n29_4);
DFFARX1 I_40(n19_4,blif_clk_net_1_r_4,n6_4,ACVQN1_5_r_4,);
not I_41(P6_5_r_4,P6_5_r_internal_4);
or I_42(n_431_0_l_4,n26_4,n_572_1_r_13);
not I_43(n6_4,blif_reset_net_1_r_4);
DFFARX1 I_44(n_431_0_l_4,blif_clk_net_1_r_4,n6_4,G78_0_l_4,);
DFFARX1 I_45(G42_1_r_13,blif_clk_net_1_r_4,n6_4,ACVQN1_5_l_4,);
not I_46(n16_4,ACVQN1_5_l_4);
DFFARX1 I_47(G42_1_r_13,blif_clk_net_1_r_4,n6_4,n17_internal_4,);
not I_48(n17_4,n17_internal_4);
nor I_49(n4_1_r_4,n30_4,n31_4);
nand I_50(n19_4,n33_4,n_549_1_r_13);
DFFARX1 I_51(G78_0_l_4,blif_clk_net_1_r_4,n6_4,n15_internal_4,);
not I_52(n15_4,n15_internal_4);
DFFARX1 I_53(ACVQN1_5_l_4,blif_clk_net_1_r_4,n6_4,P6_5_r_internal_4,);
and I_54(n20_4,n16_4,n_572_1_r_13);
nor I_55(n21_4,n_452_1_r_13,ACVQN2_3_r_13);
nand I_56(n22_4,G78_0_l_4,n25_4);
nand I_57(n23_4,n24_4,n_572_1_r_13);
not I_58(n24_4,n_452_1_r_13);
not I_59(n25_4,ACVQN2_3_r_13);
and I_60(n26_4,n27_4,P6_5_r_13);
nor I_61(n27_4,n28_4,n_573_1_r_13);
not I_62(n28_4,n_549_1_r_13);
not I_63(n29_4,n30_4);
nand I_64(n30_4,n32_4,n_266_and_0_3_r_13);
nand I_65(n31_4,n25_4,n_572_1_r_13);
nor I_66(n32_4,n33_4,n_452_1_r_13);
not I_67(n33_4,ACVQN1_5_r_13);
endmodule


