module test_I3589(I1477,I1849,I1492,I2038,I1976,I1470,I3589);
input I1477,I1849,I1492,I2038,I1976,I1470;
output I3589;
wire I1486,I1801,I3521,I3504,I1495,I3538,I3487,I3388,I3405,I1489,I1510,I3572,I1518,I1480,I3555,I2103;
DFFARX1 I_0(I1470,I1518,,,I1486,);
DFFARX1 I_1(I1470,I1518,,,I1801,);
nor I_2(I3521,I3504,I1495);
and I_3(I3504,I3487,I1489);
DFFARX1 I_4(I2103,I1470,I1518,,,I1495,);
nor I_5(I3538,I1492,I1510);
not I_6(I3487,I1486);
not I_7(I3388,I1477);
or I_8(I3405,I1480,I1495);
not I_9(I1489,I1801);
DFFARX1 I_10(I1470,I1518,,,I1510,);
nand I_11(I3572,I3555,I3405);
not I_12(I1518,I1477);
DFFARX1 I_13(I1976,I1470,I1518,,,I1480,);
and I_14(I3589,I3521,I3572);
DFFARX1 I_15(I3538,I1470,I3388,,,I3555,);
or I_16(I2103,I2038,I1849);
endmodule


