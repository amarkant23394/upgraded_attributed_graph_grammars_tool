module test_I1498(I1477,I1295,I1215,I1470,I1383,I1498);
input I1477,I1295,I1215,I1470,I1383;
output I1498;
wire I1518,I1668,I1637,I1928,I2038,I2021,I1880;
not I_0(I1518,I1477);
not I_1(I1668,I1637);
not I_2(I1637,I1215);
nor I_3(I1928,I1880,I1668);
not I_4(I2038,I2021);
DFFARX1 I_5(I1295,I1470,I1518,,,I2021,);
DFFARX1 I_6(I1383,I1470,I1518,,,I1880,);
nand I_7(I1498,I2038,I1928);
endmodule


