module test_I3234(I1351,I1319,I1431,I1477,I1470,I1335,I3234);
input I1351,I1319,I1431,I1477,I1470,I1335;
output I3234;
wire I3217,I2810,I2759,I3200,I2793;
not I_0(I3217,I3200);
nand I_1(I2810,I2793,I1335);
not I_2(I2759,I1477);
nor I_3(I3234,I3217,I2810);
DFFARX1 I_4(I1431,I1470,I2759,,,I3200,);
nor I_5(I2793,I1351,I1319);
endmodule


