module test_I1988(I1444,I1560,I1215,I1294,I1639,I1301,I1988);
input I1444,I1560,I1215,I1294,I1639,I1301;
output I1988;
wire I1319,I1749,I1656,I1971,I1342,I1334,I1797,I1509,I1310,I1577,I1780;
DFFARX1 I_0(I1749,I1294,I1342,,,I1319,);
or I_1(I1749,I1639,I1560);
nand I_2(I1656,I1639,I1509);
nor I_3(I1971,I1310,I1319);
not I_4(I1342,I1301);
DFFARX1 I_5(I1797,I1294,I1342,,,I1334,);
nand I_6(I1988,I1971,I1334);
and I_7(I1797,I1780,I1656);
DFFARX1 I_8(I1294,I1342,,,I1509,);
DFFARX1 I_9(I1577,I1294,I1342,,,I1310,);
and I_10(I1577,I1509,I1444);
DFFARX1 I_11(I1215,I1294,I1342,,,I1780,);
endmodule


