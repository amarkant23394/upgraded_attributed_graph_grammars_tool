module test_final(IN_1_1_l_16,IN_2_1_l_16,IN_3_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_3_3_l_16,IN_1_6_l_16,IN_2_6_l_16,IN_3_6_l_16,IN_4_6_l_16,IN_5_6_l_16,IN_1_8_l_16,IN_2_8_l_16,IN_3_8_l_16,IN_6_8_l_16,blif_clk_net_7_r_2,blif_reset_net_7_r_2,N1371_0_r_2,N1508_0_r_2,N1372_1_r_2,N1508_1_r_2,N6147_2_r_2,N1507_6_r_2,N1508_6_r_2,G42_7_r_2,n_572_7_r_2,n_573_7_r_2,n_549_7_r_2,n_569_7_r_2,n_452_7_r_2);
input IN_1_1_l_16,IN_2_1_l_16,IN_3_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_3_3_l_16,IN_1_6_l_16,IN_2_6_l_16,IN_3_6_l_16,IN_4_6_l_16,IN_5_6_l_16,IN_1_8_l_16,IN_2_8_l_16,IN_3_8_l_16,IN_6_8_l_16,blif_clk_net_7_r_2,blif_reset_net_7_r_2;
output N1371_0_r_2,N1508_0_r_2,N1372_1_r_2,N1508_1_r_2,N6147_2_r_2,N1507_6_r_2,N1508_6_r_2,G42_7_r_2,n_572_7_r_2,n_573_7_r_2,n_549_7_r_2,n_569_7_r_2,n_452_7_r_2;
wire N1371_0_r_16,N1508_0_r_16,N1372_1_r_16,N1508_1_r_16,N6147_2_r_16,N1507_6_r_16,N1508_6_r_16,G42_7_r_16,n_572_7_r_16,n_573_7_r_16,n_549_7_r_16,n_569_7_r_16,n_452_7_r_16,N3_8_l_16,n53_16,n29_16,n4_7_r_16,n30_16,n31_16,n32_16,n33_16,n34_16,n35_16,n36_16,n37_16,n38_16,n39_16,n40_16,n41_16,n42_16,n43_16,n44_16,n45_16,n46_16,n47_16,n48_16,n49_16,n50_16,n51_16,n52_16,n4_7_l_2,n10_2,n59_2,n33_2,N3_8_l_2,n32_internal_2,n32_2,n4_7_r_2,n34_2,n35_2,n36_2,n37_2,n38_2,n39_2,n40_2,n41_2,n42_2,n43_2,n44_2,n45_2,n46_2,n47_2,n48_2,n49_2,n50_2,n51_2,n52_2,n53_2,n54_2,n55_2,n56_2,n57_2,n58_2;
nor I_0(N1371_0_r_16,n35_16,n39_16);
nor I_1(N1508_0_r_16,n39_16,n46_16);
not I_2(N1372_1_r_16,n45_16);
nor I_3(N1508_1_r_16,n53_16,n45_16);
nor I_4(N6147_2_r_16,n37_16,n38_16);
nor I_5(N1507_6_r_16,n44_16,n49_16);
nor I_6(N1508_6_r_16,n29_16,n42_16);
DFFARX1 I_7(n4_7_r_16,blif_clk_net_7_r_2,n10_2,G42_7_r_16,);
nor I_8(n_572_7_r_16,n32_16,n33_16);
nand I_9(n_573_7_r_16,n30_16,n31_16);
nand I_10(n_549_7_r_16,IN_5_6_l_16,n47_16);
nand I_11(n_569_7_r_16,n_549_7_r_16,n30_16);
nor I_12(n_452_7_r_16,n34_16,n35_16);
and I_13(N3_8_l_16,IN_6_8_l_16,n41_16);
DFFARX1 I_14(N3_8_l_16,blif_clk_net_7_r_2,n10_2,n53_16,);
not I_15(n29_16,n53_16);
nor I_16(n4_7_r_16,n35_16,n36_16);
nand I_17(n30_16,IN_1_1_l_16,IN_2_1_l_16);
not I_18(n31_16,n34_16);
nor I_19(n32_16,IN_3_1_l_16,n30_16);
not I_20(n33_16,n_549_7_r_16);
nor I_21(n34_16,IN_1_3_l_16,n48_16);
and I_22(n35_16,IN_2_6_l_16,n50_16);
not I_23(n36_16,n30_16);
nor I_24(n37_16,n31_16,n40_16);
nand I_25(n38_16,n29_16,n39_16);
not I_26(n39_16,n32_16);
nor I_27(n40_16,IN_1_8_l_16,IN_3_8_l_16);
nand I_28(n41_16,IN_2_8_l_16,IN_3_8_l_16);
nand I_29(n42_16,n35_16,n43_16);
not I_30(n43_16,n44_16);
nor I_31(n44_16,n32_16,n49_16);
nand I_32(n45_16,n36_16,n40_16);
nor I_33(n46_16,n33_16,n34_16);
nand I_34(n47_16,IN_3_6_l_16,IN_4_6_l_16);
or I_35(n48_16,IN_2_3_l_16,IN_3_3_l_16);
and I_36(n49_16,n35_16,n36_16);
and I_37(n50_16,IN_1_6_l_16,n51_16);
nand I_38(n51_16,n47_16,n52_16);
not I_39(n52_16,IN_5_6_l_16);
nor I_40(N1371_0_r_2,n32_2,n35_2);
nor I_41(N1508_0_r_2,n32_2,n55_2);
not I_42(N1372_1_r_2,n54_2);
nor I_43(N1508_1_r_2,n59_2,n54_2);
nor I_44(N6147_2_r_2,n42_2,n43_2);
nor I_45(N1507_6_r_2,n40_2,n53_2);
nor I_46(N1508_6_r_2,n33_2,n50_2);
DFFARX1 I_47(n4_7_r_2,blif_clk_net_7_r_2,n10_2,G42_7_r_2,);
nor I_48(n_572_7_r_2,n36_2,n37_2);
or I_49(n_573_7_r_2,n34_2,n35_2);
nor I_50(n_549_7_r_2,n40_2,n41_2);
nand I_51(n_569_7_r_2,n38_2,n39_2);
nor I_52(n_452_7_r_2,n59_2,n35_2);
nor I_53(n4_7_l_2,G42_7_r_16,n_452_7_r_16);
not I_54(n10_2,blif_reset_net_7_r_2);
DFFARX1 I_55(n4_7_l_2,blif_clk_net_7_r_2,n10_2,n59_2,);
not I_56(n33_2,n59_2);
and I_57(N3_8_l_2,n49_2,N6147_2_r_16);
DFFARX1 I_58(N3_8_l_2,blif_clk_net_7_r_2,n10_2,n32_internal_2,);
not I_59(n32_2,n32_internal_2);
nor I_60(n4_7_r_2,n59_2,n36_2);
not I_61(n34_2,n39_2);
nor I_62(n35_2,N1508_0_r_16,N1508_6_r_16);
nor I_63(n36_2,N1508_1_r_16,G42_7_r_16);
or I_64(n37_2,N1371_0_r_16,N1508_0_r_16);
not I_65(n38_2,n40_2);
nand I_66(n39_2,n45_2,n57_2);
nor I_67(n40_2,n47_2,n_569_7_r_16);
nor I_68(n41_2,n32_2,n36_2);
not I_69(n42_2,n53_2);
nand I_70(n43_2,n44_2,n45_2);
nand I_71(n44_2,n38_2,n46_2);
not I_72(n45_2,N1371_0_r_16);
nand I_73(n46_2,n47_2,n48_2);
nand I_74(n47_2,N1372_1_r_16,N1507_6_r_16);
or I_75(n48_2,n_572_7_r_16,N1372_1_r_16);
nand I_76(n49_2,N1508_6_r_16,N1508_1_r_16);
nand I_77(n50_2,n51_2,n52_2);
not I_78(n51_2,n47_2);
nand I_79(n52_2,n38_2,n53_2);
nor I_80(n53_2,N1508_1_r_16,N1508_0_r_16);
nand I_81(n54_2,n42_2,n56_2);
nor I_82(n55_2,n34_2,n56_2);
nor I_83(n56_2,n_572_7_r_16,N1372_1_r_16);
nand I_84(n57_2,n58_2,n_573_7_r_16);
not I_85(n58_2,N1372_1_r_16);
endmodule


