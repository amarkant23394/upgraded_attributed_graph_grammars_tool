module test_I14965_rst(I1477_rst,I14965_rst);
,I14965_rst);
input I1477_rst;
output I14965_rst;
wire ;
not I_0(I14965_rst,I1477_rst);
endmodule


