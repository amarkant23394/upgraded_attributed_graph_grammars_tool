module test_I13392(I1477,I11576,I9083,I1470,I11327,I13392);
input I1477,I11576,I9083,I1470,I11327;
output I13392;
wire I11641,I11830,I11395,I11624,I11287,I11895,I8848,I11378,I11429,I9066,I11813,I11284,I11310,I11460,I8851;
and I_0(I11641,I11624,I11576);
not I_1(I11830,I11813);
nand I_2(I11395,I11378,I8851);
nand I_3(I11624,I11327);
DFFARX1 I_4(I11895,I1470,I11310,,,I11287,);
or I_5(I11895,I11830,I11641);
nor I_6(I8848,I9083);
nand I_7(I13392,I11287,I11284);
nor I_8(I11378,I11327,I8848);
not I_9(I11429,I8848);
DFFARX1 I_10(I1470,,,I9066,);
DFFARX1 I_11(I1470,I11310,,,I11813,);
nand I_12(I11284,I11395,I11460);
not I_13(I11310,I1477);
not I_14(I11460,I11429);
or I_15(I8851,I9083,I9066);
endmodule


