module test_I6893(I5266,I7105,I1477,I5368,I5070,I5642,I6924,I1470,I6893);
input I5266,I7105,I1477,I5368,I5070,I5642,I6924,I1470;
output I6893;
wire I7122,I5085,I5067,I6907,I5512,I5097,I7139,I5076,I6975,I7269,I6992,I5105,I7286,I7156;
and I_0(I7122,I7105,I5076);
nand I_1(I6893,I7156,I7286);
nand I_2(I5085,I5512,I5266);
DFFARX1 I_3(I5642,I1470,I5105,,,I5067,);
not I_4(I6907,I1477);
DFFARX1 I_5(I1470,I5105,,,I5512,);
nand I_6(I5097,I5642,I5368);
or I_7(I7139,I7122,I5085);
DFFARX1 I_8(I1470,I5105,,,I5076,);
nor I_9(I6975,I6924,I5070);
DFFARX1 I_10(I5067,I1470,I6907,,,I7269,);
nand I_11(I6992,I6975,I5097);
not I_12(I5105,I1477);
nor I_13(I7286,I7269,I6992);
DFFARX1 I_14(I7139,I1470,I6907,,,I7156,);
endmodule


