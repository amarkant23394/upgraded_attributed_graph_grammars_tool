module test_final(IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_4_2_l_6,IN_5_2_l_6,IN_1_6_l_6,IN_2_6_l_6,IN_3_6_l_6,IN_4_6_l_6,IN_5_6_l_6,IN_1_9_l_6,IN_2_9_l_6,IN_3_9_l_6,IN_4_9_l_6,IN_5_9_l_6,blif_clk_net_7_r_5,blif_reset_net_7_r_5,N1371_0_r_5,N1508_0_r_5,N1372_1_r_5,N1508_1_r_5,N6147_2_r_5,N1507_6_r_5,N1508_6_r_5,G42_7_r_5,n_572_7_r_5,n_573_7_r_5,n_569_7_r_5,n_452_7_r_5);
input IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_4_2_l_6,IN_5_2_l_6,IN_1_6_l_6,IN_2_6_l_6,IN_3_6_l_6,IN_4_6_l_6,IN_5_6_l_6,IN_1_9_l_6,IN_2_9_l_6,IN_3_9_l_6,IN_4_9_l_6,IN_5_9_l_6,blif_clk_net_7_r_5,blif_reset_net_7_r_5;
output N1371_0_r_5,N1508_0_r_5,N1372_1_r_5,N1508_1_r_5,N6147_2_r_5,N1507_6_r_5,N1508_6_r_5,G42_7_r_5,n_572_7_r_5,n_573_7_r_5,n_569_7_r_5,n_452_7_r_5;
wire N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,I_BUFF_1_9_r_6,N1372_10_r_6,N1508_10_r_6,N3_8_r_6,n30_6,n31_6,n32_6,n33_6,n34_6,n35_6,n36_6,n37_6,n38_6,n39_6,n40_6,n41_6,n42_6,n43_6,n44_6,n45_6,n46_6,n47_6,n48_6,n49_6,n50_6,n51_6,n52_6,n53_6,n54_6,n_549_7_r_5,n4_7_r_5,n7_5,n26_5,n27_5,n28_5,n29_5,n30_5,n31_5,n32_5,n33_5,n34_5,n35_5,n36_5,n37_5,n38_5,n39_5,n40_5,n41_5,n42_5,n43_5,n44_5,n45_5,n46_5,n47_5;
nor I_0(N1371_0_r_6,n30_6,n33_6);
nor I_1(N1508_0_r_6,n33_6,n44_6);
not I_2(N1372_1_r_6,n41_6);
nor I_3(N1508_1_r_6,n40_6,n41_6);
nor I_4(N1507_6_r_6,n39_6,n45_6);
nor I_5(N1508_6_r_6,n37_6,n38_6);
nor I_6(n_42_8_r_6,n30_6,n31_6);
DFFARX1 I_7(N3_8_r_6,blif_clk_net_7_r_5,n7_5,G199_8_r_6,);
nor I_8(N6147_9_r_6,n32_6,n33_6);
nor I_9(N6134_9_r_6,I_BUFF_1_9_r_6,n35_6);
not I_10(I_BUFF_1_9_r_6,n37_6);
not I_11(N1372_10_r_6,n43_6);
nor I_12(N1508_10_r_6,n42_6,n43_6);
nor I_13(N3_8_r_6,IN_1_9_l_6,n36_6);
nor I_14(n30_6,IN_5_9_l_6,n53_6);
not I_15(n31_6,n36_6);
nor I_16(n32_6,I_BUFF_1_9_r_6,n34_6);
not I_17(n33_6,IN_1_9_l_6);
not I_18(n34_6,n35_6);
nand I_19(n35_6,IN_2_6_l_6,n49_6);
nand I_20(n36_6,IN_5_6_l_6,n51_6);
nand I_21(n37_6,IN_2_9_l_6,n54_6);
or I_22(n38_6,n35_6,n39_6);
nor I_23(n39_6,n40_6,n45_6);
and I_24(n40_6,n46_6,n47_6);
nand I_25(n41_6,n30_6,n31_6);
nor I_26(n42_6,n34_6,n40_6);
nand I_27(n43_6,IN_1_9_l_6,n30_6);
nor I_28(n44_6,n31_6,n40_6);
nor I_29(n45_6,n35_6,n36_6);
nor I_30(n46_6,IN_1_2_l_6,IN_2_2_l_6);
or I_31(n47_6,IN_5_2_l_6,n48_6);
nor I_32(n48_6,IN_3_2_l_6,IN_4_2_l_6);
and I_33(n49_6,IN_1_6_l_6,n50_6);
nand I_34(n50_6,n51_6,n52_6);
nand I_35(n51_6,IN_3_6_l_6,IN_4_6_l_6);
not I_36(n52_6,IN_5_6_l_6);
nor I_37(n53_6,IN_3_9_l_6,IN_4_9_l_6);
or I_38(n54_6,IN_3_9_l_6,IN_4_9_l_6);
nor I_39(N1371_0_r_5,n28_5,n46_5);
nand I_40(N1508_0_r_5,n26_5,n43_5);
not I_41(N1372_1_r_5,n43_5);
nor I_42(N1508_1_r_5,n30_5,n43_5);
nor I_43(N6147_2_r_5,n29_5,n32_5);
nor I_44(N1507_6_r_5,n26_5,n44_5);
nor I_45(N1508_6_r_5,n27_5,n37_5);
DFFARX1 I_46(n4_7_r_5,blif_clk_net_7_r_5,n7_5,G42_7_r_5,);
and I_47(n_572_7_r_5,n27_5,n28_5);
nand I_48(n_573_7_r_5,n26_5,n27_5);
nand I_49(n_549_7_r_5,N1372_10_r_6,N1508_0_r_6);
nand I_50(n_569_7_r_5,n_549_7_r_5,n26_5);
not I_51(n_452_7_r_5,n29_5);
nor I_52(n4_7_r_5,n30_5,n31_5);
not I_53(n7_5,blif_reset_net_7_r_5);
not I_54(n26_5,n35_5);
nand I_55(n27_5,n40_5,n41_5);
nand I_56(n28_5,N1508_6_r_6,n_42_8_r_6);
nand I_57(n29_5,n27_5,n33_5);
nor I_58(n30_5,n45_5,N1371_0_r_6);
not I_59(n31_5,n_549_7_r_5);
nor I_60(n32_5,n34_5,n35_5);
not I_61(n33_5,n30_5);
nor I_62(n34_5,n31_5,n36_5);
nor I_63(n35_5,n28_5,N1372_1_r_6);
not I_64(n36_5,n28_5);
nand I_65(n37_5,n36_5,n38_5);
nand I_66(n38_5,n26_5,n39_5);
nand I_67(n39_5,n30_5,n31_5);
nor I_68(n40_5,N1508_1_r_6,N1507_6_r_6);
or I_69(n41_5,n42_5,N1508_0_r_6);
nor I_70(n42_5,G199_8_r_6,N6147_9_r_6);
nand I_71(n43_5,n36_5,n46_5);
nor I_72(n44_5,n_549_7_r_5,n33_5);
or I_73(n45_5,N1371_0_r_6,N1508_10_r_6);
and I_74(n46_5,n31_5,n47_5);
or I_75(n47_5,N1372_1_r_6,N6134_9_r_6);
endmodule


