module test_I16214(I1477,I1470,I16435,I16214);
input I1477,I1470,I16435;
output I16214;
wire I14338,I14362,I16452,I16257,I14341,I16291,I16469,I16240,I16274,I16503,I14537,I14370,I14332;
DFFARX1 I_0(I1470,I14370,,,I14338,);
DFFARX1 I_1(I1470,I14370,,,I14362,);
nand I_2(I16214,I16291,I16503);
and I_3(I16452,I16435,I14362);
nand I_4(I16257,I14341,I14338);
DFFARX1 I_5(I1470,I14370,,,I14341,);
DFFARX1 I_6(I16274,I1470,I16240,,,I16291,);
DFFARX1 I_7(I16452,I1470,I16240,,,I16469,);
not I_8(I16240,I1477);
and I_9(I16274,I16257,I14332);
not I_10(I16503,I16469);
DFFARX1 I_11(I1470,I14370,,,I14537,);
not I_12(I14370,I1477);
DFFARX1 I_13(I14537,I1470,I14370,,,I14332,);
endmodule


