module test_I2912(I1415,I1311,I2912);
input I1415,I1311;
output I2912;
wire I2895;
nor I_0(I2912,I2895,I1311);
not I_1(I2895,I1415);
endmodule


