module test_I7105(I1477,I3380,I1470,I5563,I3815,I5642,I7105);
input I1477,I3380,I1470,I5563,I3815,I5642;
output I7105;
wire I5659,I5156,I3388,I5079,I3359,I3371,I5088,I5139,I7088,I5105;
or I_0(I5659,I5642,I5563);
nand I_1(I5156,I5139,I3371);
not I_2(I3388,I1477);
DFFARX1 I_3(I5156,I1470,I5105,,,I5079,);
nor I_4(I7105,I7088,I5079);
DFFARX1 I_5(I1470,I3388,,,I3359,);
DFFARX1 I_6(I3815,I1470,I3388,,,I3371,);
DFFARX1 I_7(I5659,I1470,I5105,,,I5088,);
nor I_8(I5139,I3380,I3359);
not I_9(I7088,I5088);
not I_10(I5105,I1477);
endmodule


