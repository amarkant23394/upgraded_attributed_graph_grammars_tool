module test_final(G18_1_l_3,G15_1_l_3,IN_1_1_l_3,IN_4_1_l_3,IN_5_1_l_3,IN_7_1_l_3,IN_9_1_l_3,IN_10_1_l_3,IN_1_3_l_3,IN_2_3_l_3,IN_4_3_l_3,blif_clk_net_1_r_15,blif_reset_net_1_r_15,G42_1_r_15,n_572_1_r_15,n_573_1_r_15,n_549_1_r_15,n_569_1_r_15,ACVQN2_3_r_15,n_266_and_0_3_r_15,G199_4_r_15,G214_4_r_15);
input G18_1_l_3,G15_1_l_3,IN_1_1_l_3,IN_4_1_l_3,IN_5_1_l_3,IN_7_1_l_3,IN_9_1_l_3,IN_10_1_l_3,IN_1_3_l_3,IN_2_3_l_3,IN_4_3_l_3,blif_clk_net_1_r_15,blif_reset_net_1_r_15;
output G42_1_r_15,n_572_1_r_15,n_573_1_r_15,n_549_1_r_15,n_569_1_r_15,ACVQN2_3_r_15,n_266_and_0_3_r_15,G199_4_r_15,G214_4_r_15;
wire G42_1_r_3,n_572_1_r_3,n_573_1_r_3,n_549_1_r_3,n_569_1_r_3,n_452_1_r_3,n_42_2_r_3,G199_2_r_3,ACVQN2_3_r_3,n_266_and_0_3_r_3,n4_1_l_3,G42_1_l_3,n22_3,n40_3,n25_internal_3,n25_3,n4_1_r_3,N3_2_r_3,n_572_1_l_3,ACVQN1_3_r_3,n26_3,n27_3,n28_3,n29_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3,n_452_1_r_15,n4_1_l_15,n4_15,G42_1_l_15,n15_15,n17_internal_15,n17_15,n30_15,n_572_1_l_15,n14_internal_15,n14_15,N1_4_r_15,n_573_1_l_15,n18_15,n19_15,n20_15,n21_15,n22_15,n23_15,n24_15,n25_15,n26_15,n27_15,n28_15,n29_15;
DFFARX1 I_0(n4_1_r_3,blif_clk_net_1_r_15,n4_15,G42_1_r_3,);
nor I_1(n_572_1_r_3,G42_1_l_3,n28_3);
nand I_2(n_573_1_r_3,n26_3,n27_3);
nor I_3(n_549_1_r_3,n40_3,n32_3);
nand I_4(n_569_1_r_3,n27_3,n31_3);
and I_5(n_452_1_r_3,G18_1_l_3,n26_3);
nor I_6(n_42_2_r_3,n_572_1_l_3,n34_3);
DFFARX1 I_7(N3_2_r_3,blif_clk_net_1_r_15,n4_15,G199_2_r_3,);
DFFARX1 I_8(n_572_1_l_3,blif_clk_net_1_r_15,n4_15,ACVQN2_3_r_3,);
nor I_9(n_266_and_0_3_r_3,n25_3,n35_3);
nor I_10(n4_1_l_3,G18_1_l_3,IN_1_1_l_3);
DFFARX1 I_11(n4_1_l_3,blif_clk_net_1_r_15,n4_15,G42_1_l_3,);
not I_12(n22_3,G42_1_l_3);
DFFARX1 I_13(IN_1_3_l_3,blif_clk_net_1_r_15,n4_15,n40_3,);
DFFARX1 I_14(IN_2_3_l_3,blif_clk_net_1_r_15,n4_15,n25_internal_3,);
not I_15(n25_3,n25_internal_3);
nor I_16(n4_1_r_3,n40_3,n36_3);
nor I_17(N3_2_r_3,n26_3,n37_3);
nor I_18(n_572_1_l_3,G15_1_l_3,IN_7_1_l_3);
DFFARX1 I_19(G42_1_l_3,blif_clk_net_1_r_15,n4_15,ACVQN1_3_r_3,);
nor I_20(n26_3,IN_5_1_l_3,IN_9_1_l_3);
not I_21(n27_3,IN_10_1_l_3);
nor I_22(n28_3,IN_10_1_l_3,n29_3);
nor I_23(n29_3,G15_1_l_3,n30_3);
not I_24(n30_3,IN_4_1_l_3);
nor I_25(n31_3,IN_9_1_l_3,n40_3);
nor I_26(n32_3,n25_3,n33_3);
nand I_27(n33_3,IN_4_3_l_3,n22_3);
or I_28(n34_3,IN_9_1_l_3,IN_10_1_l_3);
nand I_29(n35_3,IN_4_3_l_3,ACVQN1_3_r_3);
nor I_30(n36_3,G18_1_l_3,IN_5_1_l_3);
nor I_31(n37_3,n38_3,n39_3);
not I_32(n38_3,n_572_1_l_3);
nand I_33(n39_3,n27_3,n30_3);
DFFARX1 I_34(n_452_1_r_15,blif_clk_net_1_r_15,n4_15,G42_1_r_15,);
and I_35(n_572_1_r_15,n17_15,n19_15);
nand I_36(n_573_1_r_15,n15_15,n18_15);
nor I_37(n_549_1_r_15,n21_15,n22_15);
nand I_38(n_569_1_r_15,n15_15,n20_15);
nor I_39(n_452_1_r_15,n23_15,n24_15);
DFFARX1 I_40(G42_1_l_15,blif_clk_net_1_r_15,n4_15,ACVQN2_3_r_15,);
nor I_41(n_266_and_0_3_r_15,n17_15,n14_15);
DFFARX1 I_42(N1_4_r_15,blif_clk_net_1_r_15,n4_15,G199_4_r_15,);
DFFARX1 I_43(n_573_1_l_15,blif_clk_net_1_r_15,n4_15,G214_4_r_15,);
nor I_44(n4_1_l_15,G42_1_r_3,n_42_2_r_3);
not I_45(n4_15,blif_reset_net_1_r_15);
DFFARX1 I_46(n4_1_l_15,blif_clk_net_1_r_15,n4_15,G42_1_l_15,);
not I_47(n15_15,G42_1_l_15);
DFFARX1 I_48(n_573_1_r_3,blif_clk_net_1_r_15,n4_15,n17_internal_15,);
not I_49(n17_15,n17_internal_15);
DFFARX1 I_50(n_452_1_r_3,blif_clk_net_1_r_15,n4_15,n30_15,);
nor I_51(n_572_1_l_15,n_572_1_r_3,n_266_and_0_3_r_3);
DFFARX1 I_52(n_572_1_l_15,blif_clk_net_1_r_15,n4_15,n14_internal_15,);
not I_53(n14_15,n14_internal_15);
nand I_54(N1_4_r_15,n25_15,n26_15);
or I_55(n_573_1_l_15,n_549_1_r_3,G199_2_r_3);
nor I_56(n18_15,n_569_1_r_3,G199_2_r_3);
nand I_57(n19_15,n27_15,n28_15);
nand I_58(n20_15,n30_15,ACVQN2_3_r_3);
not I_59(n21_15,n20_15);
and I_60(n22_15,n17_15,n_572_1_l_15);
nor I_61(n23_15,n_549_1_r_3,n_42_2_r_3);
or I_62(n24_15,n_569_1_r_3,G199_2_r_3);
or I_63(n25_15,n_573_1_l_15,n_42_2_r_3);
nand I_64(n26_15,n19_15,n23_15);
not I_65(n27_15,n_569_1_r_3);
nand I_66(n28_15,n29_15,G42_1_r_3);
not I_67(n29_15,n_266_and_0_3_r_3);
endmodule


