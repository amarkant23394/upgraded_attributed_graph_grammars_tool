module Benchmark_testing45000(I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1804,I1812,I1820,I1828,I1836,I1844,I1852,I1860,I1868,I1876,I1884,I1892,I1900,I1908,I1916,I1924,I1932,I1940,I1948,I1956,I1964,I1972,I1980,I1988,I1996,I2004,I2012,I2020,I2028,I2036,I2044,I2052,I2060,I2068,I2076,I2084,I2092,I2100,I2108,I2116,I2124,I2132,I2140,I2148,I2156,I2164,I2172,I2180,I2188,I2196,I2204,I2212,I2220,I2228,I2236,I2244,I2252,I2260,I2268,I2276,I2284,I2292,I2300,I2308,I2316,I2324,I2332,I2340,I2348,I2356,I2364,I2372,I2380,I2388,I2396,I2404,I2412,I2420,I2428,I2436,I2444,I2452,I2460,I2468,I2476,I2484,I2492,I2500,I2508,I2516,I2524,I2532,I2540,I2548,I2556,I2564,I2572,I2580,I2588,I2596,I2604,I2612,I2620,I2628,I2636,I2644,I2652,I2660,I2668,I2676,I2684,I2692,I2700,I2708,I2716,I2724,I2732,I2740,I2748,I2756,I2764,I2772,I2780,I2788,I2796,I2804,I2812,I2820,I2828,I2836,I2844,I2852,I2860,I2868,I2876,I2884,I2892,I2900,I2908,I2916,I2924,I2932,I2940,I2948,I2956,I2964,I2972,I2980,I2988,I2996,I3004,I3012,I3020,I3028,I3035,I3042,I124143,I124119,I124131,I124125,I124140,I124134,I124128,I124122,I124137,I170855,I170879,I170861,I170864,I170852,I170870,I170873,I170858,I170867,I170876,I184557,I184581,I184563,I184566,I184554,I184572,I184575,I184560,I184569,I184578,I191408,I191432,I191414,I191417,I191405,I191423,I191426,I191411,I191420,I191429,I216704,I216728,I216710,I216713,I216701,I216719,I216722,I216707,I216716,I216725,I241888,I241867,I241861,I241876,I241864,I241879,I241870,I241873,I241885,I241882,I247872,I247851,I247845,I247860,I247848,I247863,I247854,I247857,I247869,I247866,I254400,I254379,I254373,I254388,I254376,I254391,I254382,I254385,I254397,I254394,I392071,I392074,I392056,I392065,I392077,I392068,I392059,I392062,I392080,I414035,I414038,I414020,I414029,I414041,I414032,I414023,I414026,I414044,I432466,I432469,I432460,I432451,I432454,I432463,I432448,I432457,I447222,I447225,I447216,I447207,I447210,I447219,I447204,I447213,I489657,I489660,I489636,I489648,I489663,I489651,I489645,I489639,I489642,I489654,I494825,I494828,I494804,I494816,I494831,I494819,I494813,I494807,I494810,I494822,I557725,I557707,I557710,I557719,I557722,I557716,I557704,I557713,I571750,I571732,I571735,I571744,I571747,I571741,I571729,I571738,I608719,I608707,I608728,I608704,I608725,I608716,I608722,I608713,I608710,I631839,I631827,I631848,I631824,I631845,I631836,I631842,I631833,I631830,I700201,I700216,I700198,I700210,I700225,I700222,I700219,I700213,I700207,I700204);
input I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1804,I1812,I1820,I1828,I1836,I1844,I1852,I1860,I1868,I1876,I1884,I1892,I1900,I1908,I1916,I1924,I1932,I1940,I1948,I1956,I1964,I1972,I1980,I1988,I1996,I2004,I2012,I2020,I2028,I2036,I2044,I2052,I2060,I2068,I2076,I2084,I2092,I2100,I2108,I2116,I2124,I2132,I2140,I2148,I2156,I2164,I2172,I2180,I2188,I2196,I2204,I2212,I2220,I2228,I2236,I2244,I2252,I2260,I2268,I2276,I2284,I2292,I2300,I2308,I2316,I2324,I2332,I2340,I2348,I2356,I2364,I2372,I2380,I2388,I2396,I2404,I2412,I2420,I2428,I2436,I2444,I2452,I2460,I2468,I2476,I2484,I2492,I2500,I2508,I2516,I2524,I2532,I2540,I2548,I2556,I2564,I2572,I2580,I2588,I2596,I2604,I2612,I2620,I2628,I2636,I2644,I2652,I2660,I2668,I2676,I2684,I2692,I2700,I2708,I2716,I2724,I2732,I2740,I2748,I2756,I2764,I2772,I2780,I2788,I2796,I2804,I2812,I2820,I2828,I2836,I2844,I2852,I2860,I2868,I2876,I2884,I2892,I2900,I2908,I2916,I2924,I2932,I2940,I2948,I2956,I2964,I2972,I2980,I2988,I2996,I3004,I3012,I3020,I3028,I3035,I3042;
output I124143,I124119,I124131,I124125,I124140,I124134,I124128,I124122,I124137,I170855,I170879,I170861,I170864,I170852,I170870,I170873,I170858,I170867,I170876,I184557,I184581,I184563,I184566,I184554,I184572,I184575,I184560,I184569,I184578,I191408,I191432,I191414,I191417,I191405,I191423,I191426,I191411,I191420,I191429,I216704,I216728,I216710,I216713,I216701,I216719,I216722,I216707,I216716,I216725,I241888,I241867,I241861,I241876,I241864,I241879,I241870,I241873,I241885,I241882,I247872,I247851,I247845,I247860,I247848,I247863,I247854,I247857,I247869,I247866,I254400,I254379,I254373,I254388,I254376,I254391,I254382,I254385,I254397,I254394,I392071,I392074,I392056,I392065,I392077,I392068,I392059,I392062,I392080,I414035,I414038,I414020,I414029,I414041,I414032,I414023,I414026,I414044,I432466,I432469,I432460,I432451,I432454,I432463,I432448,I432457,I447222,I447225,I447216,I447207,I447210,I447219,I447204,I447213,I489657,I489660,I489636,I489648,I489663,I489651,I489645,I489639,I489642,I489654,I494825,I494828,I494804,I494816,I494831,I494819,I494813,I494807,I494810,I494822,I557725,I557707,I557710,I557719,I557722,I557716,I557704,I557713,I571750,I571732,I571735,I571744,I571747,I571741,I571729,I571738,I608719,I608707,I608728,I608704,I608725,I608716,I608722,I608713,I608710,I631839,I631827,I631848,I631824,I631845,I631836,I631842,I631833,I631830,I700201,I700216,I700198,I700210,I700225,I700222,I700219,I700213,I700207,I700204;
wire I1364,I1372,I1380,I1388,I1396,I1404,I1412,I1420,I1428,I1436,I1444,I1452,I1460,I1468,I1476,I1484,I1492,I1500,I1508,I1516,I1524,I1532,I1540,I1548,I1556,I1564,I1572,I1580,I1588,I1596,I1604,I1612,I1620,I1628,I1636,I1644,I1652,I1660,I1668,I1676,I1684,I1692,I1700,I1708,I1716,I1724,I1732,I1740,I1748,I1756,I1764,I1772,I1780,I1788,I1796,I1804,I1812,I1820,I1828,I1836,I1844,I1852,I1860,I1868,I1876,I1884,I1892,I1900,I1908,I1916,I1924,I1932,I1940,I1948,I1956,I1964,I1972,I1980,I1988,I1996,I2004,I2012,I2020,I2028,I2036,I2044,I2052,I2060,I2068,I2076,I2084,I2092,I2100,I2108,I2116,I2124,I2132,I2140,I2148,I2156,I2164,I2172,I2180,I2188,I2196,I2204,I2212,I2220,I2228,I2236,I2244,I2252,I2260,I2268,I2276,I2284,I2292,I2300,I2308,I2316,I2324,I2332,I2340,I2348,I2356,I2364,I2372,I2380,I2388,I2396,I2404,I2412,I2420,I2428,I2436,I2444,I2452,I2460,I2468,I2476,I2484,I2492,I2500,I2508,I2516,I2524,I2532,I2540,I2548,I2556,I2564,I2572,I2580,I2588,I2596,I2604,I2612,I2620,I2628,I2636,I2644,I2652,I2660,I2668,I2676,I2684,I2692,I2700,I2708,I2716,I2724,I2732,I2740,I2748,I2756,I2764,I2772,I2780,I2788,I2796,I2804,I2812,I2820,I2828,I2836,I2844,I2852,I2860,I2868,I2876,I2884,I2892,I2900,I2908,I2916,I2924,I2932,I2940,I2948,I2956,I2964,I2972,I2980,I2988,I2996,I3004,I3012,I3020,I3028,I3035,I3042,I3074,I213027,I3100,I3108,I213018,I3125,I3066,I213021,I3165,I3173,I3190,I213015,I3207,I213024,I3224,I3241,I3045,I3272,I3289,I3306,I213012,I213030,I3048,I3337,I3354,I3371,I213036,I3388,I3405,I3422,I3057,I3453,I213033,I3470,I3487,I3063,I3518,I3060,I3549,I213039,I3575,I3583,I3600,I3054,I3051,I3669,I116387,I3695,I3703,I3720,I3661,I116393,I3760,I3768,I3785,I116402,I3802,I116396,I3819,I3836,I3640,I3867,I3884,I3901,I116399,I116405,I3643,I3932,I3949,I116408,I3966,I116384,I3983,I4000,I4017,I3652,I4048,I116390,I4065,I4082,I3658,I4113,I3655,I4144,I4170,I4178,I4195,I3649,I3646,I4264,I731153,I4290,I4298,I731144,I4315,I4256,I731147,I4355,I4363,I4380,I731159,I4397,I731150,I4414,I4431,I4235,I4462,I4479,I4496,I731138,I4238,I4527,I4544,I731162,I4561,I731141,I4578,I4595,I4612,I4247,I4643,I731156,I4660,I4677,I4253,I4708,I4250,I4739,I731165,I4765,I4773,I4790,I4244,I4241,I4859,I270714,I4885,I4893,I270696,I4910,I4851,I270708,I4950,I4958,I4975,I270693,I4992,I270702,I5009,I5026,I4830,I5057,I5074,I5091,I270699,I270720,I4833,I5122,I5139,I270711,I5156,I270717,I5173,I5190,I5207,I4842,I5238,I5255,I5272,I4848,I5303,I4845,I5334,I270705,I5360,I5368,I5385,I4839,I4836,I5454,I639919,I5480,I5488,I5505,I5446,I639934,I5545,I5553,I5570,I639931,I5587,I639940,I5604,I5621,I5425,I5652,I5669,I5686,I639928,I639937,I5428,I5717,I5734,I639925,I5751,I639916,I5768,I5785,I5802,I5437,I5833,I639922,I5850,I5867,I5443,I5898,I5440,I5929,I5955,I5963,I5980,I5434,I5431,I6049,I393814,I6075,I6083,I393793,I6100,I6041,I393802,I6140,I6148,I6165,I393808,I6182,I393805,I6199,I6216,I6020,I6247,I6264,I6281,I393796,I393790,I6023,I6312,I6329,I393811,I6346,I6363,I6380,I6397,I6032,I6428,I393799,I6445,I6462,I6038,I6493,I6035,I6524,I6550,I6558,I6575,I6029,I6026,I6644,I572293,I6670,I6678,I6695,I6636,I572308,I6735,I6743,I6760,I572305,I6777,I572314,I6794,I6811,I6615,I6842,I6859,I6876,I572302,I572311,I6618,I6907,I6924,I572299,I6941,I572290,I6958,I6975,I6992,I6627,I7023,I572296,I7040,I7057,I6633,I7088,I6630,I7119,I7145,I7153,I7170,I6624,I6621,I7239,I429295,I7265,I7273,I429286,I7290,I7231,I429292,I7330,I7338,I7355,I7372,I429298,I7389,I7406,I7210,I7437,I7454,I7471,I429307,I429304,I7213,I7502,I7519,I7536,I429289,I7553,I7570,I7587,I7222,I7618,I7635,I7652,I7228,I7683,I7225,I7714,I429301,I7740,I7748,I7765,I7219,I7216,I7837,I118770,I7863,I7880,I7888,I7905,I118788,I118773,I7922,I118776,I7948,I7829,I7820,I118764,I7993,I8001,I118767,I8018,I7817,I118779,I8058,I8066,I7823,I7811,I8111,I118785,I118782,I8128,I8154,I8162,I7805,I8193,I8210,I8227,I8244,I8261,I7826,I8292,I7814,I7808,I8364,I74210,I8390,I8407,I8415,I8432,I74225,I8449,I74228,I8475,I8356,I8347,I74222,I8520,I8528,I74231,I8545,I8344,I74207,I8585,I8593,I8350,I8338,I8638,I74213,I8655,I74216,I8681,I8689,I8332,I8720,I8737,I74219,I8754,I8771,I8788,I8353,I8819,I8341,I8335,I8891,I137810,I8917,I8934,I8942,I8959,I137828,I137813,I8976,I137816,I9002,I8883,I8874,I137804,I9047,I9055,I137807,I9072,I8871,I137819,I9112,I9120,I8877,I8865,I9165,I137825,I137822,I9182,I9208,I9216,I8859,I9247,I9264,I9281,I9298,I9315,I8880,I9346,I8868,I8862,I9418,I459861,I9444,I9461,I9469,I9486,I459852,I459873,I9503,I459855,I9529,I9410,I9401,I9574,I9582,I459870,I9599,I9398,I459864,I9639,I9647,I9404,I9392,I9692,I459858,I459867,I9709,I9735,I9743,I9386,I9774,I9791,I9808,I9825,I9842,I9407,I9873,I9395,I9389,I9945,I436146,I9971,I9988,I9996,I10013,I436137,I436158,I10030,I436140,I10056,I9937,I9928,I10101,I10109,I436155,I10126,I9925,I436149,I10166,I10174,I9931,I9919,I10219,I436143,I436152,I10236,I10262,I10270,I9913,I10301,I10318,I10335,I10352,I10369,I9934,I10400,I9922,I9916,I10472,I121745,I10498,I10515,I10523,I10540,I121763,I121748,I10557,I121751,I10583,I10464,I10455,I121739,I10628,I10636,I121742,I10653,I10452,I121754,I10693,I10701,I10458,I10446,I10746,I121760,I121757,I10763,I10789,I10797,I10440,I10828,I10845,I10862,I10879,I10896,I10461,I10927,I10449,I10443,I10999,I705553,I11025,I11042,I11050,I11067,I705556,I705562,I11084,I705571,I11110,I10991,I10982,I705574,I11155,I11163,I705565,I11180,I10979,I11220,I11228,I10985,I10973,I11273,I705580,I705559,I11290,I705568,I11316,I11324,I10967,I11355,I11372,I705577,I11389,I11406,I11423,I10988,I11454,I10976,I10970,I11526,I703768,I11552,I11569,I11577,I11594,I703771,I703777,I11611,I703786,I11637,I11518,I11509,I703789,I11682,I11690,I703780,I11707,I11506,I11747,I11755,I11512,I11500,I11800,I703795,I703774,I11817,I703783,I11843,I11851,I11494,I11882,I11899,I703792,I11916,I11933,I11950,I11515,I11981,I11503,I11497,I12053,I119365,I12079,I12096,I12104,I12121,I119383,I119368,I12138,I119371,I12164,I12045,I12036,I119359,I12209,I12217,I119362,I12234,I12033,I119374,I12274,I12282,I12039,I12027,I12327,I119380,I119377,I12344,I12370,I12378,I12021,I12409,I12426,I12443,I12460,I12477,I12042,I12508,I12030,I12024,I12580,I616242,I12606,I12623,I12631,I12648,I616230,I616221,I12665,I616218,I12691,I12572,I12563,I616224,I12736,I12744,I616236,I12761,I12560,I616233,I12801,I12809,I12566,I12554,I12854,I616227,I12871,I616239,I12897,I12905,I12548,I12936,I12953,I12970,I12987,I13004,I12569,I13035,I12557,I12551,I13107,I734708,I13133,I13150,I13158,I13175,I734711,I734717,I13192,I734726,I13218,I13099,I13090,I734729,I13263,I13271,I734720,I13288,I13087,I13328,I13336,I13093,I13081,I13381,I734735,I734714,I13398,I734723,I13424,I13432,I13075,I13463,I13480,I734732,I13497,I13514,I13531,I13096,I13562,I13084,I13078,I13634,I406512,I13660,I13677,I13685,I13702,I406527,I406530,I13719,I406509,I13745,I13626,I13617,I406515,I13790,I13798,I406521,I13815,I13614,I13855,I13863,I13620,I13608,I13908,I406524,I406506,I13925,I406518,I13951,I13959,I13602,I13990,I14007,I14024,I14041,I14058,I13623,I14089,I13611,I13605,I14161,I261989,I14187,I14204,I14212,I14229,I261992,I14246,I262013,I14272,I14153,I14144,I262001,I14317,I14325,I262004,I14342,I14141,I262010,I14382,I14390,I14147,I14135,I14435,I262007,I261995,I14452,I261998,I14478,I14486,I14129,I14517,I14534,I262016,I14551,I14568,I14585,I14150,I14616,I14138,I14132,I14688,I511624,I14714,I14731,I14739,I14756,I511600,I511627,I14773,I511612,I14799,I14680,I14671,I511618,I14844,I14852,I511603,I14869,I14668,I511621,I14909,I14917,I14674,I14662,I14962,I511606,I511609,I14979,I15005,I15013,I14656,I15044,I15061,I511615,I15078,I15095,I15112,I14677,I15143,I14665,I14659,I15215,I59981,I15241,I15258,I15266,I15283,I59996,I15300,I59999,I15326,I15207,I15198,I59993,I15371,I15379,I60002,I15396,I15195,I59978,I15436,I15444,I15201,I15189,I15489,I59984,I15506,I59987,I15532,I15540,I15183,I15571,I15588,I59990,I15605,I15622,I15639,I15204,I15670,I15192,I15186,I15742,I684063,I15768,I15785,I15793,I15810,I684066,I684060,I15827,I684069,I15853,I15734,I15725,I684057,I15898,I15906,I684072,I15923,I15722,I684048,I15963,I15971,I15728,I15716,I16016,I684051,I16033,I16059,I16067,I15710,I16098,I16115,I684054,I16132,I16149,I16166,I15731,I16197,I15719,I15713,I16269,I674237,I16295,I16312,I16320,I16337,I674240,I674234,I16354,I674243,I16380,I16261,I16252,I674231,I16425,I16433,I674246,I16450,I16249,I674222,I16490,I16498,I16255,I16243,I16543,I674225,I16560,I16586,I16594,I16237,I16625,I16642,I674228,I16659,I16676,I16693,I16258,I16724,I16246,I16240,I16796,I178784,I16822,I16839,I16847,I16864,I178781,I178775,I16881,I178769,I16907,I16788,I16779,I178757,I16952,I16960,I178766,I16977,I16776,I178763,I17017,I17025,I16782,I16770,I17070,I178760,I178778,I17087,I17113,I17121,I16764,I17152,I17169,I178772,I17186,I17203,I17220,I16785,I17251,I16773,I16767,I17323,I190378,I17349,I17366,I17374,I17391,I190375,I190369,I17408,I190363,I17434,I17315,I17306,I190351,I17479,I17487,I190360,I17504,I17303,I190357,I17544,I17552,I17309,I17297,I17597,I190354,I190372,I17614,I17640,I17648,I17291,I17679,I17696,I190366,I17713,I17730,I17747,I17312,I17778,I17300,I17294,I17850,I127100,I17876,I17893,I17901,I17918,I127118,I127103,I17935,I127106,I17961,I17842,I17833,I127094,I18006,I18014,I127097,I18031,I17830,I127109,I18071,I18079,I17836,I17824,I18124,I127115,I127112,I18141,I18167,I18175,I17818,I18206,I18223,I18240,I18257,I18274,I17839,I18305,I17827,I17821,I18377,I421390,I18403,I18420,I18428,I18445,I421381,I421402,I18462,I421384,I18488,I18369,I18360,I18533,I18541,I421399,I18558,I18357,I421393,I18598,I18606,I18363,I18351,I18651,I421387,I421396,I18668,I18694,I18702,I18345,I18733,I18750,I18767,I18784,I18801,I18366,I18832,I18354,I18348,I18904,I467239,I18930,I18947,I18955,I18972,I467230,I467251,I18989,I467233,I19015,I18896,I18887,I19060,I19068,I467248,I19085,I18884,I467242,I19125,I19133,I18890,I18878,I19178,I467236,I467245,I19195,I19221,I19229,I18872,I19260,I19277,I19294,I19311,I19328,I18893,I19359,I18881,I18875,I19431,I441943,I19457,I19474,I19482,I19499,I441934,I441955,I19516,I441937,I19542,I19423,I19414,I19587,I19595,I441952,I19612,I19411,I441946,I19652,I19660,I19417,I19405,I19705,I441940,I441949,I19722,I19748,I19756,I19399,I19787,I19804,I19821,I19838,I19855,I19420,I19886,I19408,I19402,I19958,I275589,I19984,I20001,I20009,I20026,I275592,I20043,I275613,I20069,I19950,I19941,I275601,I20114,I20122,I275604,I20139,I19938,I275610,I20179,I20187,I19944,I19932,I20232,I275607,I275595,I20249,I275598,I20275,I20283,I19926,I20314,I20331,I275616,I20348,I20365,I20382,I19947,I20413,I19935,I19929,I20485,I258181,I20511,I20528,I20536,I20553,I258184,I20570,I258205,I20596,I20477,I20468,I258193,I20641,I20649,I258196,I20666,I20465,I258202,I20706,I20714,I20471,I20459,I20759,I258199,I258187,I20776,I258190,I20802,I20810,I20453,I20841,I20858,I258208,I20875,I20892,I20909,I20474,I20940,I20462,I20456,I21012,I605260,I21038,I21055,I21063,I21080,I605248,I605239,I21097,I605236,I21123,I21004,I20995,I605242,I21168,I21176,I605254,I21193,I20992,I605251,I21233,I21241,I20998,I20986,I21286,I605245,I21303,I605257,I21329,I21337,I20980,I21368,I21385,I21402,I21419,I21436,I21001,I21467,I20989,I20983,I21539,I584452,I21565,I21582,I21590,I21607,I584440,I584431,I21624,I584428,I21650,I21531,I21522,I584434,I21695,I21703,I584446,I21720,I21519,I584443,I21760,I21768,I21525,I21513,I21813,I584437,I21830,I584449,I21856,I21864,I21507,I21895,I21912,I21929,I21946,I21963,I21528,I21994,I21516,I21510,I22066,I160866,I22092,I22109,I22117,I22134,I160863,I160857,I22151,I160851,I22177,I22058,I22049,I160839,I22222,I22230,I160848,I22247,I22046,I160845,I22287,I22295,I22052,I22040,I22340,I160842,I160860,I22357,I22383,I22391,I22034,I22422,I22439,I160854,I22456,I22473,I22490,I22055,I22521,I22043,I22037,I22593,I165082,I22619,I22636,I22644,I22661,I165079,I165073,I22678,I165067,I22704,I22585,I22576,I165055,I22749,I22757,I165064,I22774,I22573,I165061,I22814,I22822,I22579,I22567,I22867,I165058,I165076,I22884,I22910,I22918,I22561,I22949,I22966,I165070,I22983,I23000,I23017,I22582,I23048,I22570,I22564,I23120,I481908,I23146,I23163,I23171,I23188,I481884,I481911,I23205,I481896,I23231,I23112,I23103,I481902,I23276,I23284,I481887,I23301,I23100,I481905,I23341,I23349,I23106,I23094,I23394,I481890,I481893,I23411,I23437,I23445,I23088,I23476,I23493,I481899,I23510,I23527,I23544,I23109,I23575,I23097,I23091,I23647,I292445,I23673,I23690,I23698,I23715,I292451,I292439,I23732,I292436,I23758,I23639,I23630,I292448,I23803,I23811,I292442,I23828,I23627,I292460,I23868,I23876,I23633,I23621,I23921,I292454,I292457,I23938,I23964,I23972,I23615,I24003,I24020,I24037,I24054,I24071,I23636,I24102,I23624,I23618,I24174,I272869,I24200,I24217,I24225,I24242,I272872,I24259,I272893,I24285,I24166,I24157,I272881,I24330,I24338,I272884,I24355,I24154,I272890,I24395,I24403,I24160,I24148,I24448,I272887,I272875,I24465,I272878,I24491,I24499,I24142,I24530,I24547,I272896,I24564,I24581,I24598,I24163,I24629,I24151,I24145,I24701,I671925,I24727,I24744,I24752,I24769,I671928,I671922,I24786,I671931,I24812,I24693,I24684,I671919,I24857,I24865,I671934,I24882,I24681,I671910,I24922,I24930,I24687,I24675,I24975,I671913,I24992,I25018,I25026,I24669,I25057,I25074,I671916,I25091,I25108,I25125,I24690,I25156,I24678,I24672,I25228,I277221,I25254,I25271,I25279,I25296,I277224,I25313,I277245,I25339,I25220,I25211,I277233,I25384,I25392,I277236,I25409,I25208,I277242,I25449,I25457,I25214,I25202,I25502,I277239,I277227,I25519,I277230,I25545,I25553,I25196,I25584,I25601,I277248,I25618,I25635,I25652,I25217,I25683,I25205,I25199,I25755,I585608,I25781,I25798,I25806,I25823,I585596,I585587,I25840,I585584,I25866,I25747,I25738,I585590,I25911,I25919,I585602,I25936,I25735,I585599,I25976,I25984,I25741,I25729,I26029,I585593,I26046,I585605,I26072,I26080,I25723,I26111,I26128,I26145,I26162,I26179,I25744,I26210,I25732,I25726,I26282,I239685,I26308,I26325,I26333,I26350,I239688,I26367,I239709,I26393,I26274,I26265,I239697,I26438,I26446,I239700,I26463,I26262,I239706,I26503,I26511,I26268,I26256,I26556,I239703,I239691,I26573,I239694,I26599,I26607,I26250,I26638,I26655,I239712,I26672,I26689,I26706,I26271,I26737,I26259,I26253,I26809,I26835,I26852,I26860,I26877,I26894,I26920,I26801,I26792,I26965,I26973,I26990,I26789,I27030,I27038,I26795,I26783,I27083,I27100,I27126,I27134,I26777,I27165,I27182,I27199,I27216,I27233,I26798,I27264,I26786,I26780,I27336,I345822,I27362,I27379,I27387,I27404,I345837,I345840,I27421,I345819,I27447,I27328,I27319,I345825,I27492,I27500,I345831,I27517,I27316,I27557,I27565,I27322,I27310,I27610,I345834,I345816,I27627,I345828,I27653,I27661,I27304,I27692,I27709,I27726,I27743,I27760,I27325,I27791,I27313,I27307,I27863,I281140,I27889,I27906,I27914,I27931,I281146,I281134,I27948,I281131,I27974,I27855,I27846,I281143,I28019,I28027,I281137,I28044,I27843,I281155,I28084,I28092,I27849,I27837,I28137,I281149,I281152,I28154,I28180,I28188,I27831,I28219,I28236,I28253,I28270,I28287,I27852,I28318,I27840,I27834,I28390,I225687,I28416,I28433,I28441,I28458,I225684,I225678,I28475,I225672,I28501,I28382,I28373,I225660,I28546,I28554,I225669,I28571,I28370,I225666,I28611,I28619,I28376,I28364,I28664,I225663,I225681,I28681,I28707,I28715,I28358,I28746,I28763,I225675,I28780,I28797,I28814,I28379,I28845,I28367,I28361,I28917,I111041,I28943,I28951,I28968,I111035,I111029,I28985,I111050,I29011,I111047,I29028,I29036,I111044,I29053,I28885,I29084,I29101,I28897,I29141,I28906,I29163,I111032,I29180,I111053,I29206,I29223,I28909,I29245,I28894,I29276,I111038,I29293,I29310,I29327,I28903,I29358,I28891,I28900,I28888,I29444,I465658,I29470,I29478,I29495,I465655,I465670,I29512,I465652,I29538,I465649,I29555,I29563,I29580,I29412,I29611,I29628,I29424,I29668,I29433,I29690,I465664,I29707,I465667,I29733,I29750,I29436,I29772,I29421,I29803,I465661,I29820,I29837,I29854,I29430,I29885,I29418,I29427,I29415,I29971,I301319,I29997,I30005,I30022,I301331,I301316,I30039,I301310,I30065,I301325,I30082,I30090,I301313,I30107,I29939,I30138,I30155,I29951,I301322,I30195,I29960,I30217,I301328,I301334,I30234,I30260,I30277,I29963,I30299,I29948,I30330,I30347,I30364,I30381,I29957,I30412,I29945,I29954,I29942,I30498,I457753,I30524,I30532,I30549,I457750,I457765,I30566,I457747,I30592,I457744,I30609,I30617,I30634,I30466,I30665,I30682,I30478,I30722,I30487,I30744,I457759,I30761,I457762,I30787,I30804,I30490,I30826,I30475,I30857,I457756,I30874,I30891,I30908,I30484,I30939,I30472,I30481,I30469,I31025,I521299,I31051,I31059,I31076,I521317,I521311,I31093,I521290,I31119,I521308,I31136,I31144,I521293,I31161,I30993,I31192,I31209,I31005,I521305,I31249,I31014,I31271,I521314,I521302,I31288,I521296,I31314,I31331,I31017,I31353,I31002,I31384,I31401,I31418,I31435,I31011,I31466,I30999,I31008,I30996,I31552,I483185,I31578,I31586,I31603,I483203,I483197,I31620,I483176,I31646,I483194,I31663,I31671,I483179,I31688,I31520,I31719,I31736,I31532,I483191,I31776,I31541,I31798,I483200,I483188,I31815,I483182,I31841,I31858,I31544,I31880,I31529,I31911,I31928,I31945,I31962,I31538,I31993,I31526,I31535,I31523,I32079,I594260,I32105,I32113,I32130,I594275,I594254,I32147,I594257,I32173,I594278,I32190,I32198,I32215,I32047,I32246,I32263,I32059,I32303,I32068,I32325,I594266,I594263,I32342,I594269,I32368,I32385,I32071,I32407,I32056,I32438,I594272,I32455,I32472,I32489,I32065,I32520,I32053,I32062,I32050,I32606,I469874,I32632,I32640,I32657,I469871,I469886,I32674,I469868,I32700,I469865,I32717,I32725,I32742,I32574,I32773,I32790,I32586,I32830,I32595,I32852,I469880,I32869,I469883,I32895,I32912,I32598,I32934,I32583,I32965,I469877,I32982,I32999,I33016,I32592,I33047,I32580,I32589,I32577,I33133,I33159,I33167,I33184,I33201,I33227,I33244,I33252,I33269,I33101,I33300,I33317,I33113,I33357,I33122,I33379,I33396,I33422,I33439,I33125,I33461,I33110,I33492,I33509,I33526,I33543,I33119,I33574,I33107,I33116,I33104,I33660,I216201,I33686,I33694,I33711,I216183,I216198,I33728,I216174,I33754,I216177,I33771,I33779,I216192,I33796,I33628,I33827,I33844,I33640,I216195,I33884,I33649,I33906,I216186,I33923,I216180,I33949,I33966,I33652,I33988,I33637,I34019,I216189,I34036,I34053,I34070,I33646,I34101,I33634,I33643,I33631,I34187,I450902,I34213,I34221,I34238,I450899,I450914,I34255,I450896,I34281,I450893,I34298,I34306,I34323,I34155,I34354,I34371,I34167,I34411,I34176,I34433,I450908,I34450,I450911,I34476,I34493,I34179,I34515,I34164,I34546,I450905,I34563,I34580,I34597,I34173,I34628,I34161,I34170,I34158,I34714,I105091,I34740,I34748,I34765,I105085,I105079,I34782,I105100,I34808,I105097,I34825,I34833,I105094,I34850,I34682,I34881,I34898,I34694,I34938,I34703,I34960,I105082,I34977,I105103,I35003,I35020,I34706,I35042,I34691,I35073,I105088,I35090,I35107,I35124,I34700,I35155,I34688,I34697,I34685,I35241,I139601,I35267,I35275,I35292,I139595,I139589,I35309,I139610,I35335,I139607,I35352,I35360,I139604,I35377,I35209,I35408,I35425,I35221,I35465,I35230,I35487,I139592,I35504,I139613,I35530,I35547,I35233,I35569,I35218,I35600,I139598,I35617,I35634,I35651,I35227,I35682,I35215,I35224,I35212,I35768,I416344,I35794,I35802,I35819,I416335,I416353,I35836,I416332,I35862,I35879,I35887,I416338,I35904,I35736,I35935,I35952,I35748,I35992,I35757,I36014,I416350,I416341,I36031,I416356,I36057,I36074,I35760,I36096,I35745,I36127,I416347,I36144,I36161,I36178,I35754,I36209,I35742,I35751,I35739,I36295,I323283,I36321,I36329,I36346,I323295,I323280,I36363,I323274,I36389,I323289,I36406,I36414,I323277,I36431,I36263,I36462,I36479,I36275,I323286,I36519,I36284,I36541,I323292,I323298,I36558,I36584,I36601,I36287,I36623,I36272,I36654,I36671,I36688,I36705,I36281,I36736,I36269,I36278,I36266,I36822,I356810,I36848,I36856,I36873,I356801,I356819,I36890,I356798,I36916,I36933,I36941,I356804,I36958,I36790,I36989,I37006,I36802,I37046,I36811,I37068,I356816,I356807,I37085,I356822,I37111,I37128,I36814,I37150,I36799,I37181,I356813,I37198,I37215,I37232,I36808,I37263,I36796,I36805,I36793,I37349,I540679,I37375,I37383,I37400,I540697,I540691,I37417,I540670,I37443,I540688,I37460,I37468,I540673,I37485,I37317,I37516,I37533,I37329,I540685,I37573,I37338,I37595,I540694,I540682,I37612,I540676,I37638,I37655,I37341,I37677,I37326,I37708,I37725,I37742,I37759,I37335,I37790,I37323,I37332,I37320,I37876,I554902,I37902,I37910,I37927,I554899,I554905,I37944,I37970,I37987,I37995,I38012,I37844,I38043,I38060,I37856,I554908,I38100,I37865,I38122,I554911,I554920,I38139,I554914,I38165,I38182,I37868,I38204,I37853,I38235,I554917,I38252,I38269,I38286,I37862,I38317,I37850,I37859,I37847,I38403,I80696,I38429,I38437,I38454,I80690,I80684,I38471,I80705,I38497,I80702,I38514,I38522,I80699,I38539,I38371,I38570,I38587,I38383,I38627,I38392,I38649,I80687,I38666,I80708,I38692,I38709,I38395,I38731,I38380,I38762,I80693,I38779,I38796,I38813,I38389,I38844,I38377,I38386,I38374,I38930,I38956,I38964,I38981,I38998,I39024,I39041,I39049,I39066,I38898,I39097,I39114,I38910,I39154,I38919,I39176,I39193,I39219,I39236,I38922,I39258,I38907,I39289,I39306,I39323,I39340,I38916,I39371,I38904,I38913,I38901,I39457,I446159,I39483,I39491,I39508,I446156,I446171,I39525,I446153,I39551,I446150,I39568,I39576,I39593,I39425,I39624,I39641,I39437,I39681,I39446,I39703,I446165,I39720,I446168,I39746,I39763,I39449,I39785,I39434,I39816,I446162,I39833,I39850,I39867,I39443,I39898,I39431,I39440,I39428,I39984,I189851,I40010,I40018,I40035,I189833,I189848,I40052,I189824,I40078,I189827,I40095,I40103,I189842,I40120,I39952,I40151,I40168,I39964,I189845,I40208,I39973,I40230,I189836,I40247,I189830,I40273,I40290,I39976,I40312,I39961,I40343,I189839,I40360,I40377,I40394,I39970,I40425,I39958,I39967,I39955,I40511,I659948,I40537,I40545,I40562,I659942,I659963,I40579,I659954,I40605,I659945,I40622,I40630,I659957,I40647,I40479,I40678,I40695,I40491,I40735,I40500,I40757,I659966,I659951,I40774,I40800,I40817,I40503,I40839,I40488,I40870,I659960,I40887,I40904,I40921,I40497,I40952,I40485,I40494,I40482,I41038,I41064,I41072,I41089,I41106,I41132,I41149,I41157,I41174,I41006,I41205,I41222,I41018,I41262,I41027,I41284,I41301,I41327,I41344,I41030,I41366,I41015,I41397,I41414,I41431,I41448,I41024,I41479,I41012,I41021,I41009,I41565,I609288,I41591,I41599,I41616,I609303,I609282,I41633,I609285,I41659,I609306,I41676,I41684,I41701,I41533,I41732,I41749,I41545,I41789,I41554,I41811,I609294,I609291,I41828,I609297,I41854,I41871,I41557,I41893,I41542,I41924,I609300,I41941,I41958,I41975,I41551,I42006,I41539,I41548,I41536,I42092,I650700,I42118,I42126,I42143,I650694,I650715,I42160,I650706,I42186,I650697,I42203,I42211,I650709,I42228,I42060,I42259,I42276,I42072,I42316,I42081,I42338,I650718,I650703,I42355,I42381,I42398,I42084,I42420,I42069,I42451,I650712,I42468,I42485,I42502,I42078,I42533,I42066,I42075,I42063,I42619,I552097,I42645,I42653,I42670,I552094,I552100,I42687,I42713,I42730,I42738,I42755,I42587,I42786,I42803,I42599,I552103,I42843,I42608,I42865,I552106,I552115,I42882,I552109,I42908,I42925,I42611,I42947,I42596,I42978,I552112,I42995,I43012,I43029,I42605,I43060,I42593,I42602,I42590,I43146,I223579,I43172,I43180,I43197,I223561,I223576,I43214,I223552,I43240,I223555,I43257,I43265,I223570,I43282,I43114,I43313,I43330,I43126,I223573,I43370,I43135,I43392,I223564,I43409,I223558,I43435,I43452,I43138,I43474,I43123,I43505,I223567,I43522,I43539,I43556,I43132,I43587,I43120,I43129,I43117,I43673,I331953,I43699,I43707,I43724,I331965,I331950,I43741,I331944,I43767,I331959,I43784,I43792,I331947,I43809,I43641,I43840,I43857,I43653,I331956,I43897,I43662,I43919,I331962,I331968,I43936,I43962,I43979,I43665,I44001,I43650,I44032,I44049,I44066,I44083,I43659,I44114,I43647,I43656,I43644,I44200,I240791,I44226,I44234,I44251,I240785,I240776,I44268,I240797,I44294,I240779,I44311,I44319,I240773,I44336,I44168,I44367,I44384,I44180,I44424,I44189,I44446,I240800,I240782,I44463,I240788,I44489,I44506,I44192,I44528,I44177,I44559,I240794,I44576,I44593,I44610,I44186,I44641,I44174,I44183,I44171,I44727,I431930,I44753,I44761,I44778,I431927,I431942,I44795,I431924,I44821,I431921,I44838,I44846,I44863,I44695,I44894,I44911,I44707,I44951,I44716,I44973,I431936,I44990,I431939,I45016,I45033,I44719,I45055,I44704,I45086,I431933,I45103,I45120,I45137,I44713,I45168,I44701,I44710,I44698,I45254,I688693,I45280,I45288,I45305,I688696,I688690,I45322,I688687,I45348,I688672,I45365,I45373,I688681,I45390,I45222,I45421,I45438,I45234,I45478,I45243,I45500,I688675,I688678,I45517,I688684,I45543,I45560,I45246,I45582,I45231,I45613,I45630,I45647,I45664,I45240,I45695,I45228,I45237,I45225,I45781,I536803,I45807,I45815,I45832,I536821,I536815,I45849,I536794,I45875,I536812,I45892,I45900,I536797,I45917,I45749,I45948,I45965,I45761,I536809,I46005,I45770,I46027,I536818,I536806,I46044,I536800,I46070,I46087,I45773,I46109,I45758,I46140,I46157,I46174,I46191,I45767,I46222,I45755,I45764,I45752,I46308,I730555,I46334,I46342,I46359,I730549,I730570,I46376,I730546,I46402,I730567,I46419,I46427,I730564,I46444,I46276,I46475,I46492,I46288,I730552,I46532,I46297,I46554,I730561,I730558,I46571,I730543,I46597,I46614,I46300,I46636,I46285,I46667,I46684,I46701,I46718,I46294,I46749,I46282,I46291,I46279,I46835,I597150,I46861,I46869,I46886,I597165,I597144,I46903,I597147,I46929,I597168,I46946,I46954,I46971,I46803,I47002,I47019,I46815,I47059,I46824,I47081,I597156,I597153,I47098,I597159,I47124,I47141,I46827,I47163,I46812,I47194,I597162,I47211,I47228,I47245,I46821,I47276,I46809,I46818,I46806,I47362,I326173,I47388,I47396,I47413,I326185,I326170,I47430,I326164,I47456,I326179,I47473,I47481,I326167,I47498,I47330,I47529,I47546,I47342,I326176,I47586,I47351,I47608,I326182,I326188,I47625,I47651,I47668,I47354,I47690,I47339,I47721,I47738,I47755,I47772,I47348,I47803,I47336,I47345,I47333,I47889,I204607,I47915,I47923,I47940,I204589,I204604,I47957,I204580,I47983,I204583,I48000,I48008,I204598,I48025,I47857,I48056,I48073,I47869,I204601,I48113,I47878,I48135,I204592,I48152,I204586,I48178,I48195,I47881,I48217,I47866,I48248,I204595,I48265,I48282,I48299,I47875,I48330,I47863,I47872,I47860,I48416,I172460,I48442,I48450,I48467,I172442,I172457,I48484,I172433,I48510,I172436,I48527,I48535,I172451,I48552,I48384,I48583,I48600,I48396,I172454,I48640,I48405,I48662,I172445,I48679,I172439,I48705,I48722,I48408,I48744,I48393,I48775,I172448,I48792,I48809,I48826,I48402,I48857,I48390,I48399,I48387,I48943,I76540,I48969,I48977,I48994,I76537,I76519,I49011,I76525,I49037,I76534,I49054,I49062,I76528,I49079,I48911,I49110,I49127,I48923,I76543,I49167,I48932,I49189,I76531,I76522,I49206,I49232,I49249,I48935,I49271,I48920,I49302,I76546,I49319,I49336,I49353,I48929,I49384,I48917,I48926,I48914,I49470,I174041,I49496,I49504,I49521,I174023,I174038,I49538,I174014,I49564,I174017,I49581,I49589,I174032,I49606,I49438,I49637,I49654,I49450,I174035,I49694,I49459,I49716,I174026,I49733,I174020,I49759,I49776,I49462,I49798,I49447,I49829,I174029,I49846,I49863,I49880,I49456,I49911,I49444,I49453,I49441,I49997,I326751,I50023,I50031,I50048,I326763,I326748,I50065,I326742,I50091,I326757,I50108,I50116,I326745,I50133,I49965,I50164,I50181,I49977,I326754,I50221,I49986,I50243,I326760,I326766,I50260,I50286,I50303,I49989,I50325,I49974,I50356,I50373,I50390,I50407,I49983,I50438,I49971,I49980,I49968,I50524,I731745,I50550,I50558,I50575,I731739,I731760,I50592,I731736,I50618,I731757,I50635,I50643,I731754,I50660,I50492,I50691,I50708,I50504,I731742,I50748,I50513,I50770,I731751,I731748,I50787,I731733,I50813,I50830,I50516,I50852,I50501,I50883,I50900,I50917,I50934,I50510,I50965,I50498,I50507,I50495,I51051,I390334,I51077,I51085,I51102,I390325,I390343,I51119,I390322,I51145,I51162,I51170,I390328,I51187,I51019,I51218,I51235,I51031,I51275,I51040,I51297,I390340,I390331,I51314,I390346,I51340,I51357,I51043,I51379,I51028,I51410,I390337,I51427,I51444,I51461,I51037,I51492,I51025,I51034,I51022,I51578,I51604,I51612,I51629,I51646,I51672,I51689,I51697,I51714,I51546,I51745,I51762,I51558,I51802,I51567,I51824,I51841,I51867,I51884,I51570,I51906,I51555,I51937,I51954,I51971,I51988,I51564,I52019,I51552,I51561,I51549,I52105,I52131,I52139,I52156,I52173,I52199,I52216,I52224,I52241,I52073,I52272,I52289,I52085,I52329,I52094,I52351,I52368,I52394,I52411,I52097,I52433,I52082,I52464,I52481,I52498,I52515,I52091,I52546,I52079,I52088,I52076,I52632,I491583,I52658,I52666,I52683,I491601,I491595,I52700,I491574,I52726,I491592,I52743,I52751,I491577,I52768,I52600,I52799,I52816,I52612,I491589,I52856,I52621,I52878,I491598,I491586,I52895,I491580,I52921,I52938,I52624,I52960,I52609,I52991,I53008,I53025,I53042,I52618,I53073,I52606,I52615,I52603,I53159,I53185,I53193,I53210,I53227,I53253,I53270,I53278,I53295,I53127,I53326,I53343,I53139,I53383,I53148,I53405,I53422,I53448,I53465,I53151,I53487,I53136,I53518,I53535,I53552,I53569,I53145,I53600,I53133,I53142,I53130,I53686,I463550,I53712,I53720,I53737,I463547,I463562,I53754,I463544,I53780,I463541,I53797,I53805,I53822,I53654,I53853,I53870,I53666,I53910,I53675,I53932,I463556,I53949,I463559,I53975,I53992,I53678,I54014,I53663,I54045,I463553,I54062,I54079,I54096,I53672,I54127,I53660,I53669,I53657,I54213,I194594,I54239,I54247,I54264,I194576,I194591,I54281,I194567,I54307,I194570,I54324,I54332,I194585,I54349,I54181,I54380,I54397,I54193,I194588,I54437,I54202,I54459,I194579,I54476,I194573,I54502,I54519,I54205,I54541,I54190,I54572,I194582,I54589,I54606,I54623,I54199,I54654,I54187,I54196,I54184,I54740,I89621,I54766,I54774,I54791,I89615,I89609,I54808,I89630,I54834,I89627,I54851,I54859,I89624,I54876,I54708,I54907,I54924,I54720,I54964,I54729,I54986,I89612,I55003,I89633,I55029,I55046,I54732,I55068,I54717,I55099,I89618,I55116,I55133,I55150,I54726,I55181,I54714,I54723,I54711,I55267,I390912,I55293,I55301,I55318,I390903,I390921,I55335,I390900,I55361,I55378,I55386,I390906,I55403,I55235,I55434,I55451,I55247,I55491,I55256,I55513,I390918,I390909,I55530,I390924,I55556,I55573,I55259,I55595,I55244,I55626,I390915,I55643,I55660,I55677,I55253,I55708,I55241,I55250,I55238,I55794,I278327,I55820,I55828,I55845,I278321,I278312,I55862,I278333,I55888,I278315,I55905,I55913,I278309,I55930,I55762,I55961,I55978,I55774,I56018,I55783,I56040,I278336,I278318,I56057,I278324,I56083,I56100,I55786,I56122,I55771,I56153,I278330,I56170,I56187,I56204,I55780,I56235,I55768,I55777,I55765,I56321,I740075,I56347,I56355,I56372,I740069,I740090,I56389,I740066,I56415,I740087,I56432,I56440,I740084,I56457,I56289,I56488,I56505,I56301,I740072,I56545,I56310,I56567,I740081,I740078,I56584,I740063,I56610,I56627,I56313,I56649,I56298,I56680,I56697,I56714,I56731,I56307,I56762,I56295,I56304,I56292,I56848,I211458,I56874,I56882,I56899,I211440,I211455,I56916,I211431,I56942,I211434,I56959,I56967,I211449,I56984,I56816,I57015,I57032,I56828,I211452,I57072,I56837,I57094,I211443,I57111,I211437,I57137,I57154,I56840,I57176,I56825,I57207,I211446,I57224,I57241,I57258,I56834,I57289,I56822,I56831,I56819,I57375,I297199,I57401,I57409,I57426,I297220,I297214,I57443,I297196,I57469,I57486,I57494,I297208,I57511,I57343,I57542,I57559,I57355,I297205,I57599,I57364,I57621,I297211,I297202,I57638,I57664,I57681,I57367,I57703,I57352,I57734,I297217,I57751,I57768,I57785,I57361,I57816,I57349,I57358,I57346,I57902,I134246,I57928,I57936,I57953,I134240,I134234,I57970,I134255,I57996,I134252,I58013,I58021,I134249,I58038,I57870,I58069,I58086,I57882,I58126,I57891,I58148,I134237,I58165,I134258,I58191,I58208,I57894,I58230,I57879,I58261,I134243,I58278,I58295,I58312,I57888,I58343,I57876,I57885,I57873,I58429,I438254,I58455,I58463,I58480,I438251,I438266,I58497,I438248,I58523,I438245,I58540,I58548,I58565,I58397,I58596,I58613,I58409,I58653,I58418,I58675,I438260,I58692,I438263,I58718,I58735,I58421,I58757,I58406,I58788,I438257,I58805,I58822,I58839,I58415,I58870,I58403,I58412,I58400,I58956,I729960,I58982,I58990,I59007,I729954,I729975,I59024,I729951,I59050,I729972,I59067,I59075,I729969,I59092,I58924,I59123,I59140,I58936,I729957,I59180,I58945,I59202,I729966,I729963,I59219,I729948,I59245,I59262,I58948,I59284,I58933,I59315,I59332,I59349,I59366,I58942,I59397,I58930,I58939,I58927,I59483,I399004,I59509,I59517,I59534,I398995,I399013,I59551,I398992,I59577,I59594,I59602,I398998,I59619,I59451,I59650,I59667,I59463,I59707,I59472,I59729,I399010,I399001,I59746,I399016,I59772,I59789,I59475,I59811,I59460,I59842,I399007,I59859,I59876,I59893,I59469,I59924,I59457,I59466,I59454,I60010,I109851,I60036,I60044,I60061,I109845,I109839,I60078,I109860,I60104,I109857,I60121,I60129,I109854,I60146,I60177,I60194,I60234,I60256,I109842,I60273,I109863,I60299,I60316,I60338,I60369,I109848,I60386,I60403,I60420,I60451,I60537,I269079,I60563,I60571,I60588,I269073,I269064,I60605,I269085,I60631,I269067,I60648,I60656,I269061,I60673,I60505,I60704,I60721,I60517,I60761,I60526,I60783,I269088,I269070,I60800,I269076,I60826,I60843,I60529,I60865,I60514,I60896,I269082,I60913,I60930,I60947,I60523,I60978,I60511,I60520,I60508,I61064,I356232,I61090,I61098,I61115,I356223,I356241,I61132,I356220,I61158,I61175,I61183,I356226,I61200,I61032,I61231,I61248,I61044,I61288,I61053,I61310,I356238,I356229,I61327,I356244,I61353,I61370,I61056,I61392,I61041,I61423,I356235,I61440,I61457,I61474,I61050,I61505,I61038,I61047,I61035,I61591,I180892,I61617,I61625,I61642,I180874,I180889,I61659,I180865,I61685,I180868,I61702,I61710,I180883,I61727,I61559,I61758,I61775,I61571,I180886,I61815,I61580,I61837,I180877,I61854,I180871,I61880,I61897,I61583,I61919,I61568,I61950,I180880,I61967,I61984,I62001,I61577,I62032,I61565,I61574,I61562,I62118,I180365,I62144,I62152,I62169,I180347,I180362,I62186,I180338,I62212,I180341,I62229,I62237,I180356,I62254,I62086,I62285,I62302,I62098,I180359,I62342,I62107,I62364,I180350,I62381,I180344,I62407,I62424,I62110,I62446,I62095,I62477,I180353,I62494,I62511,I62528,I62104,I62559,I62092,I62101,I62089,I62645,I175095,I62671,I62679,I62696,I175077,I175092,I62713,I175068,I62739,I175071,I62756,I62764,I175086,I62781,I62613,I62812,I62829,I62625,I175089,I62869,I62634,I62891,I175080,I62908,I175074,I62934,I62951,I62637,I62973,I62622,I63004,I175083,I63021,I63038,I63055,I62631,I63086,I62619,I62628,I62616,I63172,I529697,I63198,I63206,I63223,I529715,I529709,I63240,I529688,I63266,I529706,I63283,I63291,I529691,I63308,I63140,I63339,I63356,I63152,I529703,I63396,I63161,I63418,I529712,I529700,I63435,I529694,I63461,I63478,I63164,I63500,I63149,I63531,I63548,I63565,I63582,I63158,I63613,I63146,I63155,I63143,I63699,I516777,I63725,I63733,I63750,I516795,I516789,I63767,I516768,I63793,I516786,I63810,I63818,I516771,I63835,I63667,I63866,I63883,I63679,I516783,I63923,I63688,I63945,I516792,I516780,I63962,I516774,I63988,I64005,I63691,I64027,I63676,I64058,I64075,I64092,I64109,I63685,I64140,I63673,I63682,I63670,I64226,I738885,I64252,I64260,I64277,I738879,I738900,I64294,I738876,I64320,I738897,I64337,I64345,I738894,I64362,I64194,I64393,I64410,I64206,I738882,I64450,I64215,I64472,I738891,I738888,I64489,I738873,I64515,I64532,I64218,I64554,I64203,I64585,I64602,I64619,I64636,I64212,I64667,I64200,I64209,I64197,I64753,I382820,I64779,I64787,I64804,I382811,I382829,I64821,I382808,I64847,I64864,I64872,I382814,I64889,I64721,I64920,I64937,I64733,I64977,I64742,I64999,I382826,I382817,I65016,I382832,I65042,I65059,I64745,I65081,I64730,I65112,I382823,I65129,I65146,I65163,I64739,I65194,I64727,I64736,I64724,I65280,I300163,I65306,I65314,I65331,I300175,I300160,I65348,I300154,I65374,I300169,I65391,I65399,I300157,I65416,I65248,I65447,I65464,I65260,I300166,I65504,I65269,I65526,I300172,I300178,I65543,I65569,I65586,I65272,I65608,I65257,I65639,I65656,I65673,I65690,I65266,I65721,I65254,I65263,I65251,I65807,I378774,I65833,I65841,I65858,I378765,I378783,I65875,I378762,I65901,I65918,I65926,I378768,I65943,I65775,I65974,I65991,I65787,I66031,I65796,I66053,I378780,I378771,I66070,I378786,I66096,I66113,I65799,I66135,I65784,I66166,I378777,I66183,I66200,I66217,I65793,I66248,I65781,I65790,I65778,I66334,I613334,I66360,I66368,I66385,I613349,I613328,I66402,I613331,I66428,I613352,I66445,I66453,I66470,I66302,I66501,I66518,I66314,I66558,I66323,I66580,I613340,I613337,I66597,I613343,I66623,I66640,I66326,I66662,I66311,I66693,I613346,I66710,I66727,I66744,I66320,I66775,I66308,I66317,I66305,I66861,I117586,I66887,I66895,I66912,I117580,I117574,I66929,I117595,I66955,I117592,I66972,I66980,I117589,I66997,I66829,I67028,I67045,I66841,I67085,I66850,I67107,I117577,I67124,I117598,I67150,I67167,I66853,I67189,I66838,I67220,I117583,I67237,I67254,I67271,I66847,I67302,I66835,I66844,I66832,I67388,I368370,I67414,I67422,I67439,I368361,I368379,I67456,I368358,I67482,I67499,I67507,I368364,I67524,I67356,I67555,I67572,I67368,I67612,I67377,I67634,I368376,I368367,I67651,I368382,I67677,I67694,I67380,I67716,I67365,I67747,I368373,I67764,I67781,I67798,I67374,I67829,I67362,I67371,I67359,I67915,I694979,I67941,I67949,I67966,I694985,I695003,I67983,I695000,I68009,I694997,I68026,I68034,I694991,I68051,I67883,I68082,I68099,I67895,I68139,I67904,I68161,I694994,I694982,I68178,I695006,I68204,I68221,I67907,I68243,I67892,I68274,I694988,I68291,I68308,I68325,I67901,I68356,I67889,I67898,I67886,I68442,I177730,I68468,I68476,I68493,I177712,I177727,I68510,I177703,I68536,I177706,I68553,I68561,I177721,I68578,I68410,I68609,I68626,I68422,I177724,I68666,I68431,I68688,I177715,I68705,I177709,I68731,I68748,I68434,I68770,I68419,I68801,I177718,I68818,I68835,I68852,I68428,I68883,I68416,I68425,I68413,I68969,I574608,I68995,I69003,I69020,I574623,I574602,I69037,I574605,I69063,I574626,I69080,I69088,I69105,I68937,I69136,I69153,I68949,I69193,I68958,I69215,I574614,I574611,I69232,I574617,I69258,I69275,I68961,I69297,I68946,I69328,I574620,I69345,I69362,I69379,I68955,I69410,I68943,I68952,I68940,I69496,I193540,I69522,I69530,I69547,I193522,I193537,I69564,I193513,I69590,I193516,I69607,I69615,I193531,I69632,I69464,I69663,I69680,I69476,I193534,I69720,I69485,I69742,I193525,I69759,I193519,I69785,I69802,I69488,I69824,I69473,I69855,I193528,I69872,I69889,I69906,I69482,I69937,I69470,I69479,I69467,I70023,I131271,I70049,I70057,I70074,I131265,I131259,I70091,I131280,I70117,I131277,I70134,I70142,I131274,I70159,I69991,I70190,I70207,I70003,I70247,I70012,I70269,I131262,I70286,I131283,I70312,I70329,I70015,I70351,I70000,I70382,I131268,I70399,I70416,I70433,I70009,I70464,I69997,I70006,I69994,I70550,I652332,I70576,I70584,I70601,I652326,I652347,I70618,I652338,I70644,I652329,I70661,I70669,I652341,I70686,I70518,I70717,I70734,I70530,I70774,I70539,I70796,I652350,I652335,I70813,I70839,I70856,I70542,I70878,I70527,I70909,I652344,I70926,I70943,I70960,I70536,I70991,I70524,I70533,I70521,I71077,I592526,I71103,I71111,I71128,I592541,I592520,I71145,I592523,I71171,I592544,I71188,I71196,I71213,I71045,I71244,I71261,I71057,I71301,I71066,I71323,I592532,I592529,I71340,I592535,I71366,I71383,I71069,I71405,I71054,I71436,I592538,I71453,I71470,I71487,I71063,I71518,I71051,I71060,I71048,I71604,I199337,I71630,I71638,I71655,I199319,I199334,I71672,I199310,I71698,I199313,I71715,I71723,I199328,I71740,I71572,I71771,I71788,I71584,I199331,I71828,I71593,I71850,I199322,I71867,I199316,I71893,I71910,I71596,I71932,I71581,I71963,I199325,I71980,I71997,I72014,I71590,I72045,I71578,I71587,I71575,I72131,I348718,I72157,I72165,I72182,I348709,I348727,I72199,I348706,I72225,I72242,I72250,I348712,I72267,I72099,I72298,I72315,I72111,I72355,I72120,I72377,I348724,I348715,I72394,I348730,I72420,I72437,I72123,I72459,I72108,I72490,I348721,I72507,I72524,I72541,I72117,I72572,I72105,I72114,I72102,I72658,I533573,I72684,I72692,I72709,I533591,I533585,I72726,I533564,I72752,I533582,I72769,I72777,I533567,I72794,I72626,I72825,I72842,I72638,I533579,I72882,I72647,I72904,I533588,I533576,I72921,I533570,I72947,I72964,I72650,I72986,I72635,I73017,I73034,I73051,I73068,I72644,I73099,I72632,I72641,I72629,I73185,I152434,I73211,I73219,I73236,I152416,I152431,I73253,I152407,I73279,I152410,I73296,I73304,I152425,I73321,I73153,I73352,I73369,I73165,I152428,I73409,I73174,I73431,I152419,I73448,I152413,I73474,I73491,I73177,I73513,I73162,I73544,I152422,I73561,I73578,I73595,I73171,I73626,I73159,I73168,I73156,I73712,I248407,I73738,I73746,I73763,I248401,I248392,I73780,I248413,I73806,I248395,I73823,I73831,I248389,I73848,I73680,I73879,I73896,I73692,I73936,I73701,I73958,I248416,I248398,I73975,I248404,I74001,I74018,I73704,I74040,I73689,I74071,I248410,I74088,I74105,I74122,I73698,I74153,I73686,I73695,I73683,I74239,I441416,I74265,I74273,I74290,I441413,I441428,I74307,I441410,I74333,I441407,I74350,I74358,I74375,I74406,I74423,I74463,I74485,I441422,I74502,I441425,I74528,I74545,I74567,I74598,I441419,I74615,I74632,I74649,I74680,I74769,I287688,I74795,I74803,I287694,I74829,I74837,I287676,I74854,I287700,I74871,I74746,I74902,I287691,I74740,I74933,I287682,I74950,I74967,I287685,I287679,I74984,I75001,I75018,I74755,I74752,I74758,I75077,I75094,I75111,I287697,I75137,I74737,I75168,I75176,I74761,I75207,I75224,I75241,I74743,I75272,I75289,I74734,I74749,I75364,I130688,I75390,I75398,I130682,I75424,I75432,I130667,I75449,I130676,I75466,I75341,I75497,I130664,I75335,I75528,I130670,I75545,I75562,I130673,I130685,I75579,I75596,I75613,I75350,I75347,I75353,I75672,I75689,I75706,I130679,I75732,I75332,I75763,I75771,I75356,I75802,I75819,I75836,I75338,I75867,I75884,I75329,I75344,I75959,I107483,I75985,I75993,I107477,I76019,I76027,I107462,I76044,I107471,I76061,I75936,I76092,I107459,I75930,I76123,I107465,I76140,I76157,I107468,I107480,I76174,I76191,I76208,I75945,I75942,I75948,I76267,I76284,I76301,I107474,I76327,I75927,I76358,I76366,I75951,I76397,I76414,I76431,I75933,I76462,I76479,I75924,I75939,I76554,I249501,I76580,I76588,I249495,I76614,I76622,I249492,I76639,I249483,I76656,I76687,I249486,I76718,I249489,I76735,I76752,I249477,I249504,I76769,I76786,I76803,I76862,I76879,I76896,I249480,I76922,I76953,I76961,I249498,I76992,I77009,I77026,I77057,I77074,I77149,I494164,I77175,I77183,I494185,I77209,I77217,I494167,I77234,I494158,I77251,I77126,I77282,I494170,I77120,I77313,I494161,I77330,I77347,I494179,I494182,I77364,I77381,I77398,I77135,I77132,I77138,I77457,I77474,I77491,I494173,I494176,I77517,I77117,I77548,I77556,I77141,I77587,I77604,I77621,I77123,I77652,I77669,I77114,I77129,I77744,I374138,I77770,I77778,I374159,I77804,I77812,I77829,I374150,I77846,I77721,I77877,I374147,I77715,I77908,I374156,I77925,I77942,I374141,I77959,I77976,I77993,I77730,I77727,I77733,I78052,I78069,I78086,I374162,I374144,I78112,I77712,I78143,I78151,I374153,I77736,I78182,I78199,I78216,I77718,I78247,I78264,I77709,I77724,I78339,I342926,I78365,I78373,I342947,I78399,I78407,I78424,I342938,I78441,I78316,I78472,I342935,I78310,I78503,I342944,I78520,I78537,I342929,I78554,I78571,I78588,I78325,I78322,I78328,I78647,I78664,I78681,I342950,I342932,I78707,I78307,I78738,I78746,I342941,I78331,I78777,I78794,I78811,I78313,I78842,I78859,I78304,I78319,I78931,I698434,I78957,I78974,I78923,I78996,I698425,I79022,I79030,I79047,I698419,I79064,I698413,I79081,I79098,I698440,I79115,I79132,I698437,I79149,I78899,I79180,I79197,I79214,I79231,I78911,I78905,I79276,I698422,I78920,I78914,I79321,I79338,I698428,I79355,I698431,I79372,I698416,I79398,I79406,I78908,I78902,I79460,I79468,I78917,I79526,I576914,I79552,I79569,I79518,I79591,I79617,I79625,I79642,I576917,I79659,I576929,I79676,I79693,I576935,I79710,I576926,I79727,I576932,I79744,I79494,I79775,I79792,I79809,I79826,I79506,I79500,I79871,I576923,I79515,I79509,I79916,I79933,I576920,I79950,I576938,I79967,I79993,I80001,I79503,I79497,I80055,I80063,I79512,I80121,I509677,I80147,I80164,I80113,I80186,I509686,I80212,I80220,I80237,I509674,I80254,I509665,I80271,I80288,I509671,I80305,I509689,I80322,I509662,I80339,I80089,I80370,I80387,I80404,I80421,I80101,I80095,I80466,I509668,I80110,I80104,I80511,I80528,I509680,I80545,I80562,I509683,I80588,I80596,I80098,I80092,I80650,I80658,I80107,I80716,I673647,I80742,I80759,I80781,I673659,I80807,I80815,I80832,I673653,I80849,I673665,I80866,I80883,I673650,I80900,I673662,I80917,I673644,I80934,I80965,I80982,I80999,I81016,I81061,I673656,I81106,I81123,I81140,I81157,I673668,I81183,I81191,I81245,I81253,I81311,I235901,I81337,I81354,I81303,I81376,I235889,I81402,I81410,I81427,I235898,I81444,I235895,I81461,I81478,I235886,I81495,I235892,I81512,I235877,I81529,I81279,I81560,I81577,I81594,I81611,I81291,I81285,I81656,I81300,I81294,I81701,I81718,I235883,I81735,I235880,I81752,I235904,I81778,I81786,I81288,I81282,I81840,I81848,I81297,I81906,I188243,I81932,I81949,I81898,I81971,I188258,I81997,I82005,I82022,I188255,I82039,I82056,I82073,I188252,I82090,I188267,I82107,I188264,I82124,I81874,I82155,I82172,I82189,I82206,I81886,I81880,I82251,I188261,I81895,I81889,I82296,I82313,I188249,I82330,I188270,I82347,I188246,I82373,I82381,I81883,I81877,I82435,I82443,I81892,I82501,I424022,I82527,I82544,I82493,I82566,I424016,I82592,I82600,I82617,I424034,I82634,I82651,I82668,I82685,I424028,I82702,I424019,I82719,I82469,I82750,I82767,I82784,I82801,I82481,I82475,I82846,I424031,I82490,I82484,I82891,I82908,I424037,I82925,I82942,I424025,I82968,I82976,I82478,I82472,I83030,I83038,I82487,I83096,I363168,I83122,I83139,I83088,I83161,I363165,I83187,I83195,I83212,I363171,I83229,I363156,I83246,I83263,I363159,I83280,I363180,I83297,I363177,I83314,I83064,I83345,I83362,I83379,I83396,I83076,I83070,I83441,I83085,I83079,I83486,I83503,I363162,I83520,I363174,I83537,I83563,I83571,I83073,I83067,I83625,I83633,I83082,I83691,I83717,I83734,I83683,I83756,I83782,I83790,I83807,I83824,I83841,I83858,I83875,I83892,I83909,I83659,I83940,I83957,I83974,I83991,I83671,I83665,I84036,I83680,I83674,I84081,I84098,I84115,I84132,I84158,I84166,I83668,I83662,I84220,I84228,I83677,I84286,I693323,I84312,I84329,I84278,I84351,I693296,I84377,I84385,I84402,I693320,I84419,I693317,I84436,I84453,I84470,I693314,I84487,I693302,I84504,I84254,I84535,I84552,I84569,I84586,I84266,I84260,I84631,I693308,I84275,I84269,I84676,I84693,I693311,I84710,I693299,I84727,I693305,I84753,I84761,I84263,I84257,I84815,I84823,I84272,I84881,I530995,I84907,I84924,I84873,I84946,I531004,I84972,I84980,I84997,I530992,I85014,I530983,I85031,I85048,I530989,I85065,I531007,I85082,I530980,I85099,I84849,I85130,I85147,I85164,I85181,I84861,I84855,I85226,I530986,I84870,I84864,I85271,I85288,I530998,I85305,I85322,I531001,I85348,I85356,I84858,I84852,I85410,I85418,I84867,I85476,I503217,I85502,I85519,I85468,I85541,I503226,I85567,I85575,I85592,I503214,I85609,I503205,I85626,I85643,I503211,I85660,I503229,I85677,I503202,I85694,I85444,I85725,I85742,I85759,I85776,I85456,I85450,I85821,I503208,I85465,I85459,I85866,I85883,I503220,I85900,I85917,I503223,I85943,I85951,I85453,I85447,I86005,I86013,I85462,I86071,I325023,I86097,I86114,I86063,I86136,I325014,I86162,I86170,I86187,I325032,I86204,I325029,I86221,I86238,I325008,I86255,I325011,I86272,I325020,I86289,I86039,I86320,I86337,I86354,I86371,I86051,I86045,I86416,I325026,I86060,I86054,I86461,I86478,I86495,I325017,I86512,I86538,I86546,I86048,I86042,I86600,I86608,I86057,I86666,I632402,I86692,I86709,I86658,I86731,I86757,I86765,I86782,I632405,I86799,I632417,I86816,I86833,I632423,I86850,I632414,I86867,I632420,I86884,I86634,I86915,I86932,I86949,I86966,I86646,I86640,I87011,I632411,I86655,I86649,I87056,I87073,I632408,I87090,I632426,I87107,I87133,I87141,I86643,I86637,I87195,I87203,I86652,I87261,I155042,I87287,I87304,I87253,I87326,I155057,I87352,I87360,I87377,I155054,I87394,I87411,I87428,I155051,I87445,I155066,I87462,I155063,I87479,I87229,I87510,I87527,I87544,I87561,I87241,I87235,I87606,I155060,I87250,I87244,I87651,I87668,I155048,I87685,I155069,I87702,I155045,I87728,I87736,I87238,I87232,I87790,I87798,I87247,I87856,I728184,I87882,I87899,I87848,I87921,I728175,I87947,I87955,I87972,I728169,I87989,I728163,I88006,I88023,I728190,I88040,I88057,I728187,I88074,I87824,I88105,I88122,I88139,I88156,I87836,I87830,I88201,I728172,I87845,I87839,I88246,I88263,I728178,I88280,I728181,I88297,I728166,I88323,I88331,I87833,I87827,I88385,I88393,I87842,I88451,I88477,I88494,I88443,I88516,I88542,I88550,I88567,I88584,I88601,I88618,I88635,I88652,I88669,I88419,I88700,I88717,I88734,I88751,I88431,I88425,I88796,I88440,I88434,I88841,I88858,I88875,I88892,I88918,I88926,I88428,I88422,I88980,I88988,I88437,I89046,I89072,I89089,I89038,I89111,I89137,I89145,I89162,I89179,I89196,I89213,I89230,I89247,I89264,I89014,I89295,I89312,I89329,I89346,I89026,I89020,I89391,I89035,I89029,I89436,I89453,I89470,I89487,I89513,I89521,I89023,I89017,I89575,I89583,I89032,I89641,I709739,I89667,I89684,I89706,I709730,I89732,I89740,I89757,I709724,I89774,I709718,I89791,I89808,I709745,I89825,I89842,I709742,I89859,I89890,I89907,I89924,I89941,I89986,I709727,I90031,I90048,I709733,I90065,I709736,I90082,I709721,I90108,I90116,I90170,I90178,I90236,I744249,I90262,I90279,I90228,I90301,I744240,I90327,I90335,I90352,I744234,I90369,I744228,I90386,I90403,I744255,I90420,I90437,I744252,I90454,I90204,I90485,I90502,I90519,I90536,I90216,I90210,I90581,I744237,I90225,I90219,I90626,I90643,I744243,I90660,I744246,I90677,I744231,I90703,I90711,I90213,I90207,I90765,I90773,I90222,I90831,I499987,I90857,I90874,I90823,I90896,I499996,I90922,I90930,I90947,I499984,I90964,I499975,I90981,I90998,I499981,I91015,I499999,I91032,I499972,I91049,I90799,I91080,I91097,I91114,I91131,I90811,I90805,I91176,I499978,I90820,I90814,I91221,I91238,I499990,I91255,I91272,I499993,I91298,I91306,I90808,I90802,I91360,I91368,I90817,I91426,I675959,I91452,I91469,I91418,I91491,I675971,I91517,I91525,I91542,I675965,I91559,I675977,I91576,I91593,I675962,I91610,I675974,I91627,I675956,I91644,I91394,I91675,I91692,I91709,I91726,I91406,I91400,I91771,I675968,I91415,I91409,I91816,I91833,I91850,I91867,I675980,I91893,I91901,I91403,I91397,I91955,I91963,I91412,I92021,I92047,I92064,I92013,I92086,I92112,I92120,I92137,I92154,I92171,I92188,I92205,I92222,I92239,I91989,I92270,I92287,I92304,I92321,I92001,I91995,I92366,I92010,I92004,I92411,I92428,I92445,I92462,I92488,I92496,I91998,I91992,I92550,I92558,I92007,I92616,I479961,I92642,I92659,I92608,I92681,I479970,I92707,I92715,I92732,I479958,I92749,I479949,I92766,I92783,I479955,I92800,I479973,I92817,I479946,I92834,I92584,I92865,I92882,I92899,I92916,I92596,I92590,I92961,I479952,I92605,I92599,I93006,I93023,I479964,I93040,I93057,I479967,I93083,I93091,I92593,I92587,I93145,I93153,I92602,I93211,I547609,I93237,I93254,I93203,I93276,I547618,I93302,I93310,I93327,I547612,I93344,I547606,I93361,I93378,I547621,I93395,I93412,I547615,I93429,I93179,I93460,I93477,I93494,I93511,I93191,I93185,I93556,I93200,I93194,I93601,I93618,I547627,I93635,I547624,I93652,I93678,I93686,I93188,I93182,I93740,I93748,I93197,I93806,I334849,I93832,I93849,I93798,I93871,I334840,I93897,I93905,I93922,I334858,I93939,I334855,I93956,I93973,I334834,I93990,I334837,I94007,I334846,I94024,I93774,I94055,I94072,I94089,I94106,I93786,I93780,I94151,I334852,I93795,I93789,I94196,I94213,I94230,I334843,I94247,I94273,I94281,I93783,I93777,I94335,I94343,I93792,I94401,I357966,I94427,I94444,I94393,I94466,I357963,I94492,I94500,I94517,I357969,I94534,I357954,I94551,I94568,I357957,I94585,I357978,I94602,I357975,I94619,I94369,I94650,I94667,I94684,I94701,I94381,I94375,I94746,I94390,I94384,I94791,I94808,I357960,I94825,I357972,I94842,I94868,I94876,I94378,I94372,I94930,I94938,I94387,I94996,I219336,I95022,I95039,I94988,I95061,I219351,I95087,I95095,I95112,I219348,I95129,I95146,I95163,I219345,I95180,I219360,I95197,I219357,I95214,I94964,I95245,I95262,I95279,I95296,I94976,I94970,I95341,I219354,I94985,I94979,I95386,I95403,I219342,I95420,I219363,I95437,I219339,I95463,I95471,I94973,I94967,I95525,I95533,I94982,I95591,I722234,I95617,I95634,I95583,I95656,I722225,I95682,I95690,I95707,I722219,I95724,I722213,I95741,I95758,I722240,I95775,I95792,I722237,I95809,I95559,I95840,I95857,I95874,I95891,I95571,I95565,I95936,I722222,I95580,I95574,I95981,I95998,I722228,I96015,I722231,I96032,I722216,I96058,I96066,I95568,I95562,I96120,I96128,I95577,I96186,I161893,I96212,I96229,I96178,I96251,I161908,I96277,I96285,I96302,I161905,I96319,I96336,I96353,I161902,I96370,I161917,I96387,I161914,I96404,I96154,I96435,I96452,I96469,I96486,I96166,I96160,I96531,I161911,I96175,I96169,I96576,I96593,I161899,I96610,I161920,I96627,I161896,I96653,I96661,I96163,I96157,I96715,I96723,I96172,I96781,I162947,I96807,I96824,I96773,I96846,I162962,I96872,I96880,I96897,I162959,I96914,I96931,I96948,I162956,I96965,I162971,I96982,I162968,I96999,I96749,I97030,I97047,I97064,I97081,I96761,I96755,I97126,I162965,I96770,I96764,I97171,I97188,I162953,I97205,I162974,I97222,I162950,I97248,I97256,I96758,I96752,I97310,I97318,I96767,I97376,I666488,I97402,I97419,I97368,I97441,I666473,I97467,I97475,I97492,I666491,I97509,I97526,I97543,I666494,I97560,I666485,I97577,I666482,I97594,I97344,I97625,I97642,I97659,I97676,I97356,I97350,I97721,I666479,I97365,I97359,I97766,I97783,I666470,I97800,I666476,I97817,I97843,I97851,I97353,I97347,I97905,I97913,I97362,I97971,I633558,I97997,I98014,I97963,I98036,I98062,I98070,I98087,I633561,I98104,I633573,I98121,I98138,I633579,I98155,I633570,I98172,I633576,I98189,I97939,I98220,I98237,I98254,I98271,I97951,I97945,I98316,I633567,I97960,I97954,I98361,I98378,I633564,I98395,I633582,I98412,I98438,I98446,I97948,I97942,I98500,I98508,I97957,I98566,I617374,I98592,I98609,I98558,I98631,I98657,I98665,I98682,I617377,I98699,I617389,I98716,I98733,I617395,I98750,I617386,I98767,I617392,I98784,I98534,I98815,I98832,I98849,I98866,I98546,I98540,I98911,I617383,I98555,I98549,I98956,I98973,I617380,I98990,I617398,I99007,I99033,I99041,I98543,I98537,I99095,I99103,I98552,I99161,I531641,I99187,I99204,I99153,I99226,I531650,I99252,I99260,I99277,I531638,I99294,I531629,I99311,I99328,I531635,I99345,I531653,I99362,I531626,I99379,I99129,I99410,I99427,I99444,I99461,I99141,I99135,I99506,I531632,I99150,I99144,I99551,I99568,I531644,I99585,I99602,I531647,I99628,I99636,I99138,I99132,I99690,I99698,I99147,I99756,I593676,I99782,I99799,I99748,I99821,I99847,I99855,I99872,I593679,I99889,I593691,I99906,I99923,I593697,I99940,I593688,I99957,I593694,I99974,I99724,I100005,I100022,I100039,I100056,I99736,I99730,I100101,I593685,I99745,I99739,I100146,I100163,I593682,I100180,I593700,I100197,I100223,I100231,I99733,I99727,I100285,I100293,I99742,I100351,I100377,I100394,I100343,I100416,I100442,I100450,I100467,I100484,I100501,I100518,I100535,I100552,I100569,I100319,I100600,I100617,I100634,I100651,I100331,I100325,I100696,I100340,I100334,I100741,I100758,I100775,I100792,I100818,I100826,I100328,I100322,I100880,I100888,I100337,I100946,I409986,I100972,I100989,I100938,I101011,I409983,I101037,I101045,I101062,I409989,I101079,I409974,I101096,I101113,I409977,I101130,I409998,I101147,I409995,I101164,I100914,I101195,I101212,I101229,I101246,I100926,I100920,I101291,I100935,I100929,I101336,I101353,I409980,I101370,I409992,I101387,I101413,I101421,I100923,I100917,I101475,I101483,I100932,I101541,I351608,I101567,I101584,I101533,I101606,I351605,I101632,I101640,I101657,I351611,I101674,I351596,I101691,I101708,I351599,I101725,I351620,I101742,I351617,I101759,I101509,I101790,I101807,I101824,I101841,I101521,I101515,I101886,I101530,I101524,I101931,I101948,I351602,I101965,I351614,I101982,I102008,I102016,I101518,I101512,I102070,I102078,I101527,I102136,I396114,I102162,I102179,I102128,I102201,I396111,I102227,I102235,I102252,I396117,I102269,I396102,I102286,I102303,I396105,I102320,I396126,I102337,I396123,I102354,I102104,I102385,I102402,I102419,I102436,I102116,I102110,I102481,I102125,I102119,I102526,I102543,I396108,I102560,I396120,I102577,I102603,I102611,I102113,I102107,I102665,I102673,I102122,I102731,I445629,I102757,I102774,I102723,I102796,I445623,I102822,I102830,I102847,I445641,I102864,I102881,I102898,I102915,I445635,I102932,I445626,I102949,I102699,I102980,I102997,I103014,I103031,I102711,I102705,I103076,I445638,I102720,I102714,I103121,I103138,I445644,I103155,I103172,I445632,I103198,I103206,I102708,I102702,I103260,I103268,I102717,I103326,I103352,I103369,I103318,I103391,I103417,I103425,I103442,I103459,I103476,I103493,I103510,I103527,I103544,I103294,I103575,I103592,I103609,I103626,I103306,I103300,I103671,I103315,I103309,I103716,I103733,I103750,I103767,I103793,I103801,I103303,I103297,I103855,I103863,I103312,I103921,I261469,I103947,I103964,I103913,I103986,I261457,I104012,I104020,I104037,I261466,I104054,I261463,I104071,I104088,I261454,I104105,I261460,I104122,I261445,I104139,I103889,I104170,I104187,I104204,I104221,I103901,I103895,I104266,I103910,I103904,I104311,I104328,I261451,I104345,I261448,I104362,I261472,I104388,I104396,I103898,I103892,I104450,I104458,I103907,I104516,I104542,I104559,I104508,I104581,I104607,I104615,I104632,I104649,I104666,I104683,I104700,I104717,I104734,I104484,I104765,I104782,I104799,I104816,I104496,I104490,I104861,I104505,I104499,I104906,I104923,I104940,I104957,I104983,I104991,I104493,I104487,I105045,I105053,I104502,I105111,I245693,I105137,I105154,I105176,I245681,I105202,I105210,I105227,I245690,I105244,I245687,I105261,I105278,I245678,I105295,I245684,I105312,I245669,I105329,I105360,I105377,I105394,I105411,I105456,I105501,I105518,I245675,I105535,I245672,I105552,I245696,I105578,I105586,I105640,I105648,I105706,I105732,I105749,I105698,I105771,I105797,I105805,I105822,I105839,I105856,I105873,I105890,I105907,I105924,I105674,I105955,I105972,I105989,I106006,I105686,I105680,I106051,I105695,I105689,I106096,I106113,I106130,I106147,I106173,I106181,I105683,I105677,I106235,I106243,I105692,I106301,I106327,I106344,I106293,I106366,I106392,I106400,I106417,I106434,I106451,I106468,I106485,I106502,I106519,I106269,I106550,I106567,I106584,I106601,I106281,I106275,I106646,I106290,I106284,I106691,I106708,I106725,I106742,I106768,I106776,I106278,I106272,I106830,I106838,I106287,I106896,I567805,I106922,I106939,I106888,I106961,I567814,I106987,I106995,I107012,I567808,I107029,I567802,I107046,I107063,I567817,I107080,I107097,I567811,I107114,I106864,I107145,I107162,I107179,I107196,I106876,I106870,I107241,I106885,I106879,I107286,I107303,I567823,I107320,I567820,I107337,I107363,I107371,I106873,I106867,I107425,I107433,I106882,I107491,I415188,I107517,I107534,I107556,I415185,I107582,I107590,I107607,I415191,I107624,I415176,I107641,I107658,I415179,I107675,I415200,I107692,I415197,I107709,I107740,I107757,I107774,I107791,I107836,I107881,I107898,I415182,I107915,I415194,I107932,I107958,I107966,I108020,I108028,I108086,I411720,I108112,I108129,I108078,I108151,I411717,I108177,I108185,I108202,I411723,I108219,I411708,I108236,I108253,I411711,I108270,I411732,I108287,I411729,I108304,I108054,I108335,I108352,I108369,I108386,I108066,I108060,I108431,I108075,I108069,I108476,I108493,I411714,I108510,I411726,I108527,I108553,I108561,I108063,I108057,I108615,I108623,I108072,I108681,I271805,I108707,I108724,I108673,I108746,I271793,I108772,I108780,I108797,I271802,I108814,I271799,I108831,I108848,I271790,I108865,I271796,I108882,I271781,I108899,I108649,I108930,I108947,I108964,I108981,I108661,I108655,I109026,I108670,I108664,I109071,I109088,I271787,I109105,I271784,I109122,I271808,I109148,I109156,I108658,I108652,I109210,I109218,I108667,I109276,I680005,I109302,I109319,I109268,I109341,I680017,I109367,I109375,I109392,I680011,I109409,I680023,I109426,I109443,I680008,I109460,I680020,I109477,I680002,I109494,I109244,I109525,I109542,I109559,I109576,I109256,I109250,I109621,I680014,I109265,I109259,I109666,I109683,I109700,I109717,I680026,I109743,I109751,I109253,I109247,I109805,I109813,I109262,I109871,I231005,I109897,I109914,I109936,I230993,I109962,I109970,I109987,I231002,I110004,I230999,I110021,I110038,I230990,I110055,I230996,I110072,I230981,I110089,I110120,I110137,I110154,I110171,I110216,I110261,I110278,I230987,I110295,I230984,I110312,I231008,I110338,I110346,I110400,I110408,I110466,I662680,I110492,I110509,I110458,I110531,I662665,I110557,I110565,I110582,I662683,I110599,I110616,I110633,I662686,I110650,I662677,I110667,I662674,I110684,I110434,I110715,I110732,I110749,I110766,I110446,I110440,I110811,I662671,I110455,I110449,I110856,I110873,I662662,I110890,I662668,I110907,I110933,I110941,I110443,I110437,I110995,I111003,I110452,I111061,I597722,I111087,I111104,I111126,I111152,I111160,I111177,I597725,I111194,I597737,I111211,I111228,I597743,I111245,I597734,I111262,I597740,I111279,I111310,I111327,I111344,I111361,I111406,I597731,I111451,I111468,I597728,I111485,I597746,I111502,I111528,I111536,I111590,I111598,I111656,I546487,I111682,I111699,I111648,I111721,I546496,I111747,I111755,I111772,I546490,I111789,I546484,I111806,I111823,I546499,I111840,I111857,I546493,I111874,I111624,I111905,I111922,I111939,I111956,I111636,I111630,I112001,I111645,I111639,I112046,I112063,I546505,I112080,I546502,I112097,I112123,I112131,I111633,I111627,I112185,I112193,I111642,I112251,I562756,I112277,I112294,I112243,I112316,I562765,I112342,I112350,I112367,I562759,I112384,I562753,I112401,I112418,I562768,I112435,I112452,I562762,I112469,I112219,I112500,I112517,I112534,I112551,I112231,I112225,I112596,I112240,I112234,I112641,I112658,I562774,I112675,I562771,I112692,I112718,I112726,I112228,I112222,I112780,I112788,I112237,I112846,I520013,I112872,I112889,I112838,I112911,I520022,I112937,I112945,I112962,I520010,I112979,I520001,I112996,I113013,I520007,I113030,I520025,I113047,I519998,I113064,I112814,I113095,I113112,I113129,I113146,I112826,I112820,I113191,I520004,I112835,I112829,I113236,I113253,I520016,I113270,I113287,I520019,I113313,I113321,I112823,I112817,I113375,I113383,I112832,I113441,I558829,I113467,I113484,I113433,I113506,I558838,I113532,I113540,I113557,I558832,I113574,I558826,I113591,I113608,I558841,I113625,I113642,I558835,I113659,I113409,I113690,I113707,I113724,I113741,I113421,I113415,I113786,I113430,I113424,I113831,I113848,I558847,I113865,I558844,I113882,I113908,I113916,I113418,I113412,I113970,I113978,I113427,I114036,I114062,I114079,I114028,I114101,I114127,I114135,I114152,I114169,I114186,I114203,I114220,I114237,I114254,I114004,I114285,I114302,I114319,I114336,I114016,I114010,I114381,I114025,I114019,I114426,I114443,I114460,I114477,I114503,I114511,I114013,I114007,I114565,I114573,I114022,I114631,I635292,I114657,I114674,I114623,I114696,I114722,I114730,I114747,I635295,I114764,I635307,I114781,I114798,I635313,I114815,I635304,I114832,I635310,I114849,I114599,I114880,I114897,I114914,I114931,I114611,I114605,I114976,I635301,I114620,I114614,I115021,I115038,I635298,I115055,I635316,I115072,I115098,I115106,I114608,I114602,I115160,I115168,I114617,I115226,I623732,I115252,I115269,I115218,I115291,I115317,I115325,I115342,I623735,I115359,I623747,I115376,I115393,I623753,I115410,I623744,I115427,I623750,I115444,I115194,I115475,I115492,I115509,I115526,I115206,I115200,I115571,I623741,I115215,I115209,I115616,I115633,I623738,I115650,I623756,I115667,I115693,I115701,I115203,I115197,I115755,I115763,I115212,I115821,I426657,I115847,I115864,I115813,I115886,I426651,I115912,I115920,I115937,I426669,I115954,I115971,I115988,I116005,I426663,I116022,I426654,I116039,I115789,I116070,I116087,I116104,I116121,I115801,I115795,I116166,I426666,I115810,I115804,I116211,I116228,I426672,I116245,I116262,I426660,I116288,I116296,I115798,I115792,I116350,I116358,I115807,I116416,I327913,I116442,I116459,I116481,I327904,I116507,I116515,I116532,I327922,I116549,I327919,I116566,I116583,I327898,I116600,I327901,I116617,I327910,I116634,I116665,I116682,I116699,I116716,I116761,I327916,I116806,I116823,I116840,I327907,I116857,I116883,I116891,I116945,I116953,I117011,I396692,I117037,I117054,I117003,I117076,I396689,I117102,I117110,I117127,I396695,I117144,I396680,I117161,I117178,I396683,I117195,I396704,I117212,I396701,I117229,I116979,I117260,I117277,I117294,I117311,I116991,I116985,I117356,I117000,I116994,I117401,I117418,I396686,I117435,I396698,I117452,I117478,I117486,I116988,I116982,I117540,I117548,I116997,I117606,I366636,I117632,I117649,I117671,I366633,I117697,I117705,I117722,I366639,I117739,I366624,I117756,I117773,I366627,I117790,I366648,I117807,I366645,I117824,I117855,I117872,I117889,I117906,I117951,I117996,I118013,I366630,I118030,I366642,I118047,I118073,I118081,I118135,I118143,I118201,I564439,I118227,I118244,I118193,I118266,I564448,I118292,I118300,I118317,I564442,I118334,I564436,I118351,I118368,I564451,I118385,I118402,I564445,I118419,I118169,I118450,I118467,I118484,I118501,I118181,I118175,I118546,I118190,I118184,I118591,I118608,I564457,I118625,I564454,I118642,I118668,I118676,I118178,I118172,I118730,I118738,I118187,I118796,I236445,I118822,I118839,I118861,I236433,I118887,I118895,I118912,I236442,I118929,I236439,I118946,I118963,I236430,I118980,I236436,I118997,I236421,I119014,I119045,I119062,I119079,I119096,I119141,I119186,I119203,I236427,I119220,I236424,I119237,I236448,I119263,I119271,I119325,I119333,I119391,I583272,I119417,I119434,I119456,I119482,I119490,I119507,I583275,I119524,I583287,I119541,I119558,I583293,I119575,I583284,I119592,I583290,I119609,I119640,I119657,I119674,I119691,I119736,I583281,I119781,I119798,I583278,I119815,I583296,I119832,I119858,I119866,I119920,I119928,I119986,I384554,I120012,I120029,I119978,I120051,I384551,I120077,I120085,I120102,I384557,I120119,I384542,I120136,I120153,I384545,I120170,I384566,I120187,I384563,I120204,I119954,I120235,I120252,I120269,I120286,I119966,I119960,I120331,I119975,I119969,I120376,I120393,I384548,I120410,I384560,I120427,I120453,I120461,I119963,I119957,I120515,I120523,I119972,I120581,I629512,I120607,I120624,I120573,I120646,I120672,I120680,I120697,I629515,I120714,I629527,I120731,I120748,I629533,I120765,I629524,I120782,I629530,I120799,I120549,I120830,I120847,I120864,I120881,I120561,I120555,I120926,I629521,I120570,I120564,I120971,I120988,I629518,I121005,I629536,I121022,I121048,I121056,I120558,I120552,I121110,I121118,I120567,I121176,I121202,I121219,I121168,I121241,I121267,I121275,I121292,I121309,I121326,I121343,I121360,I121377,I121394,I121144,I121425,I121442,I121459,I121476,I121156,I121150,I121521,I121165,I121159,I121566,I121583,I121600,I121617,I121643,I121651,I121153,I121147,I121705,I121713,I121162,I121771,I726399,I121797,I121814,I121836,I726390,I121862,I121870,I121887,I726384,I121904,I726378,I121921,I121938,I726405,I121955,I121972,I726402,I121989,I122020,I122037,I122054,I122071,I122116,I726387,I122161,I122178,I726393,I122195,I726396,I122212,I726381,I122238,I122246,I122300,I122308,I122366,I122392,I122409,I122358,I122431,I122457,I122465,I122482,I122499,I122516,I122533,I122550,I122567,I122584,I122334,I122615,I122632,I122649,I122666,I122346,I122340,I122711,I122355,I122349,I122756,I122773,I122790,I122807,I122833,I122841,I122343,I122337,I122895,I122903,I122352,I122961,I122987,I123004,I122953,I123026,I123052,I123060,I123077,I123094,I123111,I123128,I123145,I123162,I123179,I122929,I123210,I123227,I123244,I123261,I122941,I122935,I123306,I122950,I122944,I123351,I123368,I123385,I123402,I123428,I123436,I122938,I122932,I123490,I123498,I122947,I123556,I548170,I123582,I123599,I123548,I123621,I548179,I123647,I123655,I123672,I548173,I123689,I548167,I123706,I123723,I548182,I123740,I123757,I548176,I123774,I123524,I123805,I123822,I123839,I123856,I123536,I123530,I123901,I123545,I123539,I123946,I123963,I548188,I123980,I548185,I123997,I124023,I124031,I123533,I123527,I124085,I124093,I123542,I124151,I317509,I124177,I124194,I124216,I317500,I124242,I124250,I124267,I317518,I124284,I317515,I124301,I124318,I317494,I124335,I317497,I124352,I317506,I124369,I124400,I124417,I124434,I124451,I124496,I317512,I124541,I124558,I124575,I317503,I124592,I124618,I124626,I124680,I124688,I124746,I618530,I124772,I124789,I124738,I124811,I124837,I124845,I124862,I618533,I124879,I618545,I124896,I124913,I618551,I124930,I618542,I124947,I618548,I124964,I124714,I124995,I125012,I125029,I125046,I124726,I124720,I125091,I618539,I124735,I124729,I125136,I125153,I618536,I125170,I618554,I125187,I125213,I125221,I124723,I124717,I125275,I125283,I124732,I125341,I349874,I125367,I125384,I125333,I125406,I349871,I125432,I125440,I125457,I349877,I125474,I349862,I125491,I125508,I349865,I125525,I349886,I125542,I349883,I125559,I125309,I125590,I125607,I125624,I125641,I125321,I125315,I125686,I125330,I125324,I125731,I125748,I349868,I125765,I349880,I125782,I125808,I125816,I125318,I125312,I125870,I125878,I125327,I125936,I125962,I125979,I125928,I126001,I126027,I126035,I126052,I126069,I126086,I126103,I126120,I126137,I126154,I125904,I126185,I126202,I126219,I126236,I125916,I125910,I126281,I125925,I125919,I126326,I126343,I126360,I126377,I126403,I126411,I125913,I125907,I126465,I126473,I125922,I126531,I402472,I126557,I126574,I126523,I126596,I402469,I126622,I126630,I126647,I402475,I126664,I402460,I126681,I126698,I402463,I126715,I402484,I126732,I402481,I126749,I126499,I126780,I126797,I126814,I126831,I126511,I126505,I126876,I126520,I126514,I126921,I126938,I402466,I126955,I402478,I126972,I126998,I127006,I126508,I126502,I127060,I127068,I126517,I127126,I367214,I127152,I127169,I127191,I367211,I127217,I127225,I127242,I367217,I127259,I367202,I127276,I127293,I367205,I127310,I367226,I127327,I367223,I127344,I127375,I127392,I127409,I127426,I127471,I127516,I127533,I367208,I127550,I367220,I127567,I127593,I127601,I127655,I127663,I127721,I227768,I127747,I127764,I127713,I127786,I227783,I127812,I127820,I127837,I227780,I127854,I127871,I127888,I227777,I127905,I227792,I127922,I227789,I127939,I127689,I127970,I127987,I128004,I128021,I127701,I127695,I128066,I227786,I127710,I127704,I128111,I128128,I227774,I128145,I227795,I128162,I227771,I128188,I128196,I127698,I127692,I128250,I128258,I127707,I128316,I128342,I128359,I128308,I128381,I128407,I128415,I128432,I128449,I128466,I128483,I128500,I128517,I128534,I128284,I128565,I128582,I128599,I128616,I128296,I128290,I128661,I128305,I128299,I128706,I128723,I128740,I128757,I128783,I128791,I128293,I128287,I128845,I128853,I128302,I128911,I469344,I128937,I128954,I128903,I128976,I469338,I129002,I129010,I129027,I469356,I129044,I129061,I129078,I129095,I469350,I129112,I469341,I129129,I128879,I129160,I129177,I129194,I129211,I128891,I128885,I129256,I469353,I128900,I128894,I129301,I129318,I469359,I129335,I129352,I469347,I129378,I129386,I128888,I128882,I129440,I129448,I128897,I129506,I418078,I129532,I129549,I129498,I129571,I418075,I129597,I129605,I129622,I418081,I129639,I418066,I129656,I129673,I418069,I129690,I418090,I129707,I418087,I129724,I129474,I129755,I129772,I129789,I129806,I129486,I129480,I129851,I129495,I129489,I129896,I129913,I418072,I129930,I418084,I129947,I129973,I129981,I129483,I129477,I130035,I130043,I129492,I130101,I517429,I130127,I130144,I130093,I130166,I517438,I130192,I130200,I130217,I517426,I130234,I517417,I130251,I130268,I517423,I130285,I517441,I130302,I517414,I130319,I130069,I130350,I130367,I130384,I130401,I130081,I130075,I130446,I517420,I130090,I130084,I130491,I130508,I517432,I130525,I130542,I517435,I130568,I130576,I130078,I130072,I130630,I130638,I130087,I130696,I230461,I130722,I130739,I130761,I230449,I130787,I130795,I130812,I230458,I130829,I230455,I130846,I130863,I230446,I130880,I230452,I130897,I230437,I130914,I130945,I130962,I130979,I130996,I131041,I131086,I131103,I230443,I131120,I230440,I131137,I230464,I131163,I131171,I131225,I131233,I131291,I435616,I131317,I131334,I131356,I435610,I131382,I131390,I131407,I435628,I131424,I131441,I131458,I131475,I435622,I131492,I435613,I131509,I131540,I131557,I131574,I131591,I131636,I435625,I131681,I131698,I435631,I131715,I131732,I435619,I131758,I131766,I131820,I131828,I131886,I131912,I131929,I131878,I131951,I131977,I131985,I132002,I132019,I132036,I132053,I132070,I132087,I132104,I131854,I132135,I132152,I132169,I132186,I131866,I131860,I132231,I131875,I131869,I132276,I132293,I132310,I132327,I132353,I132361,I131863,I131857,I132415,I132423,I131872,I132481,I632980,I132507,I132524,I132473,I132546,I132572,I132580,I132597,I632983,I132614,I632995,I132631,I132648,I633001,I132665,I632992,I132682,I632998,I132699,I132449,I132730,I132747,I132764,I132781,I132461,I132455,I132826,I632989,I132470,I132464,I132871,I132888,I632986,I132905,I633004,I132922,I132948,I132956,I132458,I132452,I133010,I133018,I132467,I133076,I290068,I133102,I133119,I133068,I133141,I290062,I133167,I133175,I133192,I290077,I133209,I290074,I133226,I133243,I290065,I133260,I290056,I133277,I290059,I133294,I133044,I133325,I133342,I133359,I133376,I133056,I133050,I133421,I290080,I133065,I133059,I133466,I133483,I290071,I133500,I133517,I133543,I133551,I133053,I133047,I133605,I133613,I133062,I133671,I527765,I133697,I133714,I133663,I133736,I527774,I133762,I133770,I133787,I527762,I133804,I527753,I133821,I133838,I527759,I133855,I527777,I133872,I527750,I133889,I133639,I133920,I133937,I133954,I133971,I133651,I133645,I134016,I527756,I133660,I133654,I134061,I134078,I527768,I134095,I134112,I527771,I134138,I134146,I133648,I133642,I134200,I134208,I133657,I134266,I161366,I134292,I134309,I134331,I161381,I134357,I134365,I134382,I161378,I134399,I134416,I134433,I161375,I134450,I161390,I134467,I161387,I134484,I134515,I134532,I134549,I134566,I134611,I161384,I134656,I134673,I161372,I134690,I161393,I134707,I161369,I134733,I134741,I134795,I134803,I134861,I187189,I134887,I134904,I134853,I134926,I187204,I134952,I134960,I134977,I187201,I134994,I135011,I135028,I187198,I135045,I187213,I135062,I187210,I135079,I134829,I135110,I135127,I135144,I135161,I134841,I134835,I135206,I187207,I134850,I134844,I135251,I135268,I187195,I135285,I187216,I135302,I187192,I135328,I135336,I134838,I134832,I135390,I135398,I134847,I135456,I501279,I135482,I135499,I135448,I135521,I501288,I135547,I135555,I135572,I501276,I135589,I501267,I135606,I135623,I501273,I135640,I501291,I135657,I501264,I135674,I135424,I135705,I135722,I135739,I135756,I135436,I135430,I135801,I501270,I135445,I135439,I135846,I135863,I501282,I135880,I135897,I501285,I135923,I135931,I135433,I135427,I135985,I135993,I135442,I136051,I156096,I136077,I136094,I136043,I136116,I156111,I136142,I136150,I136167,I156108,I136184,I136201,I136218,I156105,I136235,I156120,I136252,I156117,I136269,I136019,I136300,I136317,I136334,I136351,I136031,I136025,I136396,I156114,I136040,I136034,I136441,I136458,I156102,I136475,I156123,I136492,I156099,I136518,I136526,I136028,I136022,I136580,I136588,I136037,I136646,I194040,I136672,I136689,I136638,I136711,I194055,I136737,I136745,I136762,I194052,I136779,I136796,I136813,I194049,I136830,I194064,I136847,I194061,I136864,I136614,I136895,I136912,I136929,I136946,I136626,I136620,I136991,I194058,I136635,I136629,I137036,I137053,I194046,I137070,I194067,I137087,I194043,I137113,I137121,I136623,I136617,I137175,I137183,I136632,I137241,I266365,I137267,I137284,I137233,I137306,I266353,I137332,I137340,I137357,I266362,I137374,I266359,I137391,I137408,I266350,I137425,I266356,I137442,I266341,I137459,I137209,I137490,I137507,I137524,I137541,I137221,I137215,I137586,I137230,I137224,I137631,I137648,I266347,I137665,I266344,I137682,I266368,I137708,I137716,I137218,I137212,I137770,I137778,I137227,I137836,I178230,I137862,I137879,I137901,I178245,I137927,I137935,I137952,I178242,I137969,I137986,I138003,I178239,I138020,I178254,I138037,I178251,I138054,I138085,I138102,I138119,I138136,I138181,I178248,I138226,I138243,I178236,I138260,I178257,I138277,I178233,I138303,I138311,I138365,I138373,I138431,I589630,I138457,I138474,I138423,I138496,I138522,I138530,I138547,I589633,I138564,I589645,I138581,I138598,I589651,I138615,I589642,I138632,I589648,I138649,I138399,I138680,I138697,I138714,I138731,I138411,I138405,I138776,I589639,I138420,I138414,I138821,I138838,I589636,I138855,I589654,I138872,I138898,I138906,I138408,I138402,I138960,I138968,I138417,I139026,I664312,I139052,I139069,I139018,I139091,I664297,I139117,I139125,I139142,I664315,I139159,I139176,I139193,I664318,I139210,I664309,I139227,I664306,I139244,I138994,I139275,I139292,I139309,I139326,I139006,I139000,I139371,I664303,I139015,I139009,I139416,I139433,I664294,I139450,I664300,I139467,I139493,I139501,I139003,I138997,I139555,I139563,I139012,I139621,I648536,I139647,I139664,I139686,I648521,I139712,I139720,I139737,I648539,I139754,I139771,I139788,I648542,I139805,I648533,I139822,I648530,I139839,I139870,I139887,I139904,I139921,I139966,I648527,I140011,I140028,I648518,I140045,I648524,I140062,I140088,I140096,I140150,I140158,I140216,I155569,I140242,I140259,I140208,I140281,I155584,I140307,I140315,I140332,I155581,I140349,I140366,I140383,I155578,I140400,I155593,I140417,I155590,I140434,I140184,I140465,I140482,I140499,I140516,I140196,I140190,I140561,I155587,I140205,I140199,I140606,I140623,I155575,I140640,I155596,I140657,I155572,I140683,I140691,I140193,I140187,I140745,I140753,I140202,I140811,I463020,I140837,I140854,I140803,I140876,I463014,I140902,I140910,I140927,I463032,I140944,I140961,I140978,I140995,I463026,I141012,I463017,I141029,I140779,I141060,I141077,I141094,I141111,I140791,I140785,I141156,I463029,I140800,I140794,I141201,I141218,I463035,I141235,I141252,I463023,I141278,I141286,I140788,I140782,I141340,I141348,I140797,I141406,I667576,I141432,I141449,I141398,I141471,I667561,I141497,I141505,I141522,I667579,I141539,I141556,I141573,I667582,I141590,I667573,I141607,I667570,I141624,I141374,I141655,I141672,I141689,I141706,I141386,I141380,I141751,I667567,I141395,I141389,I141796,I141813,I667558,I141830,I667564,I141847,I141873,I141881,I141383,I141377,I141935,I141943,I141392,I142001,I590208,I142027,I142044,I141993,I142066,I142092,I142100,I142117,I590211,I142134,I590223,I142151,I142168,I590229,I142185,I590220,I142202,I590226,I142219,I141969,I142250,I142267,I142284,I142301,I141981,I141975,I142346,I590217,I141990,I141984,I142391,I142408,I590214,I142425,I590232,I142442,I142468,I142476,I141978,I141972,I142530,I142538,I141987,I142596,I296018,I142622,I142639,I142588,I142661,I296012,I142687,I142695,I142712,I296027,I142729,I296024,I142746,I142763,I296015,I142780,I296006,I142797,I296009,I142814,I142564,I142845,I142862,I142879,I142896,I142576,I142570,I142941,I296030,I142585,I142579,I142986,I143003,I296021,I143020,I143037,I143063,I143071,I142573,I142567,I143125,I143133,I142582,I143191,I143217,I143234,I143183,I143256,I143282,I143290,I143307,I143324,I143341,I143358,I143375,I143392,I143409,I143159,I143440,I143457,I143474,I143491,I143171,I143165,I143536,I143180,I143174,I143581,I143598,I143615,I143632,I143658,I143666,I143168,I143162,I143720,I143728,I143177,I143786,I143812,I143829,I143778,I143851,I143877,I143885,I143902,I143919,I143936,I143953,I143970,I143987,I144004,I143754,I144035,I144052,I144069,I144086,I143766,I143760,I144131,I143775,I143769,I144176,I144193,I144210,I144227,I144253,I144261,I143763,I143757,I144315,I144323,I143772,I144381,I401894,I144407,I144424,I144373,I144446,I401891,I144472,I144480,I144497,I401897,I144514,I401882,I144531,I144548,I401885,I144565,I401906,I144582,I401903,I144599,I144349,I144630,I144647,I144664,I144681,I144361,I144355,I144726,I144370,I144364,I144771,I144788,I401888,I144805,I401900,I144822,I144848,I144856,I144358,I144352,I144910,I144918,I144367,I144976,I409408,I145002,I145019,I144968,I145041,I409405,I145067,I145075,I145092,I409411,I145109,I409396,I145126,I145143,I409399,I145160,I409420,I145177,I409417,I145194,I144944,I145225,I145242,I145259,I145276,I144956,I144950,I145321,I144965,I144959,I145366,I145383,I409402,I145400,I409414,I145417,I145443,I145451,I144953,I144947,I145505,I145513,I144962,I145571,I375306,I145597,I145614,I145563,I145636,I375303,I145662,I145670,I145687,I375309,I145704,I375294,I145721,I145738,I375297,I145755,I375318,I145772,I375315,I145789,I145539,I145820,I145837,I145854,I145871,I145551,I145545,I145916,I145560,I145554,I145961,I145978,I375300,I145995,I375312,I146012,I146038,I146046,I145548,I145542,I146100,I146108,I145557,I146166,I474614,I146192,I146209,I146158,I146231,I474608,I146257,I146265,I146282,I474626,I146299,I146316,I146333,I146350,I474620,I146367,I474611,I146384,I146134,I146415,I146432,I146449,I146466,I146146,I146140,I146511,I474623,I146155,I146149,I146556,I146573,I474629,I146590,I146607,I474617,I146633,I146641,I146143,I146137,I146695,I146703,I146152,I146761,I146787,I146804,I146753,I146826,I146852,I146860,I146877,I146894,I146911,I146928,I146945,I146962,I146979,I146729,I147010,I147027,I147044,I147061,I146741,I146735,I147106,I146750,I146744,I147151,I147168,I147185,I147202,I147228,I147236,I146738,I146732,I147290,I147298,I146747,I147356,I693884,I147382,I147399,I147348,I147421,I693857,I147447,I147455,I147472,I693881,I147489,I693878,I147506,I147523,I147540,I693875,I147557,I693863,I147574,I147324,I147605,I147622,I147639,I147656,I147336,I147330,I147701,I693869,I147345,I147339,I147746,I147763,I693872,I147780,I693860,I147797,I693866,I147823,I147831,I147333,I147327,I147885,I147893,I147342,I147951,I630668,I147977,I147994,I147943,I148016,I148042,I148050,I148067,I630671,I148084,I630683,I148101,I148118,I630689,I148135,I630680,I148152,I630686,I148169,I147919,I148200,I148217,I148234,I148251,I147931,I147925,I148296,I630677,I147940,I147934,I148341,I148358,I630674,I148375,I630692,I148392,I148418,I148426,I147928,I147922,I148480,I148488,I147937,I148546,I510969,I148572,I148589,I148538,I148611,I510978,I148637,I148645,I148662,I510966,I148679,I510957,I148696,I148713,I510963,I148730,I510981,I148747,I510954,I148764,I148514,I148795,I148812,I148829,I148846,I148526,I148520,I148891,I510960,I148535,I148529,I148936,I148953,I510972,I148970,I148987,I510975,I149013,I149021,I148523,I148517,I149075,I149083,I148532,I149141,I538747,I149167,I149184,I149133,I149206,I538756,I149232,I149240,I149257,I538744,I149274,I538735,I149291,I149308,I538741,I149325,I538759,I149342,I538732,I149359,I149109,I149390,I149407,I149424,I149441,I149121,I149115,I149486,I538738,I149130,I149124,I149531,I149548,I538750,I149565,I149582,I538753,I149608,I149616,I149118,I149112,I149670,I149678,I149127,I149736,I205107,I149762,I149779,I149728,I149801,I205122,I149827,I149835,I149852,I205119,I149869,I149886,I149903,I205116,I149920,I205131,I149937,I205128,I149954,I149704,I149985,I150002,I150019,I150036,I149716,I149710,I150081,I205125,I149725,I149719,I150126,I150143,I205113,I150160,I205134,I150177,I205110,I150203,I150211,I149713,I149707,I150265,I150273,I149722,I150334,I542611,I150360,I150368,I542608,I542626,I150385,I542617,I150411,I150302,I150433,I542632,I150459,I150467,I542614,I150484,I150510,I150326,I150532,I150308,I542620,I150572,I150589,I150597,I150614,I150311,I150645,I542635,I150662,I542623,I150688,I150696,I150299,I150317,I150741,I542629,I150758,I150320,I150305,I150314,I150323,I150861,I445099,I150887,I150895,I445102,I445096,I150912,I445108,I150938,I150829,I150960,I445111,I150986,I150994,I151011,I151037,I150853,I151059,I150835,I445114,I151099,I151116,I151124,I151141,I150838,I151172,I445105,I151189,I151215,I151223,I150826,I150844,I151268,I445117,I151285,I150847,I150832,I150841,I150850,I151388,I291844,I151414,I151422,I291856,I151439,I291841,I151465,I151356,I151487,I291865,I151513,I151521,I291862,I151538,I151564,I151380,I151586,I151362,I291853,I151626,I151643,I151651,I151668,I151365,I151699,I291850,I151716,I291859,I151742,I151750,I151353,I151371,I151795,I291847,I151812,I151374,I151359,I151368,I151377,I151915,I471449,I151941,I151949,I471452,I471446,I151966,I471458,I151992,I151883,I152014,I471461,I152040,I152048,I152065,I152091,I151907,I152113,I151889,I471464,I152153,I152170,I152178,I152195,I151892,I152226,I471455,I152243,I152269,I152277,I151880,I151898,I152322,I471467,I152339,I151901,I151886,I151895,I151904,I152442,I291249,I152468,I152476,I291261,I152493,I291246,I152519,I152541,I291270,I152567,I152575,I291267,I152592,I152618,I152640,I291258,I152680,I152697,I152705,I152722,I152753,I291255,I152770,I291264,I152796,I152804,I152849,I291252,I152866,I152969,I690421,I152995,I153003,I690418,I690409,I153020,I690406,I153046,I152937,I153068,I690415,I153094,I153102,I690424,I153119,I153145,I152961,I153167,I152943,I690427,I153207,I153224,I153232,I153249,I152946,I153280,I690412,I153297,I690430,I153323,I153331,I152934,I152952,I153376,I153393,I152955,I152940,I152949,I152958,I153496,I458801,I153522,I153530,I458804,I458798,I153547,I458810,I153573,I153464,I153595,I458813,I153621,I153629,I153646,I153672,I153488,I153694,I153470,I458816,I153734,I153751,I153759,I153776,I153473,I153807,I458807,I153824,I153850,I153858,I153461,I153479,I153903,I458819,I153920,I153482,I153467,I153476,I153485,I154023,I737109,I154049,I154057,I737088,I154074,I737115,I154100,I153991,I154122,I737103,I154148,I154156,I737106,I154173,I154199,I154015,I154221,I153997,I737097,I154261,I154278,I154286,I154303,I154000,I154334,I737094,I737091,I154351,I737112,I154377,I154385,I153988,I154006,I154430,I737100,I154447,I154009,I153994,I154003,I154012,I154550,I658872,I154576,I154584,I658854,I658878,I154601,I658869,I154627,I154518,I154649,I658875,I154675,I154683,I658863,I154700,I154726,I154542,I154748,I154524,I154788,I154805,I154813,I154830,I154527,I154861,I658860,I658857,I154878,I658866,I154904,I154912,I154515,I154533,I154957,I154974,I154536,I154521,I154530,I154539,I155077,I155103,I155111,I155128,I155154,I155176,I155202,I155210,I155227,I155253,I155275,I155315,I155332,I155340,I155357,I155388,I155405,I155431,I155439,I155484,I155501,I155604,I619686,I155630,I155638,I619701,I155655,I619704,I155681,I155703,I619710,I155729,I155737,I619692,I155754,I155780,I155802,I619689,I155842,I155859,I155867,I155884,I155915,I619695,I155932,I619707,I155958,I155966,I156011,I619698,I156028,I156131,I156157,I156165,I156182,I156208,I156230,I156256,I156264,I156281,I156307,I156329,I156369,I156386,I156394,I156411,I156442,I156459,I156485,I156493,I156538,I156555,I156658,I156684,I156692,I156709,I156735,I156626,I156757,I156783,I156791,I156808,I156834,I156650,I156856,I156632,I156896,I156913,I156921,I156938,I156635,I156969,I156986,I157012,I157020,I156623,I156641,I157065,I157082,I156644,I156629,I156638,I156647,I157185,I725804,I157211,I157219,I725783,I157236,I725810,I157262,I157153,I157284,I725798,I157310,I157318,I725801,I157335,I157361,I157177,I157383,I157159,I725792,I157423,I157440,I157448,I157465,I157162,I157496,I725789,I725786,I157513,I725807,I157539,I157547,I157150,I157168,I157592,I725795,I157609,I157171,I157156,I157165,I157174,I157712,I234801,I157738,I157746,I234813,I234792,I157763,I234816,I157789,I157680,I157811,I234807,I157837,I157845,I234789,I157862,I157888,I157704,I157910,I157686,I234804,I157950,I157967,I157975,I157992,I157689,I158023,I234795,I158040,I234798,I158066,I158074,I157677,I157695,I158119,I234810,I158136,I157698,I157683,I157692,I157701,I158239,I361434,I158265,I158273,I361425,I361440,I158290,I361446,I158316,I158207,I158338,I361431,I158364,I158372,I158389,I158415,I158231,I158437,I158213,I361428,I158477,I158494,I158502,I158519,I158216,I158550,I361422,I361437,I158567,I158593,I158601,I158204,I158222,I158646,I361443,I158663,I158225,I158210,I158219,I158228,I158766,I720449,I158792,I158800,I720428,I158817,I720455,I158843,I158734,I158865,I720443,I158891,I158899,I720446,I158916,I158942,I158758,I158964,I158740,I720437,I159004,I159021,I159029,I159046,I158743,I159077,I720434,I720431,I159094,I720452,I159120,I159128,I158731,I158749,I159173,I720440,I159190,I158752,I158737,I158746,I158755,I159293,I373572,I159319,I159327,I373563,I373578,I159344,I373584,I159370,I159261,I159392,I373569,I159418,I159426,I159443,I159469,I159285,I159491,I159267,I373566,I159531,I159548,I159556,I159573,I159270,I159604,I373560,I373575,I159621,I159647,I159655,I159258,I159276,I159700,I373581,I159717,I159279,I159264,I159273,I159282,I159820,I159846,I159854,I159871,I159897,I159788,I159919,I159945,I159953,I159970,I159996,I159812,I160018,I159794,I160058,I160075,I160083,I160100,I159797,I160131,I160148,I160174,I160182,I159785,I159803,I160227,I160244,I159806,I159791,I159800,I159809,I160347,I383398,I160373,I160381,I383389,I383404,I160398,I383410,I160424,I160315,I160446,I383395,I160472,I160480,I160497,I160523,I160339,I160545,I160321,I383392,I160585,I160602,I160610,I160627,I160324,I160658,I383386,I383401,I160675,I160701,I160709,I160312,I160330,I160754,I383407,I160771,I160333,I160318,I160327,I160336,I160874,I707359,I160900,I160908,I707338,I160925,I707365,I160951,I160973,I707353,I160999,I161007,I707356,I161024,I161050,I161072,I707347,I161112,I161129,I161137,I161154,I161185,I707344,I707341,I161202,I707362,I161228,I161236,I161281,I707350,I161298,I161401,I161427,I161435,I161452,I161478,I161500,I161526,I161534,I161551,I161577,I161599,I161639,I161656,I161664,I161681,I161712,I161729,I161755,I161763,I161808,I161825,I161928,I476192,I161954,I161962,I476195,I476189,I161979,I476201,I162005,I162027,I476204,I162053,I162061,I162078,I162104,I162126,I476207,I162166,I162183,I162191,I162208,I162239,I476198,I162256,I162282,I162290,I162335,I476210,I162352,I162455,I695540,I162481,I162489,I695567,I695543,I162506,I695552,I162532,I162423,I162554,I162580,I162588,I695564,I162605,I162631,I162447,I162653,I162429,I695546,I162693,I162710,I162718,I162735,I162432,I162766,I695561,I695549,I162783,I695555,I162809,I162817,I162420,I162438,I162862,I695558,I162879,I162441,I162426,I162435,I162444,I162982,I163008,I163016,I163033,I163059,I163081,I163107,I163115,I163132,I163158,I163180,I163220,I163237,I163245,I163262,I163293,I163310,I163336,I163344,I163389,I163406,I163509,I368948,I163535,I163543,I368939,I368954,I163560,I368960,I163586,I163477,I163608,I368945,I163634,I163642,I163659,I163685,I163501,I163707,I163483,I368942,I163747,I163764,I163772,I163789,I163486,I163820,I368936,I368951,I163837,I163863,I163871,I163474,I163492,I163916,I368957,I163933,I163495,I163480,I163489,I163498,I164036,I559951,I164062,I164070,I559948,I164087,I559960,I164113,I164004,I164135,I164161,I164169,I559966,I164186,I164212,I164028,I164234,I164010,I559954,I164274,I164291,I164299,I164316,I164013,I164347,I559963,I559969,I164364,I164390,I164398,I164001,I164019,I164443,I559957,I164460,I164022,I164007,I164016,I164025,I164563,I550414,I164589,I164597,I550411,I164614,I550423,I164640,I164531,I164662,I164688,I164696,I550429,I164713,I164739,I164555,I164761,I164537,I550417,I164801,I164818,I164826,I164843,I164540,I164874,I550426,I550432,I164891,I164917,I164925,I164528,I164546,I164970,I550420,I164987,I164549,I164534,I164543,I164552,I165090,I165116,I165124,I165141,I165167,I165189,I165215,I165223,I165240,I165266,I165288,I165328,I165345,I165353,I165370,I165401,I165418,I165444,I165452,I165497,I165514,I165617,I165643,I165651,I165668,I165694,I165585,I165716,I165742,I165750,I165767,I165793,I165609,I165815,I165591,I165855,I165872,I165880,I165897,I165594,I165928,I165945,I165971,I165979,I165582,I165600,I166024,I166041,I165603,I165588,I165597,I165606,I166144,I166170,I166178,I166195,I166221,I166112,I166243,I166269,I166277,I166294,I166320,I166136,I166342,I166118,I166382,I166399,I166407,I166424,I166121,I166455,I166472,I166498,I166506,I166109,I166127,I166551,I166568,I166130,I166115,I166124,I166133,I166671,I166697,I166705,I166722,I166748,I166639,I166770,I166796,I166804,I166821,I166847,I166663,I166869,I166645,I166909,I166926,I166934,I166951,I166648,I166982,I166999,I167025,I167033,I166636,I166654,I167078,I167095,I166657,I166642,I166651,I166660,I167198,I449842,I167224,I167232,I449845,I449839,I167249,I449851,I167275,I167166,I167297,I449854,I167323,I167331,I167348,I167374,I167190,I167396,I167172,I449857,I167436,I167453,I167461,I167478,I167175,I167509,I449848,I167526,I167552,I167560,I167163,I167181,I167605,I449860,I167622,I167184,I167169,I167178,I167187,I167725,I530337,I167751,I167759,I530334,I530352,I167776,I530343,I167802,I167693,I167824,I530358,I167850,I167858,I530340,I167875,I167901,I167717,I167923,I167699,I530346,I167963,I167980,I167988,I168005,I167702,I168036,I530361,I168053,I530349,I168079,I168087,I167690,I167708,I168132,I530355,I168149,I167711,I167696,I167705,I167714,I168252,I405362,I168278,I168286,I405353,I405368,I168303,I405374,I168329,I168220,I168351,I405359,I168377,I168385,I168402,I168428,I168244,I168450,I168226,I405356,I168490,I168507,I168515,I168532,I168229,I168563,I405350,I405365,I168580,I168606,I168614,I168217,I168235,I168659,I405371,I168676,I168238,I168223,I168232,I168241,I168779,I168805,I168813,I168830,I168856,I168747,I168878,I168904,I168912,I168929,I168955,I168771,I168977,I168753,I169017,I169034,I169042,I169059,I168756,I169090,I169107,I169133,I169141,I168744,I168762,I169186,I169203,I168765,I168750,I168759,I168768,I169306,I302481,I169332,I169340,I302466,I302469,I169357,I302484,I169383,I169274,I169405,I302478,I169431,I169439,I169456,I169482,I169298,I169504,I169280,I302475,I169544,I169561,I169569,I169586,I169283,I169617,I302490,I169634,I302487,I169660,I169668,I169271,I169289,I169713,I302472,I169730,I169292,I169277,I169286,I169295,I169833,I576336,I169859,I169867,I576351,I169884,I576354,I169910,I169801,I169932,I576360,I169958,I169966,I576342,I169983,I170009,I169825,I170031,I169807,I576339,I170071,I170088,I170096,I170113,I169810,I170144,I576345,I170161,I576357,I170187,I170195,I169798,I169816,I170240,I576348,I170257,I169819,I169804,I169813,I169822,I170360,I170386,I170394,I170411,I170437,I170328,I170459,I170485,I170493,I170510,I170536,I170352,I170558,I170334,I170598,I170615,I170623,I170640,I170337,I170671,I170688,I170714,I170722,I170325,I170343,I170767,I170784,I170346,I170331,I170340,I170349,I170887,I439829,I170913,I170921,I439832,I439826,I170938,I439838,I170964,I170986,I439841,I171012,I171020,I171037,I171063,I171085,I439844,I171125,I171142,I171150,I171167,I171198,I439835,I171215,I171241,I171249,I171294,I439847,I171311,I171414,I171440,I171448,I171465,I171491,I171382,I171513,I171539,I171547,I171564,I171590,I171406,I171612,I171388,I171652,I171669,I171677,I171694,I171391,I171725,I171742,I171768,I171776,I171379,I171397,I171821,I171838,I171400,I171385,I171394,I171403,I171941,I670296,I171967,I171975,I670278,I670302,I171992,I670293,I172018,I171909,I172040,I670299,I172066,I172074,I670287,I172091,I172117,I171933,I172139,I171915,I172179,I172196,I172204,I172221,I171918,I172252,I670284,I670281,I172269,I670290,I172295,I172303,I171906,I171924,I172348,I172365,I171927,I171912,I171921,I171930,I172468,I473030,I172494,I172502,I473033,I473027,I172519,I473039,I172545,I172567,I473042,I172593,I172601,I172618,I172644,I172666,I473045,I172706,I172723,I172731,I172748,I172779,I473036,I172796,I172822,I172830,I172875,I473048,I172892,I172995,I460382,I173021,I173029,I460385,I460379,I173046,I460391,I173072,I172963,I173094,I460394,I173120,I173128,I173145,I173171,I172987,I173193,I172969,I460397,I173233,I173250,I173258,I173275,I172972,I173306,I460388,I173323,I173349,I173357,I172960,I172978,I173402,I460400,I173419,I172981,I172966,I172975,I172984,I173522,I616796,I173548,I173556,I616811,I173573,I616814,I173599,I173490,I173621,I616820,I173647,I173655,I616802,I173672,I173698,I173514,I173720,I173496,I616799,I173760,I173777,I173785,I173802,I173499,I173833,I616805,I173850,I616817,I173876,I173884,I173487,I173505,I173929,I616808,I173946,I173508,I173493,I173502,I173511,I174049,I661048,I174075,I174083,I661030,I661054,I174100,I661045,I174126,I174148,I661051,I174174,I174182,I661039,I174199,I174225,I174247,I174287,I174304,I174312,I174329,I174360,I661036,I661033,I174377,I661042,I174403,I174411,I174456,I174473,I174576,I518709,I174602,I174610,I518706,I518724,I174627,I518715,I174653,I174544,I174675,I518730,I174701,I174709,I518712,I174726,I174752,I174568,I174774,I174550,I518718,I174814,I174831,I174839,I174856,I174553,I174887,I518733,I174904,I518721,I174930,I174938,I174541,I174559,I174983,I518727,I175000,I174562,I174547,I174556,I174565,I175103,I665944,I175129,I175137,I665926,I665950,I175154,I665941,I175180,I175202,I665947,I175228,I175236,I665935,I175253,I175279,I175301,I175341,I175358,I175366,I175383,I175414,I665932,I665929,I175431,I665938,I175457,I175465,I175510,I175527,I175630,I371260,I175656,I175664,I371251,I371266,I175681,I371272,I175707,I175598,I175729,I371257,I175755,I175763,I175780,I175806,I175622,I175828,I175604,I371254,I175868,I175885,I175893,I175910,I175607,I175941,I371248,I371263,I175958,I175984,I175992,I175595,I175613,I176037,I371269,I176054,I175616,I175601,I175610,I175619,I176157,I525169,I176183,I176191,I525166,I525184,I176208,I525175,I176234,I176125,I176256,I525190,I176282,I176290,I525172,I176307,I176333,I176149,I176355,I176131,I525178,I176395,I176412,I176420,I176437,I176134,I176468,I525193,I176485,I525181,I176511,I176519,I176122,I176140,I176564,I525187,I176581,I176143,I176128,I176137,I176146,I176684,I552658,I176710,I176718,I552655,I176735,I552667,I176761,I176652,I176783,I176809,I176817,I552673,I176834,I176860,I176676,I176882,I176658,I552661,I176922,I176939,I176947,I176964,I176661,I176995,I552670,I552676,I177012,I177038,I177046,I176649,I176667,I177091,I552664,I177108,I176670,I176655,I176664,I176673,I177211,I412876,I177237,I177245,I412867,I412882,I177262,I412888,I177288,I177179,I177310,I412873,I177336,I177344,I177361,I177387,I177203,I177409,I177185,I412870,I177449,I177466,I177474,I177491,I177188,I177522,I412864,I412879,I177539,I177565,I177573,I177176,I177194,I177618,I412885,I177635,I177197,I177182,I177191,I177200,I177738,I420857,I177764,I177772,I420860,I420854,I177789,I420866,I177815,I177837,I420869,I177863,I177871,I177888,I177914,I177936,I420872,I177976,I177993,I178001,I178018,I178049,I420863,I178066,I178092,I178100,I178145,I420875,I178162,I178265,I699624,I178291,I178299,I699603,I178316,I699630,I178342,I178364,I699618,I178390,I178398,I699621,I178415,I178441,I178463,I699612,I178503,I178520,I178528,I178545,I178576,I699609,I699606,I178593,I699627,I178619,I178627,I178672,I699615,I178689,I178792,I405940,I178818,I178826,I405931,I405946,I178843,I405952,I178869,I178891,I405937,I178917,I178925,I178942,I178968,I178990,I405934,I179030,I179047,I179055,I179072,I179103,I405928,I405943,I179120,I179146,I179154,I179199,I405949,I179216,I179319,I367792,I179345,I179353,I367783,I367798,I179370,I367804,I179396,I179287,I179418,I367789,I179444,I179452,I179469,I179495,I179311,I179517,I179293,I367786,I179557,I179574,I179582,I179599,I179296,I179630,I367780,I367795,I179647,I179673,I179681,I179284,I179302,I179726,I367801,I179743,I179305,I179290,I179299,I179308,I179846,I381086,I179872,I179880,I381077,I381092,I179897,I381098,I179923,I179814,I179945,I381083,I179971,I179979,I179996,I180022,I179838,I180044,I179820,I381080,I180084,I180101,I180109,I180126,I179823,I180157,I381074,I381089,I180174,I180200,I180208,I179811,I179829,I180253,I381095,I180270,I179832,I179817,I179826,I179835,I180373,I449315,I180399,I180407,I449318,I449312,I180424,I449324,I180450,I180472,I449327,I180498,I180506,I180523,I180549,I180571,I449330,I180611,I180628,I180636,I180653,I180684,I449321,I180701,I180727,I180735,I180780,I449333,I180797,I180900,I613906,I180926,I180934,I613921,I180951,I613924,I180977,I180999,I613930,I181025,I181033,I613912,I181050,I181076,I181098,I613909,I181138,I181155,I181163,I181180,I181211,I613915,I181228,I613927,I181254,I181262,I181307,I613918,I181324,I181427,I595988,I181453,I181461,I596003,I181478,I596006,I181504,I181395,I181526,I596012,I181552,I181560,I595994,I181577,I181603,I181419,I181625,I181401,I595991,I181665,I181682,I181690,I181707,I181404,I181738,I595997,I181755,I596009,I181781,I181789,I181392,I181410,I181834,I596000,I181851,I181413,I181398,I181407,I181416,I181954,I408252,I181980,I181988,I408243,I408258,I182005,I408264,I182031,I181922,I182053,I408249,I182079,I182087,I182104,I182130,I181946,I182152,I181928,I408246,I182192,I182209,I182217,I182234,I181931,I182265,I408240,I408255,I182282,I182308,I182316,I181919,I181937,I182361,I408261,I182378,I181940,I181925,I181934,I181943,I182481,I259281,I182507,I182515,I259293,I259272,I182532,I259296,I182558,I182449,I182580,I259287,I182606,I182614,I259269,I182631,I182657,I182473,I182679,I182455,I259284,I182719,I182736,I182744,I182761,I182458,I182792,I259275,I182809,I259278,I182835,I182843,I182446,I182464,I182888,I259290,I182905,I182467,I182452,I182461,I182470,I183008,I183034,I183042,I183059,I183085,I182976,I183107,I183133,I183141,I183158,I183184,I183000,I183206,I182982,I183246,I183263,I183271,I183288,I182985,I183319,I183336,I183362,I183370,I182973,I182991,I183415,I183432,I182994,I182979,I182988,I182997,I183535,I183561,I183569,I183586,I183612,I183503,I183634,I183660,I183668,I183685,I183711,I183527,I183733,I183509,I183773,I183790,I183798,I183815,I183512,I183846,I183863,I183889,I183897,I183500,I183518,I183942,I183959,I183521,I183506,I183515,I183524,I184062,I674815,I184088,I184096,I674812,I674803,I184113,I674800,I184139,I184030,I184161,I674809,I184187,I184195,I674818,I184212,I184238,I184054,I184260,I184036,I674821,I184300,I184317,I184325,I184342,I184039,I184373,I674806,I184390,I674824,I184416,I184424,I184027,I184045,I184469,I184486,I184048,I184033,I184042,I184051,I184589,I669752,I184615,I184623,I669734,I669758,I184640,I669749,I184666,I184688,I669755,I184714,I184722,I669743,I184739,I184765,I184787,I184827,I184844,I184852,I184869,I184900,I669740,I669737,I184917,I669746,I184943,I184951,I184996,I185013,I185116,I185142,I185150,I185167,I185193,I185084,I185215,I185241,I185249,I185266,I185292,I185108,I185314,I185090,I185354,I185371,I185379,I185396,I185093,I185427,I185444,I185470,I185478,I185081,I185099,I185523,I185540,I185102,I185087,I185096,I185105,I185643,I570049,I185669,I185677,I570046,I185694,I570058,I185720,I185611,I185742,I185768,I185776,I570064,I185793,I185819,I185635,I185841,I185617,I570052,I185881,I185898,I185906,I185923,I185620,I185954,I570061,I570067,I185971,I185997,I186005,I185608,I185626,I186050,I570055,I186067,I185629,I185614,I185623,I185632,I186170,I186196,I186204,I186221,I186247,I186138,I186269,I186295,I186303,I186320,I186346,I186162,I186368,I186144,I186408,I186425,I186433,I186450,I186147,I186481,I186498,I186524,I186532,I186135,I186153,I186577,I186594,I186156,I186141,I186150,I186159,I186697,I284109,I186723,I186731,I284121,I186748,I284106,I186774,I186665,I186796,I284130,I186822,I186830,I284127,I186847,I186873,I186689,I186895,I186671,I284118,I186935,I186952,I186960,I186977,I186674,I187008,I284115,I187025,I284124,I187051,I187059,I186662,I186680,I187104,I284112,I187121,I186683,I186668,I186677,I186686,I187224,I187250,I187258,I187275,I187301,I187323,I187349,I187357,I187374,I187400,I187422,I187462,I187479,I187487,I187504,I187535,I187552,I187578,I187586,I187631,I187648,I187751,I742464,I187777,I187785,I742443,I187802,I742470,I187828,I187719,I187850,I742458,I187876,I187884,I742461,I187901,I187927,I187743,I187949,I187725,I742452,I187989,I188006,I188014,I188031,I187728,I188062,I742449,I742446,I188079,I742467,I188105,I188113,I187716,I187734,I188158,I742455,I188175,I187737,I187722,I187731,I187740,I188278,I481241,I188304,I188312,I481238,I481256,I188329,I481247,I188355,I188377,I481262,I188403,I188411,I481244,I188428,I188454,I188476,I481250,I188516,I188533,I188541,I188558,I188589,I481265,I188606,I481253,I188632,I188640,I188685,I481259,I188702,I188805,I711524,I188831,I188839,I711503,I188856,I711530,I188882,I188773,I188904,I711518,I188930,I188938,I711521,I188955,I188981,I188797,I189003,I188779,I711512,I189043,I189060,I189068,I189085,I188782,I189116,I711509,I711506,I189133,I711527,I189159,I189167,I188770,I188788,I189212,I711515,I189229,I188791,I188776,I188785,I188794,I189332,I323867,I189358,I189366,I323852,I323855,I189383,I323870,I189409,I189300,I189431,I323864,I189457,I189465,I189482,I189508,I189324,I189530,I189306,I323861,I189570,I189587,I189595,I189612,I189309,I189643,I323876,I189660,I323873,I189686,I189694,I189297,I189315,I189739,I323858,I189756,I189318,I189303,I189312,I189321,I189859,I372994,I189885,I189893,I372985,I373000,I189910,I373006,I189936,I189958,I372991,I189984,I189992,I190009,I190035,I190057,I372988,I190097,I190114,I190122,I190139,I190170,I372982,I372997,I190187,I190213,I190221,I190266,I373003,I190283,I190386,I628356,I190412,I190420,I628371,I190437,I628374,I190463,I190485,I628380,I190511,I190519,I628362,I190536,I190562,I190584,I628359,I190624,I190641,I190649,I190666,I190697,I628365,I190714,I628377,I190740,I190748,I190793,I628368,I190810,I190913,I190939,I190947,I190964,I190990,I190881,I191012,I191038,I191046,I191063,I191089,I190905,I191111,I190887,I191151,I191168,I191176,I191193,I190890,I191224,I191241,I191267,I191275,I190878,I190896,I191320,I191337,I190899,I190884,I190893,I190902,I191440,I191466,I191474,I191491,I191517,I191539,I191565,I191573,I191590,I191616,I191638,I191678,I191695,I191703,I191720,I191751,I191768,I191794,I191802,I191847,I191864,I191967,I191993,I192001,I192018,I192044,I191935,I192066,I192092,I192100,I192117,I192143,I191959,I192165,I191941,I192205,I192222,I192230,I192247,I191944,I192278,I192295,I192321,I192329,I191932,I191950,I192374,I192391,I191953,I191938,I191947,I191956,I192494,I444045,I192520,I192528,I444048,I444042,I192545,I444054,I192571,I192462,I192593,I444057,I192619,I192627,I192644,I192670,I192486,I192692,I192468,I444060,I192732,I192749,I192757,I192774,I192471,I192805,I444051,I192822,I192848,I192856,I192459,I192477,I192901,I444063,I192918,I192480,I192465,I192474,I192483,I193021,I746034,I193047,I193055,I746013,I193072,I746040,I193098,I192989,I193120,I746028,I193146,I193154,I746031,I193171,I193197,I193013,I193219,I192995,I746022,I193259,I193276,I193284,I193301,I192998,I193332,I746019,I746016,I193349,I746037,I193375,I193383,I192986,I193004,I193428,I746025,I193445,I193007,I192992,I193001,I193010,I193548,I380508,I193574,I193582,I380499,I380514,I193599,I380520,I193625,I193647,I380505,I193673,I193681,I193698,I193724,I193746,I380502,I193786,I193803,I193811,I193828,I193859,I380496,I380511,I193876,I193902,I193910,I193955,I380517,I193972,I194075,I303637,I194101,I194109,I303622,I303625,I194126,I303640,I194152,I194174,I303634,I194200,I194208,I194225,I194251,I194273,I303631,I194313,I194330,I194338,I194355,I194386,I303646,I194403,I303643,I194429,I194437,I194482,I303628,I194499,I194602,I593098,I194628,I194636,I593113,I194653,I593116,I194679,I194701,I593122,I194727,I194735,I593104,I194752,I194778,I194800,I593101,I194840,I194857,I194865,I194882,I194913,I593107,I194930,I593119,I194956,I194964,I195009,I593110,I195026,I195129,I252753,I195155,I195163,I252765,I252744,I195180,I252768,I195206,I195097,I195228,I252759,I195254,I195262,I252741,I195279,I195305,I195121,I195327,I195103,I252756,I195367,I195384,I195392,I195409,I195106,I195440,I252747,I195457,I252750,I195483,I195491,I195094,I195112,I195536,I252762,I195553,I195115,I195100,I195109,I195118,I195656,I442464,I195682,I195690,I442467,I442461,I195707,I442473,I195733,I195624,I195755,I442476,I195781,I195789,I195806,I195832,I195648,I195854,I195630,I442479,I195894,I195911,I195919,I195936,I195633,I195967,I442470,I195984,I196010,I196018,I195621,I195639,I196063,I442482,I196080,I195642,I195627,I195636,I195645,I196183,I575758,I196209,I196217,I575773,I196234,I575776,I196260,I196151,I196282,I575782,I196308,I196316,I575764,I196333,I196359,I196175,I196381,I196157,I575761,I196421,I196438,I196446,I196463,I196160,I196494,I575767,I196511,I575779,I196537,I196545,I196148,I196166,I196590,I575770,I196607,I196169,I196154,I196163,I196172,I196710,I579226,I196736,I196744,I579241,I196761,I579244,I196787,I196678,I196809,I579250,I196835,I196843,I579232,I196860,I196886,I196702,I196908,I196684,I579229,I196948,I196965,I196973,I196990,I196687,I197021,I579235,I197038,I579247,I197064,I197072,I196675,I196693,I197117,I579238,I197134,I196696,I196681,I196690,I196699,I197237,I348140,I197263,I197271,I348131,I348146,I197288,I348152,I197314,I197205,I197336,I348137,I197362,I197370,I197387,I197413,I197229,I197435,I197211,I348134,I197475,I197492,I197500,I197517,I197214,I197548,I348128,I348143,I197565,I197591,I197599,I197202,I197220,I197644,I348149,I197661,I197223,I197208,I197217,I197226,I197764,I505789,I197790,I197798,I505786,I505804,I197815,I505795,I197841,I197732,I197863,I505810,I197889,I197897,I505792,I197914,I197940,I197756,I197962,I197738,I505798,I198002,I198019,I198027,I198044,I197741,I198075,I505813,I198092,I505801,I198118,I198126,I197729,I197747,I198171,I505807,I198188,I197750,I197735,I197744,I197753,I198291,I657240,I198317,I198325,I657222,I657246,I198342,I657237,I198368,I198259,I198390,I657243,I198416,I198424,I657231,I198441,I198467,I198283,I198489,I198265,I198529,I198546,I198554,I198571,I198268,I198602,I657228,I657225,I198619,I657234,I198645,I198653,I198256,I198274,I198698,I198715,I198277,I198262,I198271,I198280,I198818,I604080,I198844,I198852,I604095,I198869,I604098,I198895,I198786,I198917,I604104,I198943,I198951,I604086,I198968,I198994,I198810,I199016,I198792,I604083,I199056,I199073,I199081,I199098,I198795,I199129,I604089,I199146,I604101,I199172,I199180,I198783,I198801,I199225,I604092,I199242,I198804,I198789,I198798,I198807,I199345,I199371,I199379,I199396,I199422,I199444,I199470,I199478,I199495,I199521,I199543,I199583,I199600,I199608,I199625,I199656,I199673,I199699,I199707,I199752,I199769,I199872,I541965,I199898,I199906,I541962,I541980,I199923,I541971,I199949,I199840,I199971,I541986,I199997,I200005,I541968,I200022,I200048,I199864,I200070,I199846,I541974,I200110,I200127,I200135,I200152,I199849,I200183,I541989,I200200,I541977,I200226,I200234,I199837,I199855,I200279,I541983,I200296,I199858,I199843,I199852,I199861,I200399,I200425,I200433,I200450,I200476,I200367,I200498,I200524,I200532,I200549,I200575,I200391,I200597,I200373,I200637,I200654,I200662,I200679,I200376,I200710,I200727,I200753,I200761,I200364,I200382,I200806,I200823,I200385,I200370,I200379,I200388,I200926,I200952,I200960,I200977,I201003,I200894,I201025,I201051,I201059,I201076,I201102,I200918,I201124,I200900,I201164,I201181,I201189,I201206,I200903,I201237,I201254,I201280,I201288,I200891,I200909,I201333,I201350,I200912,I200897,I200906,I200915,I201453,I258737,I201479,I201487,I258749,I258728,I201504,I258752,I201530,I201421,I201552,I258743,I201578,I201586,I258725,I201603,I201629,I201445,I201651,I201427,I258740,I201691,I201708,I201716,I201733,I201430,I201764,I258731,I201781,I258734,I201807,I201815,I201418,I201436,I201860,I258746,I201877,I201439,I201424,I201433,I201442,I201980,I279944,I202006,I202014,I279956,I202031,I279941,I202057,I201948,I202079,I279965,I202105,I202113,I279962,I202130,I202156,I201972,I202178,I201954,I279953,I202218,I202235,I202243,I202260,I201957,I202291,I279950,I202308,I279959,I202334,I202342,I201945,I201963,I202387,I279947,I202404,I201966,I201951,I201960,I201969,I202507,I499329,I202533,I202541,I499326,I499344,I202558,I499335,I202584,I202475,I202606,I499350,I202632,I202640,I499332,I202657,I202683,I202499,I202705,I202481,I499338,I202745,I202762,I202770,I202787,I202484,I202818,I499353,I202835,I499341,I202861,I202869,I202472,I202490,I202914,I499347,I202931,I202493,I202478,I202487,I202496,I203034,I423492,I203060,I203068,I423495,I423489,I203085,I423501,I203111,I203002,I203133,I423504,I203159,I203167,I203184,I203210,I203026,I203232,I203008,I423507,I203272,I203289,I203297,I203314,I203011,I203345,I423498,I203362,I203388,I203396,I202999,I203017,I203441,I423510,I203458,I203020,I203005,I203014,I203023,I203561,I485763,I203587,I203595,I485760,I485778,I203612,I485769,I203638,I203529,I203660,I485784,I203686,I203694,I485766,I203711,I203737,I203553,I203759,I203535,I485772,I203799,I203816,I203824,I203841,I203538,I203872,I485787,I203889,I485775,I203915,I203923,I203526,I203544,I203968,I485781,I203985,I203547,I203532,I203541,I203550,I204088,I318087,I204114,I204122,I318072,I318075,I204139,I318090,I204165,I204056,I204187,I318084,I204213,I204221,I204238,I204264,I204080,I204286,I204062,I318081,I204326,I204343,I204351,I204368,I204065,I204399,I318096,I204416,I318093,I204442,I204450,I204053,I204071,I204495,I318078,I204512,I204074,I204059,I204068,I204077,I204615,I605814,I204641,I204649,I605829,I204666,I605832,I204692,I204714,I605838,I204740,I204748,I605820,I204765,I204791,I204813,I605817,I204853,I204870,I204878,I204895,I204926,I605823,I204943,I605835,I204969,I204977,I205022,I605826,I205039,I205142,I232625,I205168,I205176,I232637,I232616,I205193,I232640,I205219,I205241,I232631,I205267,I205275,I232613,I205292,I205318,I205340,I232628,I205380,I205397,I205405,I205422,I205453,I232619,I205470,I232622,I205496,I205504,I205549,I232634,I205566,I205669,I205695,I205703,I205720,I205746,I205637,I205768,I205794,I205802,I205819,I205845,I205661,I205867,I205643,I205907,I205924,I205932,I205949,I205646,I205980,I205997,I206023,I206031,I205634,I205652,I206076,I206093,I205655,I205640,I205649,I205658,I206196,I573446,I206222,I206230,I573461,I206247,I573464,I206273,I206164,I206295,I573470,I206321,I206329,I573452,I206346,I206372,I206188,I206394,I206170,I573449,I206434,I206451,I206459,I206476,I206173,I206507,I573455,I206524,I573467,I206550,I206558,I206161,I206179,I206603,I573458,I206620,I206182,I206167,I206176,I206185,I206723,I438775,I206749,I206757,I438778,I438772,I206774,I438784,I206800,I206691,I206822,I438787,I206848,I206856,I206873,I206899,I206715,I206921,I206697,I438790,I206961,I206978,I206986,I207003,I206700,I207034,I438781,I207051,I207077,I207085,I206688,I206706,I207130,I438793,I207147,I206709,I206694,I206703,I206712,I207250,I207276,I207284,I207301,I207327,I207218,I207349,I207375,I207383,I207400,I207426,I207242,I207448,I207224,I207488,I207505,I207513,I207530,I207227,I207561,I207578,I207604,I207612,I207215,I207233,I207657,I207674,I207236,I207221,I207230,I207239,I207777,I394380,I207803,I207811,I394371,I394386,I207828,I394392,I207854,I207745,I207876,I394377,I207902,I207910,I207927,I207953,I207769,I207975,I207751,I394374,I208015,I208032,I208040,I208057,I207754,I208088,I394368,I394383,I208105,I208131,I208139,I207742,I207760,I208184,I394389,I208201,I207763,I207748,I207757,I207766,I208304,I532921,I208330,I208338,I532918,I532936,I208355,I532927,I208381,I208272,I208403,I532942,I208429,I208437,I532924,I208454,I208480,I208296,I208502,I208278,I532930,I208542,I208559,I208567,I208584,I208281,I208615,I532945,I208632,I532933,I208658,I208666,I208269,I208287,I208711,I532939,I208728,I208290,I208275,I208284,I208293,I208831,I737704,I208857,I208865,I737683,I208882,I737710,I208908,I208799,I208930,I737698,I208956,I208964,I737701,I208981,I209007,I208823,I209029,I208805,I737692,I209069,I209086,I209094,I209111,I208808,I209142,I737689,I737686,I209159,I737707,I209185,I209193,I208796,I208814,I209238,I737695,I209255,I208817,I208802,I208811,I208820,I209358,I624310,I209384,I209392,I624325,I209409,I624328,I209435,I209326,I209457,I624334,I209483,I209491,I624316,I209508,I209534,I209350,I209556,I209332,I624313,I209596,I209613,I209621,I209638,I209335,I209669,I624319,I209686,I624331,I209712,I209720,I209323,I209341,I209765,I624322,I209782,I209344,I209329,I209338,I209347,I209885,I641072,I209911,I209919,I641087,I209936,I641090,I209962,I209853,I209984,I641096,I210010,I210018,I641078,I210035,I210061,I209877,I210083,I209859,I641075,I210123,I210140,I210148,I210165,I209862,I210196,I641081,I210213,I641093,I210239,I210247,I209850,I209868,I210292,I641084,I210309,I209871,I209856,I209865,I209874,I210412,I697839,I210438,I210446,I697818,I210463,I697845,I210489,I210380,I210511,I697833,I210537,I210545,I697836,I210562,I210588,I210404,I210610,I210386,I697827,I210650,I210667,I210675,I210692,I210389,I210723,I697824,I697821,I210740,I697842,I210766,I210774,I210377,I210395,I210819,I697830,I210836,I210398,I210383,I210392,I210401,I210939,I238065,I210965,I210973,I238077,I238056,I210990,I238080,I211016,I210907,I211038,I238071,I211064,I211072,I238053,I211089,I211115,I210931,I211137,I210913,I238068,I211177,I211194,I211202,I211219,I210916,I211250,I238059,I211267,I238062,I211293,I211301,I210904,I210922,I211346,I238074,I211363,I210925,I210910,I210919,I210928,I211466,I372416,I211492,I211500,I372407,I372422,I211517,I372428,I211543,I211565,I372413,I211591,I211599,I211616,I211642,I211664,I372410,I211704,I211721,I211729,I211746,I211777,I372404,I372419,I211794,I211820,I211828,I211873,I372425,I211890,I211993,I723424,I212019,I212027,I723403,I212044,I723430,I212070,I211961,I212092,I723418,I212118,I212126,I723421,I212143,I212169,I211985,I212191,I211967,I723412,I212231,I212248,I212256,I212273,I211970,I212304,I723409,I723406,I212321,I723427,I212347,I212355,I211958,I211976,I212400,I723415,I212417,I211979,I211964,I211973,I211982,I212520,I668120,I212546,I212554,I668102,I668126,I212571,I668117,I212597,I212488,I212619,I668123,I212645,I212653,I668111,I212670,I212696,I212512,I212718,I212494,I212758,I212775,I212783,I212800,I212497,I212831,I668108,I668105,I212848,I668114,I212874,I212882,I212485,I212503,I212927,I212944,I212506,I212491,I212500,I212509,I213047,I213073,I213081,I213098,I213124,I213146,I213172,I213180,I213197,I213223,I213245,I213285,I213302,I213310,I213327,I213358,I213375,I213401,I213409,I213454,I213471,I213574,I213600,I213608,I213625,I213651,I213542,I213673,I213699,I213707,I213724,I213750,I213566,I213772,I213548,I213812,I213829,I213837,I213854,I213551,I213885,I213902,I213928,I213936,I213539,I213557,I213981,I213998,I213560,I213545,I213554,I213563,I214101,I293629,I214127,I214135,I293641,I214152,I293626,I214178,I214069,I214200,I293650,I214226,I214234,I293647,I214251,I214277,I214093,I214299,I214075,I293638,I214339,I214356,I214364,I214381,I214078,I214412,I293635,I214429,I293644,I214455,I214463,I214066,I214084,I214508,I293632,I214525,I214087,I214072,I214081,I214090,I214628,I421911,I214654,I214662,I421914,I421908,I214679,I421920,I214705,I214596,I214727,I421923,I214753,I214761,I214778,I214804,I214620,I214826,I214602,I421926,I214866,I214883,I214891,I214908,I214605,I214939,I421917,I214956,I214982,I214990,I214593,I214611,I215035,I421929,I215052,I214614,I214599,I214608,I214617,I215155,I256561,I215181,I215189,I256573,I256552,I215206,I256576,I215232,I215123,I215254,I256567,I215280,I215288,I256549,I215305,I215331,I215147,I215353,I215129,I256564,I215393,I215410,I215418,I215435,I215132,I215466,I256555,I215483,I256558,I215509,I215517,I215120,I215138,I215562,I256570,I215579,I215141,I215126,I215135,I215144,I215682,I286489,I215708,I215716,I286501,I215733,I286486,I215759,I215650,I215781,I286510,I215807,I215815,I286507,I215832,I215858,I215674,I215880,I215656,I286498,I215920,I215937,I215945,I215962,I215659,I215993,I286495,I216010,I286504,I216036,I216044,I215647,I215665,I216089,I286492,I216106,I215668,I215653,I215662,I215671,I216209,I630090,I216235,I216243,I630105,I216260,I630108,I216286,I216308,I630114,I216334,I216342,I630096,I216359,I216385,I216407,I630093,I216447,I216464,I216472,I216489,I216520,I630099,I216537,I630111,I216563,I216571,I216616,I630102,I216633,I216736,I689843,I216762,I216770,I689840,I689831,I216787,I689828,I216813,I216835,I689837,I216861,I216869,I689846,I216886,I216912,I216934,I689849,I216974,I216991,I216999,I217016,I217047,I689834,I217064,I689852,I217090,I217098,I217143,I217160,I217263,I713309,I217289,I217297,I713288,I217314,I713315,I217340,I217231,I217362,I713303,I217388,I217396,I713306,I217413,I217439,I217255,I217461,I217237,I713297,I217501,I217518,I217526,I217543,I217240,I217574,I713294,I713291,I217591,I713312,I217617,I217625,I217228,I217246,I217670,I713300,I217687,I217249,I217234,I217243,I217252,I217790,I273969,I217816,I217824,I273981,I273960,I217841,I273984,I217867,I217758,I217889,I273975,I217915,I217923,I273957,I217940,I217966,I217782,I217988,I217764,I273972,I218028,I218045,I218053,I218070,I217767,I218101,I273963,I218118,I273966,I218144,I218152,I217755,I217773,I218197,I273978,I218214,I217776,I217761,I217770,I217779,I218317,I451423,I218343,I218351,I451426,I451420,I218368,I451432,I218394,I218285,I218416,I451435,I218442,I218450,I218467,I218493,I218309,I218515,I218291,I451438,I218555,I218572,I218580,I218597,I218294,I218628,I451429,I218645,I218671,I218679,I218282,I218300,I218724,I451441,I218741,I218303,I218288,I218297,I218306,I218844,I483825,I218870,I218878,I483822,I483840,I218895,I483831,I218921,I218812,I218943,I483846,I218969,I218977,I483828,I218994,I219020,I218836,I219042,I218818,I483834,I219082,I219099,I219107,I219124,I218821,I219155,I483849,I219172,I483837,I219198,I219206,I218809,I218827,I219251,I483843,I219268,I218830,I218815,I218824,I218833,I219371,I578648,I219397,I219405,I578663,I219422,I578666,I219448,I219470,I578672,I219496,I219504,I578654,I219521,I219547,I219569,I578651,I219609,I219626,I219634,I219651,I219682,I578657,I219699,I578669,I219725,I219733,I219778,I578660,I219795,I219898,I267985,I219924,I219932,I267997,I267976,I219949,I268000,I219975,I219866,I219997,I267991,I220023,I220031,I267973,I220048,I220074,I219890,I220096,I219872,I267988,I220136,I220153,I220161,I220178,I219875,I220209,I267979,I220226,I267982,I220252,I220260,I219863,I219881,I220305,I267994,I220322,I219884,I219869,I219878,I219887,I220425,I722829,I220451,I220459,I722808,I220476,I722835,I220502,I220393,I220524,I722823,I220550,I220558,I722826,I220575,I220601,I220417,I220623,I220399,I722817,I220663,I220680,I220688,I220705,I220402,I220736,I722814,I722811,I220753,I722832,I220779,I220787,I220390,I220408,I220832,I722820,I220849,I220411,I220396,I220405,I220414,I220952,I704384,I220978,I220986,I704363,I221003,I704390,I221029,I220920,I221051,I704378,I221077,I221085,I704381,I221102,I221128,I220944,I221150,I220926,I704372,I221190,I221207,I221215,I221232,I220929,I221263,I704369,I704366,I221280,I704387,I221306,I221314,I220917,I220935,I221359,I704375,I221376,I220938,I220923,I220932,I220941,I221479,I221505,I221513,I221530,I221556,I221447,I221578,I221604,I221612,I221629,I221655,I221471,I221677,I221453,I221717,I221734,I221742,I221759,I221456,I221790,I221807,I221833,I221841,I221444,I221462,I221886,I221903,I221465,I221450,I221459,I221468,I222006,I651800,I222032,I222040,I651782,I651806,I222057,I651797,I222083,I221974,I222105,I651803,I222131,I222139,I651791,I222156,I222182,I221998,I222204,I221980,I222244,I222261,I222269,I222286,I221983,I222317,I651788,I651785,I222334,I651794,I222360,I222368,I221971,I221989,I222413,I222430,I221992,I221977,I221986,I221995,I222533,I222559,I222567,I222584,I222610,I222501,I222632,I222658,I222666,I222683,I222709,I222525,I222731,I222507,I222771,I222788,I222796,I222813,I222510,I222844,I222861,I222887,I222895,I222498,I222516,I222940,I222957,I222519,I222504,I222513,I222522,I223060,I560512,I223086,I223094,I560509,I223111,I560521,I223137,I223028,I223159,I223185,I223193,I560527,I223210,I223236,I223052,I223258,I223034,I560515,I223298,I223315,I223323,I223340,I223037,I223371,I560524,I560530,I223388,I223414,I223422,I223025,I223043,I223467,I560518,I223484,I223046,I223031,I223040,I223049,I223587,I231537,I223613,I223621,I231549,I231528,I223638,I231552,I223664,I223686,I231543,I223712,I223720,I231525,I223737,I223763,I223785,I231540,I223825,I223842,I223850,I223867,I223898,I231531,I223915,I231534,I223941,I223949,I223994,I231546,I224011,I224114,I267441,I224140,I224148,I267453,I267432,I224165,I267456,I224191,I224082,I224213,I267447,I224239,I224247,I267429,I224264,I224290,I224106,I224312,I224088,I267444,I224352,I224369,I224377,I224394,I224091,I224425,I267435,I224442,I267438,I224468,I224476,I224079,I224097,I224521,I267450,I224538,I224100,I224085,I224094,I224103,I224641,I744844,I224667,I224675,I744823,I224692,I744850,I224718,I224609,I224740,I744838,I224766,I224774,I744841,I224791,I224817,I224633,I224839,I224615,I744832,I224879,I224896,I224904,I224921,I224618,I224952,I744829,I744826,I224969,I744847,I224995,I225003,I224606,I224624,I225048,I744835,I225065,I224627,I224612,I224621,I224630,I225168,I425600,I225194,I225202,I425603,I425597,I225219,I425609,I225245,I225136,I225267,I425612,I225293,I225301,I225318,I225344,I225160,I225366,I225142,I425615,I225406,I225423,I225431,I225448,I225145,I225479,I425606,I225496,I225522,I225530,I225133,I225151,I225575,I425618,I225592,I225154,I225139,I225148,I225157,I225695,I287084,I225721,I225729,I287096,I225746,I287081,I225772,I225794,I287105,I225820,I225828,I287102,I225845,I225871,I225893,I287093,I225933,I225950,I225958,I225975,I226006,I287090,I226023,I287099,I226049,I226057,I226102,I287087,I226119,I226222,I255473,I226248,I226256,I255485,I255464,I226273,I255488,I226299,I226190,I226321,I255479,I226347,I226355,I255461,I226372,I226398,I226214,I226420,I226196,I255476,I226460,I226477,I226485,I226502,I226199,I226533,I255467,I226550,I255470,I226576,I226584,I226187,I226205,I226629,I255482,I226646,I226208,I226193,I226202,I226211,I226749,I474084,I226775,I226783,I474087,I474081,I226800,I474093,I226826,I226717,I226848,I474096,I226874,I226882,I226899,I226925,I226741,I226947,I226723,I474099,I226987,I227004,I227012,I227029,I226726,I227060,I474090,I227077,I227103,I227111,I226714,I226732,I227156,I474102,I227173,I226735,I226720,I226729,I226738,I227276,I543257,I227302,I227310,I543254,I543272,I227327,I543263,I227353,I227244,I227375,I543278,I227401,I227409,I543260,I227426,I227452,I227268,I227474,I227250,I543266,I227514,I227531,I227539,I227556,I227253,I227587,I543281,I227604,I543269,I227630,I227638,I227241,I227259,I227683,I543275,I227700,I227262,I227247,I227256,I227265,I227803,I227829,I227837,I227854,I227880,I227902,I227928,I227936,I227953,I227979,I228001,I228041,I228058,I228066,I228083,I228114,I228131,I228157,I228165,I228210,I228227,I228330,I263089,I228356,I228364,I263101,I263080,I228381,I263104,I228407,I228298,I228429,I263095,I228455,I228463,I263077,I228480,I228506,I228322,I228528,I228304,I263092,I228568,I228585,I228593,I228610,I228307,I228641,I263083,I228658,I263086,I228684,I228692,I228295,I228313,I228737,I263098,I228754,I228316,I228301,I228310,I228319,I228857,I392646,I228883,I228891,I392637,I392652,I228908,I392658,I228934,I228825,I228956,I392643,I228982,I228990,I229007,I229033,I228849,I229055,I228831,I392640,I229095,I229112,I229120,I229137,I228834,I229168,I392634,I392649,I229185,I229211,I229219,I228822,I228840,I229264,I392655,I229281,I228843,I228828,I228837,I228846,I229384,I229410,I229427,I229376,I229449,I229466,I229483,I229509,I229517,I229543,I229551,I229568,I229355,I229608,I229616,I229349,I229364,I229661,I229678,I229704,I229352,I229726,I229743,I229760,I229367,I229791,I229808,I229358,I229839,I229361,I229373,I229370,I229928,I647977,I229954,I229971,I229920,I229993,I230010,I647989,I647992,I230027,I647995,I230053,I230061,I647980,I230087,I230095,I647986,I230112,I229899,I647974,I230152,I230160,I229893,I229908,I230205,I647998,I230222,I647983,I230248,I229896,I230270,I230287,I230304,I229911,I230335,I230352,I229902,I230383,I229905,I229917,I229914,I230472,I230498,I230515,I230537,I230554,I230571,I230597,I230605,I230631,I230639,I230656,I230696,I230704,I230749,I230766,I230792,I230814,I230831,I230848,I230879,I230896,I230927,I231016,I231042,I231059,I231081,I231098,I231115,I231141,I231149,I231175,I231183,I231200,I231240,I231248,I231293,I231310,I231336,I231358,I231375,I231392,I231423,I231440,I231471,I231560,I231586,I231603,I231625,I231642,I231659,I231685,I231693,I231719,I231727,I231744,I231784,I231792,I231837,I231854,I231880,I231902,I231919,I231936,I231967,I231984,I232015,I232104,I320965,I232130,I232147,I232096,I232169,I232186,I320962,I320983,I232203,I320986,I232229,I232237,I320971,I232263,I232271,I320974,I232288,I232075,I320977,I232328,I232336,I232069,I232084,I232381,I320968,I232398,I320980,I232424,I232072,I232446,I232463,I232480,I232087,I232511,I232528,I232078,I232559,I232081,I232093,I232090,I232648,I437730,I232674,I232691,I232713,I232730,I437724,I437721,I232747,I437736,I232773,I232781,I232807,I232815,I437718,I232832,I232872,I232880,I232925,I437733,I437727,I232942,I232968,I232990,I233007,I233024,I233055,I233072,I437739,I233103,I233192,I459337,I233218,I233235,I233184,I233257,I233274,I459331,I459328,I233291,I459343,I233317,I233325,I233351,I233359,I459325,I233376,I233163,I233416,I233424,I233157,I233172,I233469,I459340,I459334,I233486,I233512,I233160,I233534,I233551,I233568,I233175,I233599,I233616,I459346,I233166,I233647,I233169,I233181,I233178,I233736,I620845,I233762,I233779,I233728,I233801,I233818,I620857,I233835,I620848,I233861,I233869,I620866,I233895,I233903,I620842,I233920,I233707,I620860,I233960,I233968,I233701,I233716,I234013,I620854,I620851,I234030,I620863,I234056,I233704,I234078,I234095,I234112,I233719,I234143,I234160,I233710,I234191,I233713,I233725,I233722,I234280,I628937,I234306,I234323,I234272,I234345,I234362,I628949,I234379,I628940,I234405,I234413,I628958,I234439,I234447,I628934,I234464,I234251,I628952,I234504,I234512,I234245,I234260,I234557,I628946,I628943,I234574,I628955,I234600,I234248,I234622,I234639,I234656,I234263,I234687,I234704,I234254,I234735,I234257,I234269,I234266,I234824,I488350,I234850,I234867,I234889,I234906,I488365,I488353,I234923,I488344,I234949,I234957,I488356,I234983,I234991,I488347,I235008,I488362,I235048,I235056,I235101,I488371,I488359,I235118,I488368,I235144,I235166,I235183,I235200,I235231,I235248,I235279,I235368,I235394,I235411,I235360,I235433,I235450,I235467,I235493,I235501,I235527,I235535,I235552,I235339,I235592,I235600,I235333,I235348,I235645,I235662,I235688,I235336,I235710,I235727,I235744,I235351,I235775,I235792,I235342,I235823,I235345,I235357,I235354,I235912,I479306,I235938,I235955,I235977,I235994,I479321,I479309,I236011,I479300,I236037,I236045,I479312,I236071,I236079,I479303,I236096,I479318,I236136,I236144,I236189,I479327,I479315,I236206,I479324,I236232,I236254,I236271,I236288,I236319,I236336,I236367,I236456,I236482,I236499,I236521,I236538,I236555,I236581,I236589,I236615,I236623,I236640,I236680,I236688,I236733,I236750,I236776,I236798,I236815,I236832,I236863,I236880,I236911,I237000,I237026,I237043,I236992,I237065,I237082,I237099,I237125,I237133,I237159,I237167,I237184,I236971,I237224,I237232,I236965,I236980,I237277,I237294,I237320,I236968,I237342,I237359,I237376,I236983,I237407,I237424,I236974,I237455,I236977,I236989,I236986,I237544,I505146,I237570,I237587,I237536,I237609,I237626,I505161,I505149,I237643,I505140,I237669,I237677,I505152,I237703,I237711,I505143,I237728,I237515,I505158,I237768,I237776,I237509,I237524,I237821,I505167,I505155,I237838,I505164,I237864,I237512,I237886,I237903,I237920,I237527,I237951,I237968,I237518,I237999,I237521,I237533,I237530,I238088,I365471,I238114,I238131,I238153,I238170,I365492,I365483,I238187,I238213,I238221,I365477,I238247,I238255,I365474,I238272,I365468,I238312,I238320,I238365,I365480,I238382,I365489,I238408,I238430,I238447,I238464,I238495,I238512,I365486,I238543,I238632,I702010,I238658,I238675,I238624,I238697,I238714,I701986,I702007,I238731,I702004,I238757,I238765,I701983,I238791,I238799,I701995,I238816,I238603,I701998,I238856,I238864,I238597,I238612,I238909,I702001,I701989,I238926,I701992,I238952,I238600,I238974,I238991,I239008,I238615,I239039,I239056,I238606,I239087,I238609,I238621,I238618,I239176,I239202,I239219,I239168,I239241,I239258,I239275,I239301,I239309,I239335,I239343,I239360,I239147,I239400,I239408,I239141,I239156,I239453,I239470,I239496,I239144,I239518,I239535,I239552,I239159,I239583,I239600,I239150,I239631,I239153,I239165,I239162,I239720,I341773,I239746,I239763,I239785,I239802,I341794,I341785,I239819,I239845,I239853,I341779,I239879,I239887,I341776,I239904,I341770,I239944,I239952,I239997,I341782,I240014,I341791,I240040,I240062,I240079,I240096,I240127,I240144,I341788,I240175,I240264,I496102,I240290,I240307,I240256,I240329,I240346,I496117,I496105,I240363,I496096,I240389,I240397,I496108,I240423,I240431,I496099,I240448,I240235,I496114,I240488,I240496,I240229,I240244,I240541,I496123,I496111,I240558,I496120,I240584,I240232,I240606,I240623,I240640,I240247,I240671,I240688,I240238,I240719,I240241,I240253,I240250,I240808,I240834,I240851,I240873,I240890,I240907,I240933,I240941,I240967,I240975,I240992,I241032,I241040,I241085,I241102,I241128,I241150,I241167,I241184,I241215,I241232,I241263,I241352,I516128,I241378,I241395,I241344,I241417,I241434,I516143,I516131,I241451,I516122,I241477,I241485,I516134,I241511,I241519,I516125,I241536,I241323,I516140,I241576,I241584,I241317,I241332,I241629,I516149,I516137,I241646,I516146,I241672,I241320,I241694,I241711,I241728,I241335,I241759,I241776,I241326,I241807,I241329,I241341,I241338,I241896,I683488,I241922,I241939,I241961,I241978,I683485,I683482,I241995,I683470,I242021,I242029,I683494,I242055,I242063,I683479,I242080,I683473,I242120,I242128,I242173,I683476,I242190,I683491,I242216,I242238,I242255,I242272,I242303,I242320,I242351,I242440,I242466,I242483,I242432,I242505,I242522,I242539,I242565,I242573,I242599,I242607,I242624,I242411,I242664,I242672,I242405,I242420,I242717,I242734,I242760,I242408,I242782,I242799,I242816,I242423,I242847,I242864,I242414,I242895,I242417,I242429,I242426,I242984,I243010,I243027,I242976,I243049,I243066,I243083,I243109,I243117,I243143,I243151,I243168,I242955,I243208,I243216,I242949,I242964,I243261,I243278,I243304,I242952,I243326,I243343,I243360,I242967,I243391,I243408,I242958,I243439,I242961,I242973,I242970,I243528,I243554,I243571,I243520,I243593,I243610,I243627,I243653,I243661,I243687,I243695,I243712,I243499,I243752,I243760,I243493,I243508,I243805,I243822,I243848,I243496,I243870,I243887,I243904,I243511,I243935,I243952,I243502,I243983,I243505,I243517,I243514,I244072,I582697,I244098,I244115,I244064,I244137,I244154,I582709,I244171,I582700,I244197,I244205,I582718,I244231,I244239,I582694,I244256,I244043,I582712,I244296,I244304,I244037,I244052,I244349,I582706,I582703,I244366,I582715,I244392,I244040,I244414,I244431,I244448,I244055,I244479,I244496,I244046,I244527,I244049,I244061,I244058,I244616,I607551,I244642,I244659,I244608,I244681,I244698,I607563,I244715,I607554,I244741,I244749,I607572,I244775,I244783,I607548,I244800,I244587,I607566,I244840,I244848,I244581,I244596,I244893,I607560,I607557,I244910,I607569,I244936,I244584,I244958,I244975,I244992,I244599,I245023,I245040,I244590,I245071,I244593,I244605,I244602,I245160,I676552,I245186,I245203,I245152,I245225,I245242,I676549,I676546,I245259,I676534,I245285,I245293,I676558,I245319,I245327,I676543,I245344,I245131,I676537,I245384,I245392,I245125,I245140,I245437,I676540,I245454,I676555,I245480,I245128,I245502,I245519,I245536,I245143,I245567,I245584,I245134,I245615,I245137,I245149,I245146,I245704,I337727,I245730,I245747,I245769,I245786,I337724,I337745,I245803,I337748,I245829,I245837,I337733,I245863,I245871,I337736,I245888,I337739,I245928,I245936,I245981,I337730,I245998,I337742,I246024,I246046,I246063,I246080,I246111,I246128,I246159,I246248,I246274,I246291,I246240,I246313,I246330,I246347,I246373,I246381,I246407,I246415,I246432,I246219,I246472,I246480,I246213,I246228,I246525,I246542,I246568,I246216,I246590,I246607,I246624,I246231,I246655,I246672,I246222,I246703,I246225,I246237,I246234,I246792,I353911,I246818,I246835,I246784,I246857,I246874,I353932,I353923,I246891,I246917,I246925,I353917,I246951,I246959,I353914,I246976,I246763,I353908,I247016,I247024,I246757,I246772,I247069,I353920,I247086,I353929,I247112,I246760,I247134,I247151,I247168,I246775,I247199,I247216,I353926,I246766,I247247,I246769,I246781,I246778,I247336,I247362,I247379,I247328,I247401,I247418,I247435,I247461,I247469,I247495,I247503,I247520,I247307,I247560,I247568,I247301,I247316,I247613,I247630,I247656,I247304,I247678,I247695,I247712,I247319,I247743,I247760,I247310,I247791,I247313,I247325,I247322,I247880,I320387,I247906,I247923,I247945,I247962,I320384,I320405,I247979,I320408,I248005,I248013,I320393,I248039,I248047,I320396,I248064,I320399,I248104,I248112,I248157,I320390,I248174,I320402,I248200,I248222,I248239,I248256,I248287,I248304,I248335,I248424,I248450,I248467,I248489,I248506,I248523,I248549,I248557,I248583,I248591,I248608,I248648,I248656,I248701,I248718,I248744,I248766,I248783,I248800,I248831,I248848,I248879,I248968,I600615,I248994,I249011,I248960,I249033,I249050,I600627,I249067,I600618,I249093,I249101,I600636,I249127,I249135,I600612,I249152,I248939,I600630,I249192,I249200,I248933,I248948,I249245,I600624,I600621,I249262,I600633,I249288,I248936,I249310,I249327,I249344,I248951,I249375,I249392,I248942,I249423,I248945,I248957,I248954,I249512,I561070,I249538,I249555,I249577,I249594,I561088,I249611,I561082,I249637,I249645,I561076,I249671,I249679,I561085,I249696,I561073,I249736,I249744,I249789,I561091,I249806,I249832,I249854,I249871,I249888,I249919,I249936,I561079,I249967,I250056,I643387,I250082,I250099,I250048,I250121,I250138,I643399,I250155,I643390,I250181,I250189,I643408,I250215,I250223,I643384,I250240,I250027,I643402,I250280,I250288,I250021,I250036,I250333,I643396,I643393,I250350,I643405,I250376,I250024,I250398,I250415,I250432,I250039,I250463,I250480,I250030,I250511,I250033,I250045,I250042,I250600,I713910,I250626,I250643,I250592,I250665,I250682,I713886,I713907,I250699,I713904,I250725,I250733,I713883,I250759,I250767,I713895,I250784,I250571,I713898,I250824,I250832,I250565,I250580,I250877,I713901,I713889,I250894,I713892,I250920,I250568,I250942,I250959,I250976,I250583,I251007,I251024,I250574,I251055,I250577,I250589,I250586,I251144,I251170,I251187,I251136,I251209,I251226,I251243,I251269,I251277,I251303,I251311,I251328,I251115,I251368,I251376,I251109,I251124,I251421,I251438,I251464,I251112,I251486,I251503,I251520,I251127,I251551,I251568,I251118,I251599,I251121,I251133,I251130,I251688,I251714,I251731,I251680,I251753,I251770,I251787,I251813,I251821,I251847,I251855,I251872,I251659,I251912,I251920,I251653,I251668,I251965,I251982,I252008,I251656,I252030,I252047,I252064,I251671,I252095,I252112,I251662,I252143,I251665,I251677,I251674,I252232,I685222,I252258,I252275,I252224,I252297,I252314,I685219,I685216,I252331,I685204,I252357,I252365,I685228,I252391,I252399,I685213,I252416,I252203,I685207,I252456,I252464,I252197,I252212,I252509,I685210,I252526,I685225,I252552,I252200,I252574,I252591,I252608,I252215,I252639,I252656,I252206,I252687,I252209,I252221,I252218,I252776,I252802,I252819,I252841,I252858,I252875,I252901,I252909,I252935,I252943,I252960,I253000,I253008,I253053,I253070,I253096,I253118,I253135,I253152,I253183,I253200,I253231,I253320,I534862,I253346,I253363,I253312,I253385,I253402,I534877,I534865,I253419,I534856,I253445,I253453,I534868,I253479,I253487,I534859,I253504,I253291,I534874,I253544,I253552,I253285,I253300,I253597,I534883,I534871,I253614,I534880,I253640,I253288,I253662,I253679,I253696,I253303,I253727,I253744,I253294,I253775,I253297,I253309,I253306,I253864,I281729,I253890,I253907,I253856,I253929,I253946,I281732,I281750,I253963,I281738,I253989,I253997,I254023,I254031,I281747,I254048,I253835,I281741,I254088,I254096,I253829,I253844,I254141,I281744,I281726,I254158,I281735,I254184,I253832,I254206,I254223,I254240,I253847,I254271,I254288,I253838,I254319,I253841,I253853,I253850,I254408,I623157,I254434,I254451,I254473,I254490,I623169,I254507,I623160,I254533,I254541,I623178,I254567,I254575,I623154,I254592,I623172,I254632,I254640,I254685,I623166,I623163,I254702,I623175,I254728,I254750,I254767,I254784,I254815,I254832,I254863,I254952,I254978,I254995,I254944,I255017,I255034,I255051,I255077,I255085,I255111,I255119,I255136,I254923,I255176,I255184,I254917,I254932,I255229,I255246,I255272,I254920,I255294,I255311,I255328,I254935,I255359,I255376,I254926,I255407,I254929,I254941,I254938,I255496,I728785,I255522,I255539,I255561,I255578,I728761,I728782,I255595,I728779,I255621,I255629,I728758,I255655,I255663,I728770,I255680,I728773,I255720,I255728,I255773,I728776,I728764,I255790,I728767,I255816,I255838,I255855,I255872,I255903,I255920,I255951,I256040,I256066,I256083,I256032,I256105,I256122,I256139,I256165,I256173,I256199,I256207,I256224,I256011,I256264,I256272,I256005,I256020,I256317,I256334,I256360,I256008,I256382,I256399,I256416,I256023,I256447,I256464,I256014,I256495,I256017,I256029,I256026,I256584,I256610,I256627,I256649,I256666,I256683,I256709,I256717,I256743,I256751,I256768,I256808,I256816,I256861,I256878,I256904,I256926,I256943,I256960,I256991,I257008,I257039,I257128,I386279,I257154,I257171,I257120,I257193,I257210,I386300,I386291,I257227,I257253,I257261,I386285,I257287,I257295,I386282,I257312,I257099,I386276,I257352,I257360,I257093,I257108,I257405,I386288,I257422,I386297,I257448,I257096,I257470,I257487,I257504,I257111,I257535,I257552,I386294,I257102,I257583,I257105,I257117,I257114,I257672,I523880,I257698,I257715,I257664,I257737,I257754,I523895,I523883,I257771,I523874,I257797,I257805,I523886,I257831,I257839,I523877,I257856,I257643,I523892,I257896,I257904,I257637,I257652,I257949,I523901,I523889,I257966,I523898,I257992,I257640,I258014,I258031,I258048,I257655,I258079,I258096,I257646,I258127,I257649,I257661,I257658,I258216,I258242,I258259,I258281,I258298,I258315,I258341,I258349,I258375,I258383,I258400,I258440,I258448,I258493,I258510,I258536,I258558,I258575,I258592,I258623,I258640,I258671,I258760,I465134,I258786,I258803,I258825,I258842,I465128,I465125,I258859,I465140,I258885,I258893,I258919,I258927,I465122,I258944,I258984,I258992,I259037,I465137,I465131,I259054,I259080,I259102,I259119,I259136,I259167,I259184,I465143,I259215,I259304,I657769,I259330,I259347,I259369,I259386,I657781,I657784,I259403,I657787,I259429,I259437,I657772,I259463,I259471,I657778,I259488,I657766,I259528,I259536,I259581,I657790,I259598,I657775,I259624,I259646,I259663,I259680,I259711,I259728,I259759,I259848,I259874,I259891,I259840,I259913,I259930,I259947,I259973,I259981,I260007,I260015,I260032,I259819,I260072,I260080,I259813,I259828,I260125,I260142,I260168,I259816,I260190,I260207,I260224,I259831,I260255,I260272,I259822,I260303,I259825,I259837,I259834,I260392,I567241,I260418,I260435,I260384,I260457,I260474,I567259,I260491,I567253,I260517,I260525,I567247,I260551,I260559,I567256,I260576,I260363,I567244,I260616,I260624,I260357,I260372,I260669,I567262,I260686,I260712,I260360,I260734,I260751,I260768,I260375,I260799,I260816,I567250,I260366,I260847,I260369,I260381,I260378,I260936,I315185,I260962,I260979,I260928,I261001,I261018,I315182,I315203,I261035,I315206,I261061,I261069,I315191,I261095,I261103,I315194,I261120,I260907,I315197,I261160,I261168,I260901,I260916,I261213,I315188,I261230,I315200,I261256,I260904,I261278,I261295,I261312,I260919,I261343,I261360,I260910,I261391,I260913,I260925,I260922,I261480,I347553,I261506,I261523,I261545,I261562,I347574,I347565,I261579,I261605,I261613,I347559,I261639,I261647,I347556,I261664,I347550,I261704,I261712,I261757,I347562,I261774,I347571,I261800,I261822,I261839,I261856,I261887,I261904,I347568,I261935,I262024,I378187,I262050,I262067,I262089,I262106,I378208,I378199,I262123,I262149,I262157,I378193,I262183,I262191,I378190,I262208,I378184,I262248,I262256,I262301,I378196,I262318,I378205,I262344,I262366,I262383,I262400,I262431,I262448,I378202,I262479,I262568,I650153,I262594,I262611,I262560,I262633,I262650,I650165,I650168,I262667,I650171,I262693,I262701,I650156,I262727,I262735,I650162,I262752,I262539,I650150,I262792,I262800,I262533,I262548,I262845,I650174,I262862,I650159,I262888,I262536,I262910,I262927,I262944,I262551,I262975,I262992,I262542,I263023,I262545,I262557,I262554,I263112,I569485,I263138,I263155,I263177,I263194,I569503,I263211,I569497,I263237,I263245,I569491,I263271,I263279,I569500,I263296,I569488,I263336,I263344,I263389,I569506,I263406,I263432,I263454,I263471,I263488,I263519,I263536,I569494,I263567,I263656,I263682,I263699,I263648,I263721,I263738,I263755,I263781,I263789,I263815,I263823,I263840,I263627,I263880,I263888,I263621,I263636,I263933,I263950,I263976,I263624,I263998,I264015,I264032,I263639,I264063,I264080,I263630,I264111,I263633,I263645,I263642,I264200,I332525,I264226,I264243,I264192,I264265,I264282,I332522,I332543,I264299,I332546,I264325,I264333,I332531,I264359,I264367,I332534,I264384,I264171,I332537,I264424,I264432,I264165,I264180,I264477,I332528,I264494,I332540,I264520,I264168,I264542,I264559,I264576,I264183,I264607,I264624,I264174,I264655,I264177,I264189,I264186,I264744,I398417,I264770,I264787,I264736,I264809,I264826,I398438,I398429,I264843,I264869,I264877,I398423,I264903,I264911,I398420,I264928,I264715,I398414,I264968,I264976,I264709,I264724,I265021,I398426,I265038,I398435,I265064,I264712,I265086,I265103,I265120,I264727,I265151,I265168,I398432,I264718,I265199,I264721,I264733,I264730,I265288,I696116,I265314,I265331,I265280,I265353,I265370,I696122,I696125,I265387,I696101,I265413,I265421,I696128,I265447,I265455,I696110,I265472,I265259,I696107,I265512,I265520,I265253,I265268,I265565,I696104,I696113,I265582,I696119,I265608,I265256,I265630,I265647,I265664,I265271,I265695,I265712,I265262,I265743,I265265,I265277,I265274,I265832,I718670,I265858,I265875,I265824,I265897,I265914,I718646,I718667,I265931,I718664,I265957,I265965,I718643,I265991,I265999,I718655,I266016,I265803,I718658,I266056,I266064,I265797,I265812,I266109,I718661,I718649,I266126,I718652,I266152,I265800,I266174,I266191,I266208,I265815,I266239,I266256,I265806,I266287,I265809,I265821,I265818,I266376,I719265,I266402,I266419,I266441,I266458,I719241,I719262,I266475,I719259,I266501,I266509,I719238,I266535,I266543,I719250,I266560,I719253,I266600,I266608,I266653,I719256,I719244,I266670,I719247,I266696,I266718,I266735,I266752,I266783,I266800,I266831,I266920,I266946,I266963,I266912,I266985,I267002,I267019,I267045,I267053,I267079,I267087,I267104,I266891,I267144,I267152,I266885,I266900,I267197,I267214,I267240,I266888,I267262,I267279,I267296,I266903,I267327,I267344,I266894,I267375,I266897,I266909,I266906,I267464,I703200,I267490,I267507,I267529,I267546,I703176,I703197,I267563,I703194,I267589,I267597,I703173,I267623,I267631,I703185,I267648,I703188,I267688,I267696,I267741,I703191,I703179,I267758,I703182,I267784,I267806,I267823,I267840,I267871,I267888,I267919,I268008,I268034,I268051,I268073,I268090,I268107,I268133,I268141,I268167,I268175,I268192,I268232,I268240,I268285,I268302,I268328,I268350,I268367,I268384,I268415,I268432,I268463,I268552,I688112,I268578,I268595,I268544,I268617,I268634,I688109,I688106,I268651,I688094,I268677,I268685,I688118,I268711,I268719,I688103,I268736,I268523,I688097,I268776,I268784,I268517,I268532,I268829,I688100,I268846,I688115,I268872,I268520,I268894,I268911,I268928,I268535,I268959,I268976,I268526,I269007,I268529,I268541,I268538,I269096,I493518,I269122,I269139,I269161,I269178,I493533,I493521,I269195,I493512,I269221,I269229,I493524,I269255,I269263,I493515,I269280,I493530,I269320,I269328,I269373,I493539,I493527,I269390,I493536,I269416,I269438,I269455,I269472,I269503,I269520,I269551,I269640,I557143,I269666,I269683,I269632,I269705,I269722,I557161,I269739,I557155,I269765,I269773,I557149,I269799,I269807,I557158,I269824,I269611,I557146,I269864,I269872,I269605,I269620,I269917,I557164,I269934,I269960,I269608,I269982,I269999,I270016,I269623,I270047,I270064,I557152,I269614,I270095,I269617,I269629,I269626,I270184,I640497,I270210,I270227,I270176,I270249,I270266,I640509,I270283,I640500,I270309,I270317,I640518,I270343,I270351,I640494,I270368,I270155,I640512,I270408,I270416,I270149,I270164,I270461,I640506,I640503,I270478,I640515,I270504,I270152,I270526,I270543,I270560,I270167,I270591,I270608,I270158,I270639,I270161,I270173,I270170,I270728,I354489,I270754,I270771,I270793,I270810,I354510,I354501,I270827,I270853,I270861,I354495,I270887,I270895,I354492,I270912,I354486,I270952,I270960,I271005,I354498,I271022,I354507,I271048,I271070,I271087,I271104,I271135,I271152,I354504,I271183,I271272,I310561,I271298,I271315,I271264,I271337,I271354,I310558,I310579,I271371,I310582,I271397,I271405,I310567,I271431,I271439,I310570,I271456,I271243,I310573,I271496,I271504,I271237,I271252,I271549,I310564,I271566,I310576,I271592,I271240,I271614,I271631,I271648,I271255,I271679,I271696,I271246,I271727,I271249,I271261,I271258,I271816,I271842,I271859,I271881,I271898,I271915,I271941,I271949,I271975,I271983,I272000,I272040,I272048,I272093,I272110,I272136,I272158,I272175,I272192,I272223,I272240,I272271,I272360,I456702,I272386,I272403,I272352,I272425,I272442,I456696,I456693,I272459,I456708,I272485,I272493,I272519,I272527,I456690,I272544,I272331,I272584,I272592,I272325,I272340,I272637,I456705,I456699,I272654,I272680,I272328,I272702,I272719,I272736,I272343,I272767,I272784,I456711,I272334,I272815,I272337,I272349,I272346,I272904,I272930,I272947,I272969,I272986,I273003,I273029,I273037,I273063,I273071,I273088,I273128,I273136,I273181,I273198,I273224,I273246,I273263,I273280,I273311,I273328,I273359,I273448,I401307,I273474,I273491,I273440,I273513,I273530,I401328,I401319,I273547,I273573,I273581,I401313,I273607,I273615,I401310,I273632,I273419,I401304,I273672,I273680,I273413,I273428,I273725,I401316,I273742,I401325,I273768,I273416,I273790,I273807,I273824,I273431,I273855,I273872,I401322,I273422,I273903,I273425,I273437,I273434,I273992,I478660,I274018,I274035,I274057,I274074,I478675,I478663,I274091,I478654,I274117,I274125,I478666,I274151,I274159,I478657,I274176,I478672,I274216,I274224,I274269,I478681,I478669,I274286,I478678,I274312,I274334,I274351,I274368,I274399,I274416,I274447,I274536,I602349,I274562,I274579,I274528,I274601,I274618,I602361,I274635,I602352,I274661,I274669,I602370,I274695,I274703,I602346,I274720,I274507,I602364,I274760,I274768,I274501,I274516,I274813,I602358,I602355,I274830,I602367,I274856,I274504,I274878,I274895,I274912,I274519,I274943,I274960,I274510,I274991,I274513,I274525,I274522,I275080,I610441,I275106,I275123,I275072,I275145,I275162,I610453,I275179,I610444,I275205,I275213,I610462,I275239,I275247,I610438,I275264,I275051,I610456,I275304,I275312,I275045,I275060,I275357,I610450,I610447,I275374,I610459,I275400,I275048,I275422,I275439,I275456,I275063,I275487,I275504,I275054,I275535,I275057,I275069,I275066,I275624,I656681,I275650,I275667,I275689,I275706,I656693,I656696,I275723,I656699,I275749,I275757,I656684,I275783,I275791,I656690,I275808,I656678,I275848,I275856,I275901,I656702,I275918,I656687,I275944,I275966,I275983,I276000,I276031,I276048,I276079,I276168,I276194,I276211,I276160,I276233,I276250,I276267,I276293,I276301,I276327,I276335,I276352,I276139,I276392,I276400,I276133,I276148,I276445,I276462,I276488,I276136,I276510,I276527,I276544,I276151,I276575,I276592,I276142,I276623,I276145,I276157,I276154,I276712,I276738,I276755,I276704,I276777,I276794,I276811,I276837,I276845,I276871,I276879,I276896,I276683,I276936,I276944,I276677,I276692,I276989,I277006,I277032,I276680,I277054,I277071,I277088,I276695,I277119,I277136,I276686,I277167,I276689,I276701,I276698,I277256,I277282,I277299,I277321,I277338,I277355,I277381,I277389,I277415,I277423,I277440,I277480,I277488,I277533,I277550,I277576,I277598,I277615,I277632,I277663,I277680,I277711,I277800,I277826,I277843,I277792,I277865,I277882,I277899,I277925,I277933,I277959,I277967,I277984,I277771,I278024,I278032,I277765,I277780,I278077,I278094,I278120,I277768,I278142,I278159,I278176,I277783,I278207,I278224,I277774,I278255,I277777,I277789,I277786,I278344,I278370,I278387,I278409,I278426,I278443,I278469,I278477,I278503,I278511,I278528,I278568,I278576,I278621,I278638,I278664,I278686,I278703,I278720,I278751,I278768,I278799,I278888,I712720,I278914,I278931,I278880,I278953,I278970,I712696,I712717,I278987,I712714,I279013,I279021,I712693,I279047,I279055,I712705,I279072,I278859,I712708,I279112,I279120,I278853,I278868,I279165,I712711,I712699,I279182,I712702,I279208,I278856,I279230,I279247,I279264,I278871,I279295,I279312,I278862,I279343,I278865,I278877,I278874,I279432,I490288,I279458,I279475,I279424,I279497,I279514,I490303,I490291,I279531,I490282,I279557,I279565,I490294,I279591,I279599,I490285,I279616,I279403,I490300,I279656,I279664,I279397,I279412,I279709,I490309,I490297,I279726,I490306,I279752,I279400,I279774,I279791,I279808,I279415,I279839,I279856,I279406,I279887,I279409,I279421,I279418,I279973,I443524,I279999,I280016,I443521,I280047,I280055,I280072,I280089,I443518,I280106,I443533,I280123,I280140,I280157,I280188,I443527,I280205,I443515,I280222,I280267,I280284,I280315,I443536,I280332,I280363,I280380,I443530,I280397,I280423,I280431,I280462,I280479,I280510,I280568,I645136,I280594,I280611,I280560,I645118,I280642,I280650,I645124,I280667,I280684,I645139,I280701,I645130,I280718,I280735,I280752,I280557,I280783,I645142,I280800,I645121,I280817,I280542,I280554,I280862,I280879,I280548,I280910,I645127,I280927,I280536,I280958,I645133,I280975,I280992,I281018,I281026,I280545,I281057,I281074,I280551,I281105,I280539,I281163,I281189,I281206,I281237,I281245,I281262,I281279,I281296,I281313,I281330,I281347,I281378,I281395,I281412,I281457,I281474,I281505,I281522,I281553,I281570,I281587,I281613,I281621,I281652,I281669,I281700,I281758,I572886,I281784,I281801,I572868,I281832,I281840,I572874,I281857,I281874,I572889,I281891,I572880,I281908,I281925,I281942,I281973,I572892,I281990,I572871,I282007,I282052,I282069,I282100,I572877,I282117,I282148,I572883,I282165,I282182,I282208,I282216,I282247,I282264,I282295,I282353,I319809,I282379,I282396,I282345,I319821,I282427,I282435,I319806,I282452,I282469,I319824,I282486,I319815,I282503,I282520,I282537,I282342,I282568,I319827,I282585,I319830,I282602,I282327,I282339,I282647,I282664,I282333,I282695,I282712,I282321,I282743,I319818,I282760,I319812,I282777,I282803,I282811,I282330,I282842,I282859,I282336,I282890,I282324,I282948,I358541,I282974,I282991,I282940,I358535,I283022,I283030,I358532,I283047,I283064,I358544,I283081,I358547,I283098,I283115,I283132,I282937,I283163,I358556,I283180,I358550,I283197,I282922,I282934,I283242,I283259,I282928,I283290,I358538,I283307,I282916,I283338,I358553,I283355,I283372,I283398,I283406,I282925,I283437,I283454,I282931,I283485,I282919,I283543,I283569,I283586,I283535,I283617,I283625,I283642,I283659,I283676,I283693,I283710,I283727,I283532,I283758,I283775,I283792,I283517,I283529,I283837,I283854,I283523,I283885,I283902,I283511,I283933,I283950,I283967,I283993,I284001,I283520,I284032,I284049,I283526,I284080,I283514,I284138,I284164,I284181,I284212,I284220,I284237,I284254,I284271,I284288,I284305,I284322,I284353,I284370,I284387,I284432,I284449,I284480,I284497,I284528,I284545,I284562,I284588,I284596,I284627,I284644,I284675,I284733,I284759,I284776,I284725,I284807,I284815,I284832,I284849,I284866,I284883,I284900,I284917,I284722,I284948,I284965,I284982,I284707,I284719,I285027,I285044,I284713,I285075,I285092,I284701,I285123,I285140,I285157,I285183,I285191,I284710,I285222,I285239,I284716,I285270,I284704,I285328,I285354,I285371,I285320,I285402,I285410,I285427,I285444,I285461,I285478,I285495,I285512,I285317,I285543,I285560,I285577,I285302,I285314,I285622,I285639,I285308,I285670,I285687,I285296,I285718,I285735,I285752,I285778,I285786,I285305,I285817,I285834,I285311,I285865,I285299,I285923,I285949,I285966,I285915,I285997,I286005,I286022,I286039,I286056,I286073,I286090,I286107,I285912,I286138,I286155,I286172,I285897,I285909,I286217,I286234,I285903,I286265,I286282,I285891,I286313,I286330,I286347,I286373,I286381,I285900,I286412,I286429,I285906,I286460,I285894,I286518,I303047,I286544,I286561,I303059,I286592,I286600,I303044,I286617,I286634,I303062,I286651,I303053,I286668,I286685,I286702,I286733,I303065,I286750,I303068,I286767,I286812,I286829,I286860,I286877,I286908,I303056,I286925,I303050,I286942,I286968,I286976,I287007,I287024,I287055,I287113,I287139,I287156,I287187,I287195,I287212,I287229,I287246,I287263,I287280,I287297,I287328,I287345,I287362,I287407,I287424,I287455,I287472,I287503,I287520,I287537,I287563,I287571,I287602,I287619,I287650,I287708,I717453,I287734,I287751,I717459,I287782,I287790,I717474,I287807,I287824,I717465,I287841,I717462,I287858,I287875,I287892,I287923,I287940,I717477,I287957,I288002,I288019,I288050,I717471,I288067,I288098,I717456,I288115,I717468,I288132,I717480,I288158,I288166,I288197,I288214,I288245,I288303,I288329,I288346,I288295,I288377,I288385,I288402,I288419,I288436,I288453,I288470,I288487,I288292,I288518,I288535,I288552,I288277,I288289,I288597,I288614,I288283,I288645,I288662,I288271,I288693,I288710,I288727,I288753,I288761,I288280,I288792,I288809,I288286,I288840,I288274,I288898,I522597,I288924,I288941,I288890,I522585,I288972,I288980,I522582,I288997,I289014,I522594,I289031,I522591,I289048,I289065,I289082,I288887,I289113,I522600,I289130,I522603,I289147,I288872,I288884,I289192,I289209,I288878,I289240,I522606,I289257,I288866,I289288,I522609,I289305,I522588,I289322,I289348,I289356,I288875,I289387,I289404,I288881,I289435,I288869,I289493,I289519,I289536,I289485,I289567,I289575,I289592,I289609,I289626,I289643,I289660,I289677,I289482,I289708,I289725,I289742,I289467,I289479,I289787,I289804,I289473,I289835,I289852,I289461,I289883,I289900,I289917,I289943,I289951,I289470,I289982,I289999,I289476,I290030,I289464,I290088,I382239,I290114,I290131,I382233,I290162,I290170,I382230,I290187,I290204,I382242,I290221,I382245,I290238,I290255,I290272,I290303,I382254,I290320,I382248,I290337,I290382,I290399,I290430,I382236,I290447,I290478,I382251,I290495,I290512,I290538,I290546,I290577,I290594,I290625,I290683,I290709,I290726,I290675,I290757,I290765,I290782,I290799,I290816,I290833,I290850,I290867,I290672,I290898,I290915,I290932,I290657,I290669,I290977,I290994,I290663,I291025,I291042,I290651,I291073,I291090,I291107,I291133,I291141,I290660,I291172,I291189,I290666,I291220,I290654,I291278,I612190,I291304,I291321,I612172,I291352,I291360,I612178,I291377,I291394,I612193,I291411,I612184,I291428,I291445,I291462,I291493,I612196,I291510,I612175,I291527,I291572,I291589,I291620,I612181,I291637,I291668,I612187,I291685,I291702,I291728,I291736,I291767,I291784,I291815,I291873,I746608,I291899,I291916,I746614,I291947,I291955,I746629,I291972,I291989,I746620,I292006,I746617,I292023,I292040,I292057,I292088,I292105,I746632,I292122,I292167,I292184,I292215,I746626,I292232,I292263,I746611,I292280,I746623,I292297,I746635,I292323,I292331,I292362,I292379,I292410,I292468,I432984,I292494,I292511,I432981,I292542,I292550,I292567,I292584,I432978,I292601,I432993,I292618,I292635,I292652,I292683,I432987,I292700,I432975,I292717,I292762,I292779,I292810,I432996,I292827,I292858,I292875,I432990,I292892,I292918,I292926,I292957,I292974,I293005,I293063,I735303,I293089,I293106,I293055,I735309,I293137,I293145,I735324,I293162,I293179,I735315,I293196,I735312,I293213,I293230,I293247,I293052,I293278,I293295,I735327,I293312,I293037,I293049,I293357,I293374,I293043,I293405,I735321,I293422,I293031,I293453,I735306,I293470,I735318,I293487,I735330,I293513,I293521,I293040,I293552,I293569,I293046,I293600,I293034,I293658,I507093,I293684,I293701,I507081,I293732,I293740,I507078,I293757,I293774,I507090,I293791,I507087,I293808,I293825,I293842,I293873,I507096,I293890,I507099,I293907,I293952,I293969,I294000,I507102,I294017,I294048,I507105,I294065,I507084,I294082,I294108,I294116,I294147,I294164,I294195,I294253,I697223,I294279,I294296,I294245,I697229,I294327,I294335,I697244,I294352,I294369,I697235,I294386,I697232,I294403,I294420,I294437,I294242,I294468,I294485,I697247,I294502,I294227,I294239,I294547,I294564,I294233,I294595,I697241,I294612,I294221,I294643,I697226,I294660,I697238,I294677,I697250,I294703,I294711,I294230,I294742,I294759,I294236,I294790,I294224,I294848,I539393,I294874,I294891,I294840,I539381,I294922,I294930,I539378,I294947,I294964,I539390,I294981,I539387,I294998,I295015,I295032,I294837,I295063,I539396,I295080,I539399,I295097,I294822,I294834,I295142,I295159,I294828,I295190,I539402,I295207,I294816,I295238,I539405,I295255,I539384,I295272,I295298,I295306,I294825,I295337,I295354,I294831,I295385,I294819,I295443,I587336,I295469,I295486,I295435,I587318,I295517,I295525,I587324,I295542,I295559,I587339,I295576,I587330,I295593,I295610,I295627,I295432,I295658,I587342,I295675,I587321,I295692,I295417,I295429,I295737,I295754,I295423,I295785,I587327,I295802,I295411,I295833,I587333,I295850,I295867,I295893,I295901,I295420,I295932,I295949,I295426,I295980,I295414,I296038,I513553,I296064,I296081,I513541,I296112,I296120,I513538,I296137,I296154,I513550,I296171,I513547,I296188,I296205,I296222,I296253,I513556,I296270,I513559,I296287,I296332,I296349,I296380,I513562,I296397,I296428,I513565,I296445,I513544,I296462,I296488,I296496,I296527,I296544,I296575,I296633,I404781,I296659,I296676,I296625,I404775,I296707,I296715,I404772,I296732,I296749,I404784,I296766,I404787,I296783,I296800,I296817,I296622,I296848,I404796,I296865,I404790,I296882,I296607,I296619,I296927,I296944,I296613,I296975,I404778,I296992,I296601,I297023,I404793,I297040,I297057,I297083,I297091,I296610,I297122,I297139,I296616,I297170,I296604,I297228,I422971,I297254,I297271,I422968,I297302,I297310,I297327,I297344,I422965,I297361,I422980,I297378,I297395,I297412,I297443,I422974,I297460,I422962,I297477,I297522,I297539,I297570,I422983,I297587,I297618,I297635,I422977,I297652,I297678,I297686,I297717,I297734,I297765,I297823,I626062,I297849,I297866,I297815,I626044,I297897,I297905,I626050,I297922,I297939,I626065,I297956,I626056,I297973,I297990,I298007,I297812,I298038,I626068,I298055,I626047,I298072,I297797,I297809,I298117,I298134,I297803,I298165,I626053,I298182,I297791,I298213,I626059,I298230,I298247,I298273,I298281,I297800,I298312,I298329,I297806,I298360,I297794,I298418,I299579,I298444,I298461,I298410,I299591,I298492,I298500,I299576,I298517,I298534,I299594,I298551,I299585,I298568,I298585,I298602,I298407,I298633,I299597,I298650,I299600,I298667,I298392,I298404,I298712,I298729,I298398,I298760,I298777,I298386,I298808,I299588,I298825,I299582,I298842,I298868,I298876,I298395,I298907,I298924,I298401,I298955,I298389,I299013,I299039,I299056,I299005,I299087,I299095,I299112,I299129,I299146,I299163,I299180,I299197,I299002,I299228,I299245,I299262,I298987,I298999,I299307,I299324,I298993,I299355,I299372,I298981,I299403,I299420,I299437,I299463,I299471,I298990,I299502,I299519,I298996,I299550,I298984,I299608,I385698,I299634,I299642,I385710,I299668,I299676,I385701,I299693,I385704,I299710,I299727,I385707,I299744,I299775,I299792,I299809,I299826,I385713,I299871,I299916,I385719,I299933,I299950,I299981,I299998,I385716,I300015,I385722,I300041,I300049,I300094,I300111,I300128,I300186,I634714,I300212,I300220,I634720,I300246,I300254,I300271,I634717,I300288,I300305,I634735,I300322,I300353,I300370,I300387,I634738,I300404,I300449,I300494,I634723,I300511,I300528,I300559,I634729,I300576,I634726,I300593,I634732,I300619,I300627,I300672,I300689,I300706,I300764,I300790,I300798,I300824,I300832,I300849,I300866,I300883,I300900,I300750,I300931,I300948,I300965,I300982,I300747,I300738,I301027,I300741,I300735,I301072,I301089,I301106,I300744,I301137,I301154,I301171,I301197,I301205,I300732,I300756,I301250,I301267,I301284,I300753,I301342,I468817,I301368,I301376,I301402,I301410,I468814,I301427,I468829,I301444,I301461,I468823,I301478,I301509,I301526,I301543,I468820,I301560,I468811,I301605,I301650,I468832,I301667,I301684,I301715,I301732,I301749,I468826,I301775,I301783,I301828,I301845,I301862,I301920,I637026,I301946,I301954,I637032,I301980,I301988,I302005,I637029,I302022,I302039,I637047,I302056,I301906,I302087,I302104,I302121,I637050,I302138,I301903,I301894,I302183,I301897,I301891,I302228,I637035,I302245,I302262,I301900,I302293,I637041,I302310,I637038,I302327,I637044,I302353,I302361,I301888,I301912,I302406,I302423,I302440,I301909,I302498,I302524,I302532,I302558,I302566,I302583,I302600,I302617,I302634,I302665,I302682,I302699,I302716,I302761,I302806,I302823,I302840,I302871,I302888,I302905,I302931,I302939,I302984,I303001,I303018,I303076,I653976,I303102,I303110,I653970,I303136,I303144,I653979,I303161,I653958,I303178,I303195,I653967,I303212,I303243,I303260,I303277,I653982,I303294,I653961,I303339,I303384,I653964,I303401,I303418,I303449,I653973,I303466,I303483,I303509,I303517,I303562,I303579,I303596,I303654,I303680,I303688,I303714,I303722,I303739,I303756,I303773,I303790,I303821,I303838,I303855,I303872,I303917,I303962,I303979,I303996,I304027,I304044,I304061,I304087,I304095,I304140,I304157,I304174,I304232,I344660,I304258,I304266,I344672,I304292,I304300,I344663,I304317,I344666,I304334,I304351,I344669,I304368,I304218,I304399,I304416,I304433,I304450,I344675,I304215,I304206,I304495,I304209,I304203,I304540,I344681,I304557,I304574,I304212,I304605,I304622,I344678,I304639,I344684,I304665,I304673,I304200,I304224,I304718,I304735,I304752,I304221,I304810,I654520,I304836,I304844,I654514,I304870,I304878,I654523,I304895,I654502,I304912,I304929,I654511,I304946,I304796,I304977,I304994,I305011,I654526,I305028,I654505,I304793,I304784,I305073,I304787,I304781,I305118,I654508,I305135,I305152,I304790,I305183,I654517,I305200,I305217,I305243,I305251,I304778,I304802,I305296,I305313,I305330,I304799,I305388,I305414,I305422,I305448,I305456,I305473,I305490,I305507,I305524,I305374,I305555,I305572,I305589,I305606,I305371,I305362,I305651,I305365,I305359,I305696,I305713,I305730,I305368,I305761,I305778,I305795,I305821,I305829,I305356,I305380,I305874,I305891,I305908,I305377,I305966,I416910,I305992,I306000,I416922,I306026,I306034,I416913,I306051,I416916,I306068,I306085,I416919,I306102,I305952,I306133,I306150,I306167,I306184,I416925,I305949,I305940,I306229,I305943,I305937,I306274,I416931,I306291,I306308,I305946,I306339,I306356,I416928,I306373,I416934,I306399,I306407,I305934,I305958,I306452,I306469,I306486,I305955,I306544,I306570,I306578,I306604,I306612,I306629,I306646,I306663,I306680,I306530,I306711,I306728,I306745,I306762,I306527,I306518,I306807,I306521,I306515,I306852,I306869,I306886,I306524,I306917,I306934,I306951,I306977,I306985,I306512,I306536,I307030,I307047,I307064,I306533,I307122,I502562,I307148,I307156,I502559,I307182,I307190,I502556,I307207,I502583,I307224,I307241,I502571,I307258,I307108,I307289,I307306,I307323,I502577,I307340,I502568,I307105,I307096,I307385,I307099,I307093,I307430,I502565,I307447,I307464,I307102,I307495,I502580,I307512,I502574,I307529,I307555,I307563,I307090,I307114,I307608,I307625,I307642,I307111,I307700,I716858,I307726,I307734,I307760,I307768,I716882,I307785,I716864,I307802,I307819,I716879,I307836,I307686,I307867,I307884,I307901,I716861,I307918,I716870,I307683,I307674,I307963,I307677,I307671,I308008,I716867,I308025,I308042,I307680,I308073,I716876,I308090,I716885,I308107,I716873,I308133,I308141,I307668,I307692,I308186,I308203,I308220,I307689,I308278,I379918,I308304,I308312,I379930,I308338,I308346,I379921,I308363,I379924,I308380,I308397,I379927,I308414,I308264,I308445,I308462,I308479,I308496,I379933,I308261,I308252,I308541,I308255,I308249,I308586,I379939,I308603,I308620,I308258,I308651,I308668,I379936,I308685,I379942,I308711,I308719,I308246,I308270,I308764,I308781,I308798,I308267,I308856,I678280,I308882,I308890,I678292,I308916,I308924,I678283,I308941,I678271,I308958,I308975,I678268,I308992,I308842,I309023,I309040,I309057,I678274,I309074,I308839,I308830,I309119,I308833,I308827,I309164,I678289,I309181,I309198,I308836,I309229,I678277,I309246,I309263,I678286,I309289,I309297,I308824,I308848,I309342,I309359,I309376,I308845,I309434,I309460,I309468,I309494,I309502,I309519,I309536,I309553,I309570,I309420,I309601,I309618,I309635,I309652,I309417,I309408,I309697,I309411,I309405,I309742,I309759,I309776,I309414,I309807,I309824,I309841,I309867,I309875,I309402,I309426,I309920,I309937,I309954,I309423,I310012,I478014,I310038,I310046,I478011,I310072,I310080,I478008,I310097,I478035,I310114,I310131,I478023,I310148,I309998,I310179,I310196,I310213,I478029,I310230,I478020,I309995,I309986,I310275,I309989,I309983,I310320,I478017,I310337,I310354,I309992,I310385,I478032,I310402,I478026,I310419,I310445,I310453,I309980,I310004,I310498,I310515,I310532,I310001,I310590,I721618,I310616,I310624,I310650,I310658,I721642,I310675,I721624,I310692,I310709,I721639,I310726,I310757,I310774,I310791,I721621,I310808,I721630,I310853,I310898,I721627,I310915,I310932,I310963,I721636,I310980,I721645,I310997,I721633,I311023,I311031,I311076,I311093,I311110,I311168,I506438,I311194,I311202,I506435,I311228,I311236,I506432,I311253,I506459,I311270,I311287,I506447,I311304,I311154,I311335,I311352,I311369,I506453,I311386,I506444,I311151,I311142,I311431,I311145,I311139,I311476,I506441,I311493,I311510,I311148,I311541,I506456,I311558,I506450,I311575,I311601,I311609,I311136,I311160,I311654,I311671,I311688,I311157,I311746,I490934,I311772,I311780,I490931,I311806,I311814,I490928,I311831,I490955,I311848,I311865,I490943,I311882,I311732,I311913,I311930,I311947,I490949,I311964,I490940,I311729,I311720,I312009,I311723,I311717,I312054,I490937,I312071,I312088,I311726,I312119,I490952,I312136,I490946,I312153,I312179,I312187,I311714,I311738,I312232,I312249,I312266,I311735,I312324,I312350,I312358,I312384,I312392,I312409,I312426,I312443,I312460,I312310,I312491,I312508,I312525,I312542,I312307,I312298,I312587,I312301,I312295,I312632,I312649,I312666,I312304,I312697,I312714,I312731,I312757,I312765,I312292,I312316,I312810,I312827,I312844,I312313,I312902,I312928,I312936,I312962,I312970,I312987,I313004,I313021,I313038,I312888,I313069,I313086,I313103,I313120,I312885,I312876,I313165,I312879,I312873,I313210,I313227,I313244,I312882,I313275,I313292,I313309,I313335,I313343,I312870,I312894,I313388,I313405,I313422,I312891,I313480,I313506,I313514,I313540,I313548,I313565,I313582,I313599,I313616,I313466,I313647,I313664,I313681,I313698,I313463,I313454,I313743,I313457,I313451,I313788,I313805,I313822,I313460,I313853,I313870,I313887,I313913,I313921,I313448,I313472,I313966,I313983,I314000,I313469,I314058,I415754,I314084,I314092,I415766,I314118,I314126,I415757,I314143,I415760,I314160,I314177,I415763,I314194,I314044,I314225,I314242,I314259,I314276,I415769,I314041,I314032,I314321,I314035,I314029,I314366,I415775,I314383,I314400,I314038,I314431,I314448,I415772,I314465,I415778,I314491,I314499,I314026,I314050,I314544,I314561,I314578,I314047,I314636,I314662,I314670,I314696,I314704,I314721,I314738,I314755,I314772,I314622,I314803,I314820,I314837,I314854,I314619,I314610,I314899,I314613,I314607,I314944,I314961,I314978,I314616,I315009,I315026,I315043,I315069,I315077,I314604,I314628,I315122,I315139,I315156,I314625,I315214,I665400,I315240,I315248,I665394,I315274,I315282,I665403,I315299,I665382,I315316,I315333,I665391,I315350,I315381,I315398,I315415,I665406,I315432,I665385,I315477,I315522,I665388,I315539,I315556,I315587,I665397,I315604,I315621,I315647,I315655,I315700,I315717,I315734,I315792,I359688,I315818,I315826,I359700,I315852,I315860,I359691,I315877,I359694,I315894,I315911,I359697,I315928,I315778,I315959,I315976,I315993,I316010,I359703,I315775,I315766,I316055,I315769,I315763,I316100,I359709,I316117,I316134,I315772,I316165,I316182,I359706,I316199,I359712,I316225,I316233,I315760,I315784,I316278,I316295,I316312,I315781,I316370,I343504,I316396,I316404,I343516,I316430,I316438,I343507,I316455,I343510,I316472,I316489,I343513,I316506,I316356,I316537,I316554,I316571,I316588,I343519,I316353,I316344,I316633,I316347,I316341,I316678,I343525,I316695,I316712,I316350,I316743,I316760,I343522,I316777,I343528,I316803,I316811,I316338,I316362,I316856,I316873,I316890,I316359,I316948,I627778,I316974,I316982,I627784,I317008,I317016,I317033,I627781,I317050,I317067,I627799,I317084,I316934,I317115,I317132,I317149,I627802,I317166,I316931,I316922,I317211,I316925,I316919,I317256,I627787,I317273,I317290,I316928,I317321,I627793,I317338,I627790,I317355,I627796,I317381,I317389,I316916,I316940,I317434,I317451,I317468,I316937,I317526,I419222,I317552,I317560,I419234,I317586,I317594,I419225,I317611,I419228,I317628,I317645,I419231,I317662,I317693,I317710,I317727,I317744,I419237,I317789,I317834,I419243,I317851,I317868,I317899,I317916,I419240,I317933,I419246,I317959,I317967,I318012,I318029,I318046,I318104,I318130,I318138,I318164,I318172,I318189,I318206,I318223,I318240,I318271,I318288,I318305,I318322,I318367,I318412,I318429,I318446,I318477,I318494,I318511,I318537,I318545,I318590,I318607,I318624,I318682,I318708,I318716,I318742,I318750,I318767,I318784,I318801,I318818,I318668,I318849,I318866,I318883,I318900,I318665,I318656,I318945,I318659,I318653,I318990,I319007,I319024,I318662,I319055,I319072,I319089,I319115,I319123,I318650,I318674,I319168,I319185,I319202,I318671,I319260,I362578,I319286,I319294,I362590,I319320,I319328,I362581,I319345,I362584,I319362,I319379,I362587,I319396,I319246,I319427,I319444,I319461,I319478,I362593,I319243,I319234,I319523,I319237,I319231,I319568,I362599,I319585,I319602,I319240,I319633,I319650,I362596,I319667,I362602,I319693,I319701,I319228,I319252,I319746,I319763,I319780,I319249,I319838,I353330,I319864,I319872,I353342,I319898,I319906,I353333,I319923,I353336,I319940,I319957,I353339,I319974,I320005,I320022,I320039,I320056,I353345,I320101,I320146,I353351,I320163,I320180,I320211,I320228,I353348,I320245,I353354,I320271,I320279,I320324,I320341,I320358,I320416,I320442,I320450,I320476,I320484,I320501,I320518,I320535,I320552,I320583,I320600,I320617,I320634,I320679,I320724,I320741,I320758,I320789,I320806,I320823,I320849,I320857,I320902,I320919,I320936,I320994,I339458,I321020,I321028,I339470,I321054,I321062,I339461,I321079,I339464,I321096,I321113,I339467,I321130,I321161,I321178,I321195,I321212,I339473,I321257,I321302,I339479,I321319,I321336,I321367,I321384,I339476,I321401,I339482,I321427,I321435,I321480,I321497,I321514,I321572,I321598,I321606,I321632,I321640,I321657,I321674,I321691,I321708,I321558,I321739,I321756,I321773,I321790,I321555,I321546,I321835,I321549,I321543,I321880,I321897,I321914,I321552,I321945,I321962,I321979,I322005,I322013,I321540,I321564,I322058,I322075,I322092,I321561,I322150,I582116,I322176,I322184,I582122,I322210,I322218,I322235,I582119,I322252,I322269,I582137,I322286,I322136,I322317,I322334,I322351,I582140,I322368,I322133,I322124,I322413,I322127,I322121,I322458,I582125,I322475,I322492,I322130,I322523,I582131,I322540,I582128,I322557,I582134,I322583,I322591,I322118,I322142,I322636,I322653,I322670,I322139,I322728,I422441,I322754,I322762,I322788,I322796,I422438,I322813,I422453,I322830,I322847,I422447,I322864,I322714,I322895,I322912,I322929,I422444,I322946,I422435,I322711,I322702,I322991,I322705,I322699,I323036,I422456,I323053,I323070,I322708,I323101,I323118,I323135,I422450,I323161,I323169,I322696,I322720,I323214,I323231,I323248,I322717,I323306,I435089,I323332,I323340,I323366,I323374,I435086,I323391,I435101,I323408,I323425,I435095,I323442,I323473,I323490,I323507,I435092,I323524,I435083,I323569,I323614,I435104,I323631,I323648,I323679,I323696,I323713,I435098,I323739,I323747,I323792,I323809,I323826,I323884,I515482,I323910,I323918,I515479,I323944,I323952,I515476,I323969,I515503,I323986,I324003,I515491,I324020,I324051,I324068,I324085,I515497,I324102,I515488,I324147,I324192,I515485,I324209,I324226,I324257,I515500,I324274,I515494,I324291,I324317,I324325,I324370,I324387,I324404,I324462,I434562,I324488,I324496,I324522,I324530,I434559,I324547,I434574,I324564,I324581,I434568,I324598,I324448,I324629,I324646,I324663,I434565,I324680,I434556,I324445,I324436,I324725,I324439,I324433,I324770,I434577,I324787,I324804,I324442,I324835,I324852,I324869,I434571,I324895,I324903,I324430,I324454,I324948,I324965,I324982,I324451,I325040,I349284,I325066,I325074,I349296,I325100,I325108,I349287,I325125,I349290,I325142,I325159,I349293,I325176,I325207,I325224,I325241,I325258,I349299,I325303,I325348,I349305,I325365,I325382,I325413,I325430,I349302,I325447,I349308,I325473,I325481,I325526,I325543,I325560,I325618,I456169,I325644,I325652,I325678,I325686,I456166,I325703,I456181,I325720,I325737,I456175,I325754,I325604,I325785,I325802,I325819,I456172,I325836,I456163,I325601,I325592,I325881,I325595,I325589,I325926,I456184,I325943,I325960,I325598,I325991,I326008,I326025,I456178,I326051,I326059,I325586,I325610,I326104,I326121,I326138,I325607,I326196,I341192,I326222,I326230,I341204,I326256,I326264,I341195,I326281,I341198,I326298,I326315,I341201,I326332,I326363,I326380,I326397,I326414,I341207,I326459,I326504,I341213,I326521,I326538,I326569,I326586,I341210,I326603,I341216,I326629,I326637,I326682,I326699,I326716,I326774,I326800,I326808,I326834,I326842,I326859,I326876,I326893,I326910,I326941,I326958,I326975,I326992,I327037,I327082,I327099,I327116,I327147,I327164,I327181,I327207,I327215,I327260,I327277,I327294,I327352,I470925,I327378,I327386,I327412,I327420,I470922,I327437,I470937,I327454,I327471,I470931,I327488,I327338,I327519,I327536,I327553,I470928,I327570,I470919,I327335,I327326,I327615,I327329,I327323,I327660,I470940,I327677,I327694,I327332,I327725,I327742,I327759,I470934,I327785,I327793,I327320,I327344,I327838,I327855,I327872,I327341,I327930,I587896,I327956,I327964,I587902,I327990,I327998,I328015,I587899,I328032,I328049,I587917,I328066,I328097,I328114,I328131,I587920,I328148,I328193,I328238,I587905,I328255,I328272,I328303,I587911,I328320,I587908,I328337,I587914,I328363,I328371,I328416,I328433,I328450,I328508,I359110,I328534,I328542,I359122,I328568,I328576,I359113,I328593,I359116,I328610,I328627,I359119,I328644,I328494,I328675,I328692,I328709,I328726,I359125,I328491,I328482,I328771,I328485,I328479,I328816,I359131,I328833,I328850,I328488,I328881,I328898,I359128,I328915,I359134,I328941,I328949,I328476,I328500,I328994,I329011,I329028,I328497,I329086,I329112,I329120,I329146,I329154,I329171,I329188,I329205,I329222,I329072,I329253,I329270,I329287,I329304,I329069,I329060,I329349,I329063,I329057,I329394,I329411,I329428,I329066,I329459,I329476,I329493,I329519,I329527,I329054,I329078,I329572,I329589,I329606,I329075,I329664,I329690,I329698,I329724,I329732,I329749,I329766,I329783,I329800,I329650,I329831,I329848,I329865,I329882,I329647,I329638,I329927,I329641,I329635,I329972,I329989,I330006,I329644,I330037,I330054,I330071,I330097,I330105,I329632,I329656,I330150,I330167,I330184,I329653,I330242,I680592,I330268,I330276,I680604,I330302,I330310,I680595,I330327,I680583,I330344,I330361,I680580,I330378,I330228,I330409,I330426,I330443,I680586,I330460,I330225,I330216,I330505,I330219,I330213,I330550,I680601,I330567,I330584,I330222,I330615,I680589,I330632,I330649,I680598,I330675,I330683,I330210,I330234,I330728,I330745,I330762,I330231,I330820,I561652,I330846,I330854,I561643,I330880,I330888,I561637,I330905,I561649,I330922,I330939,I561640,I330956,I330806,I330987,I331004,I331021,I561646,I331038,I561631,I330803,I330794,I331083,I330797,I330791,I331128,I331145,I331162,I330800,I331193,I561634,I331210,I331227,I331253,I331261,I330788,I330812,I331306,I331323,I331340,I330809,I331398,I634136,I331424,I331432,I634142,I331458,I331466,I331483,I634139,I331500,I331517,I634157,I331534,I331384,I331565,I331582,I331599,I634160,I331616,I331381,I331372,I331661,I331375,I331369,I331706,I634145,I331723,I331740,I331378,I331771,I634151,I331788,I634148,I331805,I634154,I331831,I331839,I331366,I331390,I331884,I331901,I331918,I331387,I331976,I332002,I332010,I332036,I332044,I332061,I332078,I332095,I332112,I332143,I332160,I332177,I332194,I332239,I332284,I332301,I332318,I332349,I332366,I332383,I332409,I332417,I332462,I332479,I332496,I332554,I508376,I332580,I332588,I508373,I332614,I332622,I508370,I332639,I508397,I332656,I332673,I508385,I332690,I332721,I332738,I332755,I508391,I332772,I508382,I332817,I332862,I508379,I332879,I332896,I332927,I508394,I332944,I508388,I332961,I332987,I332995,I333040,I333057,I333074,I333132,I437197,I333158,I333166,I333192,I333200,I437194,I333217,I437209,I333234,I333251,I437203,I333268,I333118,I333299,I333316,I333333,I437200,I333350,I437191,I333115,I333106,I333395,I333109,I333103,I333440,I437212,I333457,I333474,I333112,I333505,I333522,I333539,I437206,I333565,I333573,I333100,I333124,I333618,I333635,I333652,I333121,I333710,I466709,I333736,I333744,I333770,I333778,I466706,I333795,I466721,I333812,I333829,I466715,I333846,I333696,I333877,I333894,I333911,I466712,I333928,I466703,I333693,I333684,I333973,I333687,I333681,I334018,I466724,I334035,I334052,I333690,I334083,I334100,I334117,I466718,I334143,I334151,I333678,I333702,I334196,I334213,I334230,I333699,I334288,I424549,I334314,I334322,I334348,I334356,I424546,I334373,I424561,I334390,I334407,I424555,I334424,I334274,I334455,I334472,I334489,I424552,I334506,I424543,I334271,I334262,I334551,I334265,I334259,I334596,I424564,I334613,I334630,I334268,I334661,I334678,I334695,I424558,I334721,I334729,I334256,I334280,I334774,I334791,I334808,I334277,I334866,I376450,I334892,I334900,I376462,I334926,I334934,I376453,I334951,I376456,I334968,I334985,I376459,I335002,I335033,I335050,I335067,I335084,I376465,I335129,I335174,I376471,I335191,I335208,I335239,I335256,I376468,I335273,I376474,I335299,I335307,I335352,I335369,I335386,I335444,I335470,I335478,I335504,I335512,I335529,I335546,I335563,I335580,I335430,I335611,I335628,I335645,I335662,I335427,I335418,I335707,I335421,I335415,I335752,I335769,I335786,I335424,I335817,I335834,I335851,I335877,I335885,I335412,I335436,I335930,I335947,I335964,I335433,I336022,I743633,I336048,I336056,I336082,I336090,I743657,I336107,I743639,I336124,I336141,I743654,I336158,I336008,I336189,I336206,I336223,I743636,I336240,I743645,I336005,I335996,I336285,I335999,I335993,I336330,I743642,I336347,I336364,I336002,I336395,I743651,I336412,I743660,I336429,I743648,I336455,I336463,I335990,I336014,I336508,I336525,I336542,I336011,I336600,I568384,I336626,I336634,I568375,I336660,I336668,I568369,I336685,I568381,I336702,I336719,I568372,I336736,I336586,I336767,I336784,I336801,I568378,I336818,I568363,I336583,I336574,I336863,I336577,I336571,I336908,I336925,I336942,I336580,I336973,I568366,I336990,I337007,I337033,I337041,I336568,I336592,I337086,I337103,I337120,I336589,I337178,I635870,I337204,I337212,I635876,I337238,I337246,I337263,I635873,I337280,I337297,I635891,I337314,I337164,I337345,I337362,I337379,I635894,I337396,I337161,I337152,I337441,I337155,I337149,I337486,I635879,I337503,I337520,I337158,I337551,I635885,I337568,I635882,I337585,I635888,I337611,I337619,I337146,I337170,I337664,I337681,I337698,I337167,I337756,I337782,I337790,I337816,I337824,I337841,I337858,I337875,I337892,I337923,I337940,I337957,I337974,I338019,I338064,I338081,I338098,I338129,I338146,I338163,I338189,I338197,I338242,I338259,I338276,I338334,I563881,I338360,I338368,I338385,I563878,I563896,I338402,I563893,I338428,I338436,I563875,I338462,I338470,I338487,I338504,I338521,I338317,I563887,I338561,I338569,I338586,I338603,I338620,I338320,I338651,I563890,I338668,I338694,I338702,I338302,I338733,I338311,I338764,I338781,I338323,I338812,I563884,I338314,I338305,I338308,I338326,I338912,I338938,I338946,I338963,I338980,I339006,I339014,I339040,I339048,I339065,I339082,I339099,I338895,I339139,I339147,I339164,I339181,I339198,I338898,I339229,I339246,I339272,I339280,I338880,I339311,I338889,I339342,I339359,I338901,I339390,I338892,I338883,I338886,I338904,I339490,I575198,I339516,I339524,I339541,I575180,I575192,I339558,I575195,I339584,I339592,I575189,I575186,I339618,I339626,I339643,I339660,I339677,I575204,I339717,I339725,I339742,I339759,I339776,I339807,I575183,I339824,I339850,I339858,I339889,I339920,I339937,I339968,I575201,I340068,I685782,I340094,I340102,I340119,I685806,I685788,I340136,I685794,I340162,I340170,I685800,I685785,I340196,I340204,I340221,I340238,I340255,I340051,I685797,I340295,I340303,I340320,I340337,I340354,I340054,I340385,I685803,I685791,I340402,I340428,I340436,I340036,I340467,I340045,I340498,I340515,I340057,I340546,I340048,I340039,I340042,I340060,I340646,I340672,I340680,I340697,I340714,I340740,I340748,I340774,I340782,I340799,I340816,I340833,I340629,I340873,I340881,I340898,I340915,I340932,I340632,I340963,I340980,I341006,I341014,I340614,I341045,I340623,I341076,I341093,I340635,I341124,I340626,I340617,I340620,I340638,I341224,I341250,I341258,I341275,I341292,I341318,I341326,I341352,I341360,I341377,I341394,I341411,I341451,I341459,I341476,I341493,I341510,I341541,I341558,I341584,I341592,I341623,I341654,I341671,I341702,I341802,I341828,I341836,I341853,I341870,I341896,I341904,I341930,I341938,I341955,I341972,I341989,I342029,I342037,I342054,I342071,I342088,I342119,I342136,I342162,I342170,I342201,I342232,I342249,I342280,I342380,I608144,I342406,I342414,I342431,I608126,I608138,I342448,I608141,I342474,I342482,I608135,I608132,I342508,I342516,I342533,I342550,I342567,I342363,I608150,I342607,I342615,I342632,I342649,I342666,I342366,I342697,I608129,I342714,I342740,I342748,I342348,I342779,I342357,I342810,I342827,I342369,I342858,I608147,I342360,I342351,I342354,I342372,I342958,I606410,I342984,I342992,I343009,I606392,I606404,I343026,I606407,I343052,I343060,I606401,I606398,I343086,I343094,I343111,I343128,I343145,I606416,I343185,I343193,I343210,I343227,I343244,I343275,I606395,I343292,I343318,I343326,I343357,I343388,I343405,I343436,I606413,I343536,I436679,I343562,I343570,I343587,I436667,I436685,I343604,I436682,I343630,I343638,I436673,I436670,I343664,I343672,I343689,I343706,I343723,I436664,I343763,I343771,I343788,I343805,I343822,I343853,I343870,I343896,I343904,I343935,I343966,I343983,I344014,I436676,I344114,I344140,I344148,I344165,I344182,I344208,I344216,I344242,I344250,I344267,I344284,I344301,I344097,I344341,I344349,I344366,I344383,I344400,I344100,I344431,I344448,I344474,I344482,I344082,I344513,I344091,I344544,I344561,I344103,I344592,I344094,I344085,I344088,I344106,I344692,I344718,I344726,I344743,I344760,I344786,I344794,I344820,I344828,I344845,I344862,I344879,I344919,I344927,I344944,I344961,I344978,I345009,I345026,I345052,I345060,I345091,I345122,I345139,I345170,I345270,I655046,I345296,I345304,I345321,I655049,I655058,I345338,I655061,I345364,I345372,I655070,I655052,I345398,I345406,I345423,I345440,I345457,I345253,I345497,I345505,I345522,I345539,I345556,I345256,I345587,I655067,I345604,I655064,I345630,I345638,I345238,I345669,I345247,I345700,I345717,I345259,I345748,I655055,I345250,I345241,I345244,I345262,I345848,I345874,I345882,I345899,I345916,I345942,I345950,I345976,I345984,I346001,I346018,I346035,I346075,I346083,I346100,I346117,I346134,I346165,I346182,I346208,I346216,I346247,I346278,I346295,I346326,I346426,I346452,I346460,I346477,I346494,I346520,I346528,I346554,I346562,I346579,I346596,I346613,I346409,I346653,I346661,I346678,I346695,I346712,I346412,I346743,I346760,I346786,I346794,I346394,I346825,I346403,I346856,I346873,I346415,I346904,I346406,I346397,I346400,I346418,I347004,I347030,I347038,I347055,I347072,I347098,I347106,I347132,I347140,I347157,I347174,I347191,I346987,I347231,I347239,I347256,I347273,I347290,I346990,I347321,I347338,I347364,I347372,I346972,I347403,I346981,I347434,I347451,I346993,I347482,I346984,I346975,I346978,I346996,I347582,I347608,I347616,I347633,I347650,I347676,I347684,I347710,I347718,I347735,I347752,I347769,I347809,I347817,I347834,I347851,I347868,I347899,I347916,I347942,I347950,I347981,I348012,I348029,I348060,I348160,I497412,I348186,I348194,I348211,I497388,I497403,I348228,I497415,I348254,I348262,I497400,I497391,I348288,I348296,I348313,I348330,I348347,I348387,I348395,I348412,I348429,I348446,I348477,I497406,I497397,I348494,I497409,I348520,I348528,I348559,I348590,I348607,I348638,I497394,I348738,I348764,I348772,I348789,I348806,I348832,I348840,I348866,I348874,I348891,I348908,I348925,I348965,I348973,I348990,I349007,I349024,I349055,I349072,I349098,I349106,I349137,I349168,I349185,I349216,I349316,I349342,I349350,I349367,I349384,I349410,I349418,I349444,I349452,I349469,I349486,I349503,I349543,I349551,I349568,I349585,I349602,I349633,I349650,I349676,I349684,I349715,I349746,I349763,I349794,I349894,I536172,I349920,I349928,I349945,I536148,I536163,I349962,I536175,I349988,I349996,I536160,I536151,I350022,I350030,I350047,I350064,I350081,I350121,I350129,I350146,I350163,I350180,I350211,I536166,I536157,I350228,I536169,I350254,I350262,I350293,I350324,I350341,I350372,I536154,I350472,I431409,I350498,I350506,I350523,I431397,I431415,I350540,I431412,I350566,I350574,I431403,I431400,I350600,I350608,I350625,I350642,I350659,I350455,I431394,I350699,I350707,I350724,I350741,I350758,I350458,I350789,I350806,I350832,I350840,I350440,I350871,I350449,I350902,I350919,I350461,I350950,I431406,I350452,I350443,I350446,I350464,I351050,I719860,I351076,I351084,I351101,I719845,I719833,I351118,I719848,I351144,I351152,I719851,I351178,I351186,I351203,I351220,I351237,I351033,I719839,I351277,I351285,I351302,I351319,I351336,I351036,I351367,I719836,I719842,I351384,I719857,I351410,I351418,I351018,I351449,I351027,I351480,I351497,I351039,I351528,I719854,I351030,I351021,I351024,I351042,I351628,I351654,I351662,I351679,I351696,I351722,I351730,I351756,I351764,I351781,I351798,I351815,I351855,I351863,I351880,I351897,I351914,I351945,I351962,I351988,I351996,I352027,I352058,I352075,I352106,I352206,I352232,I352240,I352257,I352274,I352300,I352308,I352334,I352342,I352359,I352376,I352393,I352189,I352433,I352441,I352458,I352475,I352492,I352192,I352523,I352540,I352566,I352574,I352174,I352605,I352183,I352636,I352653,I352195,I352684,I352186,I352177,I352180,I352198,I352784,I681736,I352810,I352818,I352835,I681760,I681742,I352852,I681748,I352878,I352886,I681754,I681739,I352912,I352920,I352937,I352954,I352971,I352767,I681751,I353011,I353019,I353036,I353053,I353070,I352770,I353101,I681757,I681745,I353118,I353144,I353152,I352752,I353183,I352761,I353214,I353231,I352773,I353262,I352764,I352755,I352758,I352776,I353362,I353388,I353396,I353413,I353430,I353456,I353464,I353490,I353498,I353515,I353532,I353549,I353589,I353597,I353614,I353631,I353648,I353679,I353696,I353722,I353730,I353761,I353792,I353809,I353840,I353940,I353966,I353974,I353991,I354008,I354034,I354042,I354068,I354076,I354093,I354110,I354127,I354167,I354175,I354192,I354209,I354226,I354257,I354274,I354300,I354308,I354339,I354370,I354387,I354418,I354518,I547051,I354544,I354552,I354569,I547048,I547066,I354586,I547063,I354612,I354620,I547045,I354646,I354654,I354671,I354688,I354705,I547057,I354745,I354753,I354770,I354787,I354804,I354835,I547060,I354852,I354878,I354886,I354917,I354948,I354965,I354996,I547054,I355096,I355122,I355130,I355147,I355164,I355190,I355198,I355224,I355232,I355249,I355266,I355283,I355079,I355323,I355331,I355348,I355365,I355382,I355082,I355413,I355430,I355456,I355464,I355064,I355495,I355073,I355526,I355543,I355085,I355574,I355076,I355067,I355070,I355088,I355674,I485138,I355700,I355708,I355725,I485114,I485129,I355742,I485141,I355768,I355776,I485126,I485117,I355802,I355810,I355827,I355844,I355861,I355657,I355901,I355909,I355926,I355943,I355960,I355660,I355991,I485132,I485123,I356008,I485135,I356034,I356042,I355642,I356073,I355651,I356104,I356121,I355663,I356152,I485120,I355654,I355645,I355648,I355666,I356252,I356278,I356286,I356303,I356320,I356346,I356354,I356380,I356388,I356405,I356422,I356439,I356479,I356487,I356504,I356521,I356538,I356569,I356586,I356612,I356620,I356651,I356682,I356699,I356730,I356830,I739495,I356856,I356864,I356881,I739480,I739468,I356898,I739483,I356924,I356932,I739486,I356958,I356966,I356983,I357000,I357017,I739474,I357057,I357065,I357082,I357099,I357116,I357147,I739471,I739477,I357164,I739492,I357190,I357198,I357229,I357260,I357277,I357308,I739489,I357408,I622016,I357434,I357442,I357459,I621998,I622010,I357476,I622013,I357502,I357510,I622007,I622004,I357536,I357544,I357561,I357578,I357595,I357391,I622022,I357635,I357643,I357660,I357677,I357694,I357394,I357725,I622001,I357742,I357768,I357776,I357376,I357807,I357385,I357838,I357855,I357397,I357886,I622019,I357388,I357379,I357382,I357400,I357986,I358012,I358020,I358037,I358054,I358080,I358088,I358114,I358122,I358139,I358156,I358173,I358213,I358221,I358238,I358255,I358272,I358303,I358320,I358346,I358354,I358385,I358416,I358433,I358464,I358564,I358590,I358598,I358615,I358632,I358658,I358666,I358692,I358700,I358717,I358734,I358751,I358791,I358799,I358816,I358833,I358850,I358881,I358898,I358924,I358932,I358963,I358994,I359011,I359042,I359142,I472515,I359168,I359176,I359193,I472503,I472521,I359210,I472518,I359236,I359244,I472509,I472506,I359270,I359278,I359295,I359312,I359329,I472500,I359369,I359377,I359394,I359411,I359428,I359459,I359476,I359502,I359510,I359541,I359572,I359589,I359620,I472512,I359720,I359746,I359754,I359771,I359788,I359814,I359822,I359848,I359856,I359873,I359890,I359907,I359947,I359955,I359972,I359989,I360006,I360037,I360054,I360080,I360088,I360119,I360150,I360167,I360198,I360298,I360324,I360332,I360349,I360366,I360392,I360400,I360426,I360434,I360451,I360468,I360485,I360281,I360525,I360533,I360550,I360567,I360584,I360284,I360615,I360632,I360658,I360666,I360266,I360697,I360275,I360728,I360745,I360287,I360776,I360278,I360269,I360272,I360290,I360876,I672488,I360902,I360910,I360927,I672512,I672494,I360944,I672500,I360970,I360978,I672506,I672491,I361004,I361012,I361029,I361046,I361063,I360859,I672503,I361103,I361111,I361128,I361145,I361162,I360862,I361193,I672509,I672497,I361210,I361236,I361244,I360844,I361275,I360853,I361306,I361323,I360865,I361354,I360856,I360847,I360850,I360868,I361454,I624906,I361480,I361488,I361505,I624888,I624900,I361522,I624903,I361548,I361556,I624897,I624894,I361582,I361590,I361607,I361624,I361641,I624912,I361681,I361689,I361706,I361723,I361740,I361771,I624891,I361788,I361814,I361822,I361853,I361884,I361901,I361932,I624909,I362032,I426139,I362058,I362066,I362083,I426127,I426145,I362100,I426142,I362126,I362134,I426133,I426130,I362160,I362168,I362185,I362202,I362219,I362015,I426124,I362259,I362267,I362284,I362301,I362318,I362018,I362349,I362366,I362392,I362400,I362000,I362431,I362009,I362462,I362479,I362021,I362510,I426136,I362012,I362003,I362006,I362024,I362610,I715100,I362636,I362644,I362661,I715085,I715073,I362678,I715088,I362704,I362712,I715091,I362738,I362746,I362763,I362780,I362797,I715079,I362837,I362845,I362862,I362879,I362896,I362927,I715076,I715082,I362944,I715097,I362970,I362978,I363009,I363040,I363057,I363088,I715094,I363188,I363214,I363222,I363239,I363256,I363282,I363290,I363316,I363324,I363341,I363358,I363375,I363415,I363423,I363440,I363457,I363474,I363505,I363522,I363548,I363556,I363587,I363618,I363635,I363666,I363766,I363792,I363800,I363817,I363834,I363860,I363868,I363894,I363902,I363919,I363936,I363953,I363749,I363993,I364001,I364018,I364035,I364052,I363752,I364083,I364100,I364126,I364134,I363734,I364165,I363743,I364196,I364213,I363755,I364244,I363746,I363737,I363740,I363758,I364344,I364370,I364378,I364395,I364412,I364438,I364446,I364472,I364480,I364497,I364514,I364531,I364327,I364571,I364579,I364596,I364613,I364630,I364330,I364661,I364678,I364704,I364712,I364312,I364743,I364321,I364774,I364791,I364333,I364822,I364324,I364315,I364318,I364336,I364922,I364948,I364956,I364973,I364990,I365016,I365024,I365050,I365058,I365075,I365092,I365109,I364905,I365149,I365157,I365174,I365191,I365208,I364908,I365239,I365256,I365282,I365290,I364890,I365321,I364899,I365352,I365369,I364911,I365400,I364902,I364893,I364896,I364914,I365500,I365526,I365534,I365551,I365568,I365594,I365602,I365628,I365636,I365653,I365670,I365687,I365727,I365735,I365752,I365769,I365786,I365817,I365834,I365860,I365868,I365899,I365930,I365947,I365978,I366078,I425085,I366104,I366112,I366129,I425073,I425091,I366146,I425088,I366172,I366180,I425079,I425076,I366206,I366214,I366231,I366248,I366265,I366061,I425070,I366305,I366313,I366330,I366347,I366364,I366064,I366395,I366412,I366438,I366446,I366046,I366477,I366055,I366508,I366525,I366067,I366556,I425082,I366058,I366049,I366052,I366070,I366656,I366682,I366690,I366707,I366724,I366750,I366758,I366784,I366792,I366809,I366826,I366843,I366883,I366891,I366908,I366925,I366942,I366973,I366990,I367016,I367024,I367055,I367086,I367103,I367134,I367234,I367260,I367268,I367285,I367302,I367328,I367336,I367362,I367370,I367387,I367404,I367421,I367461,I367469,I367486,I367503,I367520,I367551,I367568,I367594,I367602,I367633,I367664,I367681,I367712,I367812,I367838,I367846,I367863,I367880,I367906,I367914,I367940,I367948,I367965,I367982,I367999,I368039,I368047,I368064,I368081,I368098,I368129,I368146,I368172,I368180,I368211,I368242,I368259,I368290,I368390,I701415,I368416,I368424,I368441,I701400,I701388,I368458,I701403,I368484,I368492,I701406,I368518,I368526,I368543,I368560,I368577,I701394,I368617,I368625,I368642,I368659,I368676,I368707,I701391,I701397,I368724,I701412,I368750,I368758,I368789,I368820,I368837,I368868,I701409,I368968,I368994,I369002,I369019,I369036,I369062,I369070,I369096,I369104,I369121,I369138,I369155,I369195,I369203,I369220,I369237,I369254,I369285,I369302,I369328,I369336,I369367,I369398,I369415,I369446,I369546,I369572,I369580,I369597,I369614,I369640,I369648,I369674,I369682,I369699,I369716,I369733,I369529,I369773,I369781,I369798,I369815,I369832,I369532,I369863,I369880,I369906,I369914,I369514,I369945,I369523,I369976,I369993,I369535,I370024,I369526,I369517,I369520,I369538,I370124,I370150,I370158,I370175,I370192,I370218,I370226,I370252,I370260,I370277,I370294,I370311,I370107,I370351,I370359,I370376,I370393,I370410,I370110,I370441,I370458,I370484,I370492,I370092,I370523,I370101,I370554,I370571,I370113,I370602,I370104,I370095,I370098,I370116,I370702,I370728,I370736,I370753,I370770,I370796,I370804,I370830,I370838,I370855,I370872,I370889,I370685,I370929,I370937,I370954,I370971,I370988,I370688,I371019,I371036,I371062,I371070,I370670,I371101,I370679,I371132,I371149,I370691,I371180,I370682,I370673,I370676,I370694,I371280,I371306,I371314,I371331,I371348,I371374,I371382,I371408,I371416,I371433,I371450,I371467,I371507,I371515,I371532,I371549,I371566,I371597,I371614,I371640,I371648,I371679,I371710,I371727,I371758,I371858,I681158,I371884,I371892,I371909,I681182,I681164,I371926,I681170,I371952,I371960,I681176,I681161,I371986,I371994,I372011,I372028,I372045,I371841,I681173,I372085,I372093,I372110,I372127,I372144,I371844,I372175,I681179,I681167,I372192,I372218,I372226,I371826,I372257,I371835,I372288,I372305,I371847,I372336,I371838,I371829,I371832,I371850,I372436,I652870,I372462,I372470,I372487,I652873,I652882,I372504,I652885,I372530,I372538,I652894,I652876,I372564,I372572,I372589,I372606,I372623,I372663,I372671,I372688,I372705,I372722,I372753,I652891,I372770,I652888,I372796,I372804,I372835,I372866,I372883,I372914,I652879,I373014,I373040,I373048,I373065,I373082,I373108,I373116,I373142,I373150,I373167,I373184,I373201,I373241,I373249,I373266,I373283,I373300,I373331,I373348,I373374,I373382,I373413,I373444,I373461,I373492,I373592,I745445,I373618,I373626,I373643,I745430,I745418,I373660,I745433,I373686,I373694,I745436,I373720,I373728,I373745,I373762,I373779,I745424,I373819,I373827,I373844,I373861,I373878,I373909,I745421,I745427,I373926,I745442,I373952,I373960,I373991,I374022,I374039,I374070,I745439,I374170,I520668,I374196,I374204,I374221,I520644,I520659,I374238,I520671,I374264,I374272,I520656,I520647,I374298,I374306,I374323,I374340,I374357,I374397,I374405,I374422,I374439,I374456,I374487,I520662,I520653,I374504,I520665,I374530,I374538,I374569,I374600,I374617,I374648,I520650,I374748,I374774,I374782,I374799,I374816,I374842,I374850,I374876,I374884,I374901,I374918,I374935,I374731,I374975,I374983,I375000,I375017,I375034,I374734,I375065,I375082,I375108,I375116,I374716,I375147,I374725,I375178,I375195,I374737,I375226,I374728,I374719,I374722,I374740,I375326,I375352,I375360,I375377,I375394,I375420,I375428,I375454,I375462,I375479,I375496,I375513,I375553,I375561,I375578,I375595,I375612,I375643,I375660,I375686,I375694,I375725,I375756,I375773,I375804,I375904,I375930,I375938,I375955,I375972,I375998,I376006,I376032,I376040,I376057,I376074,I376091,I375887,I376131,I376139,I376156,I376173,I376190,I375890,I376221,I376238,I376264,I376272,I375872,I376303,I375881,I376334,I376351,I375893,I376382,I375884,I375875,I375878,I375896,I376482,I376508,I376516,I376533,I376550,I376576,I376584,I376610,I376618,I376635,I376652,I376669,I376709,I376717,I376734,I376751,I376768,I376799,I376816,I376842,I376850,I376881,I376912,I376929,I376960,I377060,I519376,I377086,I377094,I377111,I519352,I519367,I377128,I519379,I377154,I377162,I519364,I519355,I377188,I377196,I377213,I377230,I377247,I377043,I377287,I377295,I377312,I377329,I377346,I377046,I377377,I519370,I519361,I377394,I519373,I377420,I377428,I377028,I377459,I377037,I377490,I377507,I377049,I377538,I519358,I377040,I377031,I377034,I377052,I377638,I448273,I377664,I377672,I377689,I448261,I448279,I377706,I448276,I377732,I377740,I448267,I448264,I377766,I377774,I377791,I377808,I377825,I377621,I448258,I377865,I377873,I377890,I377907,I377924,I377624,I377955,I377972,I377998,I378006,I377606,I378037,I377615,I378068,I378085,I377627,I378116,I448270,I377618,I377609,I377612,I377630,I378216,I627218,I378242,I378250,I378267,I627200,I627212,I378284,I627215,I378310,I378318,I627209,I627206,I378344,I378352,I378369,I378386,I378403,I627224,I378443,I378451,I378468,I378485,I378502,I378533,I627203,I378550,I378576,I378584,I378615,I378646,I378663,I378694,I627221,I378794,I543924,I378820,I378828,I378845,I543900,I543915,I378862,I543927,I378888,I378896,I543912,I543903,I378922,I378930,I378947,I378964,I378981,I379021,I379029,I379046,I379063,I379080,I379111,I543918,I543909,I379128,I543921,I379154,I379162,I379193,I379224,I379241,I379272,I543906,I379372,I428774,I379398,I379406,I379423,I428762,I428780,I379440,I428777,I379466,I379474,I428768,I428765,I379500,I379508,I379525,I379542,I379559,I379355,I428759,I379599,I379607,I379624,I379641,I379658,I379358,I379689,I379706,I379732,I379740,I379340,I379771,I379349,I379802,I379819,I379361,I379850,I428771,I379352,I379343,I379346,I379364,I379950,I379976,I379984,I380001,I380018,I380044,I380052,I380078,I380086,I380103,I380120,I380137,I380177,I380185,I380202,I380219,I380236,I380267,I380284,I380310,I380318,I380349,I380380,I380397,I380428,I380528,I380554,I380562,I380579,I380596,I380622,I380630,I380656,I380664,I380681,I380698,I380715,I380755,I380763,I380780,I380797,I380814,I380845,I380862,I380888,I380896,I380927,I380958,I380975,I381006,I381106,I734140,I381132,I381140,I381157,I734125,I734113,I381174,I734128,I381200,I381208,I734131,I381234,I381242,I381259,I381276,I381293,I734119,I381333,I381341,I381358,I381375,I381392,I381423,I734116,I734122,I381440,I734137,I381466,I381474,I381505,I381536,I381553,I381584,I734134,I381684,I381710,I381718,I381735,I381752,I381778,I381786,I381812,I381820,I381837,I381854,I381871,I381667,I381911,I381919,I381936,I381953,I381970,I381670,I382001,I382018,I382044,I382052,I381652,I382083,I381661,I382114,I382131,I381673,I382162,I381664,I381655,I381658,I381676,I382262,I721050,I382288,I382296,I382313,I721035,I721023,I382330,I721038,I382356,I382364,I721041,I382390,I382398,I382415,I382432,I382449,I721029,I382489,I382497,I382514,I382531,I382548,I382579,I721026,I721032,I382596,I721047,I382622,I382630,I382661,I382692,I382709,I382740,I721044,I382840,I382866,I382874,I382891,I382908,I382934,I382942,I382968,I382976,I382993,I383010,I383027,I383067,I383075,I383092,I383109,I383126,I383157,I383174,I383200,I383208,I383239,I383270,I383287,I383318,I383418,I383444,I383452,I383469,I383486,I383512,I383520,I383546,I383554,I383571,I383588,I383605,I383645,I383653,I383670,I383687,I383704,I383735,I383752,I383778,I383786,I383817,I383848,I383865,I383896,I383996,I589070,I384022,I384030,I384047,I589052,I589064,I384064,I589067,I384090,I384098,I589061,I589058,I384124,I384132,I384149,I384166,I384183,I383979,I589076,I384223,I384231,I384248,I384265,I384282,I383982,I384313,I589055,I384330,I384356,I384364,I383964,I384395,I383973,I384426,I384443,I383985,I384474,I589073,I383976,I383967,I383970,I383988,I384574,I384600,I384608,I384625,I384642,I384668,I384676,I384702,I384710,I384727,I384744,I384761,I384801,I384809,I384826,I384843,I384860,I384891,I384908,I384934,I384942,I384973,I385004,I385021,I385052,I385152,I385178,I385186,I385203,I385220,I385246,I385254,I385280,I385288,I385305,I385322,I385339,I385135,I385379,I385387,I385404,I385421,I385438,I385138,I385469,I385486,I385512,I385520,I385120,I385551,I385129,I385582,I385599,I385141,I385630,I385132,I385123,I385126,I385144,I385730,I385756,I385764,I385781,I385798,I385824,I385832,I385858,I385866,I385883,I385900,I385917,I385957,I385965,I385982,I385999,I386016,I386047,I386064,I386090,I386098,I386129,I386160,I386177,I386208,I386308,I386334,I386342,I386359,I386376,I386402,I386410,I386436,I386444,I386461,I386478,I386495,I386535,I386543,I386560,I386577,I386594,I386625,I386642,I386668,I386676,I386707,I386738,I386755,I386786,I386886,I386912,I386920,I386937,I386954,I386980,I386988,I387014,I387022,I387039,I387056,I387073,I386869,I387113,I387121,I387138,I387155,I387172,I386872,I387203,I387220,I387246,I387254,I386854,I387285,I386863,I387316,I387333,I386875,I387364,I386866,I386857,I386860,I386878,I387464,I387490,I387498,I387515,I387532,I387558,I387566,I387592,I387600,I387617,I387634,I387651,I387447,I387691,I387699,I387716,I387733,I387750,I387450,I387781,I387798,I387824,I387832,I387432,I387863,I387441,I387894,I387911,I387453,I387942,I387444,I387435,I387438,I387456,I388042,I388068,I388076,I388093,I388110,I388136,I388144,I388170,I388178,I388195,I388212,I388229,I388025,I388269,I388277,I388294,I388311,I388328,I388028,I388359,I388376,I388402,I388410,I388010,I388441,I388019,I388472,I388489,I388031,I388520,I388022,I388013,I388016,I388034,I388620,I715695,I388646,I388654,I388671,I715680,I715668,I388688,I715683,I388714,I388722,I715686,I388748,I388756,I388773,I388790,I388807,I388603,I715674,I388847,I388855,I388872,I388889,I388906,I388606,I388937,I715671,I715677,I388954,I715692,I388980,I388988,I388588,I389019,I388597,I389050,I389067,I388609,I389098,I715689,I388600,I388591,I388594,I388612,I389198,I389224,I389232,I389249,I389266,I389292,I389300,I389326,I389334,I389351,I389368,I389385,I389181,I389425,I389433,I389450,I389467,I389484,I389184,I389515,I389532,I389558,I389566,I389166,I389597,I389175,I389628,I389645,I389187,I389676,I389178,I389169,I389172,I389190,I389776,I389802,I389810,I389827,I389844,I389870,I389878,I389904,I389912,I389929,I389946,I389963,I389759,I390003,I390011,I390028,I390045,I390062,I389762,I390093,I390110,I390136,I390144,I389744,I390175,I389753,I390206,I390223,I389765,I390254,I389756,I389747,I389750,I389768,I390354,I390380,I390388,I390405,I390422,I390448,I390456,I390482,I390490,I390507,I390524,I390541,I390581,I390589,I390606,I390623,I390640,I390671,I390688,I390714,I390722,I390753,I390784,I390801,I390832,I390932,I390958,I390966,I390983,I391000,I391026,I391034,I391060,I391068,I391085,I391102,I391119,I391159,I391167,I391184,I391201,I391218,I391249,I391266,I391292,I391300,I391331,I391362,I391379,I391410,I391510,I391536,I391544,I391561,I391578,I391604,I391612,I391638,I391646,I391663,I391680,I391697,I391493,I391737,I391745,I391762,I391779,I391796,I391496,I391827,I391844,I391870,I391878,I391478,I391909,I391487,I391940,I391957,I391499,I391988,I391490,I391481,I391484,I391502,I392088,I392114,I392122,I392139,I392156,I392182,I392190,I392216,I392224,I392241,I392258,I392275,I392315,I392323,I392340,I392357,I392374,I392405,I392422,I392448,I392456,I392487,I392518,I392535,I392566,I392666,I392692,I392700,I392717,I392734,I392760,I392768,I392794,I392802,I392819,I392836,I392853,I392893,I392901,I392918,I392935,I392952,I392983,I393000,I393026,I393034,I393065,I393096,I393113,I393144,I393244,I475150,I393270,I393278,I393295,I475138,I475156,I393312,I475153,I393338,I393346,I475144,I475141,I393372,I393380,I393397,I393414,I393431,I393227,I475135,I393471,I393479,I393496,I393513,I393530,I393230,I393561,I393578,I393604,I393612,I393212,I393643,I393221,I393674,I393691,I393233,I393722,I475147,I393224,I393215,I393218,I393236,I393822,I393848,I393856,I393873,I393890,I393916,I393924,I393950,I393958,I393975,I393992,I394009,I394049,I394057,I394074,I394091,I394108,I394139,I394156,I394182,I394190,I394221,I394252,I394269,I394300,I394400,I555466,I394426,I394434,I394451,I555463,I555481,I394468,I555478,I394494,I394502,I555460,I394528,I394536,I394553,I394570,I394587,I555472,I394627,I394635,I394652,I394669,I394686,I394717,I555475,I394734,I394760,I394768,I394799,I394830,I394847,I394878,I555469,I394978,I395004,I395012,I395029,I395046,I395072,I395080,I395106,I395114,I395131,I395148,I395165,I394961,I395205,I395213,I395230,I395247,I395264,I394964,I395295,I395312,I395338,I395346,I394946,I395377,I394955,I395408,I395425,I394967,I395456,I394958,I394949,I394952,I394970,I395556,I395582,I395590,I395607,I395624,I395650,I395658,I395684,I395692,I395709,I395726,I395743,I395539,I395783,I395791,I395808,I395825,I395842,I395542,I395873,I395890,I395916,I395924,I395524,I395955,I395533,I395986,I396003,I395545,I396034,I395536,I395527,I395530,I395548,I396134,I396160,I396168,I396185,I396202,I396228,I396236,I396262,I396270,I396287,I396304,I396321,I396361,I396369,I396386,I396403,I396420,I396451,I396468,I396494,I396502,I396533,I396564,I396581,I396612,I396712,I686360,I396738,I396746,I396763,I686384,I686366,I396780,I686372,I396806,I396814,I686378,I686363,I396840,I396848,I396865,I396882,I396899,I686375,I396939,I396947,I396964,I396981,I396998,I397029,I686381,I686369,I397046,I397072,I397080,I397111,I397142,I397159,I397190,I397290,I397316,I397324,I397341,I397358,I397384,I397392,I397418,I397426,I397443,I397460,I397477,I397273,I397517,I397525,I397542,I397559,I397576,I397276,I397607,I397624,I397650,I397658,I397258,I397689,I397267,I397720,I397737,I397279,I397768,I397270,I397261,I397264,I397282,I397868,I454597,I397894,I397902,I397919,I454585,I454603,I397936,I454600,I397962,I397970,I454591,I454588,I397996,I398004,I398021,I398038,I398055,I397851,I454582,I398095,I398103,I398120,I398137,I398154,I397854,I398185,I398202,I398228,I398236,I397836,I398267,I397845,I398298,I398315,I397857,I398346,I454594,I397848,I397839,I397842,I397860,I398446,I669190,I398472,I398480,I398497,I669193,I669202,I398514,I669205,I398540,I398548,I669214,I669196,I398574,I398582,I398599,I398616,I398633,I398673,I398681,I398698,I398715,I398732,I398763,I669211,I398780,I669208,I398806,I398814,I398845,I398876,I398893,I398924,I669199,I399024,I399050,I399058,I399075,I399092,I399118,I399126,I399152,I399160,I399177,I399194,I399211,I399251,I399259,I399276,I399293,I399310,I399341,I399358,I399384,I399392,I399423,I399454,I399471,I399502,I399602,I399628,I399636,I399653,I399670,I399696,I399704,I399730,I399738,I399755,I399772,I399789,I399585,I399829,I399837,I399854,I399871,I399888,I399588,I399919,I399936,I399962,I399970,I399570,I400001,I399579,I400032,I400049,I399591,I400080,I399582,I399573,I399576,I399594,I400180,I670822,I400206,I400214,I400231,I670825,I670834,I400248,I670837,I400274,I400282,I670846,I670828,I400308,I400316,I400333,I400350,I400367,I400163,I400407,I400415,I400432,I400449,I400466,I400166,I400497,I670843,I400514,I670840,I400540,I400548,I400148,I400579,I400157,I400610,I400627,I400169,I400658,I670831,I400160,I400151,I400154,I400172,I400758,I545862,I400784,I400792,I400809,I545838,I545853,I400826,I545865,I400852,I400860,I545850,I545841,I400886,I400894,I400911,I400928,I400945,I400741,I400985,I400993,I401010,I401027,I401044,I400744,I401075,I545856,I545847,I401092,I545859,I401118,I401126,I400726,I401157,I400735,I401188,I401205,I400747,I401236,I545844,I400738,I400729,I400732,I400750,I401336,I401362,I401370,I401387,I401404,I401430,I401438,I401464,I401472,I401489,I401506,I401523,I401563,I401571,I401588,I401605,I401622,I401653,I401670,I401696,I401704,I401735,I401766,I401783,I401814,I401914,I706770,I401940,I401948,I401965,I706755,I706743,I401982,I706758,I402008,I402016,I706761,I402042,I402050,I402067,I402084,I402101,I706749,I402141,I402149,I402166,I402183,I402200,I402231,I706746,I706752,I402248,I706767,I402274,I402282,I402313,I402344,I402361,I402392,I706764,I402492,I402518,I402526,I402543,I402560,I402586,I402594,I402620,I402628,I402645,I402662,I402679,I402719,I402727,I402744,I402761,I402778,I402809,I402826,I402852,I402860,I402891,I402922,I402939,I402970,I403070,I403096,I403104,I403121,I403138,I403164,I403172,I403198,I403206,I403223,I403240,I403257,I403053,I403297,I403305,I403322,I403339,I403356,I403056,I403387,I403404,I403430,I403438,I403038,I403469,I403047,I403500,I403517,I403059,I403548,I403050,I403041,I403044,I403062,I403648,I403674,I403682,I403699,I403716,I403742,I403750,I403776,I403784,I403801,I403818,I403835,I403631,I403875,I403883,I403900,I403917,I403934,I403634,I403965,I403982,I404008,I404016,I403616,I404047,I403625,I404078,I404095,I403637,I404126,I403628,I403619,I403622,I403640,I404226,I550978,I404252,I404260,I404277,I550975,I550993,I404294,I550990,I404320,I404328,I550972,I404354,I404362,I404379,I404396,I404413,I404209,I550984,I404453,I404461,I404478,I404495,I404512,I404212,I404543,I550987,I404560,I404586,I404594,I404194,I404625,I404203,I404656,I404673,I404215,I404704,I550981,I404206,I404197,I404200,I404218,I404804,I404830,I404838,I404855,I404872,I404898,I404906,I404932,I404940,I404957,I404974,I404991,I405031,I405039,I405056,I405073,I405090,I405121,I405138,I405164,I405172,I405203,I405234,I405251,I405282,I405382,I480616,I405408,I405416,I405433,I480592,I480607,I405450,I480619,I405476,I405484,I480604,I480595,I405510,I405518,I405535,I405552,I405569,I405609,I405617,I405634,I405651,I405668,I405699,I480610,I480601,I405716,I480613,I405742,I405750,I405781,I405812,I405829,I405860,I480598,I405960,I405986,I405994,I406011,I406028,I406054,I406062,I406088,I406096,I406113,I406130,I406147,I406187,I406195,I406212,I406229,I406246,I406277,I406294,I406320,I406328,I406359,I406390,I406407,I406438,I406538,I406564,I406572,I406589,I406606,I406632,I406640,I406666,I406674,I406691,I406708,I406725,I406765,I406773,I406790,I406807,I406824,I406855,I406872,I406898,I406906,I406937,I406968,I406985,I407016,I407116,I407142,I407150,I407167,I407184,I407210,I407218,I407244,I407252,I407269,I407286,I407303,I407099,I407343,I407351,I407368,I407385,I407402,I407102,I407433,I407450,I407476,I407484,I407084,I407515,I407093,I407546,I407563,I407105,I407594,I407096,I407087,I407090,I407108,I407694,I407720,I407728,I407745,I407762,I407788,I407796,I407822,I407830,I407847,I407864,I407881,I407677,I407921,I407929,I407946,I407963,I407980,I407680,I408011,I408028,I408054,I408062,I407662,I408093,I407671,I408124,I408141,I407683,I408172,I407674,I407665,I407668,I407686,I408272,I740685,I408298,I408306,I408323,I740670,I740658,I408340,I740673,I408366,I408374,I740676,I408400,I408408,I408425,I408442,I408459,I740664,I408499,I408507,I408524,I408541,I408558,I408589,I740661,I740667,I408606,I740682,I408632,I408640,I408671,I408702,I408719,I408750,I740679,I408850,I408876,I408884,I408901,I408918,I408944,I408952,I408978,I408986,I409003,I409020,I409037,I408833,I409077,I409085,I409102,I409119,I409136,I408836,I409167,I409184,I409210,I409218,I408818,I409249,I408827,I409280,I409297,I408839,I409328,I408830,I408821,I408824,I408842,I409428,I409454,I409462,I409479,I409496,I409522,I409530,I409556,I409564,I409581,I409598,I409615,I409655,I409663,I409680,I409697,I409714,I409745,I409762,I409788,I409796,I409827,I409858,I409875,I409906,I410006,I410032,I410040,I410057,I410074,I410100,I410108,I410134,I410142,I410159,I410176,I410193,I410233,I410241,I410258,I410275,I410292,I410323,I410340,I410366,I410374,I410405,I410436,I410453,I410484,I410584,I598318,I410610,I410618,I410635,I598300,I598312,I410652,I598315,I410678,I410686,I598309,I598306,I410712,I410720,I410737,I410754,I410771,I410567,I598324,I410811,I410819,I410836,I410853,I410870,I410570,I410901,I598303,I410918,I410944,I410952,I410552,I410983,I410561,I411014,I411031,I410573,I411062,I598321,I410564,I410555,I410558,I410576,I411162,I411188,I411196,I411213,I411230,I411256,I411264,I411290,I411298,I411315,I411332,I411349,I411145,I411389,I411397,I411414,I411431,I411448,I411148,I411479,I411496,I411522,I411530,I411130,I411561,I411139,I411592,I411609,I411151,I411640,I411142,I411133,I411136,I411154,I411740,I411766,I411774,I411791,I411808,I411834,I411842,I411868,I411876,I411893,I411910,I411927,I411967,I411975,I411992,I412009,I412026,I412057,I412074,I412100,I412108,I412139,I412170,I412187,I412218,I412318,I412344,I412352,I412369,I412386,I412412,I412420,I412446,I412454,I412471,I412488,I412505,I412301,I412545,I412553,I412570,I412587,I412604,I412304,I412635,I412652,I412678,I412686,I412286,I412717,I412295,I412748,I412765,I412307,I412796,I412298,I412289,I412292,I412310,I412896,I412922,I412930,I412947,I412964,I412990,I412998,I413024,I413032,I413049,I413066,I413083,I413123,I413131,I413148,I413165,I413182,I413213,I413230,I413256,I413264,I413295,I413326,I413343,I413374,I413474,I413500,I413508,I413525,I413542,I413568,I413576,I413602,I413610,I413627,I413644,I413661,I413457,I413701,I413709,I413726,I413743,I413760,I413460,I413791,I413808,I413834,I413842,I413442,I413873,I413451,I413904,I413921,I413463,I413952,I413454,I413445,I413448,I413466,I414052,I553783,I414078,I414086,I414103,I553780,I553798,I414120,I553795,I414146,I414154,I553777,I414180,I414188,I414205,I414222,I414239,I553789,I414279,I414287,I414304,I414321,I414338,I414369,I553792,I414386,I414412,I414420,I414451,I414482,I414499,I414530,I553786,I414630,I544570,I414656,I414664,I414681,I544546,I544561,I414698,I544573,I414724,I414732,I544558,I544549,I414758,I414766,I414783,I414800,I414817,I414613,I414857,I414865,I414882,I414899,I414916,I414616,I414947,I544564,I544555,I414964,I544567,I414990,I414998,I414598,I415029,I414607,I415060,I415077,I414619,I415108,I544552,I414610,I414601,I414604,I414622,I415208,I473569,I415234,I415242,I415259,I473557,I473575,I415276,I473572,I415302,I415310,I473563,I473560,I415336,I415344,I415361,I415378,I415395,I473554,I415435,I415443,I415460,I415477,I415494,I415525,I415542,I415568,I415576,I415607,I415638,I415655,I415686,I473566,I415786,I415812,I415820,I415837,I415854,I415880,I415888,I415914,I415922,I415939,I415956,I415973,I416013,I416021,I416038,I416055,I416072,I416103,I416120,I416146,I416154,I416185,I416216,I416233,I416264,I416364,I416390,I416398,I416415,I416432,I416458,I416466,I416492,I416500,I416517,I416534,I416551,I416591,I416599,I416616,I416633,I416650,I416681,I416698,I416724,I416732,I416763,I416794,I416811,I416842,I416942,I416968,I416976,I416993,I417010,I417036,I417044,I417070,I417078,I417095,I417112,I417129,I417169,I417177,I417194,I417211,I417228,I417259,I417276,I417302,I417310,I417341,I417372,I417389,I417420,I417520,I417546,I417554,I417571,I417588,I417614,I417622,I417648,I417656,I417673,I417690,I417707,I417503,I417747,I417755,I417772,I417789,I417806,I417506,I417837,I417854,I417880,I417888,I417488,I417919,I417497,I417950,I417967,I417509,I417998,I417500,I417491,I417494,I417512,I418098,I418124,I418132,I418149,I418166,I418192,I418200,I418226,I418234,I418251,I418268,I418285,I418325,I418333,I418350,I418367,I418384,I418415,I418432,I418458,I418466,I418497,I418528,I418545,I418576,I418676,I418702,I418710,I418727,I418744,I418770,I418778,I418804,I418812,I418829,I418846,I418863,I418659,I418903,I418911,I418928,I418945,I418962,I418662,I418993,I419010,I419036,I419044,I418644,I419075,I418653,I419106,I419123,I418665,I419154,I418656,I418647,I418650,I418668,I419254,I636466,I419280,I419288,I419305,I636448,I636460,I419322,I636463,I419348,I419356,I636457,I636454,I419382,I419390,I419407,I419424,I419441,I636472,I419481,I419489,I419506,I419523,I419540,I419571,I636451,I419588,I419614,I419622,I419653,I419684,I419701,I419732,I636469,I419829,I419855,I419863,I419880,I419897,I419923,I419818,I419954,I419962,I419979,I420005,I420013,I419821,I420053,I419812,I419803,I420089,I420106,I420132,I420140,I420157,I419806,I420188,I420205,I420222,I419815,I420253,I419800,I420284,I420301,I419809,I420356,I586180,I420382,I420390,I420407,I586162,I420424,I586168,I420450,I420345,I586165,I420481,I420489,I586174,I420506,I420532,I420540,I420348,I586186,I420580,I420339,I420330,I420616,I586177,I586171,I420633,I420659,I420667,I420684,I420333,I420715,I586183,I420732,I420749,I420342,I420780,I420327,I420811,I420828,I420336,I420883,I420909,I420917,I420934,I420951,I420977,I421008,I421016,I421033,I421059,I421067,I421107,I421143,I421160,I421186,I421194,I421211,I421242,I421259,I421276,I421307,I421338,I421355,I421410,I486409,I421436,I421444,I421461,I486424,I486406,I421478,I421504,I486415,I421535,I421543,I486433,I421560,I421586,I421594,I486430,I421634,I421670,I486427,I486418,I421687,I486412,I421713,I421721,I421738,I421769,I486421,I421786,I421803,I421834,I421865,I421882,I421937,I421963,I421971,I421988,I422005,I422031,I422062,I422070,I422087,I422113,I422121,I422161,I422197,I422214,I422240,I422248,I422265,I422296,I422313,I422330,I422361,I422392,I422409,I422464,I422490,I422498,I422515,I422532,I422558,I422589,I422597,I422614,I422640,I422648,I422688,I422724,I422741,I422767,I422775,I422792,I422823,I422840,I422857,I422888,I422919,I422936,I422991,I423017,I423025,I423042,I423059,I423085,I423116,I423124,I423141,I423167,I423175,I423215,I423251,I423268,I423294,I423302,I423319,I423350,I423367,I423384,I423415,I423446,I423463,I423518,I710328,I423544,I423552,I423569,I710325,I710334,I423586,I710313,I423612,I710316,I423643,I423651,I710331,I423668,I423694,I423702,I710337,I423742,I423778,I710319,I710340,I423795,I710322,I423821,I423829,I423846,I423877,I423894,I423911,I423942,I423973,I423990,I424045,I424071,I424079,I424096,I424113,I424139,I424170,I424178,I424195,I424221,I424229,I424269,I424305,I424322,I424348,I424356,I424373,I424404,I424421,I424438,I424469,I424500,I424517,I424572,I424598,I424606,I424623,I424640,I424666,I424697,I424705,I424722,I424748,I424756,I424796,I424832,I424849,I424875,I424883,I424900,I424931,I424948,I424965,I424996,I425027,I425044,I425099,I425125,I425133,I425150,I425167,I425193,I425224,I425232,I425249,I425275,I425283,I425323,I425359,I425376,I425402,I425410,I425427,I425458,I425475,I425492,I425523,I425554,I425571,I425626,I425652,I425660,I425677,I425694,I425720,I425751,I425759,I425776,I425802,I425810,I425850,I425886,I425903,I425929,I425937,I425954,I425985,I426002,I426019,I426050,I426081,I426098,I426153,I426179,I426187,I426204,I426221,I426247,I426278,I426286,I426303,I426329,I426337,I426377,I426413,I426430,I426456,I426464,I426481,I426512,I426529,I426546,I426577,I426608,I426625,I426680,I426706,I426714,I426731,I426748,I426774,I426805,I426813,I426830,I426856,I426864,I426904,I426940,I426957,I426983,I426991,I427008,I427039,I427056,I427073,I427104,I427135,I427152,I427207,I580400,I427233,I427241,I427258,I580382,I427275,I580388,I427301,I427196,I580385,I427332,I427340,I580394,I427357,I427383,I427391,I427199,I580406,I427431,I427190,I427181,I427467,I580397,I580391,I427484,I427510,I427518,I427535,I427184,I427566,I580403,I427583,I427600,I427193,I427631,I427178,I427662,I427679,I427187,I427734,I427760,I427768,I427785,I427802,I427828,I427723,I427859,I427867,I427884,I427910,I427918,I427726,I427958,I427717,I427708,I427994,I428011,I428037,I428045,I428062,I427711,I428093,I428110,I428127,I427720,I428158,I427705,I428189,I428206,I427714,I428261,I428287,I428295,I428312,I428329,I428355,I428250,I428386,I428394,I428411,I428437,I428445,I428253,I428485,I428244,I428235,I428521,I428538,I428564,I428572,I428589,I428238,I428620,I428637,I428654,I428247,I428685,I428232,I428716,I428733,I428241,I428788,I595428,I428814,I428822,I428839,I595410,I428856,I595416,I428882,I595413,I428913,I428921,I595422,I428938,I428964,I428972,I595434,I429012,I429048,I595425,I595419,I429065,I429091,I429099,I429116,I429147,I595431,I429164,I429181,I429212,I429243,I429260,I429315,I429341,I429349,I429366,I429383,I429409,I429440,I429448,I429465,I429491,I429499,I429539,I429575,I429592,I429618,I429626,I429643,I429674,I429691,I429708,I429739,I429770,I429787,I429842,I590804,I429868,I429876,I429893,I590786,I429910,I590792,I429936,I429831,I590789,I429967,I429975,I590798,I429992,I430018,I430026,I429834,I590810,I430066,I429825,I429816,I430102,I590801,I590795,I430119,I430145,I430153,I430170,I429819,I430201,I590807,I430218,I430235,I429828,I430266,I429813,I430297,I430314,I429822,I430369,I430395,I430403,I430420,I430437,I430463,I430358,I430494,I430502,I430519,I430545,I430553,I430361,I430593,I430352,I430343,I430629,I430646,I430672,I430680,I430697,I430346,I430728,I430745,I430762,I430355,I430793,I430340,I430824,I430841,I430349,I430896,I556030,I430922,I430930,I430947,I556039,I556027,I430964,I556024,I430990,I430885,I431021,I431029,I556021,I431046,I431072,I431080,I430888,I431120,I430879,I430870,I431156,I556042,I556033,I431173,I556036,I431199,I431207,I431224,I430873,I431255,I431272,I431289,I430882,I431320,I430867,I431351,I431368,I430876,I431423,I431449,I431457,I431474,I431491,I431517,I431548,I431556,I431573,I431599,I431607,I431647,I431683,I431700,I431726,I431734,I431751,I431782,I431799,I431816,I431847,I431878,I431895,I431950,I431976,I431984,I432001,I432018,I432044,I432075,I432083,I432100,I432126,I432134,I432174,I432210,I432227,I432253,I432261,I432278,I432309,I432326,I432343,I432374,I432405,I432422,I432477,I727583,I432503,I432511,I432528,I727580,I727589,I432545,I727568,I432571,I727571,I432602,I432610,I727586,I432627,I432653,I432661,I727592,I432701,I432737,I727574,I727595,I432754,I727577,I432780,I432788,I432805,I432836,I432853,I432870,I432901,I432932,I432949,I433004,I696668,I433030,I433038,I433055,I696662,I696680,I433072,I696665,I433098,I696686,I433129,I433137,I696671,I433154,I433180,I433188,I696683,I433228,I433264,I696674,I696689,I433281,I696677,I433307,I433315,I433332,I433363,I433380,I433397,I433428,I433459,I433476,I433531,I433557,I433565,I433582,I433599,I433625,I433520,I433656,I433664,I433681,I433707,I433715,I433523,I433755,I433514,I433505,I433791,I433808,I433834,I433842,I433859,I433508,I433890,I433907,I433924,I433517,I433955,I433502,I433986,I434003,I433511,I434058,I586758,I434084,I434092,I434109,I586740,I434126,I586746,I434152,I434047,I586743,I434183,I434191,I586752,I434208,I434234,I434242,I434050,I586764,I434282,I434041,I434032,I434318,I586755,I586749,I434335,I434361,I434369,I434386,I434035,I434417,I586761,I434434,I434451,I434044,I434482,I434029,I434513,I434530,I434038,I434585,I736508,I434611,I434619,I434636,I736505,I736514,I434653,I736493,I434679,I736496,I434710,I434718,I736511,I434735,I434761,I434769,I736517,I434809,I434845,I736499,I736520,I434862,I736502,I434888,I434896,I434913,I434944,I434961,I434978,I435009,I435040,I435057,I435112,I514187,I435138,I435146,I435163,I514202,I514184,I435180,I435206,I514193,I435237,I435245,I514211,I435262,I435288,I435296,I514208,I435336,I435372,I514205,I514196,I435389,I514190,I435415,I435423,I435440,I435471,I514199,I435488,I435505,I435536,I435567,I435584,I435639,I435665,I435673,I435690,I435707,I435733,I435764,I435772,I435789,I435815,I435823,I435863,I435899,I435916,I435942,I435950,I435967,I435998,I436015,I436032,I436063,I436094,I436111,I436166,I436192,I436200,I436217,I436234,I436260,I436291,I436299,I436316,I436342,I436350,I436390,I436426,I436443,I436469,I436477,I436494,I436525,I436542,I436559,I436590,I436621,I436638,I436693,I436719,I436727,I436744,I436761,I436787,I436818,I436826,I436843,I436869,I436877,I436917,I436953,I436970,I436996,I437004,I437021,I437052,I437069,I437086,I437117,I437148,I437165,I437220,I476719,I437246,I437254,I437271,I476734,I476716,I437288,I437314,I476725,I437345,I437353,I476743,I437370,I437396,I437404,I476740,I437444,I437480,I476737,I476728,I437497,I476722,I437523,I437531,I437548,I437579,I476731,I437596,I437613,I437644,I437675,I437692,I437747,I551542,I437773,I437781,I437798,I551551,I551539,I437815,I551536,I437841,I437872,I437880,I551533,I437897,I437923,I437931,I437971,I438007,I551554,I551545,I438024,I551548,I438050,I438058,I438075,I438106,I438123,I438140,I438171,I438202,I438219,I438274,I438300,I438308,I438325,I438342,I438368,I438399,I438407,I438424,I438450,I438458,I438498,I438534,I438551,I438577,I438585,I438602,I438633,I438650,I438667,I438698,I438729,I438746,I438801,I438827,I438835,I438852,I438869,I438895,I438926,I438934,I438951,I438977,I438985,I439025,I439061,I439078,I439104,I439112,I439129,I439160,I439177,I439194,I439225,I439256,I439273,I439328,I439354,I439362,I439379,I439396,I439422,I439317,I439453,I439461,I439478,I439504,I439512,I439320,I439552,I439311,I439302,I439588,I439605,I439631,I439639,I439656,I439305,I439687,I439704,I439721,I439314,I439752,I439299,I439783,I439800,I439308,I439855,I439881,I439889,I439906,I439923,I439949,I439980,I439988,I440005,I440031,I440039,I440079,I440115,I440132,I440158,I440166,I440183,I440214,I440231,I440248,I440279,I440310,I440327,I440382,I583868,I440408,I440416,I440433,I583850,I440450,I583856,I440476,I440371,I583853,I440507,I440515,I583862,I440532,I440558,I440566,I440374,I583874,I440606,I440365,I440356,I440642,I583865,I583859,I440659,I440685,I440693,I440710,I440359,I440741,I583871,I440758,I440775,I440368,I440806,I440353,I440837,I440854,I440362,I440909,I440935,I440943,I440960,I440977,I441003,I440898,I441034,I441042,I441059,I441085,I441093,I440901,I441133,I440892,I440883,I441169,I441186,I441212,I441220,I441237,I440886,I441268,I441285,I441302,I440895,I441333,I440880,I441364,I441381,I440889,I441436,I653426,I441462,I441470,I441487,I653432,I653414,I441504,I653423,I441530,I653429,I441561,I441569,I653417,I441586,I441612,I441620,I653435,I441660,I441696,I653420,I441713,I653438,I441739,I441747,I441764,I441795,I441812,I441829,I441860,I441891,I441908,I441963,I741863,I441989,I441997,I442014,I741860,I741869,I442031,I741848,I442057,I741851,I442088,I442096,I741866,I442113,I442139,I442147,I741872,I442187,I442223,I741854,I741875,I442240,I741857,I442266,I442274,I442291,I442322,I442339,I442356,I442387,I442418,I442435,I442490,I649618,I442516,I442524,I442541,I649624,I649606,I442558,I649615,I442584,I649621,I442615,I442623,I649609,I442640,I442666,I442674,I649627,I442714,I442750,I649612,I442767,I649630,I442793,I442801,I442818,I442849,I442866,I442883,I442914,I442945,I442962,I443017,I443043,I443051,I443068,I443085,I443111,I443006,I443142,I443150,I443167,I443193,I443201,I443009,I443241,I443000,I442991,I443277,I443294,I443320,I443328,I443345,I442994,I443376,I443393,I443410,I443003,I443441,I442988,I443472,I443489,I442997,I443544,I646870,I443570,I443578,I443595,I646852,I443612,I646858,I443638,I646855,I443669,I443677,I646864,I443694,I443720,I443728,I646876,I443768,I443804,I646867,I646861,I443821,I443847,I443855,I443872,I443903,I646873,I443920,I443937,I443968,I443999,I444016,I444071,I444097,I444105,I444122,I444139,I444165,I444196,I444204,I444221,I444247,I444255,I444295,I444331,I444348,I444374,I444382,I444399,I444430,I444447,I444464,I444495,I444526,I444543,I444598,I596584,I444624,I444632,I444649,I596566,I444666,I596572,I444692,I444587,I596569,I444723,I444731,I596578,I444748,I444774,I444782,I444590,I596590,I444822,I444581,I444572,I444858,I596581,I596575,I444875,I444901,I444909,I444926,I444575,I444957,I596587,I444974,I444991,I444584,I445022,I444569,I445053,I445070,I444578,I445125,I514833,I445151,I445159,I445176,I514848,I514830,I445193,I445219,I514839,I445250,I445258,I514857,I445275,I445301,I445309,I514854,I445349,I445385,I514851,I514842,I445402,I514836,I445428,I445436,I445453,I445484,I514845,I445501,I445518,I445549,I445580,I445597,I445652,I615658,I445678,I445686,I445703,I615640,I445720,I615646,I445746,I615643,I445777,I445785,I615652,I445802,I445828,I445836,I615664,I445876,I445912,I615655,I615649,I445929,I445955,I445963,I445980,I446011,I615661,I446028,I446045,I446076,I446107,I446124,I446179,I446205,I446213,I446230,I446247,I446273,I446304,I446312,I446329,I446355,I446363,I446403,I446439,I446456,I446482,I446490,I446507,I446538,I446555,I446572,I446603,I446634,I446651,I446706,I446732,I446740,I446757,I446774,I446800,I446695,I446831,I446839,I446856,I446882,I446890,I446698,I446930,I446689,I446680,I446966,I446983,I447009,I447017,I447034,I446683,I447065,I447082,I447099,I446692,I447130,I446677,I447161,I447178,I446686,I447233,I447259,I447267,I447284,I447301,I447327,I447358,I447366,I447383,I447409,I447417,I447457,I447493,I447510,I447536,I447544,I447561,I447592,I447609,I447626,I447657,I447688,I447705,I447760,I504497,I447786,I447794,I447811,I504512,I504494,I447828,I447854,I447749,I504503,I447885,I447893,I504521,I447910,I447936,I447944,I447752,I504518,I447984,I447743,I447734,I448020,I504515,I504506,I448037,I504500,I448063,I448071,I448088,I447737,I448119,I504509,I448136,I448153,I447746,I448184,I447731,I448215,I448232,I447740,I448287,I686956,I448313,I448321,I448338,I686938,I686941,I448355,I686953,I448381,I686962,I448412,I448420,I686947,I448437,I448463,I448471,I686959,I448511,I448547,I686950,I686944,I448564,I448590,I448598,I448615,I448646,I448663,I448680,I448711,I448742,I448759,I448814,I448840,I448848,I448865,I448882,I448908,I448803,I448939,I448947,I448964,I448990,I448998,I448806,I449038,I448797,I448788,I449074,I449091,I449117,I449125,I449142,I448791,I449173,I449190,I449207,I448800,I449238,I448785,I449269,I449286,I448794,I449341,I619126,I449367,I449375,I449392,I619108,I449409,I619114,I449435,I619111,I449466,I449474,I619120,I449491,I449517,I449525,I619132,I449565,I449601,I619123,I619117,I449618,I449644,I449652,I449669,I449700,I619129,I449717,I449734,I449765,I449796,I449813,I449868,I449894,I449902,I449919,I449936,I449962,I449993,I450001,I450018,I450044,I450052,I450092,I450128,I450145,I450171,I450179,I450196,I450227,I450244,I450261,I450292,I450323,I450340,I450395,I631264,I450421,I450429,I450446,I631246,I450463,I631252,I450489,I450384,I631249,I450520,I450528,I631258,I450545,I450571,I450579,I450387,I631270,I450619,I450378,I450369,I450655,I631261,I631255,I450672,I450698,I450706,I450723,I450372,I450754,I631267,I450771,I450788,I450381,I450819,I450366,I450850,I450867,I450375,I450922,I450948,I450956,I450973,I450990,I451016,I451047,I451055,I451072,I451098,I451106,I451146,I451182,I451199,I451225,I451233,I451250,I451281,I451298,I451315,I451346,I451377,I451394,I451449,I487701,I451475,I451483,I451500,I487716,I487698,I451517,I451543,I487707,I451574,I451582,I487725,I451599,I451625,I451633,I487722,I451673,I451709,I487719,I487710,I451726,I487704,I451752,I451760,I451777,I451808,I487713,I451825,I451842,I451873,I451904,I451921,I451976,I488993,I452002,I452010,I452027,I489008,I488990,I452044,I452070,I451965,I488999,I452101,I452109,I489017,I452126,I452152,I452160,I451968,I489014,I452200,I451959,I451950,I452236,I489011,I489002,I452253,I488996,I452279,I452287,I452304,I451953,I452335,I489005,I452352,I452369,I451962,I452400,I451947,I452431,I452448,I451956,I452503,I611612,I452529,I452537,I452554,I611594,I452571,I611600,I452597,I452492,I611597,I452628,I452636,I611606,I452653,I452679,I452687,I452495,I611618,I452727,I452486,I452477,I452763,I611609,I611603,I452780,I452806,I452814,I452831,I452480,I452862,I611615,I452879,I452896,I452489,I452927,I452474,I452958,I452975,I452483,I453030,I453056,I453064,I453081,I453098,I453124,I453019,I453155,I453163,I453180,I453206,I453214,I453022,I453254,I453013,I453004,I453290,I453307,I453333,I453341,I453358,I453007,I453389,I453406,I453423,I453016,I453454,I453001,I453485,I453502,I453010,I453557,I638200,I453583,I453591,I453608,I638182,I453625,I638188,I453651,I453546,I638185,I453682,I453690,I638194,I453707,I453733,I453741,I453549,I638206,I453781,I453540,I453531,I453817,I638197,I638191,I453834,I453860,I453868,I453885,I453534,I453916,I638203,I453933,I453950,I453543,I453981,I453528,I454012,I454029,I453537,I454084,I454110,I454118,I454135,I454152,I454178,I454073,I454209,I454217,I454234,I454260,I454268,I454076,I454308,I454067,I454058,I454344,I454361,I454387,I454395,I454412,I454061,I454443,I454460,I454477,I454070,I454508,I454055,I454539,I454556,I454064,I454611,I454637,I454645,I454662,I454679,I454705,I454736,I454744,I454761,I454787,I454795,I454835,I454871,I454888,I454914,I454922,I454939,I454970,I454987,I455004,I455035,I455066,I455083,I455138,I455164,I455172,I455189,I455206,I455232,I455127,I455263,I455271,I455288,I455314,I455322,I455130,I455362,I455121,I455112,I455398,I455415,I455441,I455449,I455466,I455115,I455497,I455514,I455531,I455124,I455562,I455109,I455593,I455610,I455118,I455665,I455691,I455699,I455716,I455733,I455759,I455654,I455790,I455798,I455815,I455841,I455849,I455657,I455889,I455648,I455639,I455925,I455942,I455968,I455976,I455993,I455642,I456024,I456041,I456058,I455651,I456089,I455636,I456120,I456137,I455645,I456192,I456218,I456226,I456243,I456260,I456286,I456317,I456325,I456342,I456368,I456376,I456416,I456452,I456469,I456495,I456503,I456520,I456551,I456568,I456585,I456616,I456647,I456664,I456719,I456745,I456753,I456770,I456787,I456813,I456844,I456852,I456869,I456895,I456903,I456943,I456979,I456996,I457022,I457030,I457047,I457078,I457095,I457112,I457143,I457174,I457191,I457246,I585024,I457272,I457280,I457297,I585006,I457314,I585012,I457340,I457235,I585009,I457371,I457379,I585018,I457396,I457422,I457430,I457238,I585030,I457470,I457229,I457220,I457506,I585021,I585015,I457523,I457549,I457557,I457574,I457223,I457605,I585027,I457622,I457639,I457232,I457670,I457217,I457701,I457718,I457226,I457773,I457799,I457807,I457824,I457841,I457867,I457898,I457906,I457923,I457949,I457957,I457997,I458033,I458050,I458076,I458084,I458101,I458132,I458149,I458166,I458197,I458228,I458245,I458300,I644558,I458326,I458334,I458351,I644540,I458368,I644546,I458394,I458289,I644543,I458425,I458433,I644552,I458450,I458476,I458484,I458292,I644564,I458524,I458283,I458274,I458560,I644555,I644549,I458577,I458603,I458611,I458628,I458277,I458659,I644561,I458676,I458693,I458286,I458724,I458271,I458755,I458772,I458280,I458827,I496745,I458853,I458861,I458878,I496760,I496742,I458895,I458921,I496751,I458952,I458960,I496769,I458977,I459003,I459011,I496766,I459051,I459087,I496763,I496754,I459104,I496748,I459130,I459138,I459155,I459186,I496757,I459203,I459220,I459251,I459282,I459299,I459354,I646292,I459380,I459388,I459405,I646274,I459422,I646280,I459448,I646277,I459479,I459487,I646286,I459504,I459530,I459538,I646298,I459578,I459614,I646289,I646283,I459631,I459657,I459665,I459682,I459713,I646295,I459730,I459747,I459778,I459809,I459826,I459881,I459907,I459915,I459932,I459949,I459975,I460006,I460014,I460031,I460057,I460065,I460105,I460141,I460158,I460184,I460192,I460209,I460240,I460257,I460274,I460305,I460336,I460353,I460408,I525815,I460434,I460442,I460459,I525830,I525812,I460476,I460502,I525821,I460533,I460541,I525839,I460558,I460584,I460592,I525836,I460632,I460668,I525833,I525824,I460685,I525818,I460711,I460719,I460736,I460767,I525827,I460784,I460801,I460832,I460863,I460880,I460935,I617970,I460961,I460969,I460986,I617952,I461003,I617958,I461029,I460924,I617955,I461060,I461068,I617964,I461085,I461111,I461119,I460927,I617976,I461159,I460918,I460909,I461195,I617967,I617961,I461212,I461238,I461246,I461263,I460912,I461294,I617973,I461311,I461328,I460921,I461359,I460906,I461390,I461407,I460915,I461462,I461488,I461496,I461513,I461530,I461556,I461451,I461587,I461595,I461612,I461638,I461646,I461454,I461686,I461445,I461436,I461722,I461739,I461765,I461773,I461790,I461439,I461821,I461838,I461855,I461448,I461886,I461433,I461917,I461934,I461442,I461989,I462015,I462023,I462040,I462057,I462083,I461978,I462114,I462122,I462139,I462165,I462173,I461981,I462213,I461972,I461963,I462249,I462266,I462292,I462300,I462317,I461966,I462348,I462365,I462382,I461975,I462413,I461960,I462444,I462461,I461969,I462516,I462542,I462550,I462567,I462584,I462610,I462505,I462641,I462649,I462666,I462692,I462700,I462508,I462740,I462499,I462490,I462776,I462793,I462819,I462827,I462844,I462493,I462875,I462892,I462909,I462502,I462940,I462487,I462971,I462988,I462496,I463043,I463069,I463077,I463094,I463111,I463137,I463168,I463176,I463193,I463219,I463227,I463267,I463303,I463320,I463346,I463354,I463371,I463402,I463419,I463436,I463467,I463498,I463515,I463570,I463596,I463604,I463621,I463638,I463664,I463695,I463703,I463720,I463746,I463754,I463794,I463830,I463847,I463873,I463881,I463898,I463929,I463946,I463963,I463994,I464025,I464042,I464097,I563323,I464123,I464131,I464148,I563332,I563320,I464165,I563317,I464191,I464086,I464222,I464230,I563314,I464247,I464273,I464281,I464089,I464321,I464080,I464071,I464357,I563335,I563326,I464374,I563329,I464400,I464408,I464425,I464074,I464456,I464473,I464490,I464083,I464521,I464068,I464552,I464569,I464077,I464624,I464650,I464658,I464675,I464692,I464718,I464613,I464749,I464757,I464774,I464800,I464808,I464616,I464848,I464607,I464598,I464884,I464901,I464927,I464935,I464952,I464601,I464983,I465000,I465017,I464610,I465048,I464595,I465079,I465096,I464604,I465151,I465177,I465185,I465202,I465219,I465245,I465276,I465284,I465301,I465327,I465335,I465375,I465411,I465428,I465454,I465462,I465479,I465510,I465527,I465544,I465575,I465606,I465623,I465678,I465704,I465712,I465729,I465746,I465772,I465803,I465811,I465828,I465854,I465862,I465902,I465938,I465955,I465981,I465989,I466006,I466037,I466054,I466071,I466102,I466133,I466150,I466205,I712113,I466231,I466239,I466256,I712110,I712119,I466273,I712098,I466299,I466194,I712101,I466330,I466338,I712116,I466355,I466381,I466389,I466197,I712122,I466429,I466188,I466179,I466465,I712104,I712125,I466482,I712107,I466508,I466516,I466533,I466182,I466564,I466581,I466598,I466191,I466629,I466176,I466660,I466677,I466185,I466732,I466758,I466766,I466783,I466800,I466826,I466857,I466865,I466882,I466908,I466916,I466956,I466992,I467009,I467035,I467043,I467060,I467091,I467108,I467125,I467156,I467187,I467204,I467259,I467285,I467293,I467310,I467327,I467353,I467384,I467392,I467409,I467435,I467443,I467483,I467519,I467536,I467562,I467570,I467587,I467618,I467635,I467652,I467683,I467714,I467731,I467786,I500621,I467812,I467820,I467837,I500636,I500618,I467854,I467880,I467775,I500627,I467911,I467919,I500645,I467936,I467962,I467970,I467778,I500642,I468010,I467769,I467760,I468046,I500639,I500630,I468063,I500624,I468089,I468097,I468114,I467763,I468145,I500633,I468162,I468179,I467772,I468210,I467757,I468241,I468258,I467766,I468313,I468339,I468347,I468364,I468381,I468407,I468302,I468438,I468446,I468463,I468489,I468497,I468305,I468537,I468296,I468287,I468573,I468590,I468616,I468624,I468641,I468290,I468672,I468689,I468706,I468299,I468737,I468284,I468768,I468785,I468293,I468840,I468866,I468874,I468891,I468908,I468934,I468965,I468973,I468990,I469016,I469024,I469064,I469100,I469117,I469143,I469151,I469168,I469199,I469216,I469233,I469264,I469295,I469312,I469367,I710923,I469393,I469401,I469418,I710920,I710929,I469435,I710908,I469461,I710911,I469492,I469500,I710926,I469517,I469543,I469551,I710932,I469591,I469627,I710914,I710935,I469644,I710917,I469670,I469678,I469695,I469726,I469743,I469760,I469791,I469822,I469839,I469894,I469920,I469928,I469945,I469962,I469988,I470019,I470027,I470044,I470070,I470078,I470118,I470154,I470171,I470197,I470205,I470222,I470253,I470270,I470287,I470318,I470349,I470366,I470421,I470447,I470455,I470472,I470489,I470515,I470410,I470546,I470554,I470571,I470597,I470605,I470413,I470645,I470404,I470395,I470681,I470698,I470724,I470732,I470749,I470398,I470780,I470797,I470814,I470407,I470845,I470392,I470876,I470893,I470401,I470948,I700808,I470974,I470982,I470999,I700805,I700814,I471016,I700793,I471042,I700796,I471073,I471081,I700811,I471098,I471124,I471132,I700817,I471172,I471208,I700799,I700820,I471225,I700802,I471251,I471259,I471276,I471307,I471324,I471341,I471372,I471403,I471420,I471475,I532275,I471501,I471509,I471526,I532290,I532272,I471543,I471569,I532281,I471600,I471608,I532299,I471625,I471651,I471659,I532296,I471699,I471735,I532293,I532284,I471752,I532278,I471778,I471786,I471803,I471834,I532287,I471851,I471868,I471899,I471930,I471947,I472002,I615080,I472028,I472036,I472053,I615062,I472070,I615068,I472096,I471991,I615065,I472127,I472135,I615074,I472152,I472178,I472186,I471994,I615086,I472226,I471985,I471976,I472262,I615077,I615071,I472279,I472305,I472313,I472330,I471979,I472361,I615083,I472378,I472395,I471988,I472426,I471973,I472457,I472474,I471982,I472529,I472555,I472563,I472580,I472597,I472623,I472654,I472662,I472679,I472705,I472713,I472753,I472789,I472806,I472832,I472840,I472857,I472888,I472905,I472922,I472953,I472984,I473001,I473056,I473082,I473090,I473107,I473124,I473150,I473181,I473189,I473206,I473232,I473240,I473280,I473316,I473333,I473359,I473367,I473384,I473415,I473432,I473449,I473480,I473511,I473528,I473583,I473609,I473617,I473634,I473651,I473677,I473708,I473716,I473733,I473759,I473767,I473807,I473843,I473860,I473886,I473894,I473911,I473942,I473959,I473976,I474007,I474038,I474055,I474110,I638778,I474136,I474144,I474161,I638760,I474178,I638766,I474204,I638763,I474235,I474243,I638772,I474260,I474286,I474294,I638784,I474334,I474370,I638775,I638769,I474387,I474413,I474421,I474438,I474469,I638781,I474486,I474503,I474534,I474565,I474582,I474637,I474663,I474671,I474688,I474705,I474731,I474762,I474770,I474787,I474813,I474821,I474861,I474897,I474914,I474940,I474948,I474965,I474996,I475013,I475030,I475061,I475092,I475109,I475164,I498037,I475190,I475198,I475215,I498052,I498034,I475232,I475258,I498043,I475289,I475297,I498061,I475314,I475340,I475348,I498058,I475388,I475424,I498055,I498046,I475441,I498040,I475467,I475475,I475492,I475523,I498049,I475540,I475557,I475588,I475619,I475636,I475691,I475717,I475725,I475742,I475759,I475785,I475680,I475816,I475824,I475841,I475867,I475875,I475683,I475915,I475674,I475665,I475951,I475968,I475994,I476002,I476019,I475668,I476050,I476067,I476084,I475677,I476115,I475662,I476146,I476163,I475671,I476218,I622594,I476244,I476252,I476269,I622576,I476286,I622582,I476312,I622579,I476343,I476351,I622588,I476368,I476394,I476402,I622600,I476442,I476478,I622591,I622585,I476495,I476521,I476529,I476546,I476577,I622597,I476594,I476611,I476642,I476673,I476690,I476751,I476777,I476794,I476802,I476819,I476836,I476853,I476870,I476887,I476918,I476935,I476966,I476983,I477000,I477031,I477071,I477079,I477096,I477113,I477130,I477161,I477178,I477195,I477221,I477243,I477260,I477291,I477336,I477397,I477423,I477440,I477448,I477465,I477482,I477499,I477516,I477533,I477383,I477564,I477581,I477386,I477612,I477629,I477646,I477362,I477677,I477374,I477717,I477725,I477742,I477759,I477776,I477389,I477807,I477824,I477841,I477867,I477377,I477889,I477906,I477371,I477937,I477365,I477368,I477982,I477380,I478043,I478069,I478086,I478094,I478111,I478128,I478145,I478162,I478179,I478210,I478227,I478258,I478275,I478292,I478323,I478363,I478371,I478388,I478405,I478422,I478453,I478470,I478487,I478513,I478535,I478552,I478583,I478628,I478689,I478715,I478732,I478740,I478757,I478774,I478791,I478808,I478825,I478856,I478873,I478904,I478921,I478938,I478969,I479009,I479017,I479034,I479051,I479068,I479099,I479116,I479133,I479159,I479181,I479198,I479229,I479274,I479335,I479361,I479378,I479386,I479403,I479420,I479437,I479454,I479471,I479502,I479519,I479550,I479567,I479584,I479615,I479655,I479663,I479680,I479697,I479714,I479745,I479762,I479779,I479805,I479827,I479844,I479875,I479920,I479981,I480007,I480024,I480032,I480049,I480066,I480083,I480100,I480117,I480148,I480165,I480196,I480213,I480230,I480261,I480301,I480309,I480326,I480343,I480360,I480391,I480408,I480425,I480451,I480473,I480490,I480521,I480566,I480627,I480653,I480670,I480678,I480695,I480712,I480729,I480746,I480763,I480794,I480811,I480842,I480859,I480876,I480907,I480947,I480955,I480972,I480989,I481006,I481037,I481054,I481071,I481097,I481119,I481136,I481167,I481212,I481273,I481299,I481316,I481324,I481341,I481358,I481375,I481392,I481409,I481440,I481457,I481488,I481505,I481522,I481553,I481593,I481601,I481618,I481635,I481652,I481683,I481700,I481717,I481743,I481765,I481782,I481813,I481858,I481919,I481945,I481962,I481970,I481987,I482004,I482021,I482038,I482055,I482086,I482103,I482134,I482151,I482168,I482199,I482239,I482247,I482264,I482281,I482298,I482329,I482346,I482363,I482389,I482411,I482428,I482459,I482504,I482565,I554338,I482591,I554341,I482608,I482616,I482633,I482650,I554350,I482667,I554359,I482684,I554347,I482701,I482551,I482732,I482749,I482554,I482780,I482797,I554353,I482814,I482530,I482845,I482542,I482885,I482893,I482910,I482927,I554344,I482944,I482557,I482975,I554356,I482992,I483009,I483035,I482545,I483057,I483074,I482539,I483105,I482533,I482536,I483150,I482548,I483211,I483237,I483254,I483262,I483279,I483296,I483313,I483330,I483347,I483378,I483395,I483426,I483443,I483460,I483491,I483531,I483539,I483556,I483573,I483590,I483621,I483638,I483655,I483681,I483703,I483720,I483751,I483796,I483857,I483883,I483900,I483908,I483925,I483942,I483959,I483976,I483993,I484024,I484041,I484072,I484089,I484106,I484137,I484177,I484185,I484202,I484219,I484236,I484267,I484284,I484301,I484327,I484349,I484366,I484397,I484442,I484503,I484529,I484546,I484554,I484571,I484588,I484605,I484622,I484639,I484489,I484670,I484687,I484492,I484718,I484735,I484752,I484468,I484783,I484480,I484823,I484831,I484848,I484865,I484882,I484495,I484913,I484930,I484947,I484973,I484483,I484995,I485012,I484477,I485043,I484471,I484474,I485088,I484486,I485149,I485175,I485192,I485200,I485217,I485234,I485251,I485268,I485285,I485316,I485333,I485364,I485381,I485398,I485429,I485469,I485477,I485494,I485511,I485528,I485559,I485576,I485593,I485619,I485641,I485658,I485689,I485734,I485795,I549850,I485821,I549853,I485838,I485846,I485863,I485880,I549862,I485897,I549871,I485914,I549859,I485931,I485962,I485979,I486010,I486027,I549865,I486044,I486075,I486115,I486123,I486140,I486157,I549856,I486174,I486205,I549868,I486222,I486239,I486265,I486287,I486304,I486335,I486380,I486441,I548728,I486467,I548731,I486484,I486492,I486509,I486526,I548740,I486543,I548749,I486560,I548737,I486577,I486608,I486625,I486656,I486673,I548743,I486690,I486721,I486761,I486769,I486786,I486803,I548734,I486820,I486851,I548746,I486868,I486885,I486911,I486933,I486950,I486981,I487026,I487087,I487113,I487130,I487138,I487155,I487172,I487189,I487206,I487223,I487073,I487254,I487271,I487076,I487302,I487319,I487336,I487052,I487367,I487064,I487407,I487415,I487432,I487449,I487466,I487079,I487497,I487514,I487531,I487557,I487067,I487579,I487596,I487061,I487627,I487055,I487058,I487672,I487070,I487733,I487759,I487776,I487784,I487801,I487818,I487835,I487852,I487869,I487900,I487917,I487948,I487965,I487982,I488013,I488053,I488061,I488078,I488095,I488112,I488143,I488160,I488177,I488203,I488225,I488242,I488273,I488318,I488379,I488405,I488422,I488430,I488447,I488464,I488481,I488498,I488515,I488546,I488563,I488594,I488611,I488628,I488659,I488699,I488707,I488724,I488741,I488758,I488789,I488806,I488823,I488849,I488871,I488888,I488919,I488964,I489025,I601786,I489051,I601768,I489068,I489076,I489093,I601777,I489110,I601789,I489127,I601771,I489144,I601780,I489161,I489192,I489209,I489240,I489257,I601792,I489274,I489305,I489345,I489353,I489370,I489387,I489404,I489435,I601774,I489452,I601783,I489469,I489495,I489517,I489534,I489565,I489610,I489671,I601208,I489697,I601190,I489714,I489722,I489739,I601199,I489756,I601211,I489773,I601193,I489790,I601202,I489807,I489838,I489855,I489886,I489903,I601214,I489920,I489951,I489991,I489999,I490016,I490033,I490050,I490081,I601196,I490098,I601205,I490115,I490141,I490163,I490180,I490211,I490256,I490317,I490343,I490360,I490368,I490385,I490402,I490419,I490436,I490453,I490484,I490501,I490532,I490549,I490566,I490597,I490637,I490645,I490662,I490679,I490696,I490727,I490744,I490761,I490787,I490809,I490826,I490857,I490902,I490963,I568924,I490989,I568927,I491006,I491014,I491031,I491048,I568936,I491065,I568945,I491082,I568933,I491099,I491130,I491147,I491178,I491195,I568939,I491212,I491243,I491283,I491291,I491308,I491325,I568930,I491342,I491373,I568942,I491390,I491407,I491433,I491455,I491472,I491503,I491548,I491609,I491635,I491652,I491660,I491677,I491694,I491711,I491728,I491745,I491776,I491793,I491824,I491841,I491858,I491889,I491929,I491937,I491954,I491971,I491988,I492019,I492036,I492053,I492079,I492101,I492118,I492149,I492194,I492255,I492281,I492298,I492306,I492323,I492340,I492357,I492374,I492391,I492241,I492422,I492439,I492244,I492470,I492487,I492504,I492220,I492535,I492232,I492575,I492583,I492600,I492617,I492634,I492247,I492665,I492682,I492699,I492725,I492235,I492747,I492764,I492229,I492795,I492223,I492226,I492840,I492238,I492901,I682901,I492927,I682895,I492944,I492952,I492969,I682904,I492986,I682916,I493003,I682898,I493020,I493037,I492887,I493068,I493085,I492890,I493116,I493133,I682892,I493150,I492866,I493181,I492878,I493221,I493229,I493246,I493263,I682913,I493280,I492893,I493311,I682907,I493328,I493345,I682910,I493371,I492881,I493393,I493410,I492875,I493441,I492869,I492872,I493486,I492884,I493547,I493573,I493590,I493598,I493615,I493632,I493649,I493666,I493683,I493714,I493731,I493762,I493779,I493796,I493827,I493867,I493875,I493892,I493909,I493926,I493957,I493974,I493991,I494017,I494039,I494056,I494087,I494132,I494193,I647448,I494219,I647454,I494236,I494244,I494261,I647451,I494278,I647430,I494295,I647433,I494312,I647439,I494329,I494360,I494377,I494408,I494425,I494442,I494473,I494513,I494521,I494538,I494555,I647442,I494572,I494603,I494620,I647436,I494637,I647445,I494663,I494685,I494702,I494733,I494778,I494839,I494865,I494882,I494890,I494907,I494924,I494941,I494958,I494975,I495006,I495023,I495054,I495071,I495088,I495119,I495159,I495167,I495184,I495201,I495218,I495249,I495266,I495283,I495309,I495331,I495348,I495379,I495424,I495485,I495511,I495528,I495536,I495553,I495570,I495587,I495604,I495621,I495471,I495652,I495669,I495474,I495700,I495717,I495734,I495450,I495765,I495462,I495805,I495813,I495830,I495847,I495864,I495477,I495895,I495912,I495929,I495955,I495465,I495977,I495994,I495459,I496025,I495453,I495456,I496070,I495468,I496131,I726973,I496157,I726997,I496174,I496182,I496199,I726979,I496216,I726988,I496233,I496250,I726994,I496267,I496298,I496315,I496346,I496363,I726991,I496380,I496411,I496451,I496459,I496476,I496493,I726985,I496510,I496541,I726976,I496558,I727000,I496575,I726982,I496601,I496623,I496640,I496671,I496716,I496777,I496803,I496820,I496828,I496845,I496862,I496879,I496896,I496913,I496944,I496961,I496992,I497009,I497026,I497057,I497097,I497105,I497122,I497139,I497156,I497187,I497204,I497221,I497247,I497269,I497286,I497317,I497362,I497423,I497449,I497466,I497474,I497491,I497508,I497525,I497542,I497559,I497590,I497607,I497638,I497655,I497672,I497703,I497743,I497751,I497768,I497785,I497802,I497833,I497850,I497867,I497893,I497915,I497932,I497963,I498008,I498069,I498095,I498112,I498120,I498137,I498154,I498171,I498188,I498205,I498236,I498253,I498284,I498301,I498318,I498349,I498389,I498397,I498414,I498431,I498448,I498479,I498496,I498513,I498539,I498561,I498578,I498609,I498654,I498715,I498741,I498758,I498766,I498783,I498800,I498817,I498834,I498851,I498701,I498882,I498899,I498704,I498930,I498947,I498964,I498680,I498995,I498692,I499035,I499043,I499060,I499077,I499094,I498707,I499125,I499142,I499159,I499185,I498695,I499207,I499224,I498689,I499255,I498683,I498686,I499300,I498698,I499361,I499387,I499404,I499412,I499429,I499446,I499463,I499480,I499497,I499528,I499545,I499576,I499593,I499610,I499641,I499681,I499689,I499706,I499723,I499740,I499771,I499788,I499805,I499831,I499853,I499870,I499901,I499946,I500007,I500033,I500050,I500058,I500075,I500092,I500109,I500126,I500143,I500174,I500191,I500222,I500239,I500256,I500287,I500327,I500335,I500352,I500369,I500386,I500417,I500434,I500451,I500477,I500499,I500516,I500547,I500592,I500653,I500679,I500696,I500704,I500721,I500738,I500755,I500772,I500789,I500820,I500837,I500868,I500885,I500902,I500933,I500973,I500981,I500998,I501015,I501032,I501063,I501080,I501097,I501123,I501145,I501162,I501193,I501238,I501299,I501325,I501342,I501350,I501367,I501384,I501401,I501418,I501435,I501466,I501483,I501514,I501531,I501548,I501579,I501619,I501627,I501644,I501661,I501678,I501709,I501726,I501743,I501769,I501791,I501808,I501839,I501884,I501945,I501971,I501988,I501996,I502013,I502030,I502047,I502064,I502081,I501931,I502112,I502129,I501934,I502160,I502177,I502194,I501910,I502225,I501922,I502265,I502273,I502290,I502307,I502324,I501937,I502355,I502372,I502389,I502415,I501925,I502437,I502454,I501919,I502485,I501913,I501916,I502530,I501928,I502591,I502617,I502634,I502642,I502659,I502676,I502693,I502710,I502727,I502758,I502775,I502806,I502823,I502840,I502871,I502911,I502919,I502936,I502953,I502970,I503001,I503018,I503035,I503061,I503083,I503100,I503131,I503176,I503237,I503263,I503280,I503288,I503305,I503322,I503339,I503356,I503373,I503404,I503421,I503452,I503469,I503486,I503517,I503557,I503565,I503582,I503599,I503616,I503647,I503664,I503681,I503707,I503729,I503746,I503777,I503822,I503883,I503909,I503926,I503934,I503951,I503968,I503985,I504002,I504019,I503869,I504050,I504067,I503872,I504098,I504115,I504132,I503848,I504163,I503860,I504203,I504211,I504228,I504245,I504262,I503875,I504293,I504310,I504327,I504353,I503863,I504375,I504392,I503857,I504423,I503851,I503854,I504468,I503866,I504529,I504555,I504572,I504580,I504597,I504614,I504631,I504648,I504665,I504696,I504713,I504744,I504761,I504778,I504809,I504849,I504857,I504874,I504891,I504908,I504939,I504956,I504973,I504999,I505021,I505038,I505069,I505114,I505175,I505201,I505218,I505226,I505243,I505260,I505277,I505294,I505311,I505342,I505359,I505390,I505407,I505424,I505455,I505495,I505503,I505520,I505537,I505554,I505585,I505602,I505619,I505645,I505667,I505684,I505715,I505760,I505821,I505847,I505864,I505872,I505889,I505906,I505923,I505940,I505957,I505988,I506005,I506036,I506053,I506070,I506101,I506141,I506149,I506166,I506183,I506200,I506231,I506248,I506265,I506291,I506313,I506330,I506361,I506406,I506467,I506493,I506510,I506518,I506535,I506552,I506569,I506586,I506603,I506634,I506651,I506682,I506699,I506716,I506747,I506787,I506795,I506812,I506829,I506846,I506877,I506894,I506911,I506937,I506959,I506976,I507007,I507052,I507113,I507139,I507156,I507164,I507181,I507198,I507215,I507232,I507249,I507280,I507297,I507328,I507345,I507362,I507393,I507433,I507441,I507458,I507475,I507492,I507523,I507540,I507557,I507583,I507605,I507622,I507653,I507698,I507759,I507785,I507802,I507810,I507827,I507844,I507861,I507878,I507895,I507745,I507926,I507943,I507748,I507974,I507991,I508008,I507724,I508039,I507736,I508079,I508087,I508104,I508121,I508138,I507751,I508169,I508186,I508203,I508229,I507739,I508251,I508268,I507733,I508299,I507727,I507730,I508344,I507742,I508405,I743038,I508431,I743062,I508448,I508456,I508473,I743044,I508490,I743053,I508507,I508524,I743059,I508541,I508572,I508589,I508620,I508637,I743056,I508654,I508685,I508725,I508733,I508750,I508767,I743050,I508784,I508815,I743041,I508832,I743065,I508849,I743047,I508875,I508897,I508914,I508945,I508990,I509051,I509077,I509094,I509102,I509119,I509136,I509153,I509170,I509187,I509037,I509218,I509235,I509040,I509266,I509283,I509300,I509016,I509331,I509028,I509371,I509379,I509396,I509413,I509430,I509043,I509461,I509478,I509495,I509521,I509031,I509543,I509560,I509025,I509591,I509019,I509022,I509636,I509034,I509697,I509723,I509740,I509748,I509765,I509782,I509799,I509816,I509833,I509864,I509881,I509912,I509929,I509946,I509977,I510017,I510025,I510042,I510059,I510076,I510107,I510124,I510141,I510167,I510189,I510206,I510237,I510282,I510343,I510369,I510386,I510394,I510411,I510428,I510445,I510462,I510479,I510329,I510510,I510527,I510332,I510558,I510575,I510592,I510308,I510623,I510320,I510663,I510671,I510688,I510705,I510722,I510335,I510753,I510770,I510787,I510813,I510323,I510835,I510852,I510317,I510883,I510311,I510314,I510928,I510326,I510989,I566680,I511015,I566683,I511032,I511040,I511057,I511074,I566692,I511091,I566701,I511108,I566689,I511125,I511156,I511173,I511204,I511221,I566695,I511238,I511269,I511309,I511317,I511334,I511351,I566686,I511368,I511399,I566698,I511416,I511433,I511459,I511481,I511498,I511529,I511574,I511635,I511661,I511678,I511686,I511703,I511720,I511737,I511754,I511771,I511802,I511819,I511850,I511867,I511884,I511915,I511955,I511963,I511980,I511997,I512014,I512045,I512062,I512079,I512105,I512127,I512144,I512175,I512220,I512281,I724593,I512307,I724617,I512324,I512332,I512349,I724599,I512366,I724608,I512383,I512400,I724614,I512417,I512267,I512448,I512465,I512270,I512496,I512513,I724611,I512530,I512246,I512561,I512258,I512601,I512609,I512626,I512643,I724605,I512660,I512273,I512691,I724596,I512708,I724620,I512725,I724602,I512751,I512261,I512773,I512790,I512255,I512821,I512249,I512252,I512866,I512264,I512927,I512953,I512970,I512978,I512995,I513012,I513029,I513046,I513063,I512913,I513094,I513111,I512916,I513142,I513159,I513176,I512892,I513207,I512904,I513247,I513255,I513272,I513289,I513306,I512919,I513337,I513354,I513371,I513397,I512907,I513419,I513436,I512901,I513467,I512895,I512898,I513512,I512910,I513573,I513599,I513616,I513624,I513641,I513658,I513675,I513692,I513709,I513740,I513757,I513788,I513805,I513822,I513853,I513893,I513901,I513918,I513935,I513952,I513983,I514000,I514017,I514043,I514065,I514082,I514113,I514158,I514219,I514245,I514262,I514270,I514287,I514304,I514321,I514338,I514355,I514386,I514403,I514434,I514451,I514468,I514499,I514539,I514547,I514564,I514581,I514598,I514629,I514646,I514663,I514689,I514711,I514728,I514759,I514804,I514865,I626640,I514891,I626622,I514908,I514916,I514933,I626631,I514950,I626643,I514967,I626625,I514984,I626634,I515001,I515032,I515049,I515080,I515097,I626646,I515114,I515145,I515185,I515193,I515210,I515227,I515244,I515275,I626628,I515292,I626637,I515309,I515335,I515357,I515374,I515405,I515450,I515511,I668664,I515537,I668670,I515554,I515562,I515579,I668667,I515596,I668646,I515613,I668649,I515630,I668655,I515647,I515678,I515695,I515726,I515743,I515760,I515791,I515831,I515839,I515856,I515873,I668658,I515890,I515921,I515938,I668652,I515955,I668661,I515981,I516003,I516020,I516051,I516096,I516157,I516183,I516200,I516208,I516225,I516242,I516259,I516276,I516293,I516324,I516341,I516372,I516389,I516406,I516437,I516477,I516485,I516502,I516519,I516536,I516567,I516584,I516601,I516627,I516649,I516666,I516697,I516742,I516803,I516829,I516846,I516854,I516871,I516888,I516905,I516922,I516939,I516970,I516987,I517018,I517035,I517052,I517083,I517123,I517131,I517148,I517165,I517182,I517213,I517230,I517247,I517273,I517295,I517312,I517343,I517388,I517449,I716263,I517475,I716287,I517492,I517500,I517517,I716269,I517534,I716278,I517551,I517568,I716284,I517585,I517616,I517633,I517664,I517681,I716281,I517698,I517729,I517769,I517777,I517794,I517811,I716275,I517828,I517859,I716266,I517876,I716290,I517893,I716272,I517919,I517941,I517958,I517989,I518034,I518095,I518121,I518138,I518146,I518163,I518180,I518197,I518214,I518231,I518081,I518262,I518279,I518084,I518310,I518327,I518344,I518060,I518375,I518072,I518415,I518423,I518440,I518457,I518474,I518087,I518505,I518522,I518539,I518565,I518075,I518587,I518604,I518069,I518635,I518063,I518066,I518680,I518078,I518741,I518767,I518784,I518792,I518809,I518826,I518843,I518860,I518877,I518908,I518925,I518956,I518973,I518990,I519021,I519061,I519069,I519086,I519103,I519120,I519151,I519168,I519185,I519211,I519233,I519250,I519281,I519326,I519387,I519413,I519430,I519438,I519455,I519472,I519489,I519506,I519523,I519554,I519571,I519602,I519619,I519636,I519667,I519707,I519715,I519732,I519749,I519766,I519797,I519814,I519831,I519857,I519879,I519896,I519927,I519972,I520033,I520059,I520076,I520084,I520101,I520118,I520135,I520152,I520169,I520200,I520217,I520248,I520265,I520282,I520313,I520353,I520361,I520378,I520395,I520412,I520443,I520460,I520477,I520503,I520525,I520542,I520573,I520618,I520679,I520705,I520722,I520730,I520747,I520764,I520781,I520798,I520815,I520846,I520863,I520894,I520911,I520928,I520959,I520999,I521007,I521024,I521041,I521058,I521089,I521106,I521123,I521149,I521171,I521188,I521219,I521264,I521325,I611034,I521351,I611016,I521368,I521376,I521393,I611025,I521410,I611037,I521427,I611019,I521444,I611028,I521461,I521492,I521509,I521540,I521557,I611040,I521574,I521605,I521645,I521653,I521670,I521687,I521704,I521735,I611022,I521752,I611031,I521769,I521795,I521817,I521834,I521865,I521910,I521971,I521997,I522014,I522022,I522039,I522056,I522073,I522090,I522107,I521957,I522138,I522155,I521960,I522186,I522203,I522220,I521936,I522251,I521948,I522291,I522299,I522316,I522333,I522350,I521963,I522381,I522398,I522415,I522441,I521951,I522463,I522480,I521945,I522511,I521939,I521942,I522556,I521954,I522617,I577510,I522643,I577492,I522660,I522668,I522685,I577501,I522702,I577513,I522719,I577495,I522736,I577504,I522753,I522784,I522801,I522832,I522849,I577516,I522866,I522897,I522937,I522945,I522962,I522979,I522996,I523027,I577498,I523044,I577507,I523061,I523087,I523109,I523126,I523157,I523202,I523263,I523289,I523306,I523314,I523331,I523348,I523365,I523382,I523399,I523249,I523430,I523447,I523252,I523478,I523495,I523512,I523228,I523543,I523240,I523583,I523591,I523608,I523625,I523642,I523255,I523673,I523690,I523707,I523733,I523243,I523755,I523772,I523237,I523803,I523231,I523234,I523848,I523246,I523909,I523935,I523952,I523960,I523977,I523994,I524011,I524028,I524045,I524076,I524093,I524124,I524141,I524158,I524189,I524229,I524237,I524254,I524271,I524288,I524319,I524336,I524353,I524379,I524401,I524418,I524449,I524494,I524555,I524581,I524598,I524606,I524623,I524640,I524657,I524674,I524691,I524541,I524722,I524739,I524544,I524770,I524787,I524804,I524520,I524835,I524532,I524875,I524883,I524900,I524917,I524934,I524547,I524965,I524982,I524999,I525025,I524535,I525047,I525064,I524529,I525095,I524523,I524526,I525140,I524538,I525201,I614502,I525227,I614484,I525244,I525252,I525269,I614493,I525286,I614505,I525303,I614487,I525320,I614496,I525337,I525368,I525385,I525416,I525433,I614508,I525450,I525481,I525521,I525529,I525546,I525563,I525580,I525611,I614490,I525628,I614499,I525645,I525671,I525693,I525710,I525741,I525786,I525847,I525873,I525890,I525898,I525915,I525932,I525949,I525966,I525983,I526014,I526031,I526062,I526079,I526096,I526127,I526167,I526175,I526192,I526209,I526226,I526257,I526274,I526291,I526317,I526339,I526356,I526387,I526432,I526493,I694433,I526519,I694430,I526536,I526544,I526561,I694427,I526578,I694418,I526595,I694439,I526612,I526629,I526479,I526660,I526677,I526482,I526708,I526725,I694442,I526742,I526458,I526773,I526470,I526813,I526821,I526838,I526855,I694421,I526872,I526485,I526903,I694424,I526920,I694445,I526937,I694436,I526963,I526473,I526985,I527002,I526467,I527033,I526461,I526464,I527078,I526476,I527139,I527165,I527182,I527190,I527207,I527224,I527241,I527258,I527275,I527125,I527306,I527323,I527128,I527354,I527371,I527388,I527104,I527419,I527116,I527459,I527467,I527484,I527501,I527518,I527131,I527549,I527566,I527583,I527609,I527119,I527631,I527648,I527113,I527679,I527107,I527110,I527724,I527122,I527785,I527811,I527828,I527836,I527853,I527870,I527887,I527904,I527921,I527952,I527969,I528000,I528017,I528034,I528065,I528105,I528113,I528130,I528147,I528164,I528195,I528212,I528229,I528255,I528277,I528294,I528325,I528370,I528431,I528457,I528474,I528482,I528499,I528516,I528533,I528550,I528567,I528417,I528598,I528615,I528420,I528646,I528663,I528680,I528396,I528711,I528408,I528751,I528759,I528776,I528793,I528810,I528423,I528841,I528858,I528875,I528901,I528411,I528923,I528940,I528405,I528971,I528399,I528402,I529016,I528414,I529077,I529103,I529120,I529128,I529145,I529162,I529179,I529196,I529213,I529063,I529244,I529261,I529066,I529292,I529309,I529326,I529042,I529357,I529054,I529397,I529405,I529422,I529439,I529456,I529069,I529487,I529504,I529521,I529547,I529057,I529569,I529586,I529051,I529617,I529045,I529048,I529662,I529060,I529723,I529749,I529766,I529774,I529791,I529808,I529825,I529842,I529859,I529890,I529907,I529938,I529955,I529972,I530003,I530043,I530051,I530068,I530085,I530102,I530133,I530150,I530167,I530193,I530215,I530232,I530263,I530308,I530369,I606988,I530395,I606970,I530412,I530420,I530437,I606979,I530454,I606991,I530471,I606973,I530488,I606982,I530505,I530536,I530553,I530584,I530601,I606994,I530618,I530649,I530689,I530697,I530714,I530731,I530748,I530779,I606976,I530796,I606985,I530813,I530839,I530861,I530878,I530909,I530954,I531015,I531041,I531058,I531066,I531083,I531100,I531117,I531134,I531151,I531182,I531199,I531230,I531247,I531264,I531295,I531335,I531343,I531360,I531377,I531394,I531425,I531442,I531459,I531485,I531507,I531524,I531555,I531600,I531661,I531687,I531704,I531712,I531729,I531746,I531763,I531780,I531797,I531828,I531845,I531876,I531893,I531910,I531941,I531981,I531989,I532006,I532023,I532040,I532071,I532088,I532105,I532131,I532153,I532170,I532201,I532246,I532307,I532333,I532350,I532358,I532375,I532392,I532409,I532426,I532443,I532474,I532491,I532522,I532539,I532556,I532587,I532627,I532635,I532652,I532669,I532686,I532717,I532734,I532751,I532777,I532799,I532816,I532847,I532892,I532953,I532979,I532996,I533004,I533021,I533038,I533055,I533072,I533089,I533120,I533137,I533168,I533185,I533202,I533233,I533273,I533281,I533298,I533315,I533332,I533363,I533380,I533397,I533423,I533445,I533462,I533493,I533538,I533599,I533625,I533642,I533650,I533667,I533684,I533701,I533718,I533735,I533766,I533783,I533814,I533831,I533848,I533879,I533919,I533927,I533944,I533961,I533978,I534009,I534026,I534043,I534069,I534091,I534108,I534139,I534184,I534245,I534271,I534288,I534296,I534313,I534330,I534347,I534364,I534381,I534231,I534412,I534429,I534234,I534460,I534477,I534494,I534210,I534525,I534222,I534565,I534573,I534590,I534607,I534624,I534237,I534655,I534672,I534689,I534715,I534225,I534737,I534754,I534219,I534785,I534213,I534216,I534830,I534228,I534891,I642246,I534917,I642228,I534934,I534942,I534959,I642237,I534976,I642249,I534993,I642231,I535010,I642240,I535027,I535058,I535075,I535106,I535123,I642252,I535140,I535171,I535211,I535219,I535236,I535253,I535270,I535301,I642234,I535318,I642243,I535335,I535361,I535383,I535400,I535431,I535476,I535537,I535563,I535580,I535588,I535605,I535622,I535639,I535656,I535673,I535523,I535704,I535721,I535526,I535752,I535769,I535786,I535502,I535817,I535514,I535857,I535865,I535882,I535899,I535916,I535529,I535947,I535964,I535981,I536007,I535517,I536029,I536046,I535511,I536077,I535505,I535508,I536122,I535520,I536183,I536209,I536226,I536234,I536251,I536268,I536285,I536302,I536319,I536350,I536367,I536398,I536415,I536432,I536463,I536503,I536511,I536528,I536545,I536562,I536593,I536610,I536627,I536653,I536675,I536692,I536723,I536768,I536829,I536855,I536872,I536880,I536897,I536914,I536931,I536948,I536965,I536996,I537013,I537044,I537061,I537078,I537109,I537149,I537157,I537174,I537191,I537208,I537239,I537256,I537273,I537299,I537321,I537338,I537369,I537414,I537475,I663768,I537501,I663774,I537518,I537526,I537543,I663771,I537560,I663750,I537577,I663753,I537594,I663759,I537611,I537461,I537642,I537659,I537464,I537690,I537707,I537724,I537440,I537755,I537452,I537795,I537803,I537820,I537837,I663762,I537854,I537467,I537885,I537902,I663756,I537919,I663765,I537945,I537455,I537967,I537984,I537449,I538015,I537443,I537446,I538060,I537458,I538121,I538147,I538164,I538172,I538189,I538206,I538223,I538240,I538257,I538107,I538288,I538305,I538110,I538336,I538353,I538370,I538086,I538401,I538098,I538441,I538449,I538466,I538483,I538500,I538113,I538531,I538548,I538565,I538591,I538101,I538613,I538630,I538095,I538661,I538089,I538092,I538706,I538104,I538767,I643980,I538793,I643962,I538810,I538818,I538835,I643971,I538852,I643983,I538869,I643965,I538886,I643974,I538903,I538934,I538951,I538982,I538999,I643986,I539016,I539047,I539087,I539095,I539112,I539129,I539146,I539177,I643968,I539194,I643977,I539211,I539237,I539259,I539276,I539307,I539352,I539413,I687525,I539439,I687519,I539456,I539464,I539481,I687528,I539498,I687540,I539515,I687522,I539532,I539549,I539580,I539597,I539628,I539645,I687516,I539662,I539693,I539733,I539741,I539758,I539775,I687537,I539792,I539823,I687531,I539840,I539857,I687534,I539883,I539905,I539922,I539953,I539998,I540059,I540085,I540102,I540110,I540127,I540144,I540161,I540178,I540195,I540045,I540226,I540243,I540048,I540274,I540291,I540308,I540024,I540339,I540036,I540379,I540387,I540404,I540421,I540438,I540051,I540469,I540486,I540503,I540529,I540039,I540551,I540568,I540033,I540599,I540027,I540030,I540644,I540042,I540705,I540731,I540748,I540756,I540773,I540790,I540807,I540824,I540841,I540872,I540889,I540920,I540937,I540954,I540985,I541025,I541033,I541050,I541067,I541084,I541115,I541132,I541149,I541175,I541197,I541214,I541245,I541290,I541351,I541377,I541394,I541402,I541419,I541436,I541453,I541470,I541487,I541337,I541518,I541535,I541340,I541566,I541583,I541600,I541316,I541631,I541328,I541671,I541679,I541696,I541713,I541730,I541343,I541761,I541778,I541795,I541821,I541331,I541843,I541860,I541325,I541891,I541319,I541322,I541936,I541334,I541997,I542023,I542040,I542048,I542065,I542082,I542099,I542116,I542133,I542164,I542181,I542212,I542229,I542246,I542277,I542317,I542325,I542342,I542359,I542376,I542407,I542424,I542441,I542467,I542489,I542506,I542537,I542582,I542643,I566119,I542669,I566122,I542686,I542694,I542711,I542728,I566131,I542745,I566140,I542762,I566128,I542779,I542810,I542827,I542858,I542875,I566134,I542892,I542923,I542963,I542971,I542988,I543005,I566125,I543022,I543053,I566137,I543070,I543087,I543113,I543135,I543152,I543183,I543228,I543289,I543315,I543332,I543340,I543357,I543374,I543391,I543408,I543425,I543456,I543473,I543504,I543521,I543538,I543569,I543609,I543617,I543634,I543651,I543668,I543699,I543716,I543733,I543759,I543781,I543798,I543829,I543874,I543935,I660504,I543961,I660510,I543978,I543986,I544003,I660507,I544020,I660486,I544037,I660489,I544054,I660495,I544071,I544102,I544119,I544150,I544167,I544184,I544215,I544255,I544263,I544280,I544297,I660498,I544314,I544345,I544362,I660492,I544379,I660501,I544405,I544427,I544444,I544475,I544520,I544581,I663224,I544607,I663230,I544624,I544632,I544649,I663227,I544666,I663206,I544683,I663209,I544700,I663215,I544717,I544748,I544765,I544796,I544813,I544830,I544861,I544901,I544909,I544926,I544943,I663218,I544960,I544991,I545008,I663212,I545025,I663221,I545051,I545073,I545090,I545121,I545166,I545227,I679433,I545253,I679427,I545270,I545278,I545295,I679436,I545312,I679448,I545329,I679430,I545346,I545363,I545213,I545394,I545411,I545216,I545442,I545459,I679424,I545476,I545192,I545507,I545204,I545547,I545555,I545572,I545589,I679445,I545606,I545219,I545637,I679439,I545654,I545671,I679442,I545697,I545207,I545719,I545736,I545201,I545767,I545195,I545198,I545812,I545210,I545873,I545899,I545916,I545924,I545941,I545958,I545975,I545992,I546009,I546040,I546057,I546088,I546105,I546122,I546153,I546193,I546201,I546218,I546235,I546252,I546283,I546300,I546317,I546343,I546365,I546382,I546413,I546458,I546513,I546539,I546556,I546578,I546604,I546612,I546629,I546646,I546663,I546680,I546697,I546714,I546745,I546776,I546793,I546810,I546827,I546858,I546903,I546920,I546937,I546963,I546971,I547002,I547019,I547074,I547100,I547117,I547139,I547165,I547173,I547190,I547207,I547224,I547241,I547258,I547275,I547306,I547337,I547354,I547371,I547388,I547419,I547464,I547481,I547498,I547524,I547532,I547563,I547580,I547635,I547661,I547678,I547700,I547726,I547734,I547751,I547768,I547785,I547802,I547819,I547836,I547867,I547898,I547915,I547932,I547949,I547980,I548025,I548042,I548059,I548085,I548093,I548124,I548141,I548196,I548222,I548239,I548261,I548287,I548295,I548312,I548329,I548346,I548363,I548380,I548397,I548428,I548459,I548476,I548493,I548510,I548541,I548586,I548603,I548620,I548646,I548654,I548685,I548702,I548757,I548783,I548800,I548822,I548848,I548856,I548873,I548890,I548907,I548924,I548941,I548958,I548989,I549020,I549037,I549054,I549071,I549102,I549147,I549164,I549181,I549207,I549215,I549246,I549263,I549318,I549344,I549361,I549310,I549383,I549409,I549417,I549434,I549451,I549468,I549485,I549502,I549519,I549292,I549550,I549295,I549581,I549598,I549615,I549632,I549304,I549663,I549307,I549301,I549708,I549725,I549742,I549768,I549776,I549289,I549807,I549824,I549298,I549879,I549905,I549922,I549944,I549970,I549978,I549995,I550012,I550029,I550046,I550063,I550080,I550111,I550142,I550159,I550176,I550193,I550224,I550269,I550286,I550303,I550329,I550337,I550368,I550385,I550440,I550466,I550483,I550505,I550531,I550539,I550556,I550573,I550590,I550607,I550624,I550641,I550672,I550703,I550720,I550737,I550754,I550785,I550830,I550847,I550864,I550890,I550898,I550929,I550946,I551001,I667020,I551027,I551044,I551066,I667026,I551092,I551100,I667035,I551117,I551134,I667014,I551151,I667017,I551168,I551185,I667029,I551202,I551233,I551264,I667023,I551281,I551298,I551315,I551346,I551391,I667038,I551408,I551425,I667032,I551451,I551459,I551490,I551507,I551562,I551588,I551605,I551627,I551653,I551661,I551678,I551695,I551712,I551729,I551746,I551763,I551794,I551825,I551842,I551859,I551876,I551907,I551952,I551969,I551986,I552012,I552020,I552051,I552068,I552123,I552149,I552166,I552188,I552214,I552222,I552239,I552256,I552273,I552290,I552307,I552324,I552355,I552386,I552403,I552420,I552437,I552468,I552513,I552530,I552547,I552573,I552581,I552612,I552629,I552684,I612765,I552710,I552727,I552749,I612756,I552775,I552783,I612753,I552800,I552817,I612762,I552834,I612771,I552851,I552868,I612750,I552885,I552916,I552947,I612759,I552964,I552981,I552998,I553029,I553074,I612774,I553091,I553108,I612768,I553134,I553142,I553173,I553190,I553245,I553271,I553288,I553237,I553310,I553336,I553344,I553361,I553378,I553395,I553412,I553429,I553446,I553219,I553477,I553222,I553508,I553525,I553542,I553559,I553231,I553590,I553234,I553228,I553635,I553652,I553669,I553695,I553703,I553216,I553734,I553751,I553225,I553806,I553832,I553849,I553871,I553897,I553905,I553922,I553939,I553956,I553973,I553990,I554007,I554038,I554069,I554086,I554103,I554120,I554151,I554196,I554213,I554230,I554256,I554264,I554295,I554312,I554367,I714493,I554393,I554410,I554432,I714487,I554458,I554466,I714478,I554483,I554500,I714505,I554517,I714490,I714499,I554534,I554551,I714484,I554568,I554599,I554630,I714502,I554647,I554664,I554681,I554712,I554757,I714496,I554774,I554791,I714481,I554817,I554825,I554856,I554873,I554928,I554954,I554971,I554993,I555019,I555027,I555044,I555061,I555078,I555095,I555112,I555129,I555160,I555191,I555208,I555225,I555242,I555273,I555318,I555335,I555352,I555378,I555386,I555417,I555434,I555489,I555515,I555532,I555554,I555580,I555588,I555605,I555622,I555639,I555656,I555673,I555690,I555721,I555752,I555769,I555786,I555803,I555834,I555879,I555896,I555913,I555939,I555947,I555978,I555995,I556050,I645711,I556076,I556093,I556115,I645702,I556141,I556149,I645699,I556166,I556183,I645708,I556200,I645717,I556217,I556234,I645696,I556251,I556282,I556313,I645705,I556330,I556347,I556364,I556395,I556440,I645720,I556457,I556474,I645714,I556500,I556508,I556539,I556556,I556611,I556637,I556654,I556603,I556676,I556702,I556710,I556727,I556744,I556761,I556778,I556795,I556812,I556585,I556843,I556588,I556874,I556891,I556908,I556925,I556597,I556956,I556600,I556594,I557001,I557018,I557035,I557061,I557069,I556582,I557100,I557117,I556591,I557172,I557198,I557215,I557237,I557263,I557271,I557288,I557305,I557322,I557339,I557356,I557373,I557404,I557435,I557452,I557469,I557486,I557517,I557562,I557579,I557596,I557622,I557630,I557661,I557678,I557733,I625481,I557759,I557776,I557798,I625472,I557824,I557832,I625469,I557849,I557866,I625478,I557883,I625487,I557900,I557917,I625466,I557934,I557965,I557996,I625475,I558013,I558030,I558047,I558078,I558123,I625490,I558140,I558157,I625484,I558183,I558191,I558222,I558239,I558294,I558320,I558337,I558286,I558359,I558385,I558393,I558410,I558427,I558444,I558461,I558478,I558495,I558268,I558526,I558271,I558557,I558574,I558591,I558608,I558280,I558639,I558283,I558277,I558684,I558701,I558718,I558744,I558752,I558265,I558783,I558800,I558274,I558855,I637619,I558881,I558898,I558920,I637610,I558946,I558954,I637607,I558971,I558988,I637616,I559005,I637625,I559022,I559039,I637604,I559056,I559087,I559118,I637613,I559135,I559152,I559169,I559200,I559245,I637628,I559262,I559279,I637622,I559305,I559313,I559344,I559361,I559416,I559442,I559459,I559408,I559481,I559507,I559515,I559532,I559549,I559566,I559583,I559600,I559617,I559390,I559648,I559393,I559679,I559696,I559713,I559730,I559402,I559761,I559405,I559399,I559806,I559823,I559840,I559866,I559874,I559387,I559905,I559922,I559396,I559977,I718063,I560003,I560020,I560042,I718057,I560068,I560076,I718048,I560093,I560110,I718075,I560127,I718060,I718069,I560144,I560161,I718054,I560178,I560209,I560240,I718072,I560257,I560274,I560291,I560322,I560367,I718066,I560384,I560401,I718051,I560427,I560435,I560466,I560483,I560538,I560564,I560581,I560603,I560629,I560637,I560654,I560671,I560688,I560705,I560722,I560739,I560770,I560801,I560818,I560835,I560852,I560883,I560928,I560945,I560962,I560988,I560996,I561027,I561044,I561099,I561125,I561142,I561164,I561190,I561198,I561215,I561232,I561249,I561266,I561283,I561300,I561331,I561362,I561379,I561396,I561413,I561444,I561489,I561506,I561523,I561549,I561557,I561588,I561605,I561660,I561686,I561703,I561725,I561751,I561759,I561776,I561793,I561810,I561827,I561844,I561861,I561892,I561923,I561940,I561957,I561974,I562005,I562050,I562067,I562084,I562110,I562118,I562149,I562166,I562221,I562247,I562264,I562213,I562286,I562312,I562320,I562337,I562354,I562371,I562388,I562405,I562422,I562195,I562453,I562198,I562484,I562501,I562518,I562535,I562207,I562566,I562210,I562204,I562611,I562628,I562645,I562671,I562679,I562192,I562710,I562727,I562201,I562782,I562808,I562825,I562847,I562873,I562881,I562898,I562915,I562932,I562949,I562966,I562983,I563014,I563045,I563062,I563079,I563096,I563127,I563172,I563189,I563206,I563232,I563240,I563271,I563288,I563343,I563369,I563386,I563408,I563434,I563442,I563459,I563476,I563493,I563510,I563527,I563544,I563575,I563606,I563623,I563640,I563657,I563688,I563733,I563750,I563767,I563793,I563801,I563832,I563849,I563904,I563930,I563947,I563969,I563995,I564003,I564020,I564037,I564054,I564071,I564088,I564105,I564136,I564167,I564184,I564201,I564218,I564249,I564294,I564311,I564328,I564354,I564362,I564393,I564410,I564465,I564491,I564508,I564530,I564556,I564564,I564581,I564598,I564615,I564632,I564649,I564666,I564697,I564728,I564745,I564762,I564779,I564810,I564855,I564872,I564889,I564915,I564923,I564954,I564971,I565026,I702593,I565052,I565069,I565018,I565091,I702587,I565117,I565125,I702578,I565142,I565159,I702605,I565176,I702590,I702599,I565193,I565210,I702584,I565227,I565000,I565258,I565003,I565289,I702602,I565306,I565323,I565340,I565012,I565371,I565015,I565009,I565416,I702596,I565433,I565450,I702581,I565476,I565484,I564997,I565515,I565532,I565006,I565587,I642821,I565613,I565630,I565579,I565652,I642812,I565678,I565686,I642809,I565703,I565720,I642818,I565737,I642827,I565754,I565771,I642806,I565788,I565561,I565819,I565564,I565850,I642815,I565867,I565884,I565901,I565573,I565932,I565576,I565570,I565977,I642830,I565994,I566011,I642824,I566037,I566045,I565558,I566076,I566093,I565567,I566148,I566174,I566191,I566213,I566239,I566247,I566264,I566281,I566298,I566315,I566332,I566349,I566380,I566411,I566428,I566445,I566462,I566493,I566538,I566555,I566572,I566598,I566606,I566637,I566654,I566709,I566735,I566752,I566774,I566800,I566808,I566825,I566842,I566859,I566876,I566893,I566910,I566941,I566972,I566989,I567006,I567023,I567054,I567099,I567116,I567133,I567159,I567167,I567198,I567215,I567270,I567296,I567313,I567335,I567361,I567369,I567386,I567403,I567420,I567437,I567454,I567471,I567502,I567533,I567550,I567567,I567584,I567615,I567660,I567677,I567694,I567720,I567728,I567759,I567776,I567831,I567857,I567874,I567896,I567922,I567930,I567947,I567964,I567981,I567998,I568015,I568032,I568063,I568094,I568111,I568128,I568145,I568176,I568221,I568238,I568255,I568281,I568289,I568320,I568337,I568392,I692143,I568418,I568435,I568457,I692140,I568483,I568491,I692146,I568508,I568525,I692155,I568542,I692149,I568559,I568576,I692161,I568593,I568624,I568655,I692158,I568672,I568689,I568706,I568737,I568782,I692152,I568799,I692164,I568816,I568842,I568850,I568881,I568898,I568953,I568979,I568996,I569018,I569044,I569052,I569069,I569086,I569103,I569120,I569137,I569154,I569185,I569216,I569233,I569250,I569267,I569298,I569343,I569360,I569377,I569403,I569411,I569442,I569459,I569514,I569540,I569557,I569579,I569605,I569613,I569630,I569647,I569664,I569681,I569698,I569715,I569746,I569777,I569794,I569811,I569828,I569859,I569904,I569921,I569938,I569964,I569972,I570003,I570020,I570075,I570101,I570118,I570140,I570166,I570174,I570191,I570208,I570225,I570242,I570259,I570276,I570307,I570338,I570355,I570372,I570389,I570420,I570465,I570482,I570499,I570525,I570533,I570564,I570581,I570636,I570662,I570679,I570628,I570701,I570727,I570735,I570752,I570769,I570786,I570803,I570820,I570837,I570610,I570868,I570613,I570899,I570916,I570933,I570950,I570622,I570981,I570625,I570619,I571026,I571043,I571060,I571086,I571094,I570607,I571125,I571142,I570616,I571197,I571223,I571240,I571189,I571262,I571288,I571296,I571313,I571330,I571347,I571364,I571381,I571398,I571171,I571429,I571174,I571460,I571477,I571494,I571511,I571183,I571542,I571186,I571180,I571587,I571604,I571621,I571647,I571655,I571168,I571686,I571703,I571177,I571758,I571784,I571801,I571823,I571849,I571857,I571874,I571891,I571908,I571925,I571942,I571959,I571990,I572021,I572038,I572055,I572072,I572103,I572148,I572165,I572182,I572208,I572216,I572247,I572264,I572322,I729380,I572348,I572356,I729362,I729353,I572396,I572404,I729368,I572421,I729356,I572438,I572478,I572500,I729365,I572517,I572543,I572551,I572568,I729374,I572585,I572602,I572619,I572664,I729377,I572695,I572712,I729371,I729359,I572738,I572746,I572777,I572794,I572811,I572828,I572900,I572926,I572934,I572974,I572982,I572999,I573016,I573056,I573078,I573095,I573121,I573129,I573146,I573163,I573180,I573197,I573242,I573273,I573290,I573316,I573324,I573355,I573372,I573389,I573406,I573478,I573504,I573512,I573552,I573560,I573577,I573594,I573634,I573656,I573673,I573699,I573707,I573724,I573741,I573758,I573775,I573820,I573851,I573868,I573894,I573902,I573933,I573950,I573967,I573984,I574056,I574082,I574090,I574039,I574130,I574138,I574155,I574172,I574027,I574212,I574048,I574234,I574251,I574277,I574285,I574302,I574319,I574336,I574353,I574024,I574045,I574398,I574036,I574429,I574446,I574472,I574480,I574042,I574511,I574528,I574545,I574562,I574033,I574030,I574634,I671387,I574660,I574668,I671381,I671366,I574708,I574716,I671372,I574733,I671384,I574750,I574790,I574812,I574829,I574855,I574863,I574880,I671390,I574897,I671378,I574914,I574931,I574976,I671369,I575007,I575024,I671375,I575050,I575058,I575089,I575106,I575123,I575140,I575212,I575238,I575246,I575286,I575294,I575311,I575328,I575368,I575390,I575407,I575433,I575441,I575458,I575475,I575492,I575509,I575554,I575585,I575602,I575628,I575636,I575667,I575684,I575701,I575718,I575790,I575816,I575824,I575864,I575872,I575889,I575906,I575946,I575968,I575985,I576011,I576019,I576036,I576053,I576070,I576087,I576132,I576163,I576180,I576206,I576214,I576245,I576262,I576279,I576296,I576368,I684650,I576394,I576402,I684632,I684641,I576442,I576450,I684626,I576467,I684638,I576484,I576524,I576546,I684629,I576563,I576589,I576597,I576614,I576631,I576648,I576665,I576710,I684647,I576741,I576758,I684635,I684644,I576784,I576792,I576823,I576840,I576857,I576874,I576946,I576972,I576980,I577020,I577028,I577045,I577062,I577102,I577124,I577141,I577167,I577175,I577192,I577209,I577226,I577243,I577288,I577319,I577336,I577362,I577370,I577401,I577418,I577435,I577452,I577524,I577550,I577558,I577598,I577606,I577623,I577640,I577680,I577702,I577719,I577745,I577753,I577770,I577787,I577804,I577821,I577866,I577897,I577914,I577940,I577948,I577979,I577996,I578013,I578030,I578102,I578128,I578136,I578085,I578176,I578184,I578201,I578218,I578073,I578258,I578094,I578280,I578297,I578323,I578331,I578348,I578365,I578382,I578399,I578070,I578091,I578444,I578082,I578475,I578492,I578518,I578526,I578088,I578557,I578574,I578591,I578608,I578079,I578076,I578680,I578706,I578714,I578754,I578762,I578779,I578796,I578836,I578858,I578875,I578901,I578909,I578926,I578943,I578960,I578977,I579022,I579053,I579070,I579096,I579104,I579135,I579152,I579169,I579186,I579258,I579284,I579292,I579332,I579340,I579357,I579374,I579414,I579436,I579453,I579479,I579487,I579504,I579521,I579538,I579555,I579600,I579631,I579648,I579674,I579682,I579713,I579730,I579747,I579764,I579836,I579862,I579870,I579819,I579910,I579918,I579935,I579952,I579807,I579992,I579828,I580014,I580031,I580057,I580065,I580082,I580099,I580116,I580133,I579804,I579825,I580178,I579816,I580209,I580226,I580252,I580260,I579822,I580291,I580308,I580325,I580342,I579813,I579810,I580414,I580440,I580448,I580488,I580496,I580513,I580530,I580570,I580592,I580609,I580635,I580643,I580660,I580677,I580694,I580711,I580756,I580787,I580804,I580830,I580838,I580869,I580886,I580903,I580920,I580992,I581018,I581026,I580975,I581066,I581074,I581091,I581108,I580963,I581148,I580984,I581170,I581187,I581213,I581221,I581238,I581255,I581272,I581289,I580960,I580981,I581334,I580972,I581365,I581382,I581408,I581416,I580978,I581447,I581464,I581481,I581498,I580969,I580966,I581570,I581596,I581604,I581553,I581644,I581652,I581669,I581686,I581541,I581726,I581562,I581748,I581765,I581791,I581799,I581816,I581833,I581850,I581867,I581538,I581559,I581912,I581550,I581943,I581960,I581986,I581994,I581556,I582025,I582042,I582059,I582076,I581547,I581544,I582148,I582174,I582182,I582222,I582230,I582247,I582264,I582304,I582326,I582343,I582369,I582377,I582394,I582411,I582428,I582445,I582490,I582521,I582538,I582564,I582572,I582603,I582620,I582637,I582654,I582726,I582752,I582760,I582800,I582808,I582825,I582842,I582882,I582904,I582921,I582947,I582955,I582972,I582989,I583006,I583023,I583068,I583099,I583116,I583142,I583150,I583181,I583198,I583215,I583232,I583304,I675402,I583330,I583338,I675384,I675393,I583378,I583386,I675378,I583403,I675390,I583420,I583460,I583482,I675381,I583499,I583525,I583533,I583550,I583567,I583584,I583601,I583646,I675399,I583677,I583694,I675387,I675396,I583720,I583728,I583759,I583776,I583793,I583810,I583882,I738305,I583908,I583916,I738287,I738278,I583956,I583964,I738293,I583981,I738281,I583998,I584038,I584060,I738290,I584077,I584103,I584111,I584128,I738299,I584145,I584162,I584179,I584224,I738302,I584255,I584272,I738296,I738284,I584298,I584306,I584337,I584354,I584371,I584388,I584460,I584486,I584494,I584534,I584542,I584559,I584576,I584616,I584638,I584655,I584681,I584689,I584706,I584723,I584740,I584757,I584802,I584833,I584850,I584876,I584884,I584915,I584932,I584949,I584966,I585038,I661595,I585064,I585072,I661589,I661574,I585112,I585120,I661580,I585137,I661592,I585154,I585194,I585216,I585233,I585259,I585267,I585284,I661598,I585301,I661586,I585318,I585335,I585380,I661577,I585411,I585428,I661583,I585454,I585462,I585493,I585510,I585527,I585544,I585616,I585642,I585650,I585690,I585698,I585715,I585732,I585772,I585794,I585811,I585837,I585845,I585862,I585879,I585896,I585913,I585958,I585989,I586006,I586032,I586040,I586071,I586088,I586105,I586122,I586194,I586220,I586228,I586268,I586276,I586293,I586310,I586350,I586372,I586389,I586415,I586423,I586440,I586457,I586474,I586491,I586536,I586567,I586584,I586610,I586618,I586649,I586666,I586683,I586700,I586772,I586798,I586806,I586846,I586854,I586871,I586888,I586928,I586950,I586967,I586993,I587001,I587018,I587035,I587052,I587069,I587114,I587145,I587162,I587188,I587196,I587227,I587244,I587261,I587278,I587350,I699035,I587376,I587384,I699017,I699008,I587424,I587432,I699023,I587449,I699011,I587466,I587506,I587528,I699020,I587545,I587571,I587579,I587596,I699029,I587613,I587630,I587647,I587692,I699032,I587723,I587740,I699026,I699014,I587766,I587774,I587805,I587822,I587839,I587856,I587928,I651259,I587954,I587962,I651253,I651238,I588002,I588010,I651244,I588027,I651256,I588044,I588084,I588106,I588123,I588149,I588157,I588174,I651262,I588191,I651250,I588208,I588225,I588270,I651241,I588301,I588318,I651247,I588344,I588352,I588383,I588400,I588417,I588434,I588506,I588532,I588540,I588489,I588580,I588588,I588605,I588622,I588477,I588662,I588498,I588684,I588701,I588727,I588735,I588752,I588769,I588786,I588803,I588474,I588495,I588848,I588486,I588879,I588896,I588922,I588930,I588492,I588961,I588978,I588995,I589012,I588483,I588480,I589084,I589110,I589118,I589158,I589166,I589183,I589200,I589240,I589262,I589279,I589305,I589313,I589330,I589347,I589364,I589381,I589426,I589457,I589474,I589500,I589508,I589539,I589556,I589573,I589590,I589662,I589688,I589696,I589736,I589744,I589761,I589778,I589818,I589840,I589857,I589883,I589891,I589908,I589925,I589942,I589959,I590004,I590035,I590052,I590078,I590086,I590117,I590134,I590151,I590168,I590240,I590266,I590274,I590314,I590322,I590339,I590356,I590396,I590418,I590435,I590461,I590469,I590486,I590503,I590520,I590537,I590582,I590613,I590630,I590656,I590664,I590695,I590712,I590729,I590746,I590818,I590844,I590852,I590892,I590900,I590917,I590934,I590974,I590996,I591013,I591039,I591047,I591064,I591081,I591098,I591115,I591160,I591191,I591208,I591234,I591242,I591273,I591290,I591307,I591324,I591396,I591422,I591430,I591379,I591470,I591478,I591495,I591512,I591367,I591552,I591388,I591574,I591591,I591617,I591625,I591642,I591659,I591676,I591693,I591364,I591385,I591738,I591376,I591769,I591786,I591812,I591820,I591382,I591851,I591868,I591885,I591902,I591373,I591370,I591974,I592000,I592008,I591957,I592048,I592056,I592073,I592090,I591945,I592130,I591966,I592152,I592169,I592195,I592203,I592220,I592237,I592254,I592271,I591942,I591963,I592316,I591954,I592347,I592364,I592390,I592398,I591960,I592429,I592446,I592463,I592480,I591951,I591948,I592552,I592578,I592586,I592626,I592634,I592651,I592668,I592708,I592730,I592747,I592773,I592781,I592798,I592815,I592832,I592849,I592894,I592925,I592942,I592968,I592976,I593007,I593024,I593041,I593058,I593130,I593156,I593164,I593204,I593212,I593229,I593246,I593286,I593308,I593325,I593351,I593359,I593376,I593393,I593410,I593427,I593472,I593503,I593520,I593546,I593554,I593585,I593602,I593619,I593636,I593708,I593734,I593742,I593782,I593790,I593807,I593824,I593864,I593886,I593903,I593929,I593937,I593954,I593971,I593988,I594005,I594050,I594081,I594098,I594124,I594132,I594163,I594180,I594197,I594214,I594286,I594312,I594320,I594360,I594368,I594385,I594402,I594442,I594464,I594481,I594507,I594515,I594532,I594549,I594566,I594583,I594628,I594659,I594676,I594702,I594710,I594741,I594758,I594775,I594792,I594864,I594890,I594898,I594847,I594938,I594946,I594963,I594980,I594835,I595020,I594856,I595042,I595059,I595085,I595093,I595110,I595127,I595144,I595161,I594832,I594853,I595206,I594844,I595237,I595254,I595280,I595288,I594850,I595319,I595336,I595353,I595370,I594841,I594838,I595442,I595468,I595476,I595516,I595524,I595541,I595558,I595598,I595620,I595637,I595663,I595671,I595688,I595705,I595722,I595739,I595784,I595815,I595832,I595858,I595866,I595897,I595914,I595931,I595948,I596020,I596046,I596054,I596094,I596102,I596119,I596136,I596176,I596198,I596215,I596241,I596249,I596266,I596283,I596300,I596317,I596362,I596393,I596410,I596436,I596444,I596475,I596492,I596509,I596526,I596598,I724025,I596624,I596632,I724007,I723998,I596672,I596680,I724013,I596697,I724001,I596714,I596754,I596776,I724010,I596793,I596819,I596827,I596844,I724019,I596861,I596878,I596895,I596940,I724022,I596971,I596988,I724016,I724004,I597014,I597022,I597053,I597070,I597087,I597104,I597176,I597202,I597210,I597250,I597258,I597275,I597292,I597332,I597354,I597371,I597397,I597405,I597422,I597439,I597456,I597473,I597518,I597549,I597566,I597592,I597600,I597631,I597648,I597665,I597682,I597754,I597780,I597788,I597828,I597836,I597853,I597870,I597910,I597932,I597949,I597975,I597983,I598000,I598017,I598034,I598051,I598096,I598127,I598144,I598170,I598178,I598209,I598226,I598243,I598260,I598332,I598358,I598366,I598406,I598414,I598431,I598448,I598488,I598510,I598527,I598553,I598561,I598578,I598595,I598612,I598629,I598674,I598705,I598722,I598748,I598756,I598787,I598804,I598821,I598838,I598910,I598936,I598944,I598893,I598984,I598992,I599009,I599026,I598881,I599066,I598902,I599088,I599105,I599131,I599139,I599156,I599173,I599190,I599207,I598878,I598899,I599252,I598890,I599283,I599300,I599326,I599334,I598896,I599365,I599382,I599399,I599416,I598887,I598884,I599488,I741280,I599514,I599522,I741262,I599471,I741253,I599562,I599570,I741268,I599587,I741256,I599604,I599459,I599644,I599480,I599666,I741265,I599683,I599709,I599717,I599734,I741274,I599751,I599768,I599785,I599456,I599477,I599830,I741277,I599468,I599861,I599878,I741271,I741259,I599904,I599912,I599474,I599943,I599960,I599977,I599994,I599465,I599462,I600066,I600092,I600100,I600049,I600140,I600148,I600165,I600182,I600037,I600222,I600058,I600244,I600261,I600287,I600295,I600312,I600329,I600346,I600363,I600034,I600055,I600408,I600046,I600439,I600456,I600482,I600490,I600052,I600521,I600538,I600555,I600572,I600043,I600040,I600644,I600670,I600678,I600718,I600726,I600743,I600760,I600800,I600822,I600839,I600865,I600873,I600890,I600907,I600924,I600941,I600986,I601017,I601034,I601060,I601068,I601099,I601116,I601133,I601150,I601222,I601248,I601256,I601296,I601304,I601321,I601338,I601378,I601400,I601417,I601443,I601451,I601468,I601485,I601502,I601519,I601564,I601595,I601612,I601638,I601646,I601677,I601694,I601711,I601728,I601800,I601826,I601834,I601874,I601882,I601899,I601916,I601956,I601978,I601995,I602021,I602029,I602046,I602063,I602080,I602097,I602142,I602173,I602190,I602216,I602224,I602255,I602272,I602289,I602306,I602378,I602404,I602412,I602452,I602460,I602477,I602494,I602534,I602556,I602573,I602599,I602607,I602624,I602641,I602658,I602675,I602720,I602751,I602768,I602794,I602802,I602833,I602850,I602867,I602884,I602956,I602982,I602990,I602939,I603030,I603038,I603055,I603072,I602927,I603112,I602948,I603134,I603151,I603177,I603185,I603202,I603219,I603236,I603253,I602924,I602945,I603298,I602936,I603329,I603346,I603372,I603380,I602942,I603411,I603428,I603445,I603462,I602933,I602930,I603534,I603560,I603568,I603517,I603608,I603616,I603633,I603650,I603505,I603690,I603526,I603712,I603729,I603755,I603763,I603780,I603797,I603814,I603831,I603502,I603523,I603876,I603514,I603907,I603924,I603950,I603958,I603520,I603989,I604006,I604023,I604040,I603511,I603508,I604112,I604138,I604146,I604186,I604194,I604211,I604228,I604268,I604290,I604307,I604333,I604341,I604358,I604375,I604392,I604409,I604454,I604485,I604502,I604528,I604536,I604567,I604584,I604601,I604618,I604690,I604716,I604724,I604673,I604764,I604772,I604789,I604806,I604661,I604846,I604682,I604868,I604885,I604911,I604919,I604936,I604953,I604970,I604987,I604658,I604679,I605032,I604670,I605063,I605080,I605106,I605114,I604676,I605145,I605162,I605179,I605196,I604667,I604664,I605268,I605294,I605302,I605342,I605350,I605367,I605384,I605424,I605446,I605463,I605489,I605497,I605514,I605531,I605548,I605565,I605610,I605641,I605658,I605684,I605692,I605723,I605740,I605757,I605774,I605846,I605872,I605880,I605920,I605928,I605945,I605962,I606002,I606024,I606041,I606067,I606075,I606092,I606109,I606126,I606143,I606188,I606219,I606236,I606262,I606270,I606301,I606318,I606335,I606352,I606424,I606450,I606458,I606498,I606506,I606523,I606540,I606580,I606602,I606619,I606645,I606653,I606670,I606687,I606704,I606721,I606766,I606797,I606814,I606840,I606848,I606879,I606896,I606913,I606930,I607002,I607028,I607036,I607076,I607084,I607101,I607118,I607158,I607180,I607197,I607223,I607231,I607248,I607265,I607282,I607299,I607344,I607375,I607392,I607418,I607426,I607457,I607474,I607491,I607508,I607580,I656155,I607606,I607614,I656149,I656134,I607654,I607662,I656140,I607679,I656152,I607696,I607736,I607758,I607775,I607801,I607809,I607826,I656158,I607843,I656146,I607860,I607877,I607922,I656137,I607953,I607970,I656143,I607996,I608004,I608035,I608052,I608069,I608086,I608158,I608184,I608192,I608232,I608240,I608257,I608274,I608314,I608336,I608353,I608379,I608387,I608404,I608421,I608438,I608455,I608500,I608531,I608548,I608574,I608582,I608613,I608630,I608647,I608664,I608736,I608762,I608770,I608810,I608818,I608835,I608852,I608892,I608914,I608931,I608957,I608965,I608982,I608999,I609016,I609033,I609078,I609109,I609126,I609152,I609160,I609191,I609208,I609225,I609242,I609314,I609340,I609348,I609388,I609396,I609413,I609430,I609470,I609492,I609509,I609535,I609543,I609560,I609577,I609594,I609611,I609656,I609687,I609704,I609730,I609738,I609769,I609786,I609803,I609820,I609892,I664859,I609918,I609926,I664853,I609875,I664838,I609966,I609974,I664844,I609991,I664856,I610008,I609863,I610048,I609884,I610070,I610087,I610113,I610121,I610138,I664862,I610155,I664850,I610172,I610189,I609860,I609881,I610234,I664841,I609872,I610265,I610282,I664847,I610308,I610316,I609878,I610347,I610364,I610381,I610398,I609869,I609866,I610470,I610496,I610504,I610544,I610552,I610569,I610586,I610626,I610648,I610665,I610691,I610699,I610716,I610733,I610750,I610767,I610812,I610843,I610860,I610886,I610894,I610925,I610942,I610959,I610976,I611048,I611074,I611082,I611122,I611130,I611147,I611164,I611204,I611226,I611243,I611269,I611277,I611294,I611311,I611328,I611345,I611390,I611421,I611438,I611464,I611472,I611503,I611520,I611537,I611554,I611626,I611652,I611660,I611700,I611708,I611725,I611742,I611782,I611804,I611821,I611847,I611855,I611872,I611889,I611906,I611923,I611968,I611999,I612016,I612042,I612050,I612081,I612098,I612115,I612132,I612204,I733545,I612230,I612238,I733527,I733518,I612278,I612286,I733533,I612303,I733521,I612320,I612360,I612382,I733530,I612399,I612425,I612433,I612450,I733539,I612467,I612484,I612501,I612546,I733542,I612577,I612594,I733536,I733524,I612620,I612628,I612659,I612676,I612693,I612710,I612782,I612808,I612816,I612856,I612864,I612881,I612898,I612938,I612960,I612977,I613003,I613011,I613028,I613045,I613062,I613079,I613124,I613155,I613172,I613198,I613206,I613237,I613254,I613271,I613288,I613360,I613386,I613394,I613434,I613442,I613459,I613476,I613516,I613538,I613555,I613581,I613589,I613606,I613623,I613640,I613657,I613702,I613733,I613750,I613776,I613784,I613815,I613832,I613849,I613866,I613938,I613964,I613972,I614012,I614020,I614037,I614054,I614094,I614116,I614133,I614159,I614167,I614184,I614201,I614218,I614235,I614280,I614311,I614328,I614354,I614362,I614393,I614410,I614427,I614444,I614516,I614542,I614550,I614590,I614598,I614615,I614632,I614672,I614694,I614711,I614737,I614745,I614762,I614779,I614796,I614813,I614858,I614889,I614906,I614932,I614940,I614971,I614988,I615005,I615022,I615094,I615120,I615128,I615168,I615176,I615193,I615210,I615250,I615272,I615289,I615315,I615323,I615340,I615357,I615374,I615391,I615436,I615467,I615484,I615510,I615518,I615549,I615566,I615583,I615600,I615672,I615698,I615706,I615746,I615754,I615771,I615788,I615828,I615850,I615867,I615893,I615901,I615918,I615935,I615952,I615969,I616014,I616045,I616062,I616088,I616096,I616127,I616144,I616161,I616178,I616250,I616276,I616284,I616324,I616332,I616349,I616366,I616406,I616428,I616445,I616471,I616479,I616496,I616513,I616530,I616547,I616592,I616623,I616640,I616666,I616674,I616705,I616722,I616739,I616756,I616828,I616854,I616862,I616902,I616910,I616927,I616944,I616984,I617006,I617023,I617049,I617057,I617074,I617091,I617108,I617125,I617170,I617201,I617218,I617244,I617252,I617283,I617300,I617317,I617334,I617406,I707960,I617432,I617440,I707942,I707933,I617480,I617488,I707948,I617505,I707936,I617522,I617562,I617584,I707945,I617601,I617627,I617635,I617652,I707954,I617669,I617686,I617703,I617748,I707957,I617779,I617796,I707951,I707939,I617822,I617830,I617861,I617878,I617895,I617912,I617984,I618010,I618018,I618058,I618066,I618083,I618100,I618140,I618162,I618179,I618205,I618213,I618230,I618247,I618264,I618281,I618326,I618357,I618374,I618400,I618408,I618439,I618456,I618473,I618490,I618562,I618588,I618596,I618636,I618644,I618661,I618678,I618718,I618740,I618757,I618783,I618791,I618808,I618825,I618842,I618859,I618904,I618935,I618952,I618978,I618986,I619017,I619034,I619051,I619068,I619140,I619166,I619174,I619214,I619222,I619239,I619256,I619296,I619318,I619335,I619361,I619369,I619386,I619403,I619420,I619437,I619482,I619513,I619530,I619556,I619564,I619595,I619612,I619629,I619646,I619718,I682338,I619744,I619752,I682320,I682329,I619792,I619800,I682314,I619817,I682326,I619834,I619874,I619896,I682317,I619913,I619939,I619947,I619964,I619981,I619998,I620015,I620060,I682335,I620091,I620108,I682323,I682332,I620134,I620142,I620173,I620190,I620207,I620224,I620296,I620322,I620330,I620279,I620370,I620378,I620395,I620412,I620267,I620452,I620288,I620474,I620491,I620517,I620525,I620542,I620559,I620576,I620593,I620264,I620285,I620638,I620276,I620669,I620686,I620712,I620720,I620282,I620751,I620768,I620785,I620802,I620273,I620270,I620874,I708555,I620900,I620908,I708537,I708528,I620948,I620956,I708543,I620973,I708531,I620990,I621030,I621052,I708540,I621069,I621095,I621103,I621120,I708549,I621137,I621154,I621171,I621216,I708552,I621247,I621264,I708546,I708534,I621290,I621298,I621329,I621346,I621363,I621380,I621452,I621478,I621486,I621435,I621526,I621534,I621551,I621568,I621423,I621608,I621444,I621630,I621647,I621673,I621681,I621698,I621715,I621732,I621749,I621420,I621441,I621794,I621432,I621825,I621842,I621868,I621876,I621438,I621907,I621924,I621941,I621958,I621429,I621426,I622030,I622056,I622064,I622104,I622112,I622129,I622146,I622186,I622208,I622225,I622251,I622259,I622276,I622293,I622310,I622327,I622372,I622403,I622420,I622446,I622454,I622485,I622502,I622519,I622536,I622608,I691008,I622634,I622642,I690990,I690999,I622682,I622690,I690984,I622707,I690996,I622724,I622764,I622786,I690987,I622803,I622829,I622837,I622854,I622871,I622888,I622905,I622950,I691005,I622981,I622998,I690993,I691002,I623024,I623032,I623063,I623080,I623097,I623114,I623186,I649083,I623212,I623220,I649077,I649062,I623260,I623268,I649068,I623285,I649080,I623302,I623342,I623364,I623381,I623407,I623415,I623432,I649086,I623449,I649074,I623466,I623483,I623528,I649065,I623559,I623576,I649071,I623602,I623610,I623641,I623658,I623675,I623692,I623764,I623790,I623798,I623838,I623846,I623863,I623880,I623920,I623942,I623959,I623985,I623993,I624010,I624027,I624044,I624061,I624106,I624137,I624154,I624180,I624188,I624219,I624236,I624253,I624270,I624342,I624368,I624376,I624416,I624424,I624441,I624458,I624498,I624520,I624537,I624563,I624571,I624588,I624605,I624622,I624639,I624684,I624715,I624732,I624758,I624766,I624797,I624814,I624831,I624848,I624920,I624946,I624954,I624994,I625002,I625019,I625036,I625076,I625098,I625115,I625141,I625149,I625166,I625183,I625200,I625217,I625262,I625293,I625310,I625336,I625344,I625375,I625392,I625409,I625426,I625498,I625524,I625532,I625572,I625580,I625597,I625614,I625654,I625676,I625693,I625719,I625727,I625744,I625761,I625778,I625795,I625840,I625871,I625888,I625914,I625922,I625953,I625970,I625987,I626004,I626076,I626102,I626110,I626150,I626158,I626175,I626192,I626232,I626254,I626271,I626297,I626305,I626322,I626339,I626356,I626373,I626418,I626449,I626466,I626492,I626500,I626531,I626548,I626565,I626582,I626654,I626680,I626688,I626728,I626736,I626753,I626770,I626810,I626832,I626849,I626875,I626883,I626900,I626917,I626934,I626951,I626996,I627027,I627044,I627070,I627078,I627109,I627126,I627143,I627160,I627232,I627258,I627266,I627306,I627314,I627331,I627348,I627388,I627410,I627427,I627453,I627461,I627478,I627495,I627512,I627529,I627574,I627605,I627622,I627648,I627656,I627687,I627704,I627721,I627738,I627810,I627836,I627844,I627884,I627892,I627909,I627926,I627966,I627988,I628005,I628031,I628039,I628056,I628073,I628090,I628107,I628152,I628183,I628200,I628226,I628234,I628265,I628282,I628299,I628316,I628388,I662139,I628414,I628422,I662133,I662118,I628462,I628470,I662124,I628487,I662136,I628504,I628544,I628566,I628583,I628609,I628617,I628634,I662142,I628651,I662130,I628668,I628685,I628730,I662121,I628761,I628778,I662127,I628804,I628812,I628843,I628860,I628877,I628894,I628966,I628992,I629000,I629040,I629048,I629065,I629082,I629122,I629144,I629161,I629187,I629195,I629212,I629229,I629246,I629263,I629308,I629339,I629356,I629382,I629390,I629421,I629438,I629455,I629472,I629544,I629570,I629578,I629618,I629626,I629643,I629660,I629700,I629722,I629739,I629765,I629773,I629790,I629807,I629824,I629841,I629886,I629917,I629934,I629960,I629968,I629999,I630016,I630033,I630050,I630122,I630148,I630156,I630196,I630204,I630221,I630238,I630278,I630300,I630317,I630343,I630351,I630368,I630385,I630402,I630419,I630464,I630495,I630512,I630538,I630546,I630577,I630594,I630611,I630628,I630700,I630726,I630734,I630774,I630782,I630799,I630816,I630856,I630878,I630895,I630921,I630929,I630946,I630963,I630980,I630997,I631042,I631073,I631090,I631116,I631124,I631155,I631172,I631189,I631206,I631278,I631304,I631312,I631352,I631360,I631377,I631394,I631434,I631456,I631473,I631499,I631507,I631524,I631541,I631558,I631575,I631620,I631651,I631668,I631694,I631702,I631733,I631750,I631767,I631784,I631856,I678870,I631882,I631890,I678852,I678861,I631930,I631938,I678846,I631955,I678858,I631972,I632012,I632034,I678849,I632051,I632077,I632085,I632102,I632119,I632136,I632153,I632198,I678867,I632229,I632246,I678855,I678864,I632272,I632280,I632311,I632328,I632345,I632362,I632434,I632460,I632468,I632508,I632516,I632533,I632550,I632590,I632612,I632629,I632655,I632663,I632680,I632697,I632714,I632731,I632776,I632807,I632824,I632850,I632858,I632889,I632906,I632923,I632940,I633012,I633038,I633046,I633086,I633094,I633111,I633128,I633168,I633190,I633207,I633233,I633241,I633258,I633275,I633292,I633309,I633354,I633385,I633402,I633428,I633436,I633467,I633484,I633501,I633518,I633590,I633616,I633624,I633664,I633672,I633689,I633706,I633746,I633768,I633785,I633811,I633819,I633836,I633853,I633870,I633887,I633932,I633963,I633980,I634006,I634014,I634045,I634062,I634079,I634096,I634168,I634194,I634202,I634242,I634250,I634267,I634284,I634324,I634346,I634363,I634389,I634397,I634414,I634431,I634448,I634465,I634510,I634541,I634558,I634584,I634592,I634623,I634640,I634657,I634674,I634746,I634772,I634780,I634820,I634828,I634845,I634862,I634902,I634924,I634941,I634967,I634975,I634992,I635009,I635026,I635043,I635088,I635119,I635136,I635162,I635170,I635201,I635218,I635235,I635252,I635324,I635350,I635358,I635398,I635406,I635423,I635440,I635480,I635502,I635519,I635545,I635553,I635570,I635587,I635604,I635621,I635666,I635697,I635714,I635740,I635748,I635779,I635796,I635813,I635830,I635902,I635928,I635936,I635976,I635984,I636001,I636018,I636058,I636080,I636097,I636123,I636131,I636148,I636165,I636182,I636199,I636244,I636275,I636292,I636318,I636326,I636357,I636374,I636391,I636408,I636480,I636506,I636514,I636554,I636562,I636579,I636596,I636636,I636658,I636675,I636701,I636709,I636726,I636743,I636760,I636777,I636822,I636853,I636870,I636896,I636904,I636935,I636952,I636969,I636986,I637058,I637084,I637092,I637132,I637140,I637157,I637174,I637214,I637236,I637253,I637279,I637287,I637304,I637321,I637338,I637355,I637400,I637431,I637448,I637474,I637482,I637513,I637530,I637547,I637564,I637636,I637662,I637670,I637710,I637718,I637735,I637752,I637792,I637814,I637831,I637857,I637865,I637882,I637899,I637916,I637933,I637978,I638009,I638026,I638052,I638060,I638091,I638108,I638125,I638142,I638214,I638240,I638248,I638288,I638296,I638313,I638330,I638370,I638392,I638409,I638435,I638443,I638460,I638477,I638494,I638511,I638556,I638587,I638604,I638630,I638638,I638669,I638686,I638703,I638720,I638792,I638818,I638826,I638866,I638874,I638891,I638908,I638948,I638970,I638987,I639013,I639021,I639038,I639055,I639072,I639089,I639134,I639165,I639182,I639208,I639216,I639247,I639264,I639281,I639298,I639370,I639396,I639404,I639353,I639444,I639452,I639469,I639486,I639341,I639526,I639362,I639548,I639565,I639591,I639599,I639616,I639633,I639650,I639667,I639338,I639359,I639712,I639350,I639743,I639760,I639786,I639794,I639356,I639825,I639842,I639859,I639876,I639347,I639344,I639948,I639974,I639982,I640022,I640030,I640047,I640064,I640104,I640126,I640143,I640169,I640177,I640194,I640211,I640228,I640245,I640290,I640321,I640338,I640364,I640372,I640403,I640420,I640437,I640454,I640526,I640552,I640560,I640600,I640608,I640625,I640642,I640682,I640704,I640721,I640747,I640755,I640772,I640789,I640806,I640823,I640868,I640899,I640916,I640942,I640950,I640981,I640998,I641015,I641032,I641104,I641130,I641138,I641178,I641186,I641203,I641220,I641260,I641282,I641299,I641325,I641333,I641350,I641367,I641384,I641401,I641446,I641477,I641494,I641520,I641528,I641559,I641576,I641593,I641610,I641682,I641708,I641716,I641665,I641756,I641764,I641781,I641798,I641653,I641838,I641674,I641860,I641877,I641903,I641911,I641928,I641945,I641962,I641979,I641650,I641671,I642024,I641662,I642055,I642072,I642098,I642106,I641668,I642137,I642154,I642171,I642188,I641659,I641656,I642260,I642286,I642294,I642334,I642342,I642359,I642376,I642416,I642438,I642455,I642481,I642489,I642506,I642523,I642540,I642557,I642602,I642633,I642650,I642676,I642684,I642715,I642732,I642749,I642766,I642838,I642864,I642872,I642912,I642920,I642937,I642954,I642994,I643016,I643033,I643059,I643067,I643084,I643101,I643118,I643135,I643180,I643211,I643228,I643254,I643262,I643293,I643310,I643327,I643344,I643416,I643442,I643450,I643490,I643498,I643515,I643532,I643572,I643594,I643611,I643637,I643645,I643662,I643679,I643696,I643713,I643758,I643789,I643806,I643832,I643840,I643871,I643888,I643905,I643922,I643994,I644020,I644028,I644068,I644076,I644093,I644110,I644150,I644172,I644189,I644215,I644223,I644240,I644257,I644274,I644291,I644336,I644367,I644384,I644410,I644418,I644449,I644466,I644483,I644500,I644572,I644598,I644606,I644646,I644654,I644671,I644688,I644728,I644750,I644767,I644793,I644801,I644818,I644835,I644852,I644869,I644914,I644945,I644962,I644988,I644996,I645027,I645044,I645061,I645078,I645150,I645176,I645184,I645224,I645232,I645249,I645266,I645306,I645328,I645345,I645371,I645379,I645396,I645413,I645430,I645447,I645492,I645523,I645540,I645566,I645574,I645605,I645622,I645639,I645656,I645728,I645754,I645762,I645802,I645810,I645827,I645844,I645884,I645906,I645923,I645949,I645957,I645974,I645991,I646008,I646025,I646070,I646101,I646118,I646144,I646152,I646183,I646200,I646217,I646234,I646306,I646332,I646340,I646380,I646388,I646405,I646422,I646462,I646484,I646501,I646527,I646535,I646552,I646569,I646586,I646603,I646648,I646679,I646696,I646722,I646730,I646761,I646778,I646795,I646812,I646884,I706175,I646910,I646918,I706157,I706148,I646958,I646966,I706163,I646983,I706151,I647000,I647040,I647062,I706160,I647079,I647105,I647113,I647130,I706169,I647147,I647164,I647181,I647226,I706172,I647257,I647274,I706166,I706154,I647300,I647308,I647339,I647356,I647373,I647390,I647462,I647488,I647496,I647522,I647539,I647561,I647578,I647595,I647612,I647629,I647660,I647677,I647694,I647711,I647756,I647773,I647790,I647849,I647875,I647883,I647900,I647917,I647948,I648006,I648032,I648040,I648066,I648083,I648105,I648122,I648139,I648156,I648173,I648204,I648221,I648238,I648255,I648300,I648317,I648334,I648393,I648419,I648427,I648444,I648461,I648492,I648550,I648576,I648584,I648610,I648627,I648649,I648666,I648683,I648700,I648717,I648748,I648765,I648782,I648799,I648844,I648861,I648878,I648937,I648963,I648971,I648988,I649005,I649036,I649094,I649120,I649128,I649154,I649171,I649193,I649210,I649227,I649244,I649261,I649292,I649309,I649326,I649343,I649388,I649405,I649422,I649481,I649507,I649515,I649532,I649549,I649580,I649638,I649664,I649672,I649698,I649715,I649737,I649754,I649771,I649788,I649805,I649836,I649853,I649870,I649887,I649932,I649949,I649966,I650025,I650051,I650059,I650076,I650093,I650124,I650182,I650208,I650216,I650242,I650259,I650281,I650298,I650315,I650332,I650349,I650380,I650397,I650414,I650431,I650476,I650493,I650510,I650569,I650595,I650603,I650620,I650637,I650668,I650726,I677121,I650752,I650760,I677130,I677133,I650786,I650803,I650825,I677127,I650842,I677124,I650859,I677118,I650876,I650893,I650924,I677115,I650941,I677112,I650958,I650975,I651020,I651037,I651054,I651113,I677136,I651139,I651147,I651164,I651181,I651212,I651270,I651296,I651304,I651330,I651347,I651369,I651386,I651403,I651420,I651437,I651468,I651485,I651502,I651519,I651564,I651581,I651598,I651657,I651683,I651691,I651708,I651725,I651756,I651814,I651840,I651848,I651874,I651891,I651913,I651930,I651947,I651964,I651981,I652012,I652029,I652046,I652063,I652108,I652125,I652142,I652201,I652227,I652235,I652252,I652269,I652300,I652358,I652384,I652392,I652418,I652435,I652457,I652474,I652491,I652508,I652525,I652556,I652573,I652590,I652607,I652652,I652669,I652686,I652745,I652771,I652779,I652796,I652813,I652844,I652902,I652928,I652936,I652962,I652979,I653001,I653018,I653035,I653052,I653069,I653100,I653117,I653134,I653151,I653196,I653213,I653230,I653289,I653315,I653323,I653340,I653357,I653388,I653446,I653472,I653480,I653506,I653523,I653545,I653562,I653579,I653596,I653613,I653644,I653661,I653678,I653695,I653740,I653757,I653774,I653833,I653859,I653867,I653884,I653901,I653932,I653990,I654016,I654024,I654050,I654067,I654089,I654106,I654123,I654140,I654157,I654188,I654205,I654222,I654239,I654284,I654301,I654318,I654377,I654403,I654411,I654428,I654445,I654476,I654534,I677699,I654560,I654568,I677708,I677711,I654594,I654611,I654633,I677705,I654650,I677702,I654667,I677696,I654684,I654701,I654732,I677693,I654749,I677690,I654766,I654783,I654828,I654845,I654862,I654921,I677714,I654947,I654955,I654972,I654989,I655020,I655078,I673075,I655104,I655112,I673084,I673087,I655138,I655155,I655177,I673081,I655194,I673078,I655211,I673072,I655228,I655245,I655276,I673069,I655293,I673066,I655310,I655327,I655372,I655389,I655406,I655465,I673090,I655491,I655499,I655516,I655533,I655564,I655622,I655648,I655656,I655682,I655699,I655614,I655721,I655738,I655755,I655772,I655789,I655593,I655820,I655837,I655854,I655871,I655596,I655611,I655916,I655933,I655950,I655608,I655605,I655602,I656009,I656035,I656043,I656060,I656077,I655590,I656108,I655599,I656166,I656192,I656200,I656226,I656243,I656265,I656282,I656299,I656316,I656333,I656364,I656381,I656398,I656415,I656460,I656477,I656494,I656553,I656579,I656587,I656604,I656621,I656652,I656710,I656736,I656744,I656770,I656787,I656809,I656826,I656843,I656860,I656877,I656908,I656925,I656942,I656959,I657004,I657021,I657038,I657097,I657123,I657131,I657148,I657165,I657196,I657254,I657280,I657288,I657314,I657331,I657353,I657370,I657387,I657404,I657421,I657452,I657469,I657486,I657503,I657548,I657565,I657582,I657641,I657667,I657675,I657692,I657709,I657740,I657798,I691571,I657824,I657832,I691580,I691583,I657858,I657875,I657897,I691577,I657914,I691574,I657931,I691568,I657948,I657965,I657996,I691565,I658013,I691562,I658030,I658047,I658092,I658109,I658126,I658185,I691586,I658211,I658219,I658236,I658253,I658284,I658342,I658368,I658376,I658402,I658419,I658334,I658441,I658458,I658475,I658492,I658509,I658313,I658540,I658557,I658574,I658591,I658316,I658331,I658636,I658653,I658670,I658328,I658325,I658322,I658729,I658755,I658763,I658780,I658797,I658310,I658828,I658319,I658886,I658912,I658920,I658946,I658963,I658985,I659002,I659019,I659036,I659053,I659084,I659101,I659118,I659135,I659180,I659197,I659214,I659273,I659299,I659307,I659324,I659341,I659372,I659430,I659456,I659464,I659490,I659507,I659422,I659529,I659546,I659563,I659580,I659597,I659401,I659628,I659645,I659662,I659679,I659404,I659419,I659724,I659741,I659758,I659416,I659413,I659410,I659817,I659843,I659851,I659868,I659885,I659398,I659916,I659407,I659974,I660000,I660008,I660034,I660051,I660073,I660090,I660107,I660124,I660141,I660172,I660189,I660206,I660223,I660268,I660285,I660302,I660361,I660387,I660395,I660412,I660429,I660460,I660518,I660544,I660552,I660578,I660595,I660617,I660634,I660651,I660668,I660685,I660716,I660733,I660750,I660767,I660812,I660829,I660846,I660905,I660931,I660939,I660956,I660973,I661004,I661062,I661088,I661096,I661122,I661139,I661161,I661178,I661195,I661212,I661229,I661260,I661277,I661294,I661311,I661356,I661373,I661390,I661449,I661475,I661483,I661500,I661517,I661548,I661606,I661632,I661640,I661666,I661683,I661705,I661722,I661739,I661756,I661773,I661804,I661821,I661838,I661855,I661900,I661917,I661934,I661993,I662019,I662027,I662044,I662061,I662092,I662150,I662176,I662184,I662210,I662227,I662249,I662266,I662283,I662300,I662317,I662348,I662365,I662382,I662399,I662444,I662461,I662478,I662537,I662563,I662571,I662588,I662605,I662636,I662694,I662720,I662728,I662754,I662771,I662793,I662810,I662827,I662844,I662861,I662892,I662909,I662926,I662943,I662988,I663005,I663022,I663081,I663107,I663115,I663132,I663149,I663180,I663238,I704985,I663264,I663272,I704970,I704964,I663298,I663315,I663337,I704958,I663354,I704979,I663371,I704967,I663388,I663405,I663436,I704976,I663453,I704982,I663470,I704973,I663487,I663532,I704961,I663549,I663566,I663625,I663651,I663659,I663676,I663693,I663724,I663782,I663808,I663816,I663842,I663859,I663881,I663898,I663915,I663932,I663949,I663980,I663997,I664014,I664031,I664076,I664093,I664110,I664169,I664195,I664203,I664220,I664237,I664268,I664326,I664352,I664360,I664386,I664403,I664425,I664442,I664459,I664476,I664493,I664524,I664541,I664558,I664575,I664620,I664637,I664654,I664713,I664739,I664747,I664764,I664781,I664812,I664870,I664896,I664904,I664930,I664947,I664969,I664986,I665003,I665020,I665037,I665068,I665085,I665102,I665119,I665164,I665181,I665198,I665257,I665283,I665291,I665308,I665325,I665356,I665414,I732355,I665440,I665448,I732340,I732334,I665474,I665491,I665513,I732328,I665530,I732349,I665547,I732337,I665564,I665581,I665612,I732346,I665629,I732352,I665646,I732343,I665663,I665708,I732331,I665725,I665742,I665801,I665827,I665835,I665852,I665869,I665900,I665958,I665984,I665992,I666018,I666035,I666057,I666074,I666091,I666108,I666125,I666156,I666173,I666190,I666207,I666252,I666269,I666286,I666345,I666371,I666379,I666396,I666413,I666444,I666502,I666528,I666536,I666562,I666579,I666601,I666618,I666635,I666652,I666669,I666700,I666717,I666734,I666751,I666796,I666813,I666830,I666889,I666915,I666923,I666940,I666957,I666988,I667046,I725215,I667072,I667080,I725200,I725194,I667106,I667123,I667145,I725188,I667162,I725209,I667179,I725197,I667196,I667213,I667244,I725206,I667261,I725212,I667278,I725203,I667295,I667340,I725191,I667357,I667374,I667433,I667459,I667467,I667484,I667501,I667532,I667590,I667616,I667624,I667650,I667667,I667689,I667706,I667723,I667740,I667757,I667788,I667805,I667822,I667839,I667884,I667901,I667918,I667977,I668003,I668011,I668028,I668045,I668076,I668134,I668160,I668168,I668194,I668211,I668233,I668250,I668267,I668284,I668301,I668332,I668349,I668366,I668383,I668428,I668445,I668462,I668521,I668547,I668555,I668572,I668589,I668620,I668678,I668704,I668712,I668738,I668755,I668777,I668794,I668811,I668828,I668845,I668876,I668893,I668910,I668927,I668972,I668989,I669006,I669065,I669091,I669099,I669116,I669133,I669164,I669222,I669248,I669256,I669282,I669299,I669321,I669338,I669355,I669372,I669389,I669420,I669437,I669454,I669471,I669516,I669533,I669550,I669609,I669635,I669643,I669660,I669677,I669708,I669766,I735925,I669792,I669800,I735910,I735904,I669826,I669843,I669865,I735898,I669882,I735919,I669899,I735907,I669916,I669933,I669964,I735916,I669981,I735922,I669998,I735913,I670015,I670060,I735901,I670077,I670094,I670153,I670179,I670187,I670204,I670221,I670252,I670310,I670336,I670344,I670370,I670387,I670409,I670426,I670443,I670460,I670477,I670508,I670525,I670542,I670559,I670604,I670621,I670638,I670697,I670723,I670731,I670748,I670765,I670796,I670854,I670880,I670888,I670914,I670931,I670953,I670970,I670987,I671004,I671021,I671052,I671069,I671086,I671103,I671148,I671165,I671182,I671241,I671267,I671275,I671292,I671309,I671340,I671398,I671424,I671432,I671458,I671475,I671497,I671514,I671531,I671548,I671565,I671596,I671613,I671630,I671647,I671692,I671709,I671726,I671785,I671811,I671819,I671836,I671853,I671884,I671942,I671968,I671976,I671993,I672019,I672027,I672044,I672061,I672078,I672095,I672126,I672143,I672160,I672191,I672208,I672248,I672256,I672287,I672304,I672321,I672338,I672369,I672400,I672426,I672448,I672520,I672546,I672554,I672571,I672597,I672605,I672622,I672639,I672656,I672673,I672704,I672721,I672738,I672769,I672786,I672826,I672834,I672865,I672882,I672899,I672916,I672947,I672978,I673004,I673026,I673098,I673124,I673132,I673149,I673175,I673183,I673200,I673217,I673234,I673251,I673282,I673299,I673316,I673347,I673364,I673404,I673412,I673443,I673460,I673477,I673494,I673525,I673556,I673582,I673604,I673676,I673702,I673710,I673727,I673753,I673761,I673778,I673795,I673812,I673829,I673860,I673877,I673894,I673925,I673942,I673982,I673990,I674021,I674038,I674055,I674072,I674103,I674134,I674160,I674182,I674254,I674280,I674288,I674305,I674331,I674339,I674356,I674373,I674390,I674407,I674438,I674455,I674472,I674503,I674520,I674560,I674568,I674599,I674616,I674633,I674650,I674681,I674712,I674738,I674760,I674832,I674858,I674866,I674883,I674909,I674917,I674934,I674951,I674968,I674985,I675016,I675033,I675050,I675081,I675098,I675138,I675146,I675177,I675194,I675211,I675228,I675259,I675290,I675316,I675338,I675410,I675436,I675444,I675461,I675487,I675495,I675512,I675529,I675546,I675563,I675594,I675611,I675628,I675659,I675676,I675716,I675724,I675755,I675772,I675789,I675806,I675837,I675868,I675894,I675916,I675988,I676014,I676022,I676039,I676065,I676073,I676090,I676107,I676124,I676141,I676172,I676189,I676206,I676237,I676254,I676294,I676302,I676333,I676350,I676367,I676384,I676415,I676446,I676472,I676494,I676566,I676592,I676600,I676617,I676643,I676651,I676668,I676685,I676702,I676719,I676750,I676767,I676784,I676815,I676832,I676872,I676880,I676911,I676928,I676945,I676962,I676993,I677024,I677050,I677072,I677144,I677170,I677178,I677195,I677221,I677229,I677246,I677263,I677280,I677297,I677328,I677345,I677362,I677393,I677410,I677450,I677458,I677489,I677506,I677523,I677540,I677571,I677602,I677628,I677650,I677722,I677748,I677756,I677773,I677799,I677807,I677824,I677841,I677858,I677875,I677906,I677923,I677940,I677971,I677988,I678028,I678036,I678067,I678084,I678101,I678118,I678149,I678180,I678206,I678228,I678300,I678326,I678334,I678351,I678377,I678385,I678402,I678419,I678436,I678453,I678484,I678501,I678518,I678549,I678566,I678606,I678614,I678645,I678662,I678679,I678696,I678727,I678758,I678784,I678806,I678878,I678904,I678912,I678929,I678955,I678963,I678980,I678997,I679014,I679031,I679062,I679079,I679096,I679127,I679144,I679184,I679192,I679223,I679240,I679257,I679274,I679305,I679336,I679362,I679384,I679456,I709147,I679482,I679490,I709138,I679507,I709123,I679533,I679541,I679558,I709126,I679575,I709135,I679592,I679609,I709132,I679640,I709144,I679657,I679674,I679705,I709129,I679722,I679762,I679770,I679801,I709150,I679818,I679835,I679852,I679883,I679914,I709141,I679940,I679962,I680034,I680060,I680068,I680085,I680111,I680119,I680136,I680153,I680170,I680187,I680218,I680235,I680252,I680283,I680300,I680340,I680348,I680379,I680396,I680413,I680430,I680461,I680492,I680518,I680540,I680612,I680638,I680646,I680663,I680689,I680697,I680714,I680731,I680748,I680765,I680796,I680813,I680830,I680861,I680878,I680918,I680926,I680957,I680974,I680991,I681008,I681039,I681070,I681096,I681118,I681190,I681216,I681224,I681241,I681267,I681275,I681292,I681309,I681326,I681343,I681374,I681391,I681408,I681439,I681456,I681496,I681504,I681535,I681552,I681569,I681586,I681617,I681648,I681674,I681696,I681768,I681794,I681802,I681819,I681845,I681853,I681870,I681887,I681904,I681921,I681952,I681969,I681986,I682017,I682034,I682074,I682082,I682113,I682130,I682147,I682164,I682195,I682226,I682252,I682274,I682346,I682372,I682380,I682397,I682423,I682431,I682448,I682465,I682482,I682499,I682530,I682547,I682564,I682595,I682612,I682652,I682660,I682691,I682708,I682725,I682742,I682773,I682804,I682830,I682852,I682924,I682950,I682958,I682975,I683001,I683009,I683026,I683043,I683060,I683077,I683108,I683125,I683142,I683173,I683190,I683230,I683238,I683269,I683286,I683303,I683320,I683351,I683382,I683408,I683430,I683502,I683528,I683536,I683553,I683579,I683587,I683604,I683621,I683638,I683655,I683686,I683703,I683720,I683751,I683768,I683808,I683816,I683847,I683864,I683881,I683898,I683929,I683960,I683986,I684008,I684080,I684106,I684114,I684131,I684157,I684165,I684182,I684199,I684216,I684233,I684264,I684281,I684298,I684329,I684346,I684386,I684394,I684425,I684442,I684459,I684476,I684507,I684538,I684564,I684586,I684658,I684684,I684692,I684709,I684735,I684743,I684760,I684777,I684794,I684811,I684842,I684859,I684876,I684907,I684924,I684964,I684972,I685003,I685020,I685037,I685054,I685085,I685116,I685142,I685164,I685236,I685262,I685270,I685287,I685313,I685321,I685338,I685355,I685372,I685389,I685420,I685437,I685454,I685485,I685502,I685542,I685550,I685581,I685598,I685615,I685632,I685663,I685694,I685720,I685742,I685814,I685840,I685848,I685865,I685891,I685899,I685916,I685933,I685950,I685967,I685998,I686015,I686032,I686063,I686080,I686120,I686128,I686159,I686176,I686193,I686210,I686241,I686272,I686298,I686320,I686392,I686418,I686426,I686443,I686469,I686477,I686494,I686511,I686528,I686545,I686576,I686593,I686610,I686641,I686658,I686698,I686706,I686737,I686754,I686771,I686788,I686819,I686850,I686876,I686898,I686970,I686996,I687004,I687021,I687047,I687055,I687072,I687089,I687106,I687123,I687154,I687171,I687188,I687219,I687236,I687276,I687284,I687315,I687332,I687349,I687366,I687397,I687428,I687454,I687476,I687548,I732947,I687574,I687582,I732938,I687599,I732923,I687625,I687633,I687650,I732926,I687667,I732935,I687684,I687701,I732932,I687732,I732944,I687749,I687766,I687797,I732929,I687814,I687854,I687862,I687893,I732950,I687910,I687927,I687944,I687975,I688006,I732941,I688032,I688054,I688126,I688152,I688160,I688177,I688203,I688211,I688228,I688245,I688262,I688279,I688310,I688327,I688344,I688375,I688392,I688432,I688440,I688471,I688488,I688505,I688522,I688553,I688584,I688610,I688632,I688704,I688730,I688738,I688755,I688781,I688789,I688806,I688823,I688840,I688857,I688888,I688905,I688922,I688953,I688970,I689010,I689018,I689049,I689066,I689083,I689100,I689131,I689162,I689188,I689210,I689282,I689308,I689316,I689333,I689359,I689367,I689384,I689401,I689418,I689435,I689274,I689466,I689483,I689500,I689253,I689531,I689548,I689259,I689588,I689596,I689268,I689627,I689644,I689661,I689678,I689271,I689709,I689250,I689740,I689766,I689265,I689788,I689262,I689256,I689860,I689886,I689894,I689911,I689937,I689945,I689962,I689979,I689996,I690013,I690044,I690061,I690078,I690109,I690126,I690166,I690174,I690205,I690222,I690239,I690256,I690287,I690318,I690344,I690366,I690438,I690464,I690472,I690489,I690515,I690523,I690540,I690557,I690574,I690591,I690622,I690639,I690656,I690687,I690704,I690744,I690752,I690783,I690800,I690817,I690834,I690865,I690896,I690922,I690944,I691016,I691042,I691050,I691067,I691093,I691101,I691118,I691135,I691152,I691169,I691200,I691217,I691234,I691265,I691282,I691322,I691330,I691361,I691378,I691395,I691412,I691443,I691474,I691500,I691522,I691594,I691620,I691628,I691645,I691671,I691679,I691696,I691713,I691730,I691747,I691778,I691795,I691812,I691843,I691860,I691900,I691908,I691939,I691956,I691973,I691990,I692021,I692052,I692078,I692100,I692172,I692198,I692206,I692223,I692249,I692257,I692274,I692291,I692308,I692325,I692356,I692373,I692390,I692421,I692438,I692478,I692486,I692517,I692534,I692551,I692568,I692599,I692630,I692656,I692678,I692750,I692776,I692784,I692801,I692827,I692835,I692852,I692869,I692886,I692903,I692742,I692934,I692951,I692968,I692721,I692999,I693016,I692727,I693056,I693064,I692736,I693095,I693112,I693129,I693146,I692739,I693177,I692718,I693208,I693234,I692733,I693256,I692730,I692724,I693331,I693357,I693365,I693382,I693408,I693416,I693433,I693450,I693481,I693512,I693529,I693546,I693563,I693580,I693611,I693670,I693687,I693713,I693735,I693761,I693769,I693786,I693817,I693892,I693918,I693926,I693943,I693969,I693977,I693994,I694011,I694042,I694073,I694090,I694107,I694124,I694141,I694172,I694231,I694248,I694274,I694296,I694322,I694330,I694347,I694378,I694453,I694479,I694487,I694504,I694530,I694538,I694555,I694572,I694603,I694634,I694651,I694668,I694685,I694702,I694733,I694792,I694809,I694835,I694857,I694883,I694891,I694908,I694939,I695014,I695040,I695048,I695065,I695091,I695099,I695116,I695133,I695164,I695195,I695212,I695229,I695246,I695263,I695294,I695353,I695370,I695396,I695418,I695444,I695452,I695469,I695500,I695575,I695601,I695609,I695626,I695652,I695660,I695677,I695694,I695725,I695756,I695773,I695790,I695807,I695824,I695855,I695914,I695931,I695957,I695979,I696005,I696013,I696030,I696061,I696136,I696162,I696170,I696187,I696213,I696221,I696238,I696255,I696286,I696317,I696334,I696351,I696368,I696385,I696416,I696475,I696492,I696518,I696540,I696566,I696574,I696591,I696622,I696697,I696723,I696731,I696748,I696774,I696782,I696799,I696816,I696847,I696878,I696895,I696912,I696929,I696946,I696977,I697036,I697053,I697079,I697101,I697127,I697135,I697152,I697183,I697258,I697284,I697301,I697309,I697354,I697371,I697388,I697405,I697422,I697439,I697456,I697487,I697504,I697549,I697566,I697583,I697614,I697640,I697648,I697679,I697696,I697713,I697739,I697747,I697764,I697853,I697879,I697896,I697904,I697949,I697966,I697983,I698000,I698017,I698034,I698051,I698082,I698099,I698144,I698161,I698178,I698209,I698235,I698243,I698274,I698291,I698308,I698334,I698342,I698359,I698448,I698474,I698491,I698499,I698544,I698561,I698578,I698595,I698612,I698629,I698646,I698677,I698694,I698739,I698756,I698773,I698804,I698830,I698838,I698869,I698886,I698903,I698929,I698937,I698954,I699043,I699069,I699086,I699094,I699139,I699156,I699173,I699190,I699207,I699224,I699241,I699272,I699289,I699334,I699351,I699368,I699399,I699425,I699433,I699464,I699481,I699498,I699524,I699532,I699549,I699638,I699664,I699681,I699689,I699734,I699751,I699768,I699785,I699802,I699819,I699836,I699867,I699884,I699929,I699946,I699963,I699994,I700020,I700028,I700059,I700076,I700093,I700119,I700127,I700144,I700233,I700259,I700276,I700284,I700329,I700346,I700363,I700380,I700397,I700414,I700431,I700462,I700479,I700524,I700541,I700558,I700589,I700615,I700623,I700654,I700671,I700688,I700714,I700722,I700739,I700828,I700854,I700871,I700879,I700924,I700941,I700958,I700975,I700992,I701009,I701026,I701057,I701074,I701119,I701136,I701153,I701184,I701210,I701218,I701249,I701266,I701283,I701309,I701317,I701334,I701423,I701449,I701466,I701474,I701519,I701536,I701553,I701570,I701587,I701604,I701621,I701652,I701669,I701714,I701731,I701748,I701779,I701805,I701813,I701844,I701861,I701878,I701904,I701912,I701929,I702018,I702044,I702061,I702069,I702114,I702131,I702148,I702165,I702182,I702199,I702216,I702247,I702264,I702309,I702326,I702343,I702374,I702400,I702408,I702439,I702456,I702473,I702499,I702507,I702524,I702613,I702639,I702656,I702664,I702709,I702726,I702743,I702760,I702777,I702794,I702811,I702842,I702859,I702904,I702921,I702938,I702969,I702995,I703003,I703034,I703051,I703068,I703094,I703102,I703119,I703208,I703234,I703251,I703259,I703304,I703321,I703338,I703355,I703372,I703389,I703406,I703437,I703454,I703499,I703516,I703533,I703564,I703590,I703598,I703629,I703646,I703663,I703689,I703697,I703714,I703803,I703829,I703846,I703854,I703899,I703916,I703933,I703950,I703967,I703984,I704001,I704032,I704049,I704094,I704111,I704128,I704159,I704185,I704193,I704224,I704241,I704258,I704284,I704292,I704309,I704398,I704424,I704441,I704449,I704494,I704511,I704528,I704545,I704562,I704579,I704596,I704627,I704644,I704689,I704706,I704723,I704754,I704780,I704788,I704819,I704836,I704853,I704879,I704887,I704904,I704993,I705019,I705036,I705044,I705089,I705106,I705123,I705140,I705157,I705174,I705191,I705222,I705239,I705284,I705301,I705318,I705349,I705375,I705383,I705414,I705431,I705448,I705474,I705482,I705499,I705588,I705614,I705631,I705639,I705684,I705701,I705718,I705735,I705752,I705769,I705786,I705817,I705834,I705879,I705896,I705913,I705944,I705970,I705978,I706009,I706026,I706043,I706069,I706077,I706094,I706183,I706209,I706226,I706234,I706279,I706296,I706313,I706330,I706347,I706364,I706381,I706412,I706429,I706474,I706491,I706508,I706539,I706565,I706573,I706604,I706621,I706638,I706664,I706672,I706689,I706778,I706804,I706821,I706829,I706874,I706891,I706908,I706925,I706942,I706959,I706976,I707007,I707024,I707069,I707086,I707103,I707134,I707160,I707168,I707199,I707216,I707233,I707259,I707267,I707284,I707373,I707399,I707416,I707424,I707469,I707486,I707503,I707520,I707537,I707554,I707571,I707602,I707619,I707664,I707681,I707698,I707729,I707755,I707763,I707794,I707811,I707828,I707854,I707862,I707879,I707968,I707994,I708011,I708019,I708064,I708081,I708098,I708115,I708132,I708149,I708166,I708197,I708214,I708259,I708276,I708293,I708324,I708350,I708358,I708389,I708406,I708423,I708449,I708457,I708474,I708563,I708589,I708606,I708614,I708659,I708676,I708693,I708710,I708727,I708744,I708761,I708792,I708809,I708854,I708871,I708888,I708919,I708945,I708953,I708984,I709001,I709018,I709044,I709052,I709069,I709158,I709184,I709201,I709209,I709254,I709271,I709288,I709305,I709322,I709339,I709356,I709387,I709404,I709449,I709466,I709483,I709514,I709540,I709548,I709579,I709596,I709613,I709639,I709647,I709664,I709753,I709779,I709796,I709804,I709849,I709866,I709883,I709900,I709917,I709934,I709951,I709982,I709999,I710044,I710061,I710078,I710109,I710135,I710143,I710174,I710191,I710208,I710234,I710242,I710259,I710348,I710374,I710391,I710399,I710444,I710461,I710478,I710495,I710512,I710529,I710546,I710577,I710594,I710639,I710656,I710673,I710704,I710730,I710738,I710769,I710786,I710803,I710829,I710837,I710854,I710943,I710969,I710986,I710994,I711039,I711056,I711073,I711090,I711107,I711124,I711141,I711172,I711189,I711234,I711251,I711268,I711299,I711325,I711333,I711364,I711381,I711398,I711424,I711432,I711449,I711538,I711564,I711581,I711589,I711634,I711651,I711668,I711685,I711702,I711719,I711736,I711767,I711784,I711829,I711846,I711863,I711894,I711920,I711928,I711959,I711976,I711993,I712019,I712027,I712044,I712133,I712159,I712176,I712184,I712229,I712246,I712263,I712280,I712297,I712314,I712331,I712362,I712379,I712424,I712441,I712458,I712489,I712515,I712523,I712554,I712571,I712588,I712614,I712622,I712639,I712728,I712754,I712771,I712779,I712824,I712841,I712858,I712875,I712892,I712909,I712926,I712957,I712974,I713019,I713036,I713053,I713084,I713110,I713118,I713149,I713166,I713183,I713209,I713217,I713234,I713323,I713349,I713366,I713374,I713419,I713436,I713453,I713470,I713487,I713504,I713521,I713552,I713569,I713614,I713631,I713648,I713679,I713705,I713713,I713744,I713761,I713778,I713804,I713812,I713829,I713918,I713944,I713961,I713969,I714014,I714031,I714048,I714065,I714082,I714099,I714116,I714147,I714164,I714209,I714226,I714243,I714274,I714300,I714308,I714339,I714356,I714373,I714399,I714407,I714424,I714513,I714539,I714556,I714564,I714609,I714626,I714643,I714660,I714677,I714694,I714711,I714742,I714759,I714804,I714821,I714838,I714869,I714895,I714903,I714934,I714951,I714968,I714994,I715002,I715019,I715108,I715134,I715151,I715159,I715204,I715221,I715238,I715255,I715272,I715289,I715306,I715337,I715354,I715399,I715416,I715433,I715464,I715490,I715498,I715529,I715546,I715563,I715589,I715597,I715614,I715703,I715729,I715746,I715754,I715799,I715816,I715833,I715850,I715867,I715884,I715901,I715932,I715949,I715994,I716011,I716028,I716059,I716085,I716093,I716124,I716141,I716158,I716184,I716192,I716209,I716298,I716324,I716341,I716349,I716394,I716411,I716428,I716445,I716462,I716479,I716496,I716527,I716544,I716589,I716606,I716623,I716654,I716680,I716688,I716719,I716736,I716753,I716779,I716787,I716804,I716893,I716919,I716936,I716944,I716989,I717006,I717023,I717040,I717057,I717074,I717091,I717122,I717139,I717184,I717201,I717218,I717249,I717275,I717283,I717314,I717331,I717348,I717374,I717382,I717399,I717488,I717514,I717531,I717539,I717584,I717601,I717618,I717635,I717652,I717669,I717686,I717717,I717734,I717779,I717796,I717813,I717844,I717870,I717878,I717909,I717926,I717943,I717969,I717977,I717994,I718083,I718109,I718126,I718134,I718179,I718196,I718213,I718230,I718247,I718264,I718281,I718312,I718329,I718374,I718391,I718408,I718439,I718465,I718473,I718504,I718521,I718538,I718564,I718572,I718589,I718678,I718704,I718721,I718729,I718774,I718791,I718808,I718825,I718842,I718859,I718876,I718907,I718924,I718969,I718986,I719003,I719034,I719060,I719068,I719099,I719116,I719133,I719159,I719167,I719184,I719273,I719299,I719316,I719324,I719369,I719386,I719403,I719420,I719437,I719454,I719471,I719502,I719519,I719564,I719581,I719598,I719629,I719655,I719663,I719694,I719711,I719728,I719754,I719762,I719779,I719868,I719894,I719911,I719919,I719964,I719981,I719998,I720015,I720032,I720049,I720066,I720097,I720114,I720159,I720176,I720193,I720224,I720250,I720258,I720289,I720306,I720323,I720349,I720357,I720374,I720463,I720489,I720506,I720514,I720559,I720576,I720593,I720610,I720627,I720644,I720661,I720692,I720709,I720754,I720771,I720788,I720819,I720845,I720853,I720884,I720901,I720918,I720944,I720952,I720969,I721058,I721084,I721101,I721109,I721154,I721171,I721188,I721205,I721222,I721239,I721256,I721287,I721304,I721349,I721366,I721383,I721414,I721440,I721448,I721479,I721496,I721513,I721539,I721547,I721564,I721653,I721679,I721696,I721704,I721749,I721766,I721783,I721800,I721817,I721834,I721851,I721882,I721899,I721944,I721961,I721978,I722009,I722035,I722043,I722074,I722091,I722108,I722134,I722142,I722159,I722248,I722274,I722291,I722299,I722344,I722361,I722378,I722395,I722412,I722429,I722446,I722477,I722494,I722539,I722556,I722573,I722604,I722630,I722638,I722669,I722686,I722703,I722729,I722737,I722754,I722843,I722869,I722886,I722894,I722939,I722956,I722973,I722990,I723007,I723024,I723041,I723072,I723089,I723134,I723151,I723168,I723199,I723225,I723233,I723264,I723281,I723298,I723324,I723332,I723349,I723438,I723464,I723481,I723489,I723534,I723551,I723568,I723585,I723602,I723619,I723636,I723667,I723684,I723729,I723746,I723763,I723794,I723820,I723828,I723859,I723876,I723893,I723919,I723927,I723944,I724033,I724059,I724076,I724084,I724129,I724146,I724163,I724180,I724197,I724214,I724231,I724262,I724279,I724324,I724341,I724358,I724389,I724415,I724423,I724454,I724471,I724488,I724514,I724522,I724539,I724628,I724654,I724671,I724679,I724724,I724741,I724758,I724775,I724792,I724809,I724826,I724857,I724874,I724919,I724936,I724953,I724984,I725010,I725018,I725049,I725066,I725083,I725109,I725117,I725134,I725223,I725249,I725266,I725274,I725319,I725336,I725353,I725370,I725387,I725404,I725421,I725452,I725469,I725514,I725531,I725548,I725579,I725605,I725613,I725644,I725661,I725678,I725704,I725712,I725729,I725818,I725844,I725861,I725869,I725914,I725931,I725948,I725965,I725982,I725999,I726016,I726047,I726064,I726109,I726126,I726143,I726174,I726200,I726208,I726239,I726256,I726273,I726299,I726307,I726324,I726413,I726439,I726456,I726464,I726509,I726526,I726543,I726560,I726577,I726594,I726611,I726642,I726659,I726704,I726721,I726738,I726769,I726795,I726803,I726834,I726851,I726868,I726894,I726902,I726919,I727008,I727034,I727051,I727059,I727104,I727121,I727138,I727155,I727172,I727189,I727206,I727237,I727254,I727299,I727316,I727333,I727364,I727390,I727398,I727429,I727446,I727463,I727489,I727497,I727514,I727603,I727629,I727646,I727654,I727699,I727716,I727733,I727750,I727767,I727784,I727801,I727832,I727849,I727894,I727911,I727928,I727959,I727985,I727993,I728024,I728041,I728058,I728084,I728092,I728109,I728198,I728224,I728241,I728249,I728294,I728311,I728328,I728345,I728362,I728379,I728396,I728427,I728444,I728489,I728506,I728523,I728554,I728580,I728588,I728619,I728636,I728653,I728679,I728687,I728704,I728793,I728819,I728836,I728844,I728889,I728906,I728923,I728940,I728957,I728974,I728991,I729022,I729039,I729084,I729101,I729118,I729149,I729175,I729183,I729214,I729231,I729248,I729274,I729282,I729299,I729388,I729414,I729431,I729439,I729484,I729501,I729518,I729535,I729552,I729569,I729586,I729617,I729634,I729679,I729696,I729713,I729744,I729770,I729778,I729809,I729826,I729843,I729869,I729877,I729894,I729983,I730009,I730026,I730034,I730079,I730096,I730113,I730130,I730147,I730164,I730181,I730212,I730229,I730274,I730291,I730308,I730339,I730365,I730373,I730404,I730421,I730438,I730464,I730472,I730489,I730578,I730604,I730621,I730629,I730674,I730691,I730708,I730725,I730742,I730759,I730776,I730807,I730824,I730869,I730886,I730903,I730934,I730960,I730968,I730999,I731016,I731033,I731059,I731067,I731084,I731173,I731199,I731216,I731224,I731269,I731286,I731303,I731320,I731337,I731354,I731371,I731402,I731419,I731464,I731481,I731498,I731529,I731555,I731563,I731594,I731611,I731628,I731654,I731662,I731679,I731768,I731794,I731811,I731819,I731864,I731881,I731898,I731915,I731932,I731949,I731966,I731997,I732014,I732059,I732076,I732093,I732124,I732150,I732158,I732189,I732206,I732223,I732249,I732257,I732274,I732363,I732389,I732406,I732414,I732459,I732476,I732493,I732510,I732527,I732544,I732561,I732592,I732609,I732654,I732671,I732688,I732719,I732745,I732753,I732784,I732801,I732818,I732844,I732852,I732869,I732958,I732984,I733001,I733009,I733054,I733071,I733088,I733105,I733122,I733139,I733156,I733187,I733204,I733249,I733266,I733283,I733314,I733340,I733348,I733379,I733396,I733413,I733439,I733447,I733464,I733553,I733579,I733596,I733604,I733649,I733666,I733683,I733700,I733717,I733734,I733751,I733782,I733799,I733844,I733861,I733878,I733909,I733935,I733943,I733974,I733991,I734008,I734034,I734042,I734059,I734148,I734174,I734191,I734199,I734244,I734261,I734278,I734295,I734312,I734329,I734346,I734377,I734394,I734439,I734456,I734473,I734504,I734530,I734538,I734569,I734586,I734603,I734629,I734637,I734654,I734743,I734769,I734786,I734794,I734839,I734856,I734873,I734890,I734907,I734924,I734941,I734972,I734989,I735034,I735051,I735068,I735099,I735125,I735133,I735164,I735181,I735198,I735224,I735232,I735249,I735338,I735364,I735381,I735389,I735434,I735451,I735468,I735485,I735502,I735519,I735536,I735567,I735584,I735629,I735646,I735663,I735694,I735720,I735728,I735759,I735776,I735793,I735819,I735827,I735844,I735933,I735959,I735976,I735984,I736029,I736046,I736063,I736080,I736097,I736114,I736131,I736162,I736179,I736224,I736241,I736258,I736289,I736315,I736323,I736354,I736371,I736388,I736414,I736422,I736439,I736528,I736554,I736571,I736579,I736624,I736641,I736658,I736675,I736692,I736709,I736726,I736757,I736774,I736819,I736836,I736853,I736884,I736910,I736918,I736949,I736966,I736983,I737009,I737017,I737034,I737123,I737149,I737166,I737174,I737219,I737236,I737253,I737270,I737287,I737304,I737321,I737352,I737369,I737414,I737431,I737448,I737479,I737505,I737513,I737544,I737561,I737578,I737604,I737612,I737629,I737718,I737744,I737761,I737769,I737814,I737831,I737848,I737865,I737882,I737899,I737916,I737947,I737964,I738009,I738026,I738043,I738074,I738100,I738108,I738139,I738156,I738173,I738199,I738207,I738224,I738313,I738339,I738356,I738364,I738409,I738426,I738443,I738460,I738477,I738494,I738511,I738542,I738559,I738604,I738621,I738638,I738669,I738695,I738703,I738734,I738751,I738768,I738794,I738802,I738819,I738908,I738934,I738951,I738959,I739004,I739021,I739038,I739055,I739072,I739089,I739106,I739137,I739154,I739199,I739216,I739233,I739264,I739290,I739298,I739329,I739346,I739363,I739389,I739397,I739414,I739503,I739529,I739546,I739554,I739599,I739616,I739633,I739650,I739667,I739684,I739701,I739732,I739749,I739794,I739811,I739828,I739859,I739885,I739893,I739924,I739941,I739958,I739984,I739992,I740009,I740098,I740124,I740141,I740149,I740194,I740211,I740228,I740245,I740262,I740279,I740296,I740327,I740344,I740389,I740406,I740423,I740454,I740480,I740488,I740519,I740536,I740553,I740579,I740587,I740604,I740693,I740719,I740736,I740744,I740789,I740806,I740823,I740840,I740857,I740874,I740891,I740922,I740939,I740984,I741001,I741018,I741049,I741075,I741083,I741114,I741131,I741148,I741174,I741182,I741199,I741288,I741314,I741331,I741339,I741384,I741401,I741418,I741435,I741452,I741469,I741486,I741517,I741534,I741579,I741596,I741613,I741644,I741670,I741678,I741709,I741726,I741743,I741769,I741777,I741794,I741883,I741909,I741926,I741934,I741979,I741996,I742013,I742030,I742047,I742064,I742081,I742112,I742129,I742174,I742191,I742208,I742239,I742265,I742273,I742304,I742321,I742338,I742364,I742372,I742389,I742478,I742504,I742521,I742529,I742574,I742591,I742608,I742625,I742642,I742659,I742676,I742707,I742724,I742769,I742786,I742803,I742834,I742860,I742868,I742899,I742916,I742933,I742959,I742967,I742984,I743073,I743099,I743116,I743124,I743169,I743186,I743203,I743220,I743237,I743254,I743271,I743302,I743319,I743364,I743381,I743398,I743429,I743455,I743463,I743494,I743511,I743528,I743554,I743562,I743579,I743668,I743694,I743711,I743719,I743764,I743781,I743798,I743815,I743832,I743849,I743866,I743897,I743914,I743959,I743976,I743993,I744024,I744050,I744058,I744089,I744106,I744123,I744149,I744157,I744174,I744263,I744289,I744306,I744314,I744359,I744376,I744393,I744410,I744427,I744444,I744461,I744492,I744509,I744554,I744571,I744588,I744619,I744645,I744653,I744684,I744701,I744718,I744744,I744752,I744769,I744858,I744884,I744901,I744909,I744954,I744971,I744988,I745005,I745022,I745039,I745056,I745087,I745104,I745149,I745166,I745183,I745214,I745240,I745248,I745279,I745296,I745313,I745339,I745347,I745364,I745453,I745479,I745496,I745504,I745549,I745566,I745583,I745600,I745617,I745634,I745651,I745682,I745699,I745744,I745761,I745778,I745809,I745835,I745843,I745874,I745891,I745908,I745934,I745942,I745959,I746048,I746074,I746091,I746099,I746144,I746161,I746178,I746195,I746212,I746229,I746246,I746277,I746294,I746339,I746356,I746373,I746404,I746430,I746438,I746469,I746486,I746503,I746529,I746537,I746554,I746643,I746669,I746686,I746694,I746739,I746756,I746773,I746790,I746807,I746824,I746841,I746872,I746889,I746934,I746951,I746968,I746999,I747025,I747033,I747064,I747081,I747098,I747124,I747132,I747149;
not I_0 (I3074,I3042);
DFFARX1 I_1 (I213027,I3035,I3074,I3100,);
nand I_2 (I3108,I3100,I213018);
not I_3 (I3125,I3108);
DFFARX1 I_4 (I3125,I3035,I3074,I3066,);
DFFARX1 I_5 (I213021,I3035,I3074,I3165,);
not I_6 (I3173,I3165);
not I_7 (I3190,I213015);
not I_8 (I3207,I213024);
nand I_9 (I3224,I3173,I3207);
nor I_10 (I3241,I3224,I213015);
DFFARX1 I_11 (I3241,I3035,I3074,I3045,);
nor I_12 (I3272,I213024,I213015);
nand I_13 (I3289,I3165,I3272);
nor I_14 (I3306,I213012,I213030);
nor I_15 (I3048,I3224,I213012);
not I_16 (I3337,I213012);
not I_17 (I3354,I213012);
nand I_18 (I3371,I3354,I213036);
nand I_19 (I3388,I3190,I3371);
not I_20 (I3405,I3388);
nor I_21 (I3422,I213012,I213030);
nor I_22 (I3057,I3405,I3422);
nor I_23 (I3453,I213033,I213012);
and I_24 (I3470,I3453,I3306);
nor I_25 (I3487,I3388,I3470);
DFFARX1 I_26 (I3487,I3035,I3074,I3063,);
nor I_27 (I3518,I3108,I3470);
DFFARX1 I_28 (I3518,I3035,I3074,I3060,);
nor I_29 (I3549,I213033,I213039);
DFFARX1 I_30 (I3549,I3035,I3074,I3575,);
nor I_31 (I3583,I3575,I213024);
nand I_32 (I3600,I3583,I3190);
nand I_33 (I3054,I3600,I3289);
nand I_34 (I3051,I3583,I3337);
not I_35 (I3669,I3042);
DFFARX1 I_36 (I116387,I3035,I3669,I3695,);
nand I_37 (I3703,I3695,I116387);
not I_38 (I3720,I3703);
DFFARX1 I_39 (I3720,I3035,I3669,I3661,);
DFFARX1 I_40 (I116393,I3035,I3669,I3760,);
not I_41 (I3768,I3760);
not I_42 (I3785,I116402);
not I_43 (I3802,I116396);
nand I_44 (I3819,I3768,I3802);
nor I_45 (I3836,I3819,I116402);
DFFARX1 I_46 (I3836,I3035,I3669,I3640,);
nor I_47 (I3867,I116396,I116402);
nand I_48 (I3884,I3760,I3867);
nor I_49 (I3901,I116399,I116405);
nor I_50 (I3643,I3819,I116399);
not I_51 (I3932,I116399);
not I_52 (I3949,I116408);
nand I_53 (I3966,I3949,I116384);
nand I_54 (I3983,I3785,I3966);
not I_55 (I4000,I3983);
nor I_56 (I4017,I116408,I116405);
nor I_57 (I3652,I4000,I4017);
nor I_58 (I4048,I116390,I116408);
and I_59 (I4065,I4048,I3901);
nor I_60 (I4082,I3983,I4065);
DFFARX1 I_61 (I4082,I3035,I3669,I3658,);
nor I_62 (I4113,I3703,I4065);
DFFARX1 I_63 (I4113,I3035,I3669,I3655,);
nor I_64 (I4144,I116390,I116384);
DFFARX1 I_65 (I4144,I3035,I3669,I4170,);
nor I_66 (I4178,I4170,I116396);
nand I_67 (I4195,I4178,I3785);
nand I_68 (I3649,I4195,I3884);
nand I_69 (I3646,I4178,I3932);
not I_70 (I4264,I3042);
DFFARX1 I_71 (I731153,I3035,I4264,I4290,);
nand I_72 (I4298,I4290,I731144);
not I_73 (I4315,I4298);
DFFARX1 I_74 (I4315,I3035,I4264,I4256,);
DFFARX1 I_75 (I731147,I3035,I4264,I4355,);
not I_76 (I4363,I4355);
not I_77 (I4380,I731159);
not I_78 (I4397,I731150);
nand I_79 (I4414,I4363,I4397);
nor I_80 (I4431,I4414,I731159);
DFFARX1 I_81 (I4431,I3035,I4264,I4235,);
nor I_82 (I4462,I731150,I731159);
nand I_83 (I4479,I4355,I4462);
nor I_84 (I4496,I731138,I731138);
nor I_85 (I4238,I4414,I731138);
not I_86 (I4527,I731138);
not I_87 (I4544,I731162);
nand I_88 (I4561,I4544,I731141);
nand I_89 (I4578,I4380,I4561);
not I_90 (I4595,I4578);
nor I_91 (I4612,I731162,I731138);
nor I_92 (I4247,I4595,I4612);
nor I_93 (I4643,I731156,I731162);
and I_94 (I4660,I4643,I4496);
nor I_95 (I4677,I4578,I4660);
DFFARX1 I_96 (I4677,I3035,I4264,I4253,);
nor I_97 (I4708,I4298,I4660);
DFFARX1 I_98 (I4708,I3035,I4264,I4250,);
nor I_99 (I4739,I731156,I731165);
DFFARX1 I_100 (I4739,I3035,I4264,I4765,);
nor I_101 (I4773,I4765,I731150);
nand I_102 (I4790,I4773,I4380);
nand I_103 (I4244,I4790,I4479);
nand I_104 (I4241,I4773,I4527);
not I_105 (I4859,I3042);
DFFARX1 I_106 (I270714,I3035,I4859,I4885,);
nand I_107 (I4893,I4885,I270696);
not I_108 (I4910,I4893);
DFFARX1 I_109 (I4910,I3035,I4859,I4851,);
DFFARX1 I_110 (I270708,I3035,I4859,I4950,);
not I_111 (I4958,I4950);
not I_112 (I4975,I270693);
not I_113 (I4992,I270702);
nand I_114 (I5009,I4958,I4992);
nor I_115 (I5026,I5009,I270693);
DFFARX1 I_116 (I5026,I3035,I4859,I4830,);
nor I_117 (I5057,I270702,I270693);
nand I_118 (I5074,I4950,I5057);
nor I_119 (I5091,I270699,I270720);
nor I_120 (I4833,I5009,I270699);
not I_121 (I5122,I270699);
not I_122 (I5139,I270711);
nand I_123 (I5156,I5139,I270717);
nand I_124 (I5173,I4975,I5156);
not I_125 (I5190,I5173);
nor I_126 (I5207,I270711,I270720);
nor I_127 (I4842,I5190,I5207);
nor I_128 (I5238,I270693,I270711);
and I_129 (I5255,I5238,I5091);
nor I_130 (I5272,I5173,I5255);
DFFARX1 I_131 (I5272,I3035,I4859,I4848,);
nor I_132 (I5303,I4893,I5255);
DFFARX1 I_133 (I5303,I3035,I4859,I4845,);
nor I_134 (I5334,I270693,I270705);
DFFARX1 I_135 (I5334,I3035,I4859,I5360,);
nor I_136 (I5368,I5360,I270702);
nand I_137 (I5385,I5368,I4975);
nand I_138 (I4839,I5385,I5074);
nand I_139 (I4836,I5368,I5122);
not I_140 (I5454,I3042);
DFFARX1 I_141 (I639919,I3035,I5454,I5480,);
nand I_142 (I5488,I5480,I639919);
not I_143 (I5505,I5488);
DFFARX1 I_144 (I5505,I3035,I5454,I5446,);
DFFARX1 I_145 (I639934,I3035,I5454,I5545,);
not I_146 (I5553,I5545);
not I_147 (I5570,I639931);
not I_148 (I5587,I639940);
nand I_149 (I5604,I5553,I5587);
nor I_150 (I5621,I5604,I639931);
DFFARX1 I_151 (I5621,I3035,I5454,I5425,);
nor I_152 (I5652,I639940,I639931);
nand I_153 (I5669,I5545,I5652);
nor I_154 (I5686,I639928,I639937);
nor I_155 (I5428,I5604,I639928);
not I_156 (I5717,I639928);
not I_157 (I5734,I639925);
nand I_158 (I5751,I5734,I639916);
nand I_159 (I5768,I5570,I5751);
not I_160 (I5785,I5768);
nor I_161 (I5802,I639925,I639937);
nor I_162 (I5437,I5785,I5802);
nor I_163 (I5833,I639922,I639925);
and I_164 (I5850,I5833,I5686);
nor I_165 (I5867,I5768,I5850);
DFFARX1 I_166 (I5867,I3035,I5454,I5443,);
nor I_167 (I5898,I5488,I5850);
DFFARX1 I_168 (I5898,I3035,I5454,I5440,);
nor I_169 (I5929,I639922,I639916);
DFFARX1 I_170 (I5929,I3035,I5454,I5955,);
nor I_171 (I5963,I5955,I639940);
nand I_172 (I5980,I5963,I5570);
nand I_173 (I5434,I5980,I5669);
nand I_174 (I5431,I5963,I5717);
not I_175 (I6049,I3042);
DFFARX1 I_176 (I393814,I3035,I6049,I6075,);
nand I_177 (I6083,I6075,I393793);
not I_178 (I6100,I6083);
DFFARX1 I_179 (I6100,I3035,I6049,I6041,);
DFFARX1 I_180 (I393802,I3035,I6049,I6140,);
not I_181 (I6148,I6140);
not I_182 (I6165,I393808);
not I_183 (I6182,I393805);
nand I_184 (I6199,I6148,I6182);
nor I_185 (I6216,I6199,I393808);
DFFARX1 I_186 (I6216,I3035,I6049,I6020,);
nor I_187 (I6247,I393805,I393808);
nand I_188 (I6264,I6140,I6247);
nor I_189 (I6281,I393796,I393790);
nor I_190 (I6023,I6199,I393796);
not I_191 (I6312,I393796);
not I_192 (I6329,I393811);
nand I_193 (I6346,I6329,I393793);
nand I_194 (I6363,I6165,I6346);
not I_195 (I6380,I6363);
nor I_196 (I6397,I393811,I393790);
nor I_197 (I6032,I6380,I6397);
nor I_198 (I6428,I393799,I393811);
and I_199 (I6445,I6428,I6281);
nor I_200 (I6462,I6363,I6445);
DFFARX1 I_201 (I6462,I3035,I6049,I6038,);
nor I_202 (I6493,I6083,I6445);
DFFARX1 I_203 (I6493,I3035,I6049,I6035,);
nor I_204 (I6524,I393799,I393790);
DFFARX1 I_205 (I6524,I3035,I6049,I6550,);
nor I_206 (I6558,I6550,I393805);
nand I_207 (I6575,I6558,I6165);
nand I_208 (I6029,I6575,I6264);
nand I_209 (I6026,I6558,I6312);
not I_210 (I6644,I3042);
DFFARX1 I_211 (I572293,I3035,I6644,I6670,);
nand I_212 (I6678,I6670,I572293);
not I_213 (I6695,I6678);
DFFARX1 I_214 (I6695,I3035,I6644,I6636,);
DFFARX1 I_215 (I572308,I3035,I6644,I6735,);
not I_216 (I6743,I6735);
not I_217 (I6760,I572305);
not I_218 (I6777,I572314);
nand I_219 (I6794,I6743,I6777);
nor I_220 (I6811,I6794,I572305);
DFFARX1 I_221 (I6811,I3035,I6644,I6615,);
nor I_222 (I6842,I572314,I572305);
nand I_223 (I6859,I6735,I6842);
nor I_224 (I6876,I572302,I572311);
nor I_225 (I6618,I6794,I572302);
not I_226 (I6907,I572302);
not I_227 (I6924,I572299);
nand I_228 (I6941,I6924,I572290);
nand I_229 (I6958,I6760,I6941);
not I_230 (I6975,I6958);
nor I_231 (I6992,I572299,I572311);
nor I_232 (I6627,I6975,I6992);
nor I_233 (I7023,I572296,I572299);
and I_234 (I7040,I7023,I6876);
nor I_235 (I7057,I6958,I7040);
DFFARX1 I_236 (I7057,I3035,I6644,I6633,);
nor I_237 (I7088,I6678,I7040);
DFFARX1 I_238 (I7088,I3035,I6644,I6630,);
nor I_239 (I7119,I572296,I572290);
DFFARX1 I_240 (I7119,I3035,I6644,I7145,);
nor I_241 (I7153,I7145,I572314);
nand I_242 (I7170,I7153,I6760);
nand I_243 (I6624,I7170,I6859);
nand I_244 (I6621,I7153,I6907);
not I_245 (I7239,I3042);
DFFARX1 I_246 (I429295,I3035,I7239,I7265,);
nand I_247 (I7273,I7265,I429286);
not I_248 (I7290,I7273);
DFFARX1 I_249 (I7290,I3035,I7239,I7231,);
DFFARX1 I_250 (I429292,I3035,I7239,I7330,);
not I_251 (I7338,I7330);
not I_252 (I7355,I429286);
not I_253 (I7372,I429298);
nand I_254 (I7389,I7338,I7372);
nor I_255 (I7406,I7389,I429286);
DFFARX1 I_256 (I7406,I3035,I7239,I7210,);
nor I_257 (I7437,I429298,I429286);
nand I_258 (I7454,I7330,I7437);
nor I_259 (I7471,I429307,I429304);
nor I_260 (I7213,I7389,I429307);
not I_261 (I7502,I429307);
not I_262 (I7519,I429292);
nand I_263 (I7536,I7519,I429289);
nand I_264 (I7553,I7355,I7536);
not I_265 (I7570,I7553);
nor I_266 (I7587,I429292,I429304);
nor I_267 (I7222,I7570,I7587);
nor I_268 (I7618,I429289,I429292);
and I_269 (I7635,I7618,I7471);
nor I_270 (I7652,I7553,I7635);
DFFARX1 I_271 (I7652,I3035,I7239,I7228,);
nor I_272 (I7683,I7273,I7635);
DFFARX1 I_273 (I7683,I3035,I7239,I7225,);
nor I_274 (I7714,I429289,I429301);
DFFARX1 I_275 (I7714,I3035,I7239,I7740,);
nor I_276 (I7748,I7740,I429298);
nand I_277 (I7765,I7748,I7355);
nand I_278 (I7219,I7765,I7454);
nand I_279 (I7216,I7748,I7502);
not I_280 (I7837,I3042);
DFFARX1 I_281 (I118770,I3035,I7837,I7863,);
DFFARX1 I_282 (I7863,I3035,I7837,I7880,);
not I_283 (I7888,I7880);
nand I_284 (I7905,I118788,I118773);
and I_285 (I7922,I7905,I118776);
DFFARX1 I_286 (I7922,I3035,I7837,I7948,);
DFFARX1 I_287 (I7948,I3035,I7837,I7829,);
DFFARX1 I_288 (I7948,I3035,I7837,I7820,);
DFFARX1 I_289 (I118764,I3035,I7837,I7993,);
nand I_290 (I8001,I7993,I118767);
not I_291 (I8018,I8001);
nor I_292 (I7817,I7863,I8018);
DFFARX1 I_293 (I118779,I3035,I7837,I8058,);
not I_294 (I8066,I8058);
nor I_295 (I7823,I8066,I7888);
nand I_296 (I7811,I8066,I8001);
nand I_297 (I8111,I118785,I118782);
and I_298 (I8128,I8111,I118767);
DFFARX1 I_299 (I8128,I3035,I7837,I8154,);
nor I_300 (I8162,I8154,I7863);
DFFARX1 I_301 (I8162,I3035,I7837,I7805,);
not I_302 (I8193,I8154);
nor I_303 (I8210,I118764,I118782);
not I_304 (I8227,I8210);
nor I_305 (I8244,I8001,I8227);
nor I_306 (I8261,I8193,I8244);
DFFARX1 I_307 (I8261,I3035,I7837,I7826,);
nor I_308 (I8292,I8154,I8227);
nor I_309 (I7814,I8018,I8292);
nor I_310 (I7808,I8154,I8210);
not I_311 (I8364,I3042);
DFFARX1 I_312 (I74210,I3035,I8364,I8390,);
DFFARX1 I_313 (I8390,I3035,I8364,I8407,);
not I_314 (I8415,I8407);
nand I_315 (I8432,I74210,I74225);
and I_316 (I8449,I8432,I74228);
DFFARX1 I_317 (I8449,I3035,I8364,I8475,);
DFFARX1 I_318 (I8475,I3035,I8364,I8356,);
DFFARX1 I_319 (I8475,I3035,I8364,I8347,);
DFFARX1 I_320 (I74222,I3035,I8364,I8520,);
nand I_321 (I8528,I8520,I74231);
not I_322 (I8545,I8528);
nor I_323 (I8344,I8390,I8545);
DFFARX1 I_324 (I74207,I3035,I8364,I8585,);
not I_325 (I8593,I8585);
nor I_326 (I8350,I8593,I8415);
nand I_327 (I8338,I8593,I8528);
nand I_328 (I8638,I74207,I74213);
and I_329 (I8655,I8638,I74216);
DFFARX1 I_330 (I8655,I3035,I8364,I8681,);
nor I_331 (I8689,I8681,I8390);
DFFARX1 I_332 (I8689,I3035,I8364,I8332,);
not I_333 (I8720,I8681);
nor I_334 (I8737,I74219,I74213);
not I_335 (I8754,I8737);
nor I_336 (I8771,I8528,I8754);
nor I_337 (I8788,I8720,I8771);
DFFARX1 I_338 (I8788,I3035,I8364,I8353,);
nor I_339 (I8819,I8681,I8754);
nor I_340 (I8341,I8545,I8819);
nor I_341 (I8335,I8681,I8737);
not I_342 (I8891,I3042);
DFFARX1 I_343 (I137810,I3035,I8891,I8917,);
DFFARX1 I_344 (I8917,I3035,I8891,I8934,);
not I_345 (I8942,I8934);
nand I_346 (I8959,I137828,I137813);
and I_347 (I8976,I8959,I137816);
DFFARX1 I_348 (I8976,I3035,I8891,I9002,);
DFFARX1 I_349 (I9002,I3035,I8891,I8883,);
DFFARX1 I_350 (I9002,I3035,I8891,I8874,);
DFFARX1 I_351 (I137804,I3035,I8891,I9047,);
nand I_352 (I9055,I9047,I137807);
not I_353 (I9072,I9055);
nor I_354 (I8871,I8917,I9072);
DFFARX1 I_355 (I137819,I3035,I8891,I9112,);
not I_356 (I9120,I9112);
nor I_357 (I8877,I9120,I8942);
nand I_358 (I8865,I9120,I9055);
nand I_359 (I9165,I137825,I137822);
and I_360 (I9182,I9165,I137807);
DFFARX1 I_361 (I9182,I3035,I8891,I9208,);
nor I_362 (I9216,I9208,I8917);
DFFARX1 I_363 (I9216,I3035,I8891,I8859,);
not I_364 (I9247,I9208);
nor I_365 (I9264,I137804,I137822);
not I_366 (I9281,I9264);
nor I_367 (I9298,I9055,I9281);
nor I_368 (I9315,I9247,I9298);
DFFARX1 I_369 (I9315,I3035,I8891,I8880,);
nor I_370 (I9346,I9208,I9281);
nor I_371 (I8868,I9072,I9346);
nor I_372 (I8862,I9208,I9264);
not I_373 (I9418,I3042);
DFFARX1 I_374 (I459861,I3035,I9418,I9444,);
DFFARX1 I_375 (I9444,I3035,I9418,I9461,);
not I_376 (I9469,I9461);
nand I_377 (I9486,I459852,I459873);
and I_378 (I9503,I9486,I459855);
DFFARX1 I_379 (I9503,I3035,I9418,I9529,);
DFFARX1 I_380 (I9529,I3035,I9418,I9410,);
DFFARX1 I_381 (I9529,I3035,I9418,I9401,);
DFFARX1 I_382 (I459855,I3035,I9418,I9574,);
nand I_383 (I9582,I9574,I459870);
not I_384 (I9599,I9582);
nor I_385 (I9398,I9444,I9599);
DFFARX1 I_386 (I459864,I3035,I9418,I9639,);
not I_387 (I9647,I9639);
nor I_388 (I9404,I9647,I9469);
nand I_389 (I9392,I9647,I9582);
nand I_390 (I9692,I459858,I459867);
and I_391 (I9709,I9692,I459852);
DFFARX1 I_392 (I9709,I3035,I9418,I9735,);
nor I_393 (I9743,I9735,I9444);
DFFARX1 I_394 (I9743,I3035,I9418,I9386,);
not I_395 (I9774,I9735);
nor I_396 (I9791,I459858,I459867);
not I_397 (I9808,I9791);
nor I_398 (I9825,I9582,I9808);
nor I_399 (I9842,I9774,I9825);
DFFARX1 I_400 (I9842,I3035,I9418,I9407,);
nor I_401 (I9873,I9735,I9808);
nor I_402 (I9395,I9599,I9873);
nor I_403 (I9389,I9735,I9791);
not I_404 (I9945,I3042);
DFFARX1 I_405 (I436146,I3035,I9945,I9971,);
DFFARX1 I_406 (I9971,I3035,I9945,I9988,);
not I_407 (I9996,I9988);
nand I_408 (I10013,I436137,I436158);
and I_409 (I10030,I10013,I436140);
DFFARX1 I_410 (I10030,I3035,I9945,I10056,);
DFFARX1 I_411 (I10056,I3035,I9945,I9937,);
DFFARX1 I_412 (I10056,I3035,I9945,I9928,);
DFFARX1 I_413 (I436140,I3035,I9945,I10101,);
nand I_414 (I10109,I10101,I436155);
not I_415 (I10126,I10109);
nor I_416 (I9925,I9971,I10126);
DFFARX1 I_417 (I436149,I3035,I9945,I10166,);
not I_418 (I10174,I10166);
nor I_419 (I9931,I10174,I9996);
nand I_420 (I9919,I10174,I10109);
nand I_421 (I10219,I436143,I436152);
and I_422 (I10236,I10219,I436137);
DFFARX1 I_423 (I10236,I3035,I9945,I10262,);
nor I_424 (I10270,I10262,I9971);
DFFARX1 I_425 (I10270,I3035,I9945,I9913,);
not I_426 (I10301,I10262);
nor I_427 (I10318,I436143,I436152);
not I_428 (I10335,I10318);
nor I_429 (I10352,I10109,I10335);
nor I_430 (I10369,I10301,I10352);
DFFARX1 I_431 (I10369,I3035,I9945,I9934,);
nor I_432 (I10400,I10262,I10335);
nor I_433 (I9922,I10126,I10400);
nor I_434 (I9916,I10262,I10318);
not I_435 (I10472,I3042);
DFFARX1 I_436 (I121745,I3035,I10472,I10498,);
DFFARX1 I_437 (I10498,I3035,I10472,I10515,);
not I_438 (I10523,I10515);
nand I_439 (I10540,I121763,I121748);
and I_440 (I10557,I10540,I121751);
DFFARX1 I_441 (I10557,I3035,I10472,I10583,);
DFFARX1 I_442 (I10583,I3035,I10472,I10464,);
DFFARX1 I_443 (I10583,I3035,I10472,I10455,);
DFFARX1 I_444 (I121739,I3035,I10472,I10628,);
nand I_445 (I10636,I10628,I121742);
not I_446 (I10653,I10636);
nor I_447 (I10452,I10498,I10653);
DFFARX1 I_448 (I121754,I3035,I10472,I10693,);
not I_449 (I10701,I10693);
nor I_450 (I10458,I10701,I10523);
nand I_451 (I10446,I10701,I10636);
nand I_452 (I10746,I121760,I121757);
and I_453 (I10763,I10746,I121742);
DFFARX1 I_454 (I10763,I3035,I10472,I10789,);
nor I_455 (I10797,I10789,I10498);
DFFARX1 I_456 (I10797,I3035,I10472,I10440,);
not I_457 (I10828,I10789);
nor I_458 (I10845,I121739,I121757);
not I_459 (I10862,I10845);
nor I_460 (I10879,I10636,I10862);
nor I_461 (I10896,I10828,I10879);
DFFARX1 I_462 (I10896,I3035,I10472,I10461,);
nor I_463 (I10927,I10789,I10862);
nor I_464 (I10449,I10653,I10927);
nor I_465 (I10443,I10789,I10845);
not I_466 (I10999,I3042);
DFFARX1 I_467 (I705553,I3035,I10999,I11025,);
DFFARX1 I_468 (I11025,I3035,I10999,I11042,);
not I_469 (I11050,I11042);
nand I_470 (I11067,I705556,I705562);
and I_471 (I11084,I11067,I705571);
DFFARX1 I_472 (I11084,I3035,I10999,I11110,);
DFFARX1 I_473 (I11110,I3035,I10999,I10991,);
DFFARX1 I_474 (I11110,I3035,I10999,I10982,);
DFFARX1 I_475 (I705574,I3035,I10999,I11155,);
nand I_476 (I11163,I11155,I705565);
not I_477 (I11180,I11163);
nor I_478 (I10979,I11025,I11180);
DFFARX1 I_479 (I705553,I3035,I10999,I11220,);
not I_480 (I11228,I11220);
nor I_481 (I10985,I11228,I11050);
nand I_482 (I10973,I11228,I11163);
nand I_483 (I11273,I705580,I705559);
and I_484 (I11290,I11273,I705568);
DFFARX1 I_485 (I11290,I3035,I10999,I11316,);
nor I_486 (I11324,I11316,I11025);
DFFARX1 I_487 (I11324,I3035,I10999,I10967,);
not I_488 (I11355,I11316);
nor I_489 (I11372,I705577,I705559);
not I_490 (I11389,I11372);
nor I_491 (I11406,I11163,I11389);
nor I_492 (I11423,I11355,I11406);
DFFARX1 I_493 (I11423,I3035,I10999,I10988,);
nor I_494 (I11454,I11316,I11389);
nor I_495 (I10976,I11180,I11454);
nor I_496 (I10970,I11316,I11372);
not I_497 (I11526,I3042);
DFFARX1 I_498 (I703768,I3035,I11526,I11552,);
DFFARX1 I_499 (I11552,I3035,I11526,I11569,);
not I_500 (I11577,I11569);
nand I_501 (I11594,I703771,I703777);
and I_502 (I11611,I11594,I703786);
DFFARX1 I_503 (I11611,I3035,I11526,I11637,);
DFFARX1 I_504 (I11637,I3035,I11526,I11518,);
DFFARX1 I_505 (I11637,I3035,I11526,I11509,);
DFFARX1 I_506 (I703789,I3035,I11526,I11682,);
nand I_507 (I11690,I11682,I703780);
not I_508 (I11707,I11690);
nor I_509 (I11506,I11552,I11707);
DFFARX1 I_510 (I703768,I3035,I11526,I11747,);
not I_511 (I11755,I11747);
nor I_512 (I11512,I11755,I11577);
nand I_513 (I11500,I11755,I11690);
nand I_514 (I11800,I703795,I703774);
and I_515 (I11817,I11800,I703783);
DFFARX1 I_516 (I11817,I3035,I11526,I11843,);
nor I_517 (I11851,I11843,I11552);
DFFARX1 I_518 (I11851,I3035,I11526,I11494,);
not I_519 (I11882,I11843);
nor I_520 (I11899,I703792,I703774);
not I_521 (I11916,I11899);
nor I_522 (I11933,I11690,I11916);
nor I_523 (I11950,I11882,I11933);
DFFARX1 I_524 (I11950,I3035,I11526,I11515,);
nor I_525 (I11981,I11843,I11916);
nor I_526 (I11503,I11707,I11981);
nor I_527 (I11497,I11843,I11899);
not I_528 (I12053,I3042);
DFFARX1 I_529 (I119365,I3035,I12053,I12079,);
DFFARX1 I_530 (I12079,I3035,I12053,I12096,);
not I_531 (I12104,I12096);
nand I_532 (I12121,I119383,I119368);
and I_533 (I12138,I12121,I119371);
DFFARX1 I_534 (I12138,I3035,I12053,I12164,);
DFFARX1 I_535 (I12164,I3035,I12053,I12045,);
DFFARX1 I_536 (I12164,I3035,I12053,I12036,);
DFFARX1 I_537 (I119359,I3035,I12053,I12209,);
nand I_538 (I12217,I12209,I119362);
not I_539 (I12234,I12217);
nor I_540 (I12033,I12079,I12234);
DFFARX1 I_541 (I119374,I3035,I12053,I12274,);
not I_542 (I12282,I12274);
nor I_543 (I12039,I12282,I12104);
nand I_544 (I12027,I12282,I12217);
nand I_545 (I12327,I119380,I119377);
and I_546 (I12344,I12327,I119362);
DFFARX1 I_547 (I12344,I3035,I12053,I12370,);
nor I_548 (I12378,I12370,I12079);
DFFARX1 I_549 (I12378,I3035,I12053,I12021,);
not I_550 (I12409,I12370);
nor I_551 (I12426,I119359,I119377);
not I_552 (I12443,I12426);
nor I_553 (I12460,I12217,I12443);
nor I_554 (I12477,I12409,I12460);
DFFARX1 I_555 (I12477,I3035,I12053,I12042,);
nor I_556 (I12508,I12370,I12443);
nor I_557 (I12030,I12234,I12508);
nor I_558 (I12024,I12370,I12426);
not I_559 (I12580,I3042);
DFFARX1 I_560 (I616242,I3035,I12580,I12606,);
DFFARX1 I_561 (I12606,I3035,I12580,I12623,);
not I_562 (I12631,I12623);
nand I_563 (I12648,I616230,I616221);
and I_564 (I12665,I12648,I616218);
DFFARX1 I_565 (I12665,I3035,I12580,I12691,);
DFFARX1 I_566 (I12691,I3035,I12580,I12572,);
DFFARX1 I_567 (I12691,I3035,I12580,I12563,);
DFFARX1 I_568 (I616224,I3035,I12580,I12736,);
nand I_569 (I12744,I12736,I616236);
not I_570 (I12761,I12744);
nor I_571 (I12560,I12606,I12761);
DFFARX1 I_572 (I616233,I3035,I12580,I12801,);
not I_573 (I12809,I12801);
nor I_574 (I12566,I12809,I12631);
nand I_575 (I12554,I12809,I12744);
nand I_576 (I12854,I616227,I616221);
and I_577 (I12871,I12854,I616239);
DFFARX1 I_578 (I12871,I3035,I12580,I12897,);
nor I_579 (I12905,I12897,I12606);
DFFARX1 I_580 (I12905,I3035,I12580,I12548,);
not I_581 (I12936,I12897);
nor I_582 (I12953,I616218,I616221);
not I_583 (I12970,I12953);
nor I_584 (I12987,I12744,I12970);
nor I_585 (I13004,I12936,I12987);
DFFARX1 I_586 (I13004,I3035,I12580,I12569,);
nor I_587 (I13035,I12897,I12970);
nor I_588 (I12557,I12761,I13035);
nor I_589 (I12551,I12897,I12953);
not I_590 (I13107,I3042);
DFFARX1 I_591 (I734708,I3035,I13107,I13133,);
DFFARX1 I_592 (I13133,I3035,I13107,I13150,);
not I_593 (I13158,I13150);
nand I_594 (I13175,I734711,I734717);
and I_595 (I13192,I13175,I734726);
DFFARX1 I_596 (I13192,I3035,I13107,I13218,);
DFFARX1 I_597 (I13218,I3035,I13107,I13099,);
DFFARX1 I_598 (I13218,I3035,I13107,I13090,);
DFFARX1 I_599 (I734729,I3035,I13107,I13263,);
nand I_600 (I13271,I13263,I734720);
not I_601 (I13288,I13271);
nor I_602 (I13087,I13133,I13288);
DFFARX1 I_603 (I734708,I3035,I13107,I13328,);
not I_604 (I13336,I13328);
nor I_605 (I13093,I13336,I13158);
nand I_606 (I13081,I13336,I13271);
nand I_607 (I13381,I734735,I734714);
and I_608 (I13398,I13381,I734723);
DFFARX1 I_609 (I13398,I3035,I13107,I13424,);
nor I_610 (I13432,I13424,I13133);
DFFARX1 I_611 (I13432,I3035,I13107,I13075,);
not I_612 (I13463,I13424);
nor I_613 (I13480,I734732,I734714);
not I_614 (I13497,I13480);
nor I_615 (I13514,I13271,I13497);
nor I_616 (I13531,I13463,I13514);
DFFARX1 I_617 (I13531,I3035,I13107,I13096,);
nor I_618 (I13562,I13424,I13497);
nor I_619 (I13084,I13288,I13562);
nor I_620 (I13078,I13424,I13480);
not I_621 (I13634,I3042);
DFFARX1 I_622 (I406512,I3035,I13634,I13660,);
DFFARX1 I_623 (I13660,I3035,I13634,I13677,);
not I_624 (I13685,I13677);
nand I_625 (I13702,I406527,I406530);
and I_626 (I13719,I13702,I406509);
DFFARX1 I_627 (I13719,I3035,I13634,I13745,);
DFFARX1 I_628 (I13745,I3035,I13634,I13626,);
DFFARX1 I_629 (I13745,I3035,I13634,I13617,);
DFFARX1 I_630 (I406515,I3035,I13634,I13790,);
nand I_631 (I13798,I13790,I406521);
not I_632 (I13815,I13798);
nor I_633 (I13614,I13660,I13815);
DFFARX1 I_634 (I406509,I3035,I13634,I13855,);
not I_635 (I13863,I13855);
nor I_636 (I13620,I13863,I13685);
nand I_637 (I13608,I13863,I13798);
nand I_638 (I13908,I406524,I406506);
and I_639 (I13925,I13908,I406518);
DFFARX1 I_640 (I13925,I3035,I13634,I13951,);
nor I_641 (I13959,I13951,I13660);
DFFARX1 I_642 (I13959,I3035,I13634,I13602,);
not I_643 (I13990,I13951);
nor I_644 (I14007,I406506,I406506);
not I_645 (I14024,I14007);
nor I_646 (I14041,I13798,I14024);
nor I_647 (I14058,I13990,I14041);
DFFARX1 I_648 (I14058,I3035,I13634,I13623,);
nor I_649 (I14089,I13951,I14024);
nor I_650 (I13611,I13815,I14089);
nor I_651 (I13605,I13951,I14007);
not I_652 (I14161,I3042);
DFFARX1 I_653 (I261989,I3035,I14161,I14187,);
DFFARX1 I_654 (I14187,I3035,I14161,I14204,);
not I_655 (I14212,I14204);
nand I_656 (I14229,I261989,I261992);
and I_657 (I14246,I14229,I262013);
DFFARX1 I_658 (I14246,I3035,I14161,I14272,);
DFFARX1 I_659 (I14272,I3035,I14161,I14153,);
DFFARX1 I_660 (I14272,I3035,I14161,I14144,);
DFFARX1 I_661 (I262001,I3035,I14161,I14317,);
nand I_662 (I14325,I14317,I262004);
not I_663 (I14342,I14325);
nor I_664 (I14141,I14187,I14342);
DFFARX1 I_665 (I262010,I3035,I14161,I14382,);
not I_666 (I14390,I14382);
nor I_667 (I14147,I14390,I14212);
nand I_668 (I14135,I14390,I14325);
nand I_669 (I14435,I262007,I261995);
and I_670 (I14452,I14435,I261998);
DFFARX1 I_671 (I14452,I3035,I14161,I14478,);
nor I_672 (I14486,I14478,I14187);
DFFARX1 I_673 (I14486,I3035,I14161,I14129,);
not I_674 (I14517,I14478);
nor I_675 (I14534,I262016,I261995);
not I_676 (I14551,I14534);
nor I_677 (I14568,I14325,I14551);
nor I_678 (I14585,I14517,I14568);
DFFARX1 I_679 (I14585,I3035,I14161,I14150,);
nor I_680 (I14616,I14478,I14551);
nor I_681 (I14138,I14342,I14616);
nor I_682 (I14132,I14478,I14534);
not I_683 (I14688,I3042);
DFFARX1 I_684 (I511624,I3035,I14688,I14714,);
DFFARX1 I_685 (I14714,I3035,I14688,I14731,);
not I_686 (I14739,I14731);
nand I_687 (I14756,I511600,I511627);
and I_688 (I14773,I14756,I511612);
DFFARX1 I_689 (I14773,I3035,I14688,I14799,);
DFFARX1 I_690 (I14799,I3035,I14688,I14680,);
DFFARX1 I_691 (I14799,I3035,I14688,I14671,);
DFFARX1 I_692 (I511618,I3035,I14688,I14844,);
nand I_693 (I14852,I14844,I511603);
not I_694 (I14869,I14852);
nor I_695 (I14668,I14714,I14869);
DFFARX1 I_696 (I511621,I3035,I14688,I14909,);
not I_697 (I14917,I14909);
nor I_698 (I14674,I14917,I14739);
nand I_699 (I14662,I14917,I14852);
nand I_700 (I14962,I511606,I511609);
and I_701 (I14979,I14962,I511600);
DFFARX1 I_702 (I14979,I3035,I14688,I15005,);
nor I_703 (I15013,I15005,I14714);
DFFARX1 I_704 (I15013,I3035,I14688,I14656,);
not I_705 (I15044,I15005);
nor I_706 (I15061,I511615,I511609);
not I_707 (I15078,I15061);
nor I_708 (I15095,I14852,I15078);
nor I_709 (I15112,I15044,I15095);
DFFARX1 I_710 (I15112,I3035,I14688,I14677,);
nor I_711 (I15143,I15005,I15078);
nor I_712 (I14665,I14869,I15143);
nor I_713 (I14659,I15005,I15061);
not I_714 (I15215,I3042);
DFFARX1 I_715 (I59981,I3035,I15215,I15241,);
DFFARX1 I_716 (I15241,I3035,I15215,I15258,);
not I_717 (I15266,I15258);
nand I_718 (I15283,I59981,I59996);
and I_719 (I15300,I15283,I59999);
DFFARX1 I_720 (I15300,I3035,I15215,I15326,);
DFFARX1 I_721 (I15326,I3035,I15215,I15207,);
DFFARX1 I_722 (I15326,I3035,I15215,I15198,);
DFFARX1 I_723 (I59993,I3035,I15215,I15371,);
nand I_724 (I15379,I15371,I60002);
not I_725 (I15396,I15379);
nor I_726 (I15195,I15241,I15396);
DFFARX1 I_727 (I59978,I3035,I15215,I15436,);
not I_728 (I15444,I15436);
nor I_729 (I15201,I15444,I15266);
nand I_730 (I15189,I15444,I15379);
nand I_731 (I15489,I59978,I59984);
and I_732 (I15506,I15489,I59987);
DFFARX1 I_733 (I15506,I3035,I15215,I15532,);
nor I_734 (I15540,I15532,I15241);
DFFARX1 I_735 (I15540,I3035,I15215,I15183,);
not I_736 (I15571,I15532);
nor I_737 (I15588,I59990,I59984);
not I_738 (I15605,I15588);
nor I_739 (I15622,I15379,I15605);
nor I_740 (I15639,I15571,I15622);
DFFARX1 I_741 (I15639,I3035,I15215,I15204,);
nor I_742 (I15670,I15532,I15605);
nor I_743 (I15192,I15396,I15670);
nor I_744 (I15186,I15532,I15588);
not I_745 (I15742,I3042);
DFFARX1 I_746 (I684063,I3035,I15742,I15768,);
DFFARX1 I_747 (I15768,I3035,I15742,I15785,);
not I_748 (I15793,I15785);
nand I_749 (I15810,I684066,I684060);
and I_750 (I15827,I15810,I684069);
DFFARX1 I_751 (I15827,I3035,I15742,I15853,);
DFFARX1 I_752 (I15853,I3035,I15742,I15734,);
DFFARX1 I_753 (I15853,I3035,I15742,I15725,);
DFFARX1 I_754 (I684057,I3035,I15742,I15898,);
nand I_755 (I15906,I15898,I684072);
not I_756 (I15923,I15906);
nor I_757 (I15722,I15768,I15923);
DFFARX1 I_758 (I684048,I3035,I15742,I15963,);
not I_759 (I15971,I15963);
nor I_760 (I15728,I15971,I15793);
nand I_761 (I15716,I15971,I15906);
nand I_762 (I16016,I684051,I684051);
and I_763 (I16033,I16016,I684048);
DFFARX1 I_764 (I16033,I3035,I15742,I16059,);
nor I_765 (I16067,I16059,I15768);
DFFARX1 I_766 (I16067,I3035,I15742,I15710,);
not I_767 (I16098,I16059);
nor I_768 (I16115,I684054,I684051);
not I_769 (I16132,I16115);
nor I_770 (I16149,I15906,I16132);
nor I_771 (I16166,I16098,I16149);
DFFARX1 I_772 (I16166,I3035,I15742,I15731,);
nor I_773 (I16197,I16059,I16132);
nor I_774 (I15719,I15923,I16197);
nor I_775 (I15713,I16059,I16115);
not I_776 (I16269,I3042);
DFFARX1 I_777 (I674237,I3035,I16269,I16295,);
DFFARX1 I_778 (I16295,I3035,I16269,I16312,);
not I_779 (I16320,I16312);
nand I_780 (I16337,I674240,I674234);
and I_781 (I16354,I16337,I674243);
DFFARX1 I_782 (I16354,I3035,I16269,I16380,);
DFFARX1 I_783 (I16380,I3035,I16269,I16261,);
DFFARX1 I_784 (I16380,I3035,I16269,I16252,);
DFFARX1 I_785 (I674231,I3035,I16269,I16425,);
nand I_786 (I16433,I16425,I674246);
not I_787 (I16450,I16433);
nor I_788 (I16249,I16295,I16450);
DFFARX1 I_789 (I674222,I3035,I16269,I16490,);
not I_790 (I16498,I16490);
nor I_791 (I16255,I16498,I16320);
nand I_792 (I16243,I16498,I16433);
nand I_793 (I16543,I674225,I674225);
and I_794 (I16560,I16543,I674222);
DFFARX1 I_795 (I16560,I3035,I16269,I16586,);
nor I_796 (I16594,I16586,I16295);
DFFARX1 I_797 (I16594,I3035,I16269,I16237,);
not I_798 (I16625,I16586);
nor I_799 (I16642,I674228,I674225);
not I_800 (I16659,I16642);
nor I_801 (I16676,I16433,I16659);
nor I_802 (I16693,I16625,I16676);
DFFARX1 I_803 (I16693,I3035,I16269,I16258,);
nor I_804 (I16724,I16586,I16659);
nor I_805 (I16246,I16450,I16724);
nor I_806 (I16240,I16586,I16642);
not I_807 (I16796,I3042);
DFFARX1 I_808 (I178784,I3035,I16796,I16822,);
DFFARX1 I_809 (I16822,I3035,I16796,I16839,);
not I_810 (I16847,I16839);
nand I_811 (I16864,I178781,I178775);
and I_812 (I16881,I16864,I178769);
DFFARX1 I_813 (I16881,I3035,I16796,I16907,);
DFFARX1 I_814 (I16907,I3035,I16796,I16788,);
DFFARX1 I_815 (I16907,I3035,I16796,I16779,);
DFFARX1 I_816 (I178757,I3035,I16796,I16952,);
nand I_817 (I16960,I16952,I178766);
not I_818 (I16977,I16960);
nor I_819 (I16776,I16822,I16977);
DFFARX1 I_820 (I178763,I3035,I16796,I17017,);
not I_821 (I17025,I17017);
nor I_822 (I16782,I17025,I16847);
nand I_823 (I16770,I17025,I16960);
nand I_824 (I17070,I178760,I178778);
and I_825 (I17087,I17070,I178757);
DFFARX1 I_826 (I17087,I3035,I16796,I17113,);
nor I_827 (I17121,I17113,I16822);
DFFARX1 I_828 (I17121,I3035,I16796,I16764,);
not I_829 (I17152,I17113);
nor I_830 (I17169,I178772,I178778);
not I_831 (I17186,I17169);
nor I_832 (I17203,I16960,I17186);
nor I_833 (I17220,I17152,I17203);
DFFARX1 I_834 (I17220,I3035,I16796,I16785,);
nor I_835 (I17251,I17113,I17186);
nor I_836 (I16773,I16977,I17251);
nor I_837 (I16767,I17113,I17169);
not I_838 (I17323,I3042);
DFFARX1 I_839 (I190378,I3035,I17323,I17349,);
DFFARX1 I_840 (I17349,I3035,I17323,I17366,);
not I_841 (I17374,I17366);
nand I_842 (I17391,I190375,I190369);
and I_843 (I17408,I17391,I190363);
DFFARX1 I_844 (I17408,I3035,I17323,I17434,);
DFFARX1 I_845 (I17434,I3035,I17323,I17315,);
DFFARX1 I_846 (I17434,I3035,I17323,I17306,);
DFFARX1 I_847 (I190351,I3035,I17323,I17479,);
nand I_848 (I17487,I17479,I190360);
not I_849 (I17504,I17487);
nor I_850 (I17303,I17349,I17504);
DFFARX1 I_851 (I190357,I3035,I17323,I17544,);
not I_852 (I17552,I17544);
nor I_853 (I17309,I17552,I17374);
nand I_854 (I17297,I17552,I17487);
nand I_855 (I17597,I190354,I190372);
and I_856 (I17614,I17597,I190351);
DFFARX1 I_857 (I17614,I3035,I17323,I17640,);
nor I_858 (I17648,I17640,I17349);
DFFARX1 I_859 (I17648,I3035,I17323,I17291,);
not I_860 (I17679,I17640);
nor I_861 (I17696,I190366,I190372);
not I_862 (I17713,I17696);
nor I_863 (I17730,I17487,I17713);
nor I_864 (I17747,I17679,I17730);
DFFARX1 I_865 (I17747,I3035,I17323,I17312,);
nor I_866 (I17778,I17640,I17713);
nor I_867 (I17300,I17504,I17778);
nor I_868 (I17294,I17640,I17696);
not I_869 (I17850,I3042);
DFFARX1 I_870 (I127100,I3035,I17850,I17876,);
DFFARX1 I_871 (I17876,I3035,I17850,I17893,);
not I_872 (I17901,I17893);
nand I_873 (I17918,I127118,I127103);
and I_874 (I17935,I17918,I127106);
DFFARX1 I_875 (I17935,I3035,I17850,I17961,);
DFFARX1 I_876 (I17961,I3035,I17850,I17842,);
DFFARX1 I_877 (I17961,I3035,I17850,I17833,);
DFFARX1 I_878 (I127094,I3035,I17850,I18006,);
nand I_879 (I18014,I18006,I127097);
not I_880 (I18031,I18014);
nor I_881 (I17830,I17876,I18031);
DFFARX1 I_882 (I127109,I3035,I17850,I18071,);
not I_883 (I18079,I18071);
nor I_884 (I17836,I18079,I17901);
nand I_885 (I17824,I18079,I18014);
nand I_886 (I18124,I127115,I127112);
and I_887 (I18141,I18124,I127097);
DFFARX1 I_888 (I18141,I3035,I17850,I18167,);
nor I_889 (I18175,I18167,I17876);
DFFARX1 I_890 (I18175,I3035,I17850,I17818,);
not I_891 (I18206,I18167);
nor I_892 (I18223,I127094,I127112);
not I_893 (I18240,I18223);
nor I_894 (I18257,I18014,I18240);
nor I_895 (I18274,I18206,I18257);
DFFARX1 I_896 (I18274,I3035,I17850,I17839,);
nor I_897 (I18305,I18167,I18240);
nor I_898 (I17827,I18031,I18305);
nor I_899 (I17821,I18167,I18223);
not I_900 (I18377,I3042);
DFFARX1 I_901 (I421390,I3035,I18377,I18403,);
DFFARX1 I_902 (I18403,I3035,I18377,I18420,);
not I_903 (I18428,I18420);
nand I_904 (I18445,I421381,I421402);
and I_905 (I18462,I18445,I421384);
DFFARX1 I_906 (I18462,I3035,I18377,I18488,);
DFFARX1 I_907 (I18488,I3035,I18377,I18369,);
DFFARX1 I_908 (I18488,I3035,I18377,I18360,);
DFFARX1 I_909 (I421384,I3035,I18377,I18533,);
nand I_910 (I18541,I18533,I421399);
not I_911 (I18558,I18541);
nor I_912 (I18357,I18403,I18558);
DFFARX1 I_913 (I421393,I3035,I18377,I18598,);
not I_914 (I18606,I18598);
nor I_915 (I18363,I18606,I18428);
nand I_916 (I18351,I18606,I18541);
nand I_917 (I18651,I421387,I421396);
and I_918 (I18668,I18651,I421381);
DFFARX1 I_919 (I18668,I3035,I18377,I18694,);
nor I_920 (I18702,I18694,I18403);
DFFARX1 I_921 (I18702,I3035,I18377,I18345,);
not I_922 (I18733,I18694);
nor I_923 (I18750,I421387,I421396);
not I_924 (I18767,I18750);
nor I_925 (I18784,I18541,I18767);
nor I_926 (I18801,I18733,I18784);
DFFARX1 I_927 (I18801,I3035,I18377,I18366,);
nor I_928 (I18832,I18694,I18767);
nor I_929 (I18354,I18558,I18832);
nor I_930 (I18348,I18694,I18750);
not I_931 (I18904,I3042);
DFFARX1 I_932 (I467239,I3035,I18904,I18930,);
DFFARX1 I_933 (I18930,I3035,I18904,I18947,);
not I_934 (I18955,I18947);
nand I_935 (I18972,I467230,I467251);
and I_936 (I18989,I18972,I467233);
DFFARX1 I_937 (I18989,I3035,I18904,I19015,);
DFFARX1 I_938 (I19015,I3035,I18904,I18896,);
DFFARX1 I_939 (I19015,I3035,I18904,I18887,);
DFFARX1 I_940 (I467233,I3035,I18904,I19060,);
nand I_941 (I19068,I19060,I467248);
not I_942 (I19085,I19068);
nor I_943 (I18884,I18930,I19085);
DFFARX1 I_944 (I467242,I3035,I18904,I19125,);
not I_945 (I19133,I19125);
nor I_946 (I18890,I19133,I18955);
nand I_947 (I18878,I19133,I19068);
nand I_948 (I19178,I467236,I467245);
and I_949 (I19195,I19178,I467230);
DFFARX1 I_950 (I19195,I3035,I18904,I19221,);
nor I_951 (I19229,I19221,I18930);
DFFARX1 I_952 (I19229,I3035,I18904,I18872,);
not I_953 (I19260,I19221);
nor I_954 (I19277,I467236,I467245);
not I_955 (I19294,I19277);
nor I_956 (I19311,I19068,I19294);
nor I_957 (I19328,I19260,I19311);
DFFARX1 I_958 (I19328,I3035,I18904,I18893,);
nor I_959 (I19359,I19221,I19294);
nor I_960 (I18881,I19085,I19359);
nor I_961 (I18875,I19221,I19277);
not I_962 (I19431,I3042);
DFFARX1 I_963 (I441943,I3035,I19431,I19457,);
DFFARX1 I_964 (I19457,I3035,I19431,I19474,);
not I_965 (I19482,I19474);
nand I_966 (I19499,I441934,I441955);
and I_967 (I19516,I19499,I441937);
DFFARX1 I_968 (I19516,I3035,I19431,I19542,);
DFFARX1 I_969 (I19542,I3035,I19431,I19423,);
DFFARX1 I_970 (I19542,I3035,I19431,I19414,);
DFFARX1 I_971 (I441937,I3035,I19431,I19587,);
nand I_972 (I19595,I19587,I441952);
not I_973 (I19612,I19595);
nor I_974 (I19411,I19457,I19612);
DFFARX1 I_975 (I441946,I3035,I19431,I19652,);
not I_976 (I19660,I19652);
nor I_977 (I19417,I19660,I19482);
nand I_978 (I19405,I19660,I19595);
nand I_979 (I19705,I441940,I441949);
and I_980 (I19722,I19705,I441934);
DFFARX1 I_981 (I19722,I3035,I19431,I19748,);
nor I_982 (I19756,I19748,I19457);
DFFARX1 I_983 (I19756,I3035,I19431,I19399,);
not I_984 (I19787,I19748);
nor I_985 (I19804,I441940,I441949);
not I_986 (I19821,I19804);
nor I_987 (I19838,I19595,I19821);
nor I_988 (I19855,I19787,I19838);
DFFARX1 I_989 (I19855,I3035,I19431,I19420,);
nor I_990 (I19886,I19748,I19821);
nor I_991 (I19408,I19612,I19886);
nor I_992 (I19402,I19748,I19804);
not I_993 (I19958,I3042);
DFFARX1 I_994 (I275589,I3035,I19958,I19984,);
DFFARX1 I_995 (I19984,I3035,I19958,I20001,);
not I_996 (I20009,I20001);
nand I_997 (I20026,I275589,I275592);
and I_998 (I20043,I20026,I275613);
DFFARX1 I_999 (I20043,I3035,I19958,I20069,);
DFFARX1 I_1000 (I20069,I3035,I19958,I19950,);
DFFARX1 I_1001 (I20069,I3035,I19958,I19941,);
DFFARX1 I_1002 (I275601,I3035,I19958,I20114,);
nand I_1003 (I20122,I20114,I275604);
not I_1004 (I20139,I20122);
nor I_1005 (I19938,I19984,I20139);
DFFARX1 I_1006 (I275610,I3035,I19958,I20179,);
not I_1007 (I20187,I20179);
nor I_1008 (I19944,I20187,I20009);
nand I_1009 (I19932,I20187,I20122);
nand I_1010 (I20232,I275607,I275595);
and I_1011 (I20249,I20232,I275598);
DFFARX1 I_1012 (I20249,I3035,I19958,I20275,);
nor I_1013 (I20283,I20275,I19984);
DFFARX1 I_1014 (I20283,I3035,I19958,I19926,);
not I_1015 (I20314,I20275);
nor I_1016 (I20331,I275616,I275595);
not I_1017 (I20348,I20331);
nor I_1018 (I20365,I20122,I20348);
nor I_1019 (I20382,I20314,I20365);
DFFARX1 I_1020 (I20382,I3035,I19958,I19947,);
nor I_1021 (I20413,I20275,I20348);
nor I_1022 (I19935,I20139,I20413);
nor I_1023 (I19929,I20275,I20331);
not I_1024 (I20485,I3042);
DFFARX1 I_1025 (I258181,I3035,I20485,I20511,);
DFFARX1 I_1026 (I20511,I3035,I20485,I20528,);
not I_1027 (I20536,I20528);
nand I_1028 (I20553,I258181,I258184);
and I_1029 (I20570,I20553,I258205);
DFFARX1 I_1030 (I20570,I3035,I20485,I20596,);
DFFARX1 I_1031 (I20596,I3035,I20485,I20477,);
DFFARX1 I_1032 (I20596,I3035,I20485,I20468,);
DFFARX1 I_1033 (I258193,I3035,I20485,I20641,);
nand I_1034 (I20649,I20641,I258196);
not I_1035 (I20666,I20649);
nor I_1036 (I20465,I20511,I20666);
DFFARX1 I_1037 (I258202,I3035,I20485,I20706,);
not I_1038 (I20714,I20706);
nor I_1039 (I20471,I20714,I20536);
nand I_1040 (I20459,I20714,I20649);
nand I_1041 (I20759,I258199,I258187);
and I_1042 (I20776,I20759,I258190);
DFFARX1 I_1043 (I20776,I3035,I20485,I20802,);
nor I_1044 (I20810,I20802,I20511);
DFFARX1 I_1045 (I20810,I3035,I20485,I20453,);
not I_1046 (I20841,I20802);
nor I_1047 (I20858,I258208,I258187);
not I_1048 (I20875,I20858);
nor I_1049 (I20892,I20649,I20875);
nor I_1050 (I20909,I20841,I20892);
DFFARX1 I_1051 (I20909,I3035,I20485,I20474,);
nor I_1052 (I20940,I20802,I20875);
nor I_1053 (I20462,I20666,I20940);
nor I_1054 (I20456,I20802,I20858);
not I_1055 (I21012,I3042);
DFFARX1 I_1056 (I605260,I3035,I21012,I21038,);
DFFARX1 I_1057 (I21038,I3035,I21012,I21055,);
not I_1058 (I21063,I21055);
nand I_1059 (I21080,I605248,I605239);
and I_1060 (I21097,I21080,I605236);
DFFARX1 I_1061 (I21097,I3035,I21012,I21123,);
DFFARX1 I_1062 (I21123,I3035,I21012,I21004,);
DFFARX1 I_1063 (I21123,I3035,I21012,I20995,);
DFFARX1 I_1064 (I605242,I3035,I21012,I21168,);
nand I_1065 (I21176,I21168,I605254);
not I_1066 (I21193,I21176);
nor I_1067 (I20992,I21038,I21193);
DFFARX1 I_1068 (I605251,I3035,I21012,I21233,);
not I_1069 (I21241,I21233);
nor I_1070 (I20998,I21241,I21063);
nand I_1071 (I20986,I21241,I21176);
nand I_1072 (I21286,I605245,I605239);
and I_1073 (I21303,I21286,I605257);
DFFARX1 I_1074 (I21303,I3035,I21012,I21329,);
nor I_1075 (I21337,I21329,I21038);
DFFARX1 I_1076 (I21337,I3035,I21012,I20980,);
not I_1077 (I21368,I21329);
nor I_1078 (I21385,I605236,I605239);
not I_1079 (I21402,I21385);
nor I_1080 (I21419,I21176,I21402);
nor I_1081 (I21436,I21368,I21419);
DFFARX1 I_1082 (I21436,I3035,I21012,I21001,);
nor I_1083 (I21467,I21329,I21402);
nor I_1084 (I20989,I21193,I21467);
nor I_1085 (I20983,I21329,I21385);
not I_1086 (I21539,I3042);
DFFARX1 I_1087 (I584452,I3035,I21539,I21565,);
DFFARX1 I_1088 (I21565,I3035,I21539,I21582,);
not I_1089 (I21590,I21582);
nand I_1090 (I21607,I584440,I584431);
and I_1091 (I21624,I21607,I584428);
DFFARX1 I_1092 (I21624,I3035,I21539,I21650,);
DFFARX1 I_1093 (I21650,I3035,I21539,I21531,);
DFFARX1 I_1094 (I21650,I3035,I21539,I21522,);
DFFARX1 I_1095 (I584434,I3035,I21539,I21695,);
nand I_1096 (I21703,I21695,I584446);
not I_1097 (I21720,I21703);
nor I_1098 (I21519,I21565,I21720);
DFFARX1 I_1099 (I584443,I3035,I21539,I21760,);
not I_1100 (I21768,I21760);
nor I_1101 (I21525,I21768,I21590);
nand I_1102 (I21513,I21768,I21703);
nand I_1103 (I21813,I584437,I584431);
and I_1104 (I21830,I21813,I584449);
DFFARX1 I_1105 (I21830,I3035,I21539,I21856,);
nor I_1106 (I21864,I21856,I21565);
DFFARX1 I_1107 (I21864,I3035,I21539,I21507,);
not I_1108 (I21895,I21856);
nor I_1109 (I21912,I584428,I584431);
not I_1110 (I21929,I21912);
nor I_1111 (I21946,I21703,I21929);
nor I_1112 (I21963,I21895,I21946);
DFFARX1 I_1113 (I21963,I3035,I21539,I21528,);
nor I_1114 (I21994,I21856,I21929);
nor I_1115 (I21516,I21720,I21994);
nor I_1116 (I21510,I21856,I21912);
not I_1117 (I22066,I3042);
DFFARX1 I_1118 (I160866,I3035,I22066,I22092,);
DFFARX1 I_1119 (I22092,I3035,I22066,I22109,);
not I_1120 (I22117,I22109);
nand I_1121 (I22134,I160863,I160857);
and I_1122 (I22151,I22134,I160851);
DFFARX1 I_1123 (I22151,I3035,I22066,I22177,);
DFFARX1 I_1124 (I22177,I3035,I22066,I22058,);
DFFARX1 I_1125 (I22177,I3035,I22066,I22049,);
DFFARX1 I_1126 (I160839,I3035,I22066,I22222,);
nand I_1127 (I22230,I22222,I160848);
not I_1128 (I22247,I22230);
nor I_1129 (I22046,I22092,I22247);
DFFARX1 I_1130 (I160845,I3035,I22066,I22287,);
not I_1131 (I22295,I22287);
nor I_1132 (I22052,I22295,I22117);
nand I_1133 (I22040,I22295,I22230);
nand I_1134 (I22340,I160842,I160860);
and I_1135 (I22357,I22340,I160839);
DFFARX1 I_1136 (I22357,I3035,I22066,I22383,);
nor I_1137 (I22391,I22383,I22092);
DFFARX1 I_1138 (I22391,I3035,I22066,I22034,);
not I_1139 (I22422,I22383);
nor I_1140 (I22439,I160854,I160860);
not I_1141 (I22456,I22439);
nor I_1142 (I22473,I22230,I22456);
nor I_1143 (I22490,I22422,I22473);
DFFARX1 I_1144 (I22490,I3035,I22066,I22055,);
nor I_1145 (I22521,I22383,I22456);
nor I_1146 (I22043,I22247,I22521);
nor I_1147 (I22037,I22383,I22439);
not I_1148 (I22593,I3042);
DFFARX1 I_1149 (I165082,I3035,I22593,I22619,);
DFFARX1 I_1150 (I22619,I3035,I22593,I22636,);
not I_1151 (I22644,I22636);
nand I_1152 (I22661,I165079,I165073);
and I_1153 (I22678,I22661,I165067);
DFFARX1 I_1154 (I22678,I3035,I22593,I22704,);
DFFARX1 I_1155 (I22704,I3035,I22593,I22585,);
DFFARX1 I_1156 (I22704,I3035,I22593,I22576,);
DFFARX1 I_1157 (I165055,I3035,I22593,I22749,);
nand I_1158 (I22757,I22749,I165064);
not I_1159 (I22774,I22757);
nor I_1160 (I22573,I22619,I22774);
DFFARX1 I_1161 (I165061,I3035,I22593,I22814,);
not I_1162 (I22822,I22814);
nor I_1163 (I22579,I22822,I22644);
nand I_1164 (I22567,I22822,I22757);
nand I_1165 (I22867,I165058,I165076);
and I_1166 (I22884,I22867,I165055);
DFFARX1 I_1167 (I22884,I3035,I22593,I22910,);
nor I_1168 (I22918,I22910,I22619);
DFFARX1 I_1169 (I22918,I3035,I22593,I22561,);
not I_1170 (I22949,I22910);
nor I_1171 (I22966,I165070,I165076);
not I_1172 (I22983,I22966);
nor I_1173 (I23000,I22757,I22983);
nor I_1174 (I23017,I22949,I23000);
DFFARX1 I_1175 (I23017,I3035,I22593,I22582,);
nor I_1176 (I23048,I22910,I22983);
nor I_1177 (I22570,I22774,I23048);
nor I_1178 (I22564,I22910,I22966);
not I_1179 (I23120,I3042);
DFFARX1 I_1180 (I481908,I3035,I23120,I23146,);
DFFARX1 I_1181 (I23146,I3035,I23120,I23163,);
not I_1182 (I23171,I23163);
nand I_1183 (I23188,I481884,I481911);
and I_1184 (I23205,I23188,I481896);
DFFARX1 I_1185 (I23205,I3035,I23120,I23231,);
DFFARX1 I_1186 (I23231,I3035,I23120,I23112,);
DFFARX1 I_1187 (I23231,I3035,I23120,I23103,);
DFFARX1 I_1188 (I481902,I3035,I23120,I23276,);
nand I_1189 (I23284,I23276,I481887);
not I_1190 (I23301,I23284);
nor I_1191 (I23100,I23146,I23301);
DFFARX1 I_1192 (I481905,I3035,I23120,I23341,);
not I_1193 (I23349,I23341);
nor I_1194 (I23106,I23349,I23171);
nand I_1195 (I23094,I23349,I23284);
nand I_1196 (I23394,I481890,I481893);
and I_1197 (I23411,I23394,I481884);
DFFARX1 I_1198 (I23411,I3035,I23120,I23437,);
nor I_1199 (I23445,I23437,I23146);
DFFARX1 I_1200 (I23445,I3035,I23120,I23088,);
not I_1201 (I23476,I23437);
nor I_1202 (I23493,I481899,I481893);
not I_1203 (I23510,I23493);
nor I_1204 (I23527,I23284,I23510);
nor I_1205 (I23544,I23476,I23527);
DFFARX1 I_1206 (I23544,I3035,I23120,I23109,);
nor I_1207 (I23575,I23437,I23510);
nor I_1208 (I23097,I23301,I23575);
nor I_1209 (I23091,I23437,I23493);
not I_1210 (I23647,I3042);
DFFARX1 I_1211 (I292445,I3035,I23647,I23673,);
DFFARX1 I_1212 (I23673,I3035,I23647,I23690,);
not I_1213 (I23698,I23690);
nand I_1214 (I23715,I292451,I292439);
and I_1215 (I23732,I23715,I292436);
DFFARX1 I_1216 (I23732,I3035,I23647,I23758,);
DFFARX1 I_1217 (I23758,I3035,I23647,I23639,);
DFFARX1 I_1218 (I23758,I3035,I23647,I23630,);
DFFARX1 I_1219 (I292448,I3035,I23647,I23803,);
nand I_1220 (I23811,I23803,I292442);
not I_1221 (I23828,I23811);
nor I_1222 (I23627,I23673,I23828);
DFFARX1 I_1223 (I292460,I3035,I23647,I23868,);
not I_1224 (I23876,I23868);
nor I_1225 (I23633,I23876,I23698);
nand I_1226 (I23621,I23876,I23811);
nand I_1227 (I23921,I292454,I292457);
and I_1228 (I23938,I23921,I292439);
DFFARX1 I_1229 (I23938,I3035,I23647,I23964,);
nor I_1230 (I23972,I23964,I23673);
DFFARX1 I_1231 (I23972,I3035,I23647,I23615,);
not I_1232 (I24003,I23964);
nor I_1233 (I24020,I292436,I292457);
not I_1234 (I24037,I24020);
nor I_1235 (I24054,I23811,I24037);
nor I_1236 (I24071,I24003,I24054);
DFFARX1 I_1237 (I24071,I3035,I23647,I23636,);
nor I_1238 (I24102,I23964,I24037);
nor I_1239 (I23624,I23828,I24102);
nor I_1240 (I23618,I23964,I24020);
not I_1241 (I24174,I3042);
DFFARX1 I_1242 (I272869,I3035,I24174,I24200,);
DFFARX1 I_1243 (I24200,I3035,I24174,I24217,);
not I_1244 (I24225,I24217);
nand I_1245 (I24242,I272869,I272872);
and I_1246 (I24259,I24242,I272893);
DFFARX1 I_1247 (I24259,I3035,I24174,I24285,);
DFFARX1 I_1248 (I24285,I3035,I24174,I24166,);
DFFARX1 I_1249 (I24285,I3035,I24174,I24157,);
DFFARX1 I_1250 (I272881,I3035,I24174,I24330,);
nand I_1251 (I24338,I24330,I272884);
not I_1252 (I24355,I24338);
nor I_1253 (I24154,I24200,I24355);
DFFARX1 I_1254 (I272890,I3035,I24174,I24395,);
not I_1255 (I24403,I24395);
nor I_1256 (I24160,I24403,I24225);
nand I_1257 (I24148,I24403,I24338);
nand I_1258 (I24448,I272887,I272875);
and I_1259 (I24465,I24448,I272878);
DFFARX1 I_1260 (I24465,I3035,I24174,I24491,);
nor I_1261 (I24499,I24491,I24200);
DFFARX1 I_1262 (I24499,I3035,I24174,I24142,);
not I_1263 (I24530,I24491);
nor I_1264 (I24547,I272896,I272875);
not I_1265 (I24564,I24547);
nor I_1266 (I24581,I24338,I24564);
nor I_1267 (I24598,I24530,I24581);
DFFARX1 I_1268 (I24598,I3035,I24174,I24163,);
nor I_1269 (I24629,I24491,I24564);
nor I_1270 (I24151,I24355,I24629);
nor I_1271 (I24145,I24491,I24547);
not I_1272 (I24701,I3042);
DFFARX1 I_1273 (I671925,I3035,I24701,I24727,);
DFFARX1 I_1274 (I24727,I3035,I24701,I24744,);
not I_1275 (I24752,I24744);
nand I_1276 (I24769,I671928,I671922);
and I_1277 (I24786,I24769,I671931);
DFFARX1 I_1278 (I24786,I3035,I24701,I24812,);
DFFARX1 I_1279 (I24812,I3035,I24701,I24693,);
DFFARX1 I_1280 (I24812,I3035,I24701,I24684,);
DFFARX1 I_1281 (I671919,I3035,I24701,I24857,);
nand I_1282 (I24865,I24857,I671934);
not I_1283 (I24882,I24865);
nor I_1284 (I24681,I24727,I24882);
DFFARX1 I_1285 (I671910,I3035,I24701,I24922,);
not I_1286 (I24930,I24922);
nor I_1287 (I24687,I24930,I24752);
nand I_1288 (I24675,I24930,I24865);
nand I_1289 (I24975,I671913,I671913);
and I_1290 (I24992,I24975,I671910);
DFFARX1 I_1291 (I24992,I3035,I24701,I25018,);
nor I_1292 (I25026,I25018,I24727);
DFFARX1 I_1293 (I25026,I3035,I24701,I24669,);
not I_1294 (I25057,I25018);
nor I_1295 (I25074,I671916,I671913);
not I_1296 (I25091,I25074);
nor I_1297 (I25108,I24865,I25091);
nor I_1298 (I25125,I25057,I25108);
DFFARX1 I_1299 (I25125,I3035,I24701,I24690,);
nor I_1300 (I25156,I25018,I25091);
nor I_1301 (I24678,I24882,I25156);
nor I_1302 (I24672,I25018,I25074);
not I_1303 (I25228,I3042);
DFFARX1 I_1304 (I277221,I3035,I25228,I25254,);
DFFARX1 I_1305 (I25254,I3035,I25228,I25271,);
not I_1306 (I25279,I25271);
nand I_1307 (I25296,I277221,I277224);
and I_1308 (I25313,I25296,I277245);
DFFARX1 I_1309 (I25313,I3035,I25228,I25339,);
DFFARX1 I_1310 (I25339,I3035,I25228,I25220,);
DFFARX1 I_1311 (I25339,I3035,I25228,I25211,);
DFFARX1 I_1312 (I277233,I3035,I25228,I25384,);
nand I_1313 (I25392,I25384,I277236);
not I_1314 (I25409,I25392);
nor I_1315 (I25208,I25254,I25409);
DFFARX1 I_1316 (I277242,I3035,I25228,I25449,);
not I_1317 (I25457,I25449);
nor I_1318 (I25214,I25457,I25279);
nand I_1319 (I25202,I25457,I25392);
nand I_1320 (I25502,I277239,I277227);
and I_1321 (I25519,I25502,I277230);
DFFARX1 I_1322 (I25519,I3035,I25228,I25545,);
nor I_1323 (I25553,I25545,I25254);
DFFARX1 I_1324 (I25553,I3035,I25228,I25196,);
not I_1325 (I25584,I25545);
nor I_1326 (I25601,I277248,I277227);
not I_1327 (I25618,I25601);
nor I_1328 (I25635,I25392,I25618);
nor I_1329 (I25652,I25584,I25635);
DFFARX1 I_1330 (I25652,I3035,I25228,I25217,);
nor I_1331 (I25683,I25545,I25618);
nor I_1332 (I25205,I25409,I25683);
nor I_1333 (I25199,I25545,I25601);
not I_1334 (I25755,I3042);
DFFARX1 I_1335 (I585608,I3035,I25755,I25781,);
DFFARX1 I_1336 (I25781,I3035,I25755,I25798,);
not I_1337 (I25806,I25798);
nand I_1338 (I25823,I585596,I585587);
and I_1339 (I25840,I25823,I585584);
DFFARX1 I_1340 (I25840,I3035,I25755,I25866,);
DFFARX1 I_1341 (I25866,I3035,I25755,I25747,);
DFFARX1 I_1342 (I25866,I3035,I25755,I25738,);
DFFARX1 I_1343 (I585590,I3035,I25755,I25911,);
nand I_1344 (I25919,I25911,I585602);
not I_1345 (I25936,I25919);
nor I_1346 (I25735,I25781,I25936);
DFFARX1 I_1347 (I585599,I3035,I25755,I25976,);
not I_1348 (I25984,I25976);
nor I_1349 (I25741,I25984,I25806);
nand I_1350 (I25729,I25984,I25919);
nand I_1351 (I26029,I585593,I585587);
and I_1352 (I26046,I26029,I585605);
DFFARX1 I_1353 (I26046,I3035,I25755,I26072,);
nor I_1354 (I26080,I26072,I25781);
DFFARX1 I_1355 (I26080,I3035,I25755,I25723,);
not I_1356 (I26111,I26072);
nor I_1357 (I26128,I585584,I585587);
not I_1358 (I26145,I26128);
nor I_1359 (I26162,I25919,I26145);
nor I_1360 (I26179,I26111,I26162);
DFFARX1 I_1361 (I26179,I3035,I25755,I25744,);
nor I_1362 (I26210,I26072,I26145);
nor I_1363 (I25732,I25936,I26210);
nor I_1364 (I25726,I26072,I26128);
not I_1365 (I26282,I3042);
DFFARX1 I_1366 (I239685,I3035,I26282,I26308,);
DFFARX1 I_1367 (I26308,I3035,I26282,I26325,);
not I_1368 (I26333,I26325);
nand I_1369 (I26350,I239685,I239688);
and I_1370 (I26367,I26350,I239709);
DFFARX1 I_1371 (I26367,I3035,I26282,I26393,);
DFFARX1 I_1372 (I26393,I3035,I26282,I26274,);
DFFARX1 I_1373 (I26393,I3035,I26282,I26265,);
DFFARX1 I_1374 (I239697,I3035,I26282,I26438,);
nand I_1375 (I26446,I26438,I239700);
not I_1376 (I26463,I26446);
nor I_1377 (I26262,I26308,I26463);
DFFARX1 I_1378 (I239706,I3035,I26282,I26503,);
not I_1379 (I26511,I26503);
nor I_1380 (I26268,I26511,I26333);
nand I_1381 (I26256,I26511,I26446);
nand I_1382 (I26556,I239703,I239691);
and I_1383 (I26573,I26556,I239694);
DFFARX1 I_1384 (I26573,I3035,I26282,I26599,);
nor I_1385 (I26607,I26599,I26308);
DFFARX1 I_1386 (I26607,I3035,I26282,I26250,);
not I_1387 (I26638,I26599);
nor I_1388 (I26655,I239712,I239691);
not I_1389 (I26672,I26655);
nor I_1390 (I26689,I26446,I26672);
nor I_1391 (I26706,I26638,I26689);
DFFARX1 I_1392 (I26706,I3035,I26282,I26271,);
nor I_1393 (I26737,I26599,I26672);
nor I_1394 (I26259,I26463,I26737);
nor I_1395 (I26253,I26599,I26655);
not I_1396 (I26809,I3042);
DFFARX1 I_1397 (I3661,I3035,I26809,I26835,);
DFFARX1 I_1398 (I26835,I3035,I26809,I26852,);
not I_1399 (I26860,I26852);
nand I_1400 (I26877,I3655,I3649);
and I_1401 (I26894,I26877,I3646);
DFFARX1 I_1402 (I26894,I3035,I26809,I26920,);
DFFARX1 I_1403 (I26920,I3035,I26809,I26801,);
DFFARX1 I_1404 (I26920,I3035,I26809,I26792,);
DFFARX1 I_1405 (I3652,I3035,I26809,I26965,);
nand I_1406 (I26973,I26965,I3646);
not I_1407 (I26990,I26973);
nor I_1408 (I26789,I26835,I26990);
DFFARX1 I_1409 (I3643,I3035,I26809,I27030,);
not I_1410 (I27038,I27030);
nor I_1411 (I26795,I27038,I26860);
nand I_1412 (I26783,I27038,I26973);
nand I_1413 (I27083,I3640,I3640);
and I_1414 (I27100,I27083,I3658);
DFFARX1 I_1415 (I27100,I3035,I26809,I27126,);
nor I_1416 (I27134,I27126,I26835);
DFFARX1 I_1417 (I27134,I3035,I26809,I26777,);
not I_1418 (I27165,I27126);
nor I_1419 (I27182,I3643,I3640);
not I_1420 (I27199,I27182);
nor I_1421 (I27216,I26973,I27199);
nor I_1422 (I27233,I27165,I27216);
DFFARX1 I_1423 (I27233,I3035,I26809,I26798,);
nor I_1424 (I27264,I27126,I27199);
nor I_1425 (I26786,I26990,I27264);
nor I_1426 (I26780,I27126,I27182);
not I_1427 (I27336,I3042);
DFFARX1 I_1428 (I345822,I3035,I27336,I27362,);
DFFARX1 I_1429 (I27362,I3035,I27336,I27379,);
not I_1430 (I27387,I27379);
nand I_1431 (I27404,I345837,I345840);
and I_1432 (I27421,I27404,I345819);
DFFARX1 I_1433 (I27421,I3035,I27336,I27447,);
DFFARX1 I_1434 (I27447,I3035,I27336,I27328,);
DFFARX1 I_1435 (I27447,I3035,I27336,I27319,);
DFFARX1 I_1436 (I345825,I3035,I27336,I27492,);
nand I_1437 (I27500,I27492,I345831);
not I_1438 (I27517,I27500);
nor I_1439 (I27316,I27362,I27517);
DFFARX1 I_1440 (I345819,I3035,I27336,I27557,);
not I_1441 (I27565,I27557);
nor I_1442 (I27322,I27565,I27387);
nand I_1443 (I27310,I27565,I27500);
nand I_1444 (I27610,I345834,I345816);
and I_1445 (I27627,I27610,I345828);
DFFARX1 I_1446 (I27627,I3035,I27336,I27653,);
nor I_1447 (I27661,I27653,I27362);
DFFARX1 I_1448 (I27661,I3035,I27336,I27304,);
not I_1449 (I27692,I27653);
nor I_1450 (I27709,I345816,I345816);
not I_1451 (I27726,I27709);
nor I_1452 (I27743,I27500,I27726);
nor I_1453 (I27760,I27692,I27743);
DFFARX1 I_1454 (I27760,I3035,I27336,I27325,);
nor I_1455 (I27791,I27653,I27726);
nor I_1456 (I27313,I27517,I27791);
nor I_1457 (I27307,I27653,I27709);
not I_1458 (I27863,I3042);
DFFARX1 I_1459 (I281140,I3035,I27863,I27889,);
DFFARX1 I_1460 (I27889,I3035,I27863,I27906,);
not I_1461 (I27914,I27906);
nand I_1462 (I27931,I281146,I281134);
and I_1463 (I27948,I27931,I281131);
DFFARX1 I_1464 (I27948,I3035,I27863,I27974,);
DFFARX1 I_1465 (I27974,I3035,I27863,I27855,);
DFFARX1 I_1466 (I27974,I3035,I27863,I27846,);
DFFARX1 I_1467 (I281143,I3035,I27863,I28019,);
nand I_1468 (I28027,I28019,I281137);
not I_1469 (I28044,I28027);
nor I_1470 (I27843,I27889,I28044);
DFFARX1 I_1471 (I281155,I3035,I27863,I28084,);
not I_1472 (I28092,I28084);
nor I_1473 (I27849,I28092,I27914);
nand I_1474 (I27837,I28092,I28027);
nand I_1475 (I28137,I281149,I281152);
and I_1476 (I28154,I28137,I281134);
DFFARX1 I_1477 (I28154,I3035,I27863,I28180,);
nor I_1478 (I28188,I28180,I27889);
DFFARX1 I_1479 (I28188,I3035,I27863,I27831,);
not I_1480 (I28219,I28180);
nor I_1481 (I28236,I281131,I281152);
not I_1482 (I28253,I28236);
nor I_1483 (I28270,I28027,I28253);
nor I_1484 (I28287,I28219,I28270);
DFFARX1 I_1485 (I28287,I3035,I27863,I27852,);
nor I_1486 (I28318,I28180,I28253);
nor I_1487 (I27840,I28044,I28318);
nor I_1488 (I27834,I28180,I28236);
not I_1489 (I28390,I3042);
DFFARX1 I_1490 (I225687,I3035,I28390,I28416,);
DFFARX1 I_1491 (I28416,I3035,I28390,I28433,);
not I_1492 (I28441,I28433);
nand I_1493 (I28458,I225684,I225678);
and I_1494 (I28475,I28458,I225672);
DFFARX1 I_1495 (I28475,I3035,I28390,I28501,);
DFFARX1 I_1496 (I28501,I3035,I28390,I28382,);
DFFARX1 I_1497 (I28501,I3035,I28390,I28373,);
DFFARX1 I_1498 (I225660,I3035,I28390,I28546,);
nand I_1499 (I28554,I28546,I225669);
not I_1500 (I28571,I28554);
nor I_1501 (I28370,I28416,I28571);
DFFARX1 I_1502 (I225666,I3035,I28390,I28611,);
not I_1503 (I28619,I28611);
nor I_1504 (I28376,I28619,I28441);
nand I_1505 (I28364,I28619,I28554);
nand I_1506 (I28664,I225663,I225681);
and I_1507 (I28681,I28664,I225660);
DFFARX1 I_1508 (I28681,I3035,I28390,I28707,);
nor I_1509 (I28715,I28707,I28416);
DFFARX1 I_1510 (I28715,I3035,I28390,I28358,);
not I_1511 (I28746,I28707);
nor I_1512 (I28763,I225675,I225681);
not I_1513 (I28780,I28763);
nor I_1514 (I28797,I28554,I28780);
nor I_1515 (I28814,I28746,I28797);
DFFARX1 I_1516 (I28814,I3035,I28390,I28379,);
nor I_1517 (I28845,I28707,I28780);
nor I_1518 (I28367,I28571,I28845);
nor I_1519 (I28361,I28707,I28763);
not I_1520 (I28917,I3042);
DFFARX1 I_1521 (I111041,I3035,I28917,I28943,);
not I_1522 (I28951,I28943);
nand I_1523 (I28968,I111035,I111029);
and I_1524 (I28985,I28968,I111050);
DFFARX1 I_1525 (I28985,I3035,I28917,I29011,);
DFFARX1 I_1526 (I111047,I3035,I28917,I29028,);
and I_1527 (I29036,I29028,I111044);
nor I_1528 (I29053,I29011,I29036);
DFFARX1 I_1529 (I29053,I3035,I28917,I28885,);
nand I_1530 (I29084,I29028,I111044);
nand I_1531 (I29101,I28951,I29084);
not I_1532 (I28897,I29101);
DFFARX1 I_1533 (I111029,I3035,I28917,I29141,);
DFFARX1 I_1534 (I29141,I3035,I28917,I28906,);
nand I_1535 (I29163,I111032,I111032);
and I_1536 (I29180,I29163,I111053);
DFFARX1 I_1537 (I29180,I3035,I28917,I29206,);
DFFARX1 I_1538 (I29206,I3035,I28917,I29223,);
not I_1539 (I28909,I29223);
not I_1540 (I29245,I29206);
nand I_1541 (I28894,I29245,I29084);
nor I_1542 (I29276,I111038,I111032);
not I_1543 (I29293,I29276);
nor I_1544 (I29310,I29245,I29293);
nor I_1545 (I29327,I28951,I29310);
DFFARX1 I_1546 (I29327,I3035,I28917,I28903,);
nor I_1547 (I29358,I29011,I29293);
nor I_1548 (I28891,I29206,I29358);
nor I_1549 (I28900,I29141,I29276);
nor I_1550 (I28888,I29011,I29276);
not I_1551 (I29444,I3042);
DFFARX1 I_1552 (I465658,I3035,I29444,I29470,);
not I_1553 (I29478,I29470);
nand I_1554 (I29495,I465655,I465670);
and I_1555 (I29512,I29495,I465652);
DFFARX1 I_1556 (I29512,I3035,I29444,I29538,);
DFFARX1 I_1557 (I465649,I3035,I29444,I29555,);
and I_1558 (I29563,I29555,I465649);
nor I_1559 (I29580,I29538,I29563);
DFFARX1 I_1560 (I29580,I3035,I29444,I29412,);
nand I_1561 (I29611,I29555,I465649);
nand I_1562 (I29628,I29478,I29611);
not I_1563 (I29424,I29628);
DFFARX1 I_1564 (I465652,I3035,I29444,I29668,);
DFFARX1 I_1565 (I29668,I3035,I29444,I29433,);
nand I_1566 (I29690,I465664,I465655);
and I_1567 (I29707,I29690,I465667);
DFFARX1 I_1568 (I29707,I3035,I29444,I29733,);
DFFARX1 I_1569 (I29733,I3035,I29444,I29750,);
not I_1570 (I29436,I29750);
not I_1571 (I29772,I29733);
nand I_1572 (I29421,I29772,I29611);
nor I_1573 (I29803,I465661,I465655);
not I_1574 (I29820,I29803);
nor I_1575 (I29837,I29772,I29820);
nor I_1576 (I29854,I29478,I29837);
DFFARX1 I_1577 (I29854,I3035,I29444,I29430,);
nor I_1578 (I29885,I29538,I29820);
nor I_1579 (I29418,I29733,I29885);
nor I_1580 (I29427,I29668,I29803);
nor I_1581 (I29415,I29538,I29803);
not I_1582 (I29971,I3042);
DFFARX1 I_1583 (I301319,I3035,I29971,I29997,);
not I_1584 (I30005,I29997);
nand I_1585 (I30022,I301331,I301316);
and I_1586 (I30039,I30022,I301310);
DFFARX1 I_1587 (I30039,I3035,I29971,I30065,);
DFFARX1 I_1588 (I301325,I3035,I29971,I30082,);
and I_1589 (I30090,I30082,I301313);
nor I_1590 (I30107,I30065,I30090);
DFFARX1 I_1591 (I30107,I3035,I29971,I29939,);
nand I_1592 (I30138,I30082,I301313);
nand I_1593 (I30155,I30005,I30138);
not I_1594 (I29951,I30155);
DFFARX1 I_1595 (I301322,I3035,I29971,I30195,);
DFFARX1 I_1596 (I30195,I3035,I29971,I29960,);
nand I_1597 (I30217,I301328,I301334);
and I_1598 (I30234,I30217,I301310);
DFFARX1 I_1599 (I30234,I3035,I29971,I30260,);
DFFARX1 I_1600 (I30260,I3035,I29971,I30277,);
not I_1601 (I29963,I30277);
not I_1602 (I30299,I30260);
nand I_1603 (I29948,I30299,I30138);
nor I_1604 (I30330,I301313,I301334);
not I_1605 (I30347,I30330);
nor I_1606 (I30364,I30299,I30347);
nor I_1607 (I30381,I30005,I30364);
DFFARX1 I_1608 (I30381,I3035,I29971,I29957,);
nor I_1609 (I30412,I30065,I30347);
nor I_1610 (I29945,I30260,I30412);
nor I_1611 (I29954,I30195,I30330);
nor I_1612 (I29942,I30065,I30330);
not I_1613 (I30498,I3042);
DFFARX1 I_1614 (I457753,I3035,I30498,I30524,);
not I_1615 (I30532,I30524);
nand I_1616 (I30549,I457750,I457765);
and I_1617 (I30566,I30549,I457747);
DFFARX1 I_1618 (I30566,I3035,I30498,I30592,);
DFFARX1 I_1619 (I457744,I3035,I30498,I30609,);
and I_1620 (I30617,I30609,I457744);
nor I_1621 (I30634,I30592,I30617);
DFFARX1 I_1622 (I30634,I3035,I30498,I30466,);
nand I_1623 (I30665,I30609,I457744);
nand I_1624 (I30682,I30532,I30665);
not I_1625 (I30478,I30682);
DFFARX1 I_1626 (I457747,I3035,I30498,I30722,);
DFFARX1 I_1627 (I30722,I3035,I30498,I30487,);
nand I_1628 (I30744,I457759,I457750);
and I_1629 (I30761,I30744,I457762);
DFFARX1 I_1630 (I30761,I3035,I30498,I30787,);
DFFARX1 I_1631 (I30787,I3035,I30498,I30804,);
not I_1632 (I30490,I30804);
not I_1633 (I30826,I30787);
nand I_1634 (I30475,I30826,I30665);
nor I_1635 (I30857,I457756,I457750);
not I_1636 (I30874,I30857);
nor I_1637 (I30891,I30826,I30874);
nor I_1638 (I30908,I30532,I30891);
DFFARX1 I_1639 (I30908,I3035,I30498,I30484,);
nor I_1640 (I30939,I30592,I30874);
nor I_1641 (I30472,I30787,I30939);
nor I_1642 (I30481,I30722,I30857);
nor I_1643 (I30469,I30592,I30857);
not I_1644 (I31025,I3042);
DFFARX1 I_1645 (I521299,I3035,I31025,I31051,);
not I_1646 (I31059,I31051);
nand I_1647 (I31076,I521317,I521311);
and I_1648 (I31093,I31076,I521290);
DFFARX1 I_1649 (I31093,I3035,I31025,I31119,);
DFFARX1 I_1650 (I521308,I3035,I31025,I31136,);
and I_1651 (I31144,I31136,I521293);
nor I_1652 (I31161,I31119,I31144);
DFFARX1 I_1653 (I31161,I3035,I31025,I30993,);
nand I_1654 (I31192,I31136,I521293);
nand I_1655 (I31209,I31059,I31192);
not I_1656 (I31005,I31209);
DFFARX1 I_1657 (I521305,I3035,I31025,I31249,);
DFFARX1 I_1658 (I31249,I3035,I31025,I31014,);
nand I_1659 (I31271,I521314,I521302);
and I_1660 (I31288,I31271,I521296);
DFFARX1 I_1661 (I31288,I3035,I31025,I31314,);
DFFARX1 I_1662 (I31314,I3035,I31025,I31331,);
not I_1663 (I31017,I31331);
not I_1664 (I31353,I31314);
nand I_1665 (I31002,I31353,I31192);
nor I_1666 (I31384,I521290,I521302);
not I_1667 (I31401,I31384);
nor I_1668 (I31418,I31353,I31401);
nor I_1669 (I31435,I31059,I31418);
DFFARX1 I_1670 (I31435,I3035,I31025,I31011,);
nor I_1671 (I31466,I31119,I31401);
nor I_1672 (I30999,I31314,I31466);
nor I_1673 (I31008,I31249,I31384);
nor I_1674 (I30996,I31119,I31384);
not I_1675 (I31552,I3042);
DFFARX1 I_1676 (I483185,I3035,I31552,I31578,);
not I_1677 (I31586,I31578);
nand I_1678 (I31603,I483203,I483197);
and I_1679 (I31620,I31603,I483176);
DFFARX1 I_1680 (I31620,I3035,I31552,I31646,);
DFFARX1 I_1681 (I483194,I3035,I31552,I31663,);
and I_1682 (I31671,I31663,I483179);
nor I_1683 (I31688,I31646,I31671);
DFFARX1 I_1684 (I31688,I3035,I31552,I31520,);
nand I_1685 (I31719,I31663,I483179);
nand I_1686 (I31736,I31586,I31719);
not I_1687 (I31532,I31736);
DFFARX1 I_1688 (I483191,I3035,I31552,I31776,);
DFFARX1 I_1689 (I31776,I3035,I31552,I31541,);
nand I_1690 (I31798,I483200,I483188);
and I_1691 (I31815,I31798,I483182);
DFFARX1 I_1692 (I31815,I3035,I31552,I31841,);
DFFARX1 I_1693 (I31841,I3035,I31552,I31858,);
not I_1694 (I31544,I31858);
not I_1695 (I31880,I31841);
nand I_1696 (I31529,I31880,I31719);
nor I_1697 (I31911,I483176,I483188);
not I_1698 (I31928,I31911);
nor I_1699 (I31945,I31880,I31928);
nor I_1700 (I31962,I31586,I31945);
DFFARX1 I_1701 (I31962,I3035,I31552,I31538,);
nor I_1702 (I31993,I31646,I31928);
nor I_1703 (I31526,I31841,I31993);
nor I_1704 (I31535,I31776,I31911);
nor I_1705 (I31523,I31646,I31911);
not I_1706 (I32079,I3042);
DFFARX1 I_1707 (I594260,I3035,I32079,I32105,);
not I_1708 (I32113,I32105);
nand I_1709 (I32130,I594275,I594254);
and I_1710 (I32147,I32130,I594257);
DFFARX1 I_1711 (I32147,I3035,I32079,I32173,);
DFFARX1 I_1712 (I594278,I3035,I32079,I32190,);
and I_1713 (I32198,I32190,I594257);
nor I_1714 (I32215,I32173,I32198);
DFFARX1 I_1715 (I32215,I3035,I32079,I32047,);
nand I_1716 (I32246,I32190,I594257);
nand I_1717 (I32263,I32113,I32246);
not I_1718 (I32059,I32263);
DFFARX1 I_1719 (I594254,I3035,I32079,I32303,);
DFFARX1 I_1720 (I32303,I3035,I32079,I32068,);
nand I_1721 (I32325,I594266,I594263);
and I_1722 (I32342,I32325,I594269);
DFFARX1 I_1723 (I32342,I3035,I32079,I32368,);
DFFARX1 I_1724 (I32368,I3035,I32079,I32385,);
not I_1725 (I32071,I32385);
not I_1726 (I32407,I32368);
nand I_1727 (I32056,I32407,I32246);
nor I_1728 (I32438,I594272,I594263);
not I_1729 (I32455,I32438);
nor I_1730 (I32472,I32407,I32455);
nor I_1731 (I32489,I32113,I32472);
DFFARX1 I_1732 (I32489,I3035,I32079,I32065,);
nor I_1733 (I32520,I32173,I32455);
nor I_1734 (I32053,I32368,I32520);
nor I_1735 (I32062,I32303,I32438);
nor I_1736 (I32050,I32173,I32438);
not I_1737 (I32606,I3042);
DFFARX1 I_1738 (I469874,I3035,I32606,I32632,);
not I_1739 (I32640,I32632);
nand I_1740 (I32657,I469871,I469886);
and I_1741 (I32674,I32657,I469868);
DFFARX1 I_1742 (I32674,I3035,I32606,I32700,);
DFFARX1 I_1743 (I469865,I3035,I32606,I32717,);
and I_1744 (I32725,I32717,I469865);
nor I_1745 (I32742,I32700,I32725);
DFFARX1 I_1746 (I32742,I3035,I32606,I32574,);
nand I_1747 (I32773,I32717,I469865);
nand I_1748 (I32790,I32640,I32773);
not I_1749 (I32586,I32790);
DFFARX1 I_1750 (I469868,I3035,I32606,I32830,);
DFFARX1 I_1751 (I32830,I3035,I32606,I32595,);
nand I_1752 (I32852,I469880,I469871);
and I_1753 (I32869,I32852,I469883);
DFFARX1 I_1754 (I32869,I3035,I32606,I32895,);
DFFARX1 I_1755 (I32895,I3035,I32606,I32912,);
not I_1756 (I32598,I32912);
not I_1757 (I32934,I32895);
nand I_1758 (I32583,I32934,I32773);
nor I_1759 (I32965,I469877,I469871);
not I_1760 (I32982,I32965);
nor I_1761 (I32999,I32934,I32982);
nor I_1762 (I33016,I32640,I32999);
DFFARX1 I_1763 (I33016,I3035,I32606,I32592,);
nor I_1764 (I33047,I32700,I32982);
nor I_1765 (I32580,I32895,I33047);
nor I_1766 (I32589,I32830,I32965);
nor I_1767 (I32577,I32700,I32965);
not I_1768 (I33133,I3042);
DFFARX1 I_1769 (I1516,I3035,I33133,I33159,);
not I_1770 (I33167,I33159);
nand I_1771 (I33184,I2764,I1524);
and I_1772 (I33201,I33184,I2876);
DFFARX1 I_1773 (I33201,I3035,I33133,I33227,);
DFFARX1 I_1774 (I2588,I3035,I33133,I33244,);
and I_1775 (I33252,I33244,I2996);
nor I_1776 (I33269,I33227,I33252);
DFFARX1 I_1777 (I33269,I3035,I33133,I33101,);
nand I_1778 (I33300,I33244,I2996);
nand I_1779 (I33317,I33167,I33300);
not I_1780 (I33113,I33317);
DFFARX1 I_1781 (I1996,I3035,I33133,I33357,);
DFFARX1 I_1782 (I33357,I3035,I33133,I33122,);
nand I_1783 (I33379,I2948,I1844);
and I_1784 (I33396,I33379,I2580);
DFFARX1 I_1785 (I33396,I3035,I33133,I33422,);
DFFARX1 I_1786 (I33422,I3035,I33133,I33439,);
not I_1787 (I33125,I33439);
not I_1788 (I33461,I33422);
nand I_1789 (I33110,I33461,I33300);
nor I_1790 (I33492,I2908,I1844);
not I_1791 (I33509,I33492);
nor I_1792 (I33526,I33461,I33509);
nor I_1793 (I33543,I33167,I33526);
DFFARX1 I_1794 (I33543,I3035,I33133,I33119,);
nor I_1795 (I33574,I33227,I33509);
nor I_1796 (I33107,I33422,I33574);
nor I_1797 (I33116,I33357,I33492);
nor I_1798 (I33104,I33227,I33492);
not I_1799 (I33660,I3042);
DFFARX1 I_1800 (I216201,I3035,I33660,I33686,);
not I_1801 (I33694,I33686);
nand I_1802 (I33711,I216183,I216198);
and I_1803 (I33728,I33711,I216174);
DFFARX1 I_1804 (I33728,I3035,I33660,I33754,);
DFFARX1 I_1805 (I216177,I3035,I33660,I33771,);
and I_1806 (I33779,I33771,I216192);
nor I_1807 (I33796,I33754,I33779);
DFFARX1 I_1808 (I33796,I3035,I33660,I33628,);
nand I_1809 (I33827,I33771,I216192);
nand I_1810 (I33844,I33694,I33827);
not I_1811 (I33640,I33844);
DFFARX1 I_1812 (I216195,I3035,I33660,I33884,);
DFFARX1 I_1813 (I33884,I3035,I33660,I33649,);
nand I_1814 (I33906,I216174,I216186);
and I_1815 (I33923,I33906,I216180);
DFFARX1 I_1816 (I33923,I3035,I33660,I33949,);
DFFARX1 I_1817 (I33949,I3035,I33660,I33966,);
not I_1818 (I33652,I33966);
not I_1819 (I33988,I33949);
nand I_1820 (I33637,I33988,I33827);
nor I_1821 (I34019,I216189,I216186);
not I_1822 (I34036,I34019);
nor I_1823 (I34053,I33988,I34036);
nor I_1824 (I34070,I33694,I34053);
DFFARX1 I_1825 (I34070,I3035,I33660,I33646,);
nor I_1826 (I34101,I33754,I34036);
nor I_1827 (I33634,I33949,I34101);
nor I_1828 (I33643,I33884,I34019);
nor I_1829 (I33631,I33754,I34019);
not I_1830 (I34187,I3042);
DFFARX1 I_1831 (I450902,I3035,I34187,I34213,);
not I_1832 (I34221,I34213);
nand I_1833 (I34238,I450899,I450914);
and I_1834 (I34255,I34238,I450896);
DFFARX1 I_1835 (I34255,I3035,I34187,I34281,);
DFFARX1 I_1836 (I450893,I3035,I34187,I34298,);
and I_1837 (I34306,I34298,I450893);
nor I_1838 (I34323,I34281,I34306);
DFFARX1 I_1839 (I34323,I3035,I34187,I34155,);
nand I_1840 (I34354,I34298,I450893);
nand I_1841 (I34371,I34221,I34354);
not I_1842 (I34167,I34371);
DFFARX1 I_1843 (I450896,I3035,I34187,I34411,);
DFFARX1 I_1844 (I34411,I3035,I34187,I34176,);
nand I_1845 (I34433,I450908,I450899);
and I_1846 (I34450,I34433,I450911);
DFFARX1 I_1847 (I34450,I3035,I34187,I34476,);
DFFARX1 I_1848 (I34476,I3035,I34187,I34493,);
not I_1849 (I34179,I34493);
not I_1850 (I34515,I34476);
nand I_1851 (I34164,I34515,I34354);
nor I_1852 (I34546,I450905,I450899);
not I_1853 (I34563,I34546);
nor I_1854 (I34580,I34515,I34563);
nor I_1855 (I34597,I34221,I34580);
DFFARX1 I_1856 (I34597,I3035,I34187,I34173,);
nor I_1857 (I34628,I34281,I34563);
nor I_1858 (I34161,I34476,I34628);
nor I_1859 (I34170,I34411,I34546);
nor I_1860 (I34158,I34281,I34546);
not I_1861 (I34714,I3042);
DFFARX1 I_1862 (I105091,I3035,I34714,I34740,);
not I_1863 (I34748,I34740);
nand I_1864 (I34765,I105085,I105079);
and I_1865 (I34782,I34765,I105100);
DFFARX1 I_1866 (I34782,I3035,I34714,I34808,);
DFFARX1 I_1867 (I105097,I3035,I34714,I34825,);
and I_1868 (I34833,I34825,I105094);
nor I_1869 (I34850,I34808,I34833);
DFFARX1 I_1870 (I34850,I3035,I34714,I34682,);
nand I_1871 (I34881,I34825,I105094);
nand I_1872 (I34898,I34748,I34881);
not I_1873 (I34694,I34898);
DFFARX1 I_1874 (I105079,I3035,I34714,I34938,);
DFFARX1 I_1875 (I34938,I3035,I34714,I34703,);
nand I_1876 (I34960,I105082,I105082);
and I_1877 (I34977,I34960,I105103);
DFFARX1 I_1878 (I34977,I3035,I34714,I35003,);
DFFARX1 I_1879 (I35003,I3035,I34714,I35020,);
not I_1880 (I34706,I35020);
not I_1881 (I35042,I35003);
nand I_1882 (I34691,I35042,I34881);
nor I_1883 (I35073,I105088,I105082);
not I_1884 (I35090,I35073);
nor I_1885 (I35107,I35042,I35090);
nor I_1886 (I35124,I34748,I35107);
DFFARX1 I_1887 (I35124,I3035,I34714,I34700,);
nor I_1888 (I35155,I34808,I35090);
nor I_1889 (I34688,I35003,I35155);
nor I_1890 (I34697,I34938,I35073);
nor I_1891 (I34685,I34808,I35073);
not I_1892 (I35241,I3042);
DFFARX1 I_1893 (I139601,I3035,I35241,I35267,);
not I_1894 (I35275,I35267);
nand I_1895 (I35292,I139595,I139589);
and I_1896 (I35309,I35292,I139610);
DFFARX1 I_1897 (I35309,I3035,I35241,I35335,);
DFFARX1 I_1898 (I139607,I3035,I35241,I35352,);
and I_1899 (I35360,I35352,I139604);
nor I_1900 (I35377,I35335,I35360);
DFFARX1 I_1901 (I35377,I3035,I35241,I35209,);
nand I_1902 (I35408,I35352,I139604);
nand I_1903 (I35425,I35275,I35408);
not I_1904 (I35221,I35425);
DFFARX1 I_1905 (I139589,I3035,I35241,I35465,);
DFFARX1 I_1906 (I35465,I3035,I35241,I35230,);
nand I_1907 (I35487,I139592,I139592);
and I_1908 (I35504,I35487,I139613);
DFFARX1 I_1909 (I35504,I3035,I35241,I35530,);
DFFARX1 I_1910 (I35530,I3035,I35241,I35547,);
not I_1911 (I35233,I35547);
not I_1912 (I35569,I35530);
nand I_1913 (I35218,I35569,I35408);
nor I_1914 (I35600,I139598,I139592);
not I_1915 (I35617,I35600);
nor I_1916 (I35634,I35569,I35617);
nor I_1917 (I35651,I35275,I35634);
DFFARX1 I_1918 (I35651,I3035,I35241,I35227,);
nor I_1919 (I35682,I35335,I35617);
nor I_1920 (I35215,I35530,I35682);
nor I_1921 (I35224,I35465,I35600);
nor I_1922 (I35212,I35335,I35600);
not I_1923 (I35768,I3042);
DFFARX1 I_1924 (I416344,I3035,I35768,I35794,);
not I_1925 (I35802,I35794);
nand I_1926 (I35819,I416335,I416353);
and I_1927 (I35836,I35819,I416332);
DFFARX1 I_1928 (I35836,I3035,I35768,I35862,);
DFFARX1 I_1929 (I416335,I3035,I35768,I35879,);
and I_1930 (I35887,I35879,I416338);
nor I_1931 (I35904,I35862,I35887);
DFFARX1 I_1932 (I35904,I3035,I35768,I35736,);
nand I_1933 (I35935,I35879,I416338);
nand I_1934 (I35952,I35802,I35935);
not I_1935 (I35748,I35952);
DFFARX1 I_1936 (I416332,I3035,I35768,I35992,);
DFFARX1 I_1937 (I35992,I3035,I35768,I35757,);
nand I_1938 (I36014,I416350,I416341);
and I_1939 (I36031,I36014,I416356);
DFFARX1 I_1940 (I36031,I3035,I35768,I36057,);
DFFARX1 I_1941 (I36057,I3035,I35768,I36074,);
not I_1942 (I35760,I36074);
not I_1943 (I36096,I36057);
nand I_1944 (I35745,I36096,I35935);
nor I_1945 (I36127,I416347,I416341);
not I_1946 (I36144,I36127);
nor I_1947 (I36161,I36096,I36144);
nor I_1948 (I36178,I35802,I36161);
DFFARX1 I_1949 (I36178,I3035,I35768,I35754,);
nor I_1950 (I36209,I35862,I36144);
nor I_1951 (I35742,I36057,I36209);
nor I_1952 (I35751,I35992,I36127);
nor I_1953 (I35739,I35862,I36127);
not I_1954 (I36295,I3042);
DFFARX1 I_1955 (I323283,I3035,I36295,I36321,);
not I_1956 (I36329,I36321);
nand I_1957 (I36346,I323295,I323280);
and I_1958 (I36363,I36346,I323274);
DFFARX1 I_1959 (I36363,I3035,I36295,I36389,);
DFFARX1 I_1960 (I323289,I3035,I36295,I36406,);
and I_1961 (I36414,I36406,I323277);
nor I_1962 (I36431,I36389,I36414);
DFFARX1 I_1963 (I36431,I3035,I36295,I36263,);
nand I_1964 (I36462,I36406,I323277);
nand I_1965 (I36479,I36329,I36462);
not I_1966 (I36275,I36479);
DFFARX1 I_1967 (I323286,I3035,I36295,I36519,);
DFFARX1 I_1968 (I36519,I3035,I36295,I36284,);
nand I_1969 (I36541,I323292,I323298);
and I_1970 (I36558,I36541,I323274);
DFFARX1 I_1971 (I36558,I3035,I36295,I36584,);
DFFARX1 I_1972 (I36584,I3035,I36295,I36601,);
not I_1973 (I36287,I36601);
not I_1974 (I36623,I36584);
nand I_1975 (I36272,I36623,I36462);
nor I_1976 (I36654,I323277,I323298);
not I_1977 (I36671,I36654);
nor I_1978 (I36688,I36623,I36671);
nor I_1979 (I36705,I36329,I36688);
DFFARX1 I_1980 (I36705,I3035,I36295,I36281,);
nor I_1981 (I36736,I36389,I36671);
nor I_1982 (I36269,I36584,I36736);
nor I_1983 (I36278,I36519,I36654);
nor I_1984 (I36266,I36389,I36654);
not I_1985 (I36822,I3042);
DFFARX1 I_1986 (I356810,I3035,I36822,I36848,);
not I_1987 (I36856,I36848);
nand I_1988 (I36873,I356801,I356819);
and I_1989 (I36890,I36873,I356798);
DFFARX1 I_1990 (I36890,I3035,I36822,I36916,);
DFFARX1 I_1991 (I356801,I3035,I36822,I36933,);
and I_1992 (I36941,I36933,I356804);
nor I_1993 (I36958,I36916,I36941);
DFFARX1 I_1994 (I36958,I3035,I36822,I36790,);
nand I_1995 (I36989,I36933,I356804);
nand I_1996 (I37006,I36856,I36989);
not I_1997 (I36802,I37006);
DFFARX1 I_1998 (I356798,I3035,I36822,I37046,);
DFFARX1 I_1999 (I37046,I3035,I36822,I36811,);
nand I_2000 (I37068,I356816,I356807);
and I_2001 (I37085,I37068,I356822);
DFFARX1 I_2002 (I37085,I3035,I36822,I37111,);
DFFARX1 I_2003 (I37111,I3035,I36822,I37128,);
not I_2004 (I36814,I37128);
not I_2005 (I37150,I37111);
nand I_2006 (I36799,I37150,I36989);
nor I_2007 (I37181,I356813,I356807);
not I_2008 (I37198,I37181);
nor I_2009 (I37215,I37150,I37198);
nor I_2010 (I37232,I36856,I37215);
DFFARX1 I_2011 (I37232,I3035,I36822,I36808,);
nor I_2012 (I37263,I36916,I37198);
nor I_2013 (I36796,I37111,I37263);
nor I_2014 (I36805,I37046,I37181);
nor I_2015 (I36793,I36916,I37181);
not I_2016 (I37349,I3042);
DFFARX1 I_2017 (I540679,I3035,I37349,I37375,);
not I_2018 (I37383,I37375);
nand I_2019 (I37400,I540697,I540691);
and I_2020 (I37417,I37400,I540670);
DFFARX1 I_2021 (I37417,I3035,I37349,I37443,);
DFFARX1 I_2022 (I540688,I3035,I37349,I37460,);
and I_2023 (I37468,I37460,I540673);
nor I_2024 (I37485,I37443,I37468);
DFFARX1 I_2025 (I37485,I3035,I37349,I37317,);
nand I_2026 (I37516,I37460,I540673);
nand I_2027 (I37533,I37383,I37516);
not I_2028 (I37329,I37533);
DFFARX1 I_2029 (I540685,I3035,I37349,I37573,);
DFFARX1 I_2030 (I37573,I3035,I37349,I37338,);
nand I_2031 (I37595,I540694,I540682);
and I_2032 (I37612,I37595,I540676);
DFFARX1 I_2033 (I37612,I3035,I37349,I37638,);
DFFARX1 I_2034 (I37638,I3035,I37349,I37655,);
not I_2035 (I37341,I37655);
not I_2036 (I37677,I37638);
nand I_2037 (I37326,I37677,I37516);
nor I_2038 (I37708,I540670,I540682);
not I_2039 (I37725,I37708);
nor I_2040 (I37742,I37677,I37725);
nor I_2041 (I37759,I37383,I37742);
DFFARX1 I_2042 (I37759,I3035,I37349,I37335,);
nor I_2043 (I37790,I37443,I37725);
nor I_2044 (I37323,I37638,I37790);
nor I_2045 (I37332,I37573,I37708);
nor I_2046 (I37320,I37443,I37708);
not I_2047 (I37876,I3042);
DFFARX1 I_2048 (I554902,I3035,I37876,I37902,);
not I_2049 (I37910,I37902);
nand I_2050 (I37927,I554899,I554905);
and I_2051 (I37944,I37927,I554902);
DFFARX1 I_2052 (I37944,I3035,I37876,I37970,);
DFFARX1 I_2053 (I554905,I3035,I37876,I37987,);
and I_2054 (I37995,I37987,I554899);
nor I_2055 (I38012,I37970,I37995);
DFFARX1 I_2056 (I38012,I3035,I37876,I37844,);
nand I_2057 (I38043,I37987,I554899);
nand I_2058 (I38060,I37910,I38043);
not I_2059 (I37856,I38060);
DFFARX1 I_2060 (I554908,I3035,I37876,I38100,);
DFFARX1 I_2061 (I38100,I3035,I37876,I37865,);
nand I_2062 (I38122,I554911,I554920);
and I_2063 (I38139,I38122,I554914);
DFFARX1 I_2064 (I38139,I3035,I37876,I38165,);
DFFARX1 I_2065 (I38165,I3035,I37876,I38182,);
not I_2066 (I37868,I38182);
not I_2067 (I38204,I38165);
nand I_2068 (I37853,I38204,I38043);
nor I_2069 (I38235,I554917,I554920);
not I_2070 (I38252,I38235);
nor I_2071 (I38269,I38204,I38252);
nor I_2072 (I38286,I37910,I38269);
DFFARX1 I_2073 (I38286,I3035,I37876,I37862,);
nor I_2074 (I38317,I37970,I38252);
nor I_2075 (I37850,I38165,I38317);
nor I_2076 (I37859,I38100,I38235);
nor I_2077 (I37847,I37970,I38235);
not I_2078 (I38403,I3042);
DFFARX1 I_2079 (I80696,I3035,I38403,I38429,);
not I_2080 (I38437,I38429);
nand I_2081 (I38454,I80690,I80684);
and I_2082 (I38471,I38454,I80705);
DFFARX1 I_2083 (I38471,I3035,I38403,I38497,);
DFFARX1 I_2084 (I80702,I3035,I38403,I38514,);
and I_2085 (I38522,I38514,I80699);
nor I_2086 (I38539,I38497,I38522);
DFFARX1 I_2087 (I38539,I3035,I38403,I38371,);
nand I_2088 (I38570,I38514,I80699);
nand I_2089 (I38587,I38437,I38570);
not I_2090 (I38383,I38587);
DFFARX1 I_2091 (I80684,I3035,I38403,I38627,);
DFFARX1 I_2092 (I38627,I3035,I38403,I38392,);
nand I_2093 (I38649,I80687,I80687);
and I_2094 (I38666,I38649,I80708);
DFFARX1 I_2095 (I38666,I3035,I38403,I38692,);
DFFARX1 I_2096 (I38692,I3035,I38403,I38709,);
not I_2097 (I38395,I38709);
not I_2098 (I38731,I38692);
nand I_2099 (I38380,I38731,I38570);
nor I_2100 (I38762,I80693,I80687);
not I_2101 (I38779,I38762);
nor I_2102 (I38796,I38731,I38779);
nor I_2103 (I38813,I38437,I38796);
DFFARX1 I_2104 (I38813,I3035,I38403,I38389,);
nor I_2105 (I38844,I38497,I38779);
nor I_2106 (I38377,I38692,I38844);
nor I_2107 (I38386,I38627,I38762);
nor I_2108 (I38374,I38497,I38762);
not I_2109 (I38930,I3042);
DFFARX1 I_2110 (I10464,I3035,I38930,I38956,);
not I_2111 (I38964,I38956);
nand I_2112 (I38981,I10452,I10458);
and I_2113 (I38998,I38981,I10461);
DFFARX1 I_2114 (I38998,I3035,I38930,I39024,);
DFFARX1 I_2115 (I10443,I3035,I38930,I39041,);
and I_2116 (I39049,I39041,I10449);
nor I_2117 (I39066,I39024,I39049);
DFFARX1 I_2118 (I39066,I3035,I38930,I38898,);
nand I_2119 (I39097,I39041,I10449);
nand I_2120 (I39114,I38964,I39097);
not I_2121 (I38910,I39114);
DFFARX1 I_2122 (I10443,I3035,I38930,I39154,);
DFFARX1 I_2123 (I39154,I3035,I38930,I38919,);
nand I_2124 (I39176,I10446,I10440);
and I_2125 (I39193,I39176,I10455);
DFFARX1 I_2126 (I39193,I3035,I38930,I39219,);
DFFARX1 I_2127 (I39219,I3035,I38930,I39236,);
not I_2128 (I38922,I39236);
not I_2129 (I39258,I39219);
nand I_2130 (I38907,I39258,I39097);
nor I_2131 (I39289,I10440,I10440);
not I_2132 (I39306,I39289);
nor I_2133 (I39323,I39258,I39306);
nor I_2134 (I39340,I38964,I39323);
DFFARX1 I_2135 (I39340,I3035,I38930,I38916,);
nor I_2136 (I39371,I39024,I39306);
nor I_2137 (I38904,I39219,I39371);
nor I_2138 (I38913,I39154,I39289);
nor I_2139 (I38901,I39024,I39289);
not I_2140 (I39457,I3042);
DFFARX1 I_2141 (I446159,I3035,I39457,I39483,);
not I_2142 (I39491,I39483);
nand I_2143 (I39508,I446156,I446171);
and I_2144 (I39525,I39508,I446153);
DFFARX1 I_2145 (I39525,I3035,I39457,I39551,);
DFFARX1 I_2146 (I446150,I3035,I39457,I39568,);
and I_2147 (I39576,I39568,I446150);
nor I_2148 (I39593,I39551,I39576);
DFFARX1 I_2149 (I39593,I3035,I39457,I39425,);
nand I_2150 (I39624,I39568,I446150);
nand I_2151 (I39641,I39491,I39624);
not I_2152 (I39437,I39641);
DFFARX1 I_2153 (I446153,I3035,I39457,I39681,);
DFFARX1 I_2154 (I39681,I3035,I39457,I39446,);
nand I_2155 (I39703,I446165,I446156);
and I_2156 (I39720,I39703,I446168);
DFFARX1 I_2157 (I39720,I3035,I39457,I39746,);
DFFARX1 I_2158 (I39746,I3035,I39457,I39763,);
not I_2159 (I39449,I39763);
not I_2160 (I39785,I39746);
nand I_2161 (I39434,I39785,I39624);
nor I_2162 (I39816,I446162,I446156);
not I_2163 (I39833,I39816);
nor I_2164 (I39850,I39785,I39833);
nor I_2165 (I39867,I39491,I39850);
DFFARX1 I_2166 (I39867,I3035,I39457,I39443,);
nor I_2167 (I39898,I39551,I39833);
nor I_2168 (I39431,I39746,I39898);
nor I_2169 (I39440,I39681,I39816);
nor I_2170 (I39428,I39551,I39816);
not I_2171 (I39984,I3042);
DFFARX1 I_2172 (I189851,I3035,I39984,I40010,);
not I_2173 (I40018,I40010);
nand I_2174 (I40035,I189833,I189848);
and I_2175 (I40052,I40035,I189824);
DFFARX1 I_2176 (I40052,I3035,I39984,I40078,);
DFFARX1 I_2177 (I189827,I3035,I39984,I40095,);
and I_2178 (I40103,I40095,I189842);
nor I_2179 (I40120,I40078,I40103);
DFFARX1 I_2180 (I40120,I3035,I39984,I39952,);
nand I_2181 (I40151,I40095,I189842);
nand I_2182 (I40168,I40018,I40151);
not I_2183 (I39964,I40168);
DFFARX1 I_2184 (I189845,I3035,I39984,I40208,);
DFFARX1 I_2185 (I40208,I3035,I39984,I39973,);
nand I_2186 (I40230,I189824,I189836);
and I_2187 (I40247,I40230,I189830);
DFFARX1 I_2188 (I40247,I3035,I39984,I40273,);
DFFARX1 I_2189 (I40273,I3035,I39984,I40290,);
not I_2190 (I39976,I40290);
not I_2191 (I40312,I40273);
nand I_2192 (I39961,I40312,I40151);
nor I_2193 (I40343,I189839,I189836);
not I_2194 (I40360,I40343);
nor I_2195 (I40377,I40312,I40360);
nor I_2196 (I40394,I40018,I40377);
DFFARX1 I_2197 (I40394,I3035,I39984,I39970,);
nor I_2198 (I40425,I40078,I40360);
nor I_2199 (I39958,I40273,I40425);
nor I_2200 (I39967,I40208,I40343);
nor I_2201 (I39955,I40078,I40343);
not I_2202 (I40511,I3042);
DFFARX1 I_2203 (I659948,I3035,I40511,I40537,);
not I_2204 (I40545,I40537);
nand I_2205 (I40562,I659942,I659963);
and I_2206 (I40579,I40562,I659954);
DFFARX1 I_2207 (I40579,I3035,I40511,I40605,);
DFFARX1 I_2208 (I659945,I3035,I40511,I40622,);
and I_2209 (I40630,I40622,I659957);
nor I_2210 (I40647,I40605,I40630);
DFFARX1 I_2211 (I40647,I3035,I40511,I40479,);
nand I_2212 (I40678,I40622,I659957);
nand I_2213 (I40695,I40545,I40678);
not I_2214 (I40491,I40695);
DFFARX1 I_2215 (I659945,I3035,I40511,I40735,);
DFFARX1 I_2216 (I40735,I3035,I40511,I40500,);
nand I_2217 (I40757,I659966,I659951);
and I_2218 (I40774,I40757,I659942);
DFFARX1 I_2219 (I40774,I3035,I40511,I40800,);
DFFARX1 I_2220 (I40800,I3035,I40511,I40817,);
not I_2221 (I40503,I40817);
not I_2222 (I40839,I40800);
nand I_2223 (I40488,I40839,I40678);
nor I_2224 (I40870,I659960,I659951);
not I_2225 (I40887,I40870);
nor I_2226 (I40904,I40839,I40887);
nor I_2227 (I40921,I40545,I40904);
DFFARX1 I_2228 (I40921,I3035,I40511,I40497,);
nor I_2229 (I40952,I40605,I40887);
nor I_2230 (I40485,I40800,I40952);
nor I_2231 (I40494,I40735,I40870);
nor I_2232 (I40482,I40605,I40870);
not I_2233 (I41038,I3042);
DFFARX1 I_2234 (I13099,I3035,I41038,I41064,);
not I_2235 (I41072,I41064);
nand I_2236 (I41089,I13087,I13093);
and I_2237 (I41106,I41089,I13096);
DFFARX1 I_2238 (I41106,I3035,I41038,I41132,);
DFFARX1 I_2239 (I13078,I3035,I41038,I41149,);
and I_2240 (I41157,I41149,I13084);
nor I_2241 (I41174,I41132,I41157);
DFFARX1 I_2242 (I41174,I3035,I41038,I41006,);
nand I_2243 (I41205,I41149,I13084);
nand I_2244 (I41222,I41072,I41205);
not I_2245 (I41018,I41222);
DFFARX1 I_2246 (I13078,I3035,I41038,I41262,);
DFFARX1 I_2247 (I41262,I3035,I41038,I41027,);
nand I_2248 (I41284,I13081,I13075);
and I_2249 (I41301,I41284,I13090);
DFFARX1 I_2250 (I41301,I3035,I41038,I41327,);
DFFARX1 I_2251 (I41327,I3035,I41038,I41344,);
not I_2252 (I41030,I41344);
not I_2253 (I41366,I41327);
nand I_2254 (I41015,I41366,I41205);
nor I_2255 (I41397,I13075,I13075);
not I_2256 (I41414,I41397);
nor I_2257 (I41431,I41366,I41414);
nor I_2258 (I41448,I41072,I41431);
DFFARX1 I_2259 (I41448,I3035,I41038,I41024,);
nor I_2260 (I41479,I41132,I41414);
nor I_2261 (I41012,I41327,I41479);
nor I_2262 (I41021,I41262,I41397);
nor I_2263 (I41009,I41132,I41397);
not I_2264 (I41565,I3042);
DFFARX1 I_2265 (I609288,I3035,I41565,I41591,);
not I_2266 (I41599,I41591);
nand I_2267 (I41616,I609303,I609282);
and I_2268 (I41633,I41616,I609285);
DFFARX1 I_2269 (I41633,I3035,I41565,I41659,);
DFFARX1 I_2270 (I609306,I3035,I41565,I41676,);
and I_2271 (I41684,I41676,I609285);
nor I_2272 (I41701,I41659,I41684);
DFFARX1 I_2273 (I41701,I3035,I41565,I41533,);
nand I_2274 (I41732,I41676,I609285);
nand I_2275 (I41749,I41599,I41732);
not I_2276 (I41545,I41749);
DFFARX1 I_2277 (I609282,I3035,I41565,I41789,);
DFFARX1 I_2278 (I41789,I3035,I41565,I41554,);
nand I_2279 (I41811,I609294,I609291);
and I_2280 (I41828,I41811,I609297);
DFFARX1 I_2281 (I41828,I3035,I41565,I41854,);
DFFARX1 I_2282 (I41854,I3035,I41565,I41871,);
not I_2283 (I41557,I41871);
not I_2284 (I41893,I41854);
nand I_2285 (I41542,I41893,I41732);
nor I_2286 (I41924,I609300,I609291);
not I_2287 (I41941,I41924);
nor I_2288 (I41958,I41893,I41941);
nor I_2289 (I41975,I41599,I41958);
DFFARX1 I_2290 (I41975,I3035,I41565,I41551,);
nor I_2291 (I42006,I41659,I41941);
nor I_2292 (I41539,I41854,I42006);
nor I_2293 (I41548,I41789,I41924);
nor I_2294 (I41536,I41659,I41924);
not I_2295 (I42092,I3042);
DFFARX1 I_2296 (I650700,I3035,I42092,I42118,);
not I_2297 (I42126,I42118);
nand I_2298 (I42143,I650694,I650715);
and I_2299 (I42160,I42143,I650706);
DFFARX1 I_2300 (I42160,I3035,I42092,I42186,);
DFFARX1 I_2301 (I650697,I3035,I42092,I42203,);
and I_2302 (I42211,I42203,I650709);
nor I_2303 (I42228,I42186,I42211);
DFFARX1 I_2304 (I42228,I3035,I42092,I42060,);
nand I_2305 (I42259,I42203,I650709);
nand I_2306 (I42276,I42126,I42259);
not I_2307 (I42072,I42276);
DFFARX1 I_2308 (I650697,I3035,I42092,I42316,);
DFFARX1 I_2309 (I42316,I3035,I42092,I42081,);
nand I_2310 (I42338,I650718,I650703);
and I_2311 (I42355,I42338,I650694);
DFFARX1 I_2312 (I42355,I3035,I42092,I42381,);
DFFARX1 I_2313 (I42381,I3035,I42092,I42398,);
not I_2314 (I42084,I42398);
not I_2315 (I42420,I42381);
nand I_2316 (I42069,I42420,I42259);
nor I_2317 (I42451,I650712,I650703);
not I_2318 (I42468,I42451);
nor I_2319 (I42485,I42420,I42468);
nor I_2320 (I42502,I42126,I42485);
DFFARX1 I_2321 (I42502,I3035,I42092,I42078,);
nor I_2322 (I42533,I42186,I42468);
nor I_2323 (I42066,I42381,I42533);
nor I_2324 (I42075,I42316,I42451);
nor I_2325 (I42063,I42186,I42451);
not I_2326 (I42619,I3042);
DFFARX1 I_2327 (I552097,I3035,I42619,I42645,);
not I_2328 (I42653,I42645);
nand I_2329 (I42670,I552094,I552100);
and I_2330 (I42687,I42670,I552097);
DFFARX1 I_2331 (I42687,I3035,I42619,I42713,);
DFFARX1 I_2332 (I552100,I3035,I42619,I42730,);
and I_2333 (I42738,I42730,I552094);
nor I_2334 (I42755,I42713,I42738);
DFFARX1 I_2335 (I42755,I3035,I42619,I42587,);
nand I_2336 (I42786,I42730,I552094);
nand I_2337 (I42803,I42653,I42786);
not I_2338 (I42599,I42803);
DFFARX1 I_2339 (I552103,I3035,I42619,I42843,);
DFFARX1 I_2340 (I42843,I3035,I42619,I42608,);
nand I_2341 (I42865,I552106,I552115);
and I_2342 (I42882,I42865,I552109);
DFFARX1 I_2343 (I42882,I3035,I42619,I42908,);
DFFARX1 I_2344 (I42908,I3035,I42619,I42925,);
not I_2345 (I42611,I42925);
not I_2346 (I42947,I42908);
nand I_2347 (I42596,I42947,I42786);
nor I_2348 (I42978,I552112,I552115);
not I_2349 (I42995,I42978);
nor I_2350 (I43012,I42947,I42995);
nor I_2351 (I43029,I42653,I43012);
DFFARX1 I_2352 (I43029,I3035,I42619,I42605,);
nor I_2353 (I43060,I42713,I42995);
nor I_2354 (I42593,I42908,I43060);
nor I_2355 (I42602,I42843,I42978);
nor I_2356 (I42590,I42713,I42978);
not I_2357 (I43146,I3042);
DFFARX1 I_2358 (I223579,I3035,I43146,I43172,);
not I_2359 (I43180,I43172);
nand I_2360 (I43197,I223561,I223576);
and I_2361 (I43214,I43197,I223552);
DFFARX1 I_2362 (I43214,I3035,I43146,I43240,);
DFFARX1 I_2363 (I223555,I3035,I43146,I43257,);
and I_2364 (I43265,I43257,I223570);
nor I_2365 (I43282,I43240,I43265);
DFFARX1 I_2366 (I43282,I3035,I43146,I43114,);
nand I_2367 (I43313,I43257,I223570);
nand I_2368 (I43330,I43180,I43313);
not I_2369 (I43126,I43330);
DFFARX1 I_2370 (I223573,I3035,I43146,I43370,);
DFFARX1 I_2371 (I43370,I3035,I43146,I43135,);
nand I_2372 (I43392,I223552,I223564);
and I_2373 (I43409,I43392,I223558);
DFFARX1 I_2374 (I43409,I3035,I43146,I43435,);
DFFARX1 I_2375 (I43435,I3035,I43146,I43452,);
not I_2376 (I43138,I43452);
not I_2377 (I43474,I43435);
nand I_2378 (I43123,I43474,I43313);
nor I_2379 (I43505,I223567,I223564);
not I_2380 (I43522,I43505);
nor I_2381 (I43539,I43474,I43522);
nor I_2382 (I43556,I43180,I43539);
DFFARX1 I_2383 (I43556,I3035,I43146,I43132,);
nor I_2384 (I43587,I43240,I43522);
nor I_2385 (I43120,I43435,I43587);
nor I_2386 (I43129,I43370,I43505);
nor I_2387 (I43117,I43240,I43505);
not I_2388 (I43673,I3042);
DFFARX1 I_2389 (I331953,I3035,I43673,I43699,);
not I_2390 (I43707,I43699);
nand I_2391 (I43724,I331965,I331950);
and I_2392 (I43741,I43724,I331944);
DFFARX1 I_2393 (I43741,I3035,I43673,I43767,);
DFFARX1 I_2394 (I331959,I3035,I43673,I43784,);
and I_2395 (I43792,I43784,I331947);
nor I_2396 (I43809,I43767,I43792);
DFFARX1 I_2397 (I43809,I3035,I43673,I43641,);
nand I_2398 (I43840,I43784,I331947);
nand I_2399 (I43857,I43707,I43840);
not I_2400 (I43653,I43857);
DFFARX1 I_2401 (I331956,I3035,I43673,I43897,);
DFFARX1 I_2402 (I43897,I3035,I43673,I43662,);
nand I_2403 (I43919,I331962,I331968);
and I_2404 (I43936,I43919,I331944);
DFFARX1 I_2405 (I43936,I3035,I43673,I43962,);
DFFARX1 I_2406 (I43962,I3035,I43673,I43979,);
not I_2407 (I43665,I43979);
not I_2408 (I44001,I43962);
nand I_2409 (I43650,I44001,I43840);
nor I_2410 (I44032,I331947,I331968);
not I_2411 (I44049,I44032);
nor I_2412 (I44066,I44001,I44049);
nor I_2413 (I44083,I43707,I44066);
DFFARX1 I_2414 (I44083,I3035,I43673,I43659,);
nor I_2415 (I44114,I43767,I44049);
nor I_2416 (I43647,I43962,I44114);
nor I_2417 (I43656,I43897,I44032);
nor I_2418 (I43644,I43767,I44032);
not I_2419 (I44200,I3042);
DFFARX1 I_2420 (I240791,I3035,I44200,I44226,);
not I_2421 (I44234,I44226);
nand I_2422 (I44251,I240785,I240776);
and I_2423 (I44268,I44251,I240797);
DFFARX1 I_2424 (I44268,I3035,I44200,I44294,);
DFFARX1 I_2425 (I240779,I3035,I44200,I44311,);
and I_2426 (I44319,I44311,I240773);
nor I_2427 (I44336,I44294,I44319);
DFFARX1 I_2428 (I44336,I3035,I44200,I44168,);
nand I_2429 (I44367,I44311,I240773);
nand I_2430 (I44384,I44234,I44367);
not I_2431 (I44180,I44384);
DFFARX1 I_2432 (I240773,I3035,I44200,I44424,);
DFFARX1 I_2433 (I44424,I3035,I44200,I44189,);
nand I_2434 (I44446,I240800,I240782);
and I_2435 (I44463,I44446,I240788);
DFFARX1 I_2436 (I44463,I3035,I44200,I44489,);
DFFARX1 I_2437 (I44489,I3035,I44200,I44506,);
not I_2438 (I44192,I44506);
not I_2439 (I44528,I44489);
nand I_2440 (I44177,I44528,I44367);
nor I_2441 (I44559,I240794,I240782);
not I_2442 (I44576,I44559);
nor I_2443 (I44593,I44528,I44576);
nor I_2444 (I44610,I44234,I44593);
DFFARX1 I_2445 (I44610,I3035,I44200,I44186,);
nor I_2446 (I44641,I44294,I44576);
nor I_2447 (I44174,I44489,I44641);
nor I_2448 (I44183,I44424,I44559);
nor I_2449 (I44171,I44294,I44559);
not I_2450 (I44727,I3042);
DFFARX1 I_2451 (I431930,I3035,I44727,I44753,);
not I_2452 (I44761,I44753);
nand I_2453 (I44778,I431927,I431942);
and I_2454 (I44795,I44778,I431924);
DFFARX1 I_2455 (I44795,I3035,I44727,I44821,);
DFFARX1 I_2456 (I431921,I3035,I44727,I44838,);
and I_2457 (I44846,I44838,I431921);
nor I_2458 (I44863,I44821,I44846);
DFFARX1 I_2459 (I44863,I3035,I44727,I44695,);
nand I_2460 (I44894,I44838,I431921);
nand I_2461 (I44911,I44761,I44894);
not I_2462 (I44707,I44911);
DFFARX1 I_2463 (I431924,I3035,I44727,I44951,);
DFFARX1 I_2464 (I44951,I3035,I44727,I44716,);
nand I_2465 (I44973,I431936,I431927);
and I_2466 (I44990,I44973,I431939);
DFFARX1 I_2467 (I44990,I3035,I44727,I45016,);
DFFARX1 I_2468 (I45016,I3035,I44727,I45033,);
not I_2469 (I44719,I45033);
not I_2470 (I45055,I45016);
nand I_2471 (I44704,I45055,I44894);
nor I_2472 (I45086,I431933,I431927);
not I_2473 (I45103,I45086);
nor I_2474 (I45120,I45055,I45103);
nor I_2475 (I45137,I44761,I45120);
DFFARX1 I_2476 (I45137,I3035,I44727,I44713,);
nor I_2477 (I45168,I44821,I45103);
nor I_2478 (I44701,I45016,I45168);
nor I_2479 (I44710,I44951,I45086);
nor I_2480 (I44698,I44821,I45086);
not I_2481 (I45254,I3042);
DFFARX1 I_2482 (I688693,I3035,I45254,I45280,);
not I_2483 (I45288,I45280);
nand I_2484 (I45305,I688696,I688690);
and I_2485 (I45322,I45305,I688687);
DFFARX1 I_2486 (I45322,I3035,I45254,I45348,);
DFFARX1 I_2487 (I688672,I3035,I45254,I45365,);
and I_2488 (I45373,I45365,I688681);
nor I_2489 (I45390,I45348,I45373);
DFFARX1 I_2490 (I45390,I3035,I45254,I45222,);
nand I_2491 (I45421,I45365,I688681);
nand I_2492 (I45438,I45288,I45421);
not I_2493 (I45234,I45438);
DFFARX1 I_2494 (I688672,I3035,I45254,I45478,);
DFFARX1 I_2495 (I45478,I3035,I45254,I45243,);
nand I_2496 (I45500,I688675,I688678);
and I_2497 (I45517,I45500,I688684);
DFFARX1 I_2498 (I45517,I3035,I45254,I45543,);
DFFARX1 I_2499 (I45543,I3035,I45254,I45560,);
not I_2500 (I45246,I45560);
not I_2501 (I45582,I45543);
nand I_2502 (I45231,I45582,I45421);
nor I_2503 (I45613,I688675,I688678);
not I_2504 (I45630,I45613);
nor I_2505 (I45647,I45582,I45630);
nor I_2506 (I45664,I45288,I45647);
DFFARX1 I_2507 (I45664,I3035,I45254,I45240,);
nor I_2508 (I45695,I45348,I45630);
nor I_2509 (I45228,I45543,I45695);
nor I_2510 (I45237,I45478,I45613);
nor I_2511 (I45225,I45348,I45613);
not I_2512 (I45781,I3042);
DFFARX1 I_2513 (I536803,I3035,I45781,I45807,);
not I_2514 (I45815,I45807);
nand I_2515 (I45832,I536821,I536815);
and I_2516 (I45849,I45832,I536794);
DFFARX1 I_2517 (I45849,I3035,I45781,I45875,);
DFFARX1 I_2518 (I536812,I3035,I45781,I45892,);
and I_2519 (I45900,I45892,I536797);
nor I_2520 (I45917,I45875,I45900);
DFFARX1 I_2521 (I45917,I3035,I45781,I45749,);
nand I_2522 (I45948,I45892,I536797);
nand I_2523 (I45965,I45815,I45948);
not I_2524 (I45761,I45965);
DFFARX1 I_2525 (I536809,I3035,I45781,I46005,);
DFFARX1 I_2526 (I46005,I3035,I45781,I45770,);
nand I_2527 (I46027,I536818,I536806);
and I_2528 (I46044,I46027,I536800);
DFFARX1 I_2529 (I46044,I3035,I45781,I46070,);
DFFARX1 I_2530 (I46070,I3035,I45781,I46087,);
not I_2531 (I45773,I46087);
not I_2532 (I46109,I46070);
nand I_2533 (I45758,I46109,I45948);
nor I_2534 (I46140,I536794,I536806);
not I_2535 (I46157,I46140);
nor I_2536 (I46174,I46109,I46157);
nor I_2537 (I46191,I45815,I46174);
DFFARX1 I_2538 (I46191,I3035,I45781,I45767,);
nor I_2539 (I46222,I45875,I46157);
nor I_2540 (I45755,I46070,I46222);
nor I_2541 (I45764,I46005,I46140);
nor I_2542 (I45752,I45875,I46140);
not I_2543 (I46308,I3042);
DFFARX1 I_2544 (I730555,I3035,I46308,I46334,);
not I_2545 (I46342,I46334);
nand I_2546 (I46359,I730549,I730570);
and I_2547 (I46376,I46359,I730546);
DFFARX1 I_2548 (I46376,I3035,I46308,I46402,);
DFFARX1 I_2549 (I730567,I3035,I46308,I46419,);
and I_2550 (I46427,I46419,I730564);
nor I_2551 (I46444,I46402,I46427);
DFFARX1 I_2552 (I46444,I3035,I46308,I46276,);
nand I_2553 (I46475,I46419,I730564);
nand I_2554 (I46492,I46342,I46475);
not I_2555 (I46288,I46492);
DFFARX1 I_2556 (I730552,I3035,I46308,I46532,);
DFFARX1 I_2557 (I46532,I3035,I46308,I46297,);
nand I_2558 (I46554,I730561,I730558);
and I_2559 (I46571,I46554,I730543);
DFFARX1 I_2560 (I46571,I3035,I46308,I46597,);
DFFARX1 I_2561 (I46597,I3035,I46308,I46614,);
not I_2562 (I46300,I46614);
not I_2563 (I46636,I46597);
nand I_2564 (I46285,I46636,I46475);
nor I_2565 (I46667,I730543,I730558);
not I_2566 (I46684,I46667);
nor I_2567 (I46701,I46636,I46684);
nor I_2568 (I46718,I46342,I46701);
DFFARX1 I_2569 (I46718,I3035,I46308,I46294,);
nor I_2570 (I46749,I46402,I46684);
nor I_2571 (I46282,I46597,I46749);
nor I_2572 (I46291,I46532,I46667);
nor I_2573 (I46279,I46402,I46667);
not I_2574 (I46835,I3042);
DFFARX1 I_2575 (I597150,I3035,I46835,I46861,);
not I_2576 (I46869,I46861);
nand I_2577 (I46886,I597165,I597144);
and I_2578 (I46903,I46886,I597147);
DFFARX1 I_2579 (I46903,I3035,I46835,I46929,);
DFFARX1 I_2580 (I597168,I3035,I46835,I46946,);
and I_2581 (I46954,I46946,I597147);
nor I_2582 (I46971,I46929,I46954);
DFFARX1 I_2583 (I46971,I3035,I46835,I46803,);
nand I_2584 (I47002,I46946,I597147);
nand I_2585 (I47019,I46869,I47002);
not I_2586 (I46815,I47019);
DFFARX1 I_2587 (I597144,I3035,I46835,I47059,);
DFFARX1 I_2588 (I47059,I3035,I46835,I46824,);
nand I_2589 (I47081,I597156,I597153);
and I_2590 (I47098,I47081,I597159);
DFFARX1 I_2591 (I47098,I3035,I46835,I47124,);
DFFARX1 I_2592 (I47124,I3035,I46835,I47141,);
not I_2593 (I46827,I47141);
not I_2594 (I47163,I47124);
nand I_2595 (I46812,I47163,I47002);
nor I_2596 (I47194,I597162,I597153);
not I_2597 (I47211,I47194);
nor I_2598 (I47228,I47163,I47211);
nor I_2599 (I47245,I46869,I47228);
DFFARX1 I_2600 (I47245,I3035,I46835,I46821,);
nor I_2601 (I47276,I46929,I47211);
nor I_2602 (I46809,I47124,I47276);
nor I_2603 (I46818,I47059,I47194);
nor I_2604 (I46806,I46929,I47194);
not I_2605 (I47362,I3042);
DFFARX1 I_2606 (I326173,I3035,I47362,I47388,);
not I_2607 (I47396,I47388);
nand I_2608 (I47413,I326185,I326170);
and I_2609 (I47430,I47413,I326164);
DFFARX1 I_2610 (I47430,I3035,I47362,I47456,);
DFFARX1 I_2611 (I326179,I3035,I47362,I47473,);
and I_2612 (I47481,I47473,I326167);
nor I_2613 (I47498,I47456,I47481);
DFFARX1 I_2614 (I47498,I3035,I47362,I47330,);
nand I_2615 (I47529,I47473,I326167);
nand I_2616 (I47546,I47396,I47529);
not I_2617 (I47342,I47546);
DFFARX1 I_2618 (I326176,I3035,I47362,I47586,);
DFFARX1 I_2619 (I47586,I3035,I47362,I47351,);
nand I_2620 (I47608,I326182,I326188);
and I_2621 (I47625,I47608,I326164);
DFFARX1 I_2622 (I47625,I3035,I47362,I47651,);
DFFARX1 I_2623 (I47651,I3035,I47362,I47668,);
not I_2624 (I47354,I47668);
not I_2625 (I47690,I47651);
nand I_2626 (I47339,I47690,I47529);
nor I_2627 (I47721,I326167,I326188);
not I_2628 (I47738,I47721);
nor I_2629 (I47755,I47690,I47738);
nor I_2630 (I47772,I47396,I47755);
DFFARX1 I_2631 (I47772,I3035,I47362,I47348,);
nor I_2632 (I47803,I47456,I47738);
nor I_2633 (I47336,I47651,I47803);
nor I_2634 (I47345,I47586,I47721);
nor I_2635 (I47333,I47456,I47721);
not I_2636 (I47889,I3042);
DFFARX1 I_2637 (I204607,I3035,I47889,I47915,);
not I_2638 (I47923,I47915);
nand I_2639 (I47940,I204589,I204604);
and I_2640 (I47957,I47940,I204580);
DFFARX1 I_2641 (I47957,I3035,I47889,I47983,);
DFFARX1 I_2642 (I204583,I3035,I47889,I48000,);
and I_2643 (I48008,I48000,I204598);
nor I_2644 (I48025,I47983,I48008);
DFFARX1 I_2645 (I48025,I3035,I47889,I47857,);
nand I_2646 (I48056,I48000,I204598);
nand I_2647 (I48073,I47923,I48056);
not I_2648 (I47869,I48073);
DFFARX1 I_2649 (I204601,I3035,I47889,I48113,);
DFFARX1 I_2650 (I48113,I3035,I47889,I47878,);
nand I_2651 (I48135,I204580,I204592);
and I_2652 (I48152,I48135,I204586);
DFFARX1 I_2653 (I48152,I3035,I47889,I48178,);
DFFARX1 I_2654 (I48178,I3035,I47889,I48195,);
not I_2655 (I47881,I48195);
not I_2656 (I48217,I48178);
nand I_2657 (I47866,I48217,I48056);
nor I_2658 (I48248,I204595,I204592);
not I_2659 (I48265,I48248);
nor I_2660 (I48282,I48217,I48265);
nor I_2661 (I48299,I47923,I48282);
DFFARX1 I_2662 (I48299,I3035,I47889,I47875,);
nor I_2663 (I48330,I47983,I48265);
nor I_2664 (I47863,I48178,I48330);
nor I_2665 (I47872,I48113,I48248);
nor I_2666 (I47860,I47983,I48248);
not I_2667 (I48416,I3042);
DFFARX1 I_2668 (I172460,I3035,I48416,I48442,);
not I_2669 (I48450,I48442);
nand I_2670 (I48467,I172442,I172457);
and I_2671 (I48484,I48467,I172433);
DFFARX1 I_2672 (I48484,I3035,I48416,I48510,);
DFFARX1 I_2673 (I172436,I3035,I48416,I48527,);
and I_2674 (I48535,I48527,I172451);
nor I_2675 (I48552,I48510,I48535);
DFFARX1 I_2676 (I48552,I3035,I48416,I48384,);
nand I_2677 (I48583,I48527,I172451);
nand I_2678 (I48600,I48450,I48583);
not I_2679 (I48396,I48600);
DFFARX1 I_2680 (I172454,I3035,I48416,I48640,);
DFFARX1 I_2681 (I48640,I3035,I48416,I48405,);
nand I_2682 (I48662,I172433,I172445);
and I_2683 (I48679,I48662,I172439);
DFFARX1 I_2684 (I48679,I3035,I48416,I48705,);
DFFARX1 I_2685 (I48705,I3035,I48416,I48722,);
not I_2686 (I48408,I48722);
not I_2687 (I48744,I48705);
nand I_2688 (I48393,I48744,I48583);
nor I_2689 (I48775,I172448,I172445);
not I_2690 (I48792,I48775);
nor I_2691 (I48809,I48744,I48792);
nor I_2692 (I48826,I48450,I48809);
DFFARX1 I_2693 (I48826,I3035,I48416,I48402,);
nor I_2694 (I48857,I48510,I48792);
nor I_2695 (I48390,I48705,I48857);
nor I_2696 (I48399,I48640,I48775);
nor I_2697 (I48387,I48510,I48775);
not I_2698 (I48943,I3042);
DFFARX1 I_2699 (I76540,I3035,I48943,I48969,);
not I_2700 (I48977,I48969);
nand I_2701 (I48994,I76537,I76519);
and I_2702 (I49011,I48994,I76525);
DFFARX1 I_2703 (I49011,I3035,I48943,I49037,);
DFFARX1 I_2704 (I76534,I3035,I48943,I49054,);
and I_2705 (I49062,I49054,I76528);
nor I_2706 (I49079,I49037,I49062);
DFFARX1 I_2707 (I49079,I3035,I48943,I48911,);
nand I_2708 (I49110,I49054,I76528);
nand I_2709 (I49127,I48977,I49110);
not I_2710 (I48923,I49127);
DFFARX1 I_2711 (I76543,I3035,I48943,I49167,);
DFFARX1 I_2712 (I49167,I3035,I48943,I48932,);
nand I_2713 (I49189,I76531,I76522);
and I_2714 (I49206,I49189,I76519);
DFFARX1 I_2715 (I49206,I3035,I48943,I49232,);
DFFARX1 I_2716 (I49232,I3035,I48943,I49249,);
not I_2717 (I48935,I49249);
not I_2718 (I49271,I49232);
nand I_2719 (I48920,I49271,I49110);
nor I_2720 (I49302,I76546,I76522);
not I_2721 (I49319,I49302);
nor I_2722 (I49336,I49271,I49319);
nor I_2723 (I49353,I48977,I49336);
DFFARX1 I_2724 (I49353,I3035,I48943,I48929,);
nor I_2725 (I49384,I49037,I49319);
nor I_2726 (I48917,I49232,I49384);
nor I_2727 (I48926,I49167,I49302);
nor I_2728 (I48914,I49037,I49302);
not I_2729 (I49470,I3042);
DFFARX1 I_2730 (I174041,I3035,I49470,I49496,);
not I_2731 (I49504,I49496);
nand I_2732 (I49521,I174023,I174038);
and I_2733 (I49538,I49521,I174014);
DFFARX1 I_2734 (I49538,I3035,I49470,I49564,);
DFFARX1 I_2735 (I174017,I3035,I49470,I49581,);
and I_2736 (I49589,I49581,I174032);
nor I_2737 (I49606,I49564,I49589);
DFFARX1 I_2738 (I49606,I3035,I49470,I49438,);
nand I_2739 (I49637,I49581,I174032);
nand I_2740 (I49654,I49504,I49637);
not I_2741 (I49450,I49654);
DFFARX1 I_2742 (I174035,I3035,I49470,I49694,);
DFFARX1 I_2743 (I49694,I3035,I49470,I49459,);
nand I_2744 (I49716,I174014,I174026);
and I_2745 (I49733,I49716,I174020);
DFFARX1 I_2746 (I49733,I3035,I49470,I49759,);
DFFARX1 I_2747 (I49759,I3035,I49470,I49776,);
not I_2748 (I49462,I49776);
not I_2749 (I49798,I49759);
nand I_2750 (I49447,I49798,I49637);
nor I_2751 (I49829,I174029,I174026);
not I_2752 (I49846,I49829);
nor I_2753 (I49863,I49798,I49846);
nor I_2754 (I49880,I49504,I49863);
DFFARX1 I_2755 (I49880,I3035,I49470,I49456,);
nor I_2756 (I49911,I49564,I49846);
nor I_2757 (I49444,I49759,I49911);
nor I_2758 (I49453,I49694,I49829);
nor I_2759 (I49441,I49564,I49829);
not I_2760 (I49997,I3042);
DFFARX1 I_2761 (I326751,I3035,I49997,I50023,);
not I_2762 (I50031,I50023);
nand I_2763 (I50048,I326763,I326748);
and I_2764 (I50065,I50048,I326742);
DFFARX1 I_2765 (I50065,I3035,I49997,I50091,);
DFFARX1 I_2766 (I326757,I3035,I49997,I50108,);
and I_2767 (I50116,I50108,I326745);
nor I_2768 (I50133,I50091,I50116);
DFFARX1 I_2769 (I50133,I3035,I49997,I49965,);
nand I_2770 (I50164,I50108,I326745);
nand I_2771 (I50181,I50031,I50164);
not I_2772 (I49977,I50181);
DFFARX1 I_2773 (I326754,I3035,I49997,I50221,);
DFFARX1 I_2774 (I50221,I3035,I49997,I49986,);
nand I_2775 (I50243,I326760,I326766);
and I_2776 (I50260,I50243,I326742);
DFFARX1 I_2777 (I50260,I3035,I49997,I50286,);
DFFARX1 I_2778 (I50286,I3035,I49997,I50303,);
not I_2779 (I49989,I50303);
not I_2780 (I50325,I50286);
nand I_2781 (I49974,I50325,I50164);
nor I_2782 (I50356,I326745,I326766);
not I_2783 (I50373,I50356);
nor I_2784 (I50390,I50325,I50373);
nor I_2785 (I50407,I50031,I50390);
DFFARX1 I_2786 (I50407,I3035,I49997,I49983,);
nor I_2787 (I50438,I50091,I50373);
nor I_2788 (I49971,I50286,I50438);
nor I_2789 (I49980,I50221,I50356);
nor I_2790 (I49968,I50091,I50356);
not I_2791 (I50524,I3042);
DFFARX1 I_2792 (I731745,I3035,I50524,I50550,);
not I_2793 (I50558,I50550);
nand I_2794 (I50575,I731739,I731760);
and I_2795 (I50592,I50575,I731736);
DFFARX1 I_2796 (I50592,I3035,I50524,I50618,);
DFFARX1 I_2797 (I731757,I3035,I50524,I50635,);
and I_2798 (I50643,I50635,I731754);
nor I_2799 (I50660,I50618,I50643);
DFFARX1 I_2800 (I50660,I3035,I50524,I50492,);
nand I_2801 (I50691,I50635,I731754);
nand I_2802 (I50708,I50558,I50691);
not I_2803 (I50504,I50708);
DFFARX1 I_2804 (I731742,I3035,I50524,I50748,);
DFFARX1 I_2805 (I50748,I3035,I50524,I50513,);
nand I_2806 (I50770,I731751,I731748);
and I_2807 (I50787,I50770,I731733);
DFFARX1 I_2808 (I50787,I3035,I50524,I50813,);
DFFARX1 I_2809 (I50813,I3035,I50524,I50830,);
not I_2810 (I50516,I50830);
not I_2811 (I50852,I50813);
nand I_2812 (I50501,I50852,I50691);
nor I_2813 (I50883,I731733,I731748);
not I_2814 (I50900,I50883);
nor I_2815 (I50917,I50852,I50900);
nor I_2816 (I50934,I50558,I50917);
DFFARX1 I_2817 (I50934,I3035,I50524,I50510,);
nor I_2818 (I50965,I50618,I50900);
nor I_2819 (I50498,I50813,I50965);
nor I_2820 (I50507,I50748,I50883);
nor I_2821 (I50495,I50618,I50883);
not I_2822 (I51051,I3042);
DFFARX1 I_2823 (I390334,I3035,I51051,I51077,);
not I_2824 (I51085,I51077);
nand I_2825 (I51102,I390325,I390343);
and I_2826 (I51119,I51102,I390322);
DFFARX1 I_2827 (I51119,I3035,I51051,I51145,);
DFFARX1 I_2828 (I390325,I3035,I51051,I51162,);
and I_2829 (I51170,I51162,I390328);
nor I_2830 (I51187,I51145,I51170);
DFFARX1 I_2831 (I51187,I3035,I51051,I51019,);
nand I_2832 (I51218,I51162,I390328);
nand I_2833 (I51235,I51085,I51218);
not I_2834 (I51031,I51235);
DFFARX1 I_2835 (I390322,I3035,I51051,I51275,);
DFFARX1 I_2836 (I51275,I3035,I51051,I51040,);
nand I_2837 (I51297,I390340,I390331);
and I_2838 (I51314,I51297,I390346);
DFFARX1 I_2839 (I51314,I3035,I51051,I51340,);
DFFARX1 I_2840 (I51340,I3035,I51051,I51357,);
not I_2841 (I51043,I51357);
not I_2842 (I51379,I51340);
nand I_2843 (I51028,I51379,I51218);
nor I_2844 (I51410,I390337,I390331);
not I_2845 (I51427,I51410);
nor I_2846 (I51444,I51379,I51427);
nor I_2847 (I51461,I51085,I51444);
DFFARX1 I_2848 (I51461,I3035,I51051,I51037,);
nor I_2849 (I51492,I51145,I51427);
nor I_2850 (I51025,I51340,I51492);
nor I_2851 (I51034,I51275,I51410);
nor I_2852 (I51022,I51145,I51410);
not I_2853 (I51578,I3042);
DFFARX1 I_2854 (I1836,I3035,I51578,I51604,);
not I_2855 (I51612,I51604);
nand I_2856 (I51629,I1676,I1700);
and I_2857 (I51646,I51629,I2564);
DFFARX1 I_2858 (I51646,I3035,I51578,I51672,);
DFFARX1 I_2859 (I2444,I3035,I51578,I51689,);
and I_2860 (I51697,I51689,I2068);
nor I_2861 (I51714,I51672,I51697);
DFFARX1 I_2862 (I51714,I3035,I51578,I51546,);
nand I_2863 (I51745,I51689,I2068);
nand I_2864 (I51762,I51612,I51745);
not I_2865 (I51558,I51762);
DFFARX1 I_2866 (I2020,I3035,I51578,I51802,);
DFFARX1 I_2867 (I51802,I3035,I51578,I51567,);
nand I_2868 (I51824,I1636,I2804);
and I_2869 (I51841,I51824,I2820);
DFFARX1 I_2870 (I51841,I3035,I51578,I51867,);
DFFARX1 I_2871 (I51867,I3035,I51578,I51884,);
not I_2872 (I51570,I51884);
not I_2873 (I51906,I51867);
nand I_2874 (I51555,I51906,I51745);
nor I_2875 (I51937,I2524,I2804);
not I_2876 (I51954,I51937);
nor I_2877 (I51971,I51906,I51954);
nor I_2878 (I51988,I51612,I51971);
DFFARX1 I_2879 (I51988,I3035,I51578,I51564,);
nor I_2880 (I52019,I51672,I51954);
nor I_2881 (I51552,I51867,I52019);
nor I_2882 (I51561,I51802,I51937);
nor I_2883 (I51549,I51672,I51937);
not I_2884 (I52105,I3042);
DFFARX1 I_2885 (I16788,I3035,I52105,I52131,);
not I_2886 (I52139,I52131);
nand I_2887 (I52156,I16776,I16782);
and I_2888 (I52173,I52156,I16785);
DFFARX1 I_2889 (I52173,I3035,I52105,I52199,);
DFFARX1 I_2890 (I16767,I3035,I52105,I52216,);
and I_2891 (I52224,I52216,I16773);
nor I_2892 (I52241,I52199,I52224);
DFFARX1 I_2893 (I52241,I3035,I52105,I52073,);
nand I_2894 (I52272,I52216,I16773);
nand I_2895 (I52289,I52139,I52272);
not I_2896 (I52085,I52289);
DFFARX1 I_2897 (I16767,I3035,I52105,I52329,);
DFFARX1 I_2898 (I52329,I3035,I52105,I52094,);
nand I_2899 (I52351,I16770,I16764);
and I_2900 (I52368,I52351,I16779);
DFFARX1 I_2901 (I52368,I3035,I52105,I52394,);
DFFARX1 I_2902 (I52394,I3035,I52105,I52411,);
not I_2903 (I52097,I52411);
not I_2904 (I52433,I52394);
nand I_2905 (I52082,I52433,I52272);
nor I_2906 (I52464,I16764,I16764);
not I_2907 (I52481,I52464);
nor I_2908 (I52498,I52433,I52481);
nor I_2909 (I52515,I52139,I52498);
DFFARX1 I_2910 (I52515,I3035,I52105,I52091,);
nor I_2911 (I52546,I52199,I52481);
nor I_2912 (I52079,I52394,I52546);
nor I_2913 (I52088,I52329,I52464);
nor I_2914 (I52076,I52199,I52464);
not I_2915 (I52632,I3042);
DFFARX1 I_2916 (I491583,I3035,I52632,I52658,);
not I_2917 (I52666,I52658);
nand I_2918 (I52683,I491601,I491595);
and I_2919 (I52700,I52683,I491574);
DFFARX1 I_2920 (I52700,I3035,I52632,I52726,);
DFFARX1 I_2921 (I491592,I3035,I52632,I52743,);
and I_2922 (I52751,I52743,I491577);
nor I_2923 (I52768,I52726,I52751);
DFFARX1 I_2924 (I52768,I3035,I52632,I52600,);
nand I_2925 (I52799,I52743,I491577);
nand I_2926 (I52816,I52666,I52799);
not I_2927 (I52612,I52816);
DFFARX1 I_2928 (I491589,I3035,I52632,I52856,);
DFFARX1 I_2929 (I52856,I3035,I52632,I52621,);
nand I_2930 (I52878,I491598,I491586);
and I_2931 (I52895,I52878,I491580);
DFFARX1 I_2932 (I52895,I3035,I52632,I52921,);
DFFARX1 I_2933 (I52921,I3035,I52632,I52938,);
not I_2934 (I52624,I52938);
not I_2935 (I52960,I52921);
nand I_2936 (I52609,I52960,I52799);
nor I_2937 (I52991,I491574,I491586);
not I_2938 (I53008,I52991);
nor I_2939 (I53025,I52960,I53008);
nor I_2940 (I53042,I52666,I53025);
DFFARX1 I_2941 (I53042,I3035,I52632,I52618,);
nor I_2942 (I53073,I52726,I53008);
nor I_2943 (I52606,I52921,I53073);
nor I_2944 (I52615,I52856,I52991);
nor I_2945 (I52603,I52726,I52991);
not I_2946 (I53159,I3042);
DFFARX1 I_2947 (I24166,I3035,I53159,I53185,);
not I_2948 (I53193,I53185);
nand I_2949 (I53210,I24154,I24160);
and I_2950 (I53227,I53210,I24163);
DFFARX1 I_2951 (I53227,I3035,I53159,I53253,);
DFFARX1 I_2952 (I24145,I3035,I53159,I53270,);
and I_2953 (I53278,I53270,I24151);
nor I_2954 (I53295,I53253,I53278);
DFFARX1 I_2955 (I53295,I3035,I53159,I53127,);
nand I_2956 (I53326,I53270,I24151);
nand I_2957 (I53343,I53193,I53326);
not I_2958 (I53139,I53343);
DFFARX1 I_2959 (I24145,I3035,I53159,I53383,);
DFFARX1 I_2960 (I53383,I3035,I53159,I53148,);
nand I_2961 (I53405,I24148,I24142);
and I_2962 (I53422,I53405,I24157);
DFFARX1 I_2963 (I53422,I3035,I53159,I53448,);
DFFARX1 I_2964 (I53448,I3035,I53159,I53465,);
not I_2965 (I53151,I53465);
not I_2966 (I53487,I53448);
nand I_2967 (I53136,I53487,I53326);
nor I_2968 (I53518,I24142,I24142);
not I_2969 (I53535,I53518);
nor I_2970 (I53552,I53487,I53535);
nor I_2971 (I53569,I53193,I53552);
DFFARX1 I_2972 (I53569,I3035,I53159,I53145,);
nor I_2973 (I53600,I53253,I53535);
nor I_2974 (I53133,I53448,I53600);
nor I_2975 (I53142,I53383,I53518);
nor I_2976 (I53130,I53253,I53518);
not I_2977 (I53686,I3042);
DFFARX1 I_2978 (I463550,I3035,I53686,I53712,);
not I_2979 (I53720,I53712);
nand I_2980 (I53737,I463547,I463562);
and I_2981 (I53754,I53737,I463544);
DFFARX1 I_2982 (I53754,I3035,I53686,I53780,);
DFFARX1 I_2983 (I463541,I3035,I53686,I53797,);
and I_2984 (I53805,I53797,I463541);
nor I_2985 (I53822,I53780,I53805);
DFFARX1 I_2986 (I53822,I3035,I53686,I53654,);
nand I_2987 (I53853,I53797,I463541);
nand I_2988 (I53870,I53720,I53853);
not I_2989 (I53666,I53870);
DFFARX1 I_2990 (I463544,I3035,I53686,I53910,);
DFFARX1 I_2991 (I53910,I3035,I53686,I53675,);
nand I_2992 (I53932,I463556,I463547);
and I_2993 (I53949,I53932,I463559);
DFFARX1 I_2994 (I53949,I3035,I53686,I53975,);
DFFARX1 I_2995 (I53975,I3035,I53686,I53992,);
not I_2996 (I53678,I53992);
not I_2997 (I54014,I53975);
nand I_2998 (I53663,I54014,I53853);
nor I_2999 (I54045,I463553,I463547);
not I_3000 (I54062,I54045);
nor I_3001 (I54079,I54014,I54062);
nor I_3002 (I54096,I53720,I54079);
DFFARX1 I_3003 (I54096,I3035,I53686,I53672,);
nor I_3004 (I54127,I53780,I54062);
nor I_3005 (I53660,I53975,I54127);
nor I_3006 (I53669,I53910,I54045);
nor I_3007 (I53657,I53780,I54045);
not I_3008 (I54213,I3042);
DFFARX1 I_3009 (I194594,I3035,I54213,I54239,);
not I_3010 (I54247,I54239);
nand I_3011 (I54264,I194576,I194591);
and I_3012 (I54281,I54264,I194567);
DFFARX1 I_3013 (I54281,I3035,I54213,I54307,);
DFFARX1 I_3014 (I194570,I3035,I54213,I54324,);
and I_3015 (I54332,I54324,I194585);
nor I_3016 (I54349,I54307,I54332);
DFFARX1 I_3017 (I54349,I3035,I54213,I54181,);
nand I_3018 (I54380,I54324,I194585);
nand I_3019 (I54397,I54247,I54380);
not I_3020 (I54193,I54397);
DFFARX1 I_3021 (I194588,I3035,I54213,I54437,);
DFFARX1 I_3022 (I54437,I3035,I54213,I54202,);
nand I_3023 (I54459,I194567,I194579);
and I_3024 (I54476,I54459,I194573);
DFFARX1 I_3025 (I54476,I3035,I54213,I54502,);
DFFARX1 I_3026 (I54502,I3035,I54213,I54519,);
not I_3027 (I54205,I54519);
not I_3028 (I54541,I54502);
nand I_3029 (I54190,I54541,I54380);
nor I_3030 (I54572,I194582,I194579);
not I_3031 (I54589,I54572);
nor I_3032 (I54606,I54541,I54589);
nor I_3033 (I54623,I54247,I54606);
DFFARX1 I_3034 (I54623,I3035,I54213,I54199,);
nor I_3035 (I54654,I54307,I54589);
nor I_3036 (I54187,I54502,I54654);
nor I_3037 (I54196,I54437,I54572);
nor I_3038 (I54184,I54307,I54572);
not I_3039 (I54740,I3042);
DFFARX1 I_3040 (I89621,I3035,I54740,I54766,);
not I_3041 (I54774,I54766);
nand I_3042 (I54791,I89615,I89609);
and I_3043 (I54808,I54791,I89630);
DFFARX1 I_3044 (I54808,I3035,I54740,I54834,);
DFFARX1 I_3045 (I89627,I3035,I54740,I54851,);
and I_3046 (I54859,I54851,I89624);
nor I_3047 (I54876,I54834,I54859);
DFFARX1 I_3048 (I54876,I3035,I54740,I54708,);
nand I_3049 (I54907,I54851,I89624);
nand I_3050 (I54924,I54774,I54907);
not I_3051 (I54720,I54924);
DFFARX1 I_3052 (I89609,I3035,I54740,I54964,);
DFFARX1 I_3053 (I54964,I3035,I54740,I54729,);
nand I_3054 (I54986,I89612,I89612);
and I_3055 (I55003,I54986,I89633);
DFFARX1 I_3056 (I55003,I3035,I54740,I55029,);
DFFARX1 I_3057 (I55029,I3035,I54740,I55046,);
not I_3058 (I54732,I55046);
not I_3059 (I55068,I55029);
nand I_3060 (I54717,I55068,I54907);
nor I_3061 (I55099,I89618,I89612);
not I_3062 (I55116,I55099);
nor I_3063 (I55133,I55068,I55116);
nor I_3064 (I55150,I54774,I55133);
DFFARX1 I_3065 (I55150,I3035,I54740,I54726,);
nor I_3066 (I55181,I54834,I55116);
nor I_3067 (I54714,I55029,I55181);
nor I_3068 (I54723,I54964,I55099);
nor I_3069 (I54711,I54834,I55099);
not I_3070 (I55267,I3042);
DFFARX1 I_3071 (I390912,I3035,I55267,I55293,);
not I_3072 (I55301,I55293);
nand I_3073 (I55318,I390903,I390921);
and I_3074 (I55335,I55318,I390900);
DFFARX1 I_3075 (I55335,I3035,I55267,I55361,);
DFFARX1 I_3076 (I390903,I3035,I55267,I55378,);
and I_3077 (I55386,I55378,I390906);
nor I_3078 (I55403,I55361,I55386);
DFFARX1 I_3079 (I55403,I3035,I55267,I55235,);
nand I_3080 (I55434,I55378,I390906);
nand I_3081 (I55451,I55301,I55434);
not I_3082 (I55247,I55451);
DFFARX1 I_3083 (I390900,I3035,I55267,I55491,);
DFFARX1 I_3084 (I55491,I3035,I55267,I55256,);
nand I_3085 (I55513,I390918,I390909);
and I_3086 (I55530,I55513,I390924);
DFFARX1 I_3087 (I55530,I3035,I55267,I55556,);
DFFARX1 I_3088 (I55556,I3035,I55267,I55573,);
not I_3089 (I55259,I55573);
not I_3090 (I55595,I55556);
nand I_3091 (I55244,I55595,I55434);
nor I_3092 (I55626,I390915,I390909);
not I_3093 (I55643,I55626);
nor I_3094 (I55660,I55595,I55643);
nor I_3095 (I55677,I55301,I55660);
DFFARX1 I_3096 (I55677,I3035,I55267,I55253,);
nor I_3097 (I55708,I55361,I55643);
nor I_3098 (I55241,I55556,I55708);
nor I_3099 (I55250,I55491,I55626);
nor I_3100 (I55238,I55361,I55626);
not I_3101 (I55794,I3042);
DFFARX1 I_3102 (I278327,I3035,I55794,I55820,);
not I_3103 (I55828,I55820);
nand I_3104 (I55845,I278321,I278312);
and I_3105 (I55862,I55845,I278333);
DFFARX1 I_3106 (I55862,I3035,I55794,I55888,);
DFFARX1 I_3107 (I278315,I3035,I55794,I55905,);
and I_3108 (I55913,I55905,I278309);
nor I_3109 (I55930,I55888,I55913);
DFFARX1 I_3110 (I55930,I3035,I55794,I55762,);
nand I_3111 (I55961,I55905,I278309);
nand I_3112 (I55978,I55828,I55961);
not I_3113 (I55774,I55978);
DFFARX1 I_3114 (I278309,I3035,I55794,I56018,);
DFFARX1 I_3115 (I56018,I3035,I55794,I55783,);
nand I_3116 (I56040,I278336,I278318);
and I_3117 (I56057,I56040,I278324);
DFFARX1 I_3118 (I56057,I3035,I55794,I56083,);
DFFARX1 I_3119 (I56083,I3035,I55794,I56100,);
not I_3120 (I55786,I56100);
not I_3121 (I56122,I56083);
nand I_3122 (I55771,I56122,I55961);
nor I_3123 (I56153,I278330,I278318);
not I_3124 (I56170,I56153);
nor I_3125 (I56187,I56122,I56170);
nor I_3126 (I56204,I55828,I56187);
DFFARX1 I_3127 (I56204,I3035,I55794,I55780,);
nor I_3128 (I56235,I55888,I56170);
nor I_3129 (I55768,I56083,I56235);
nor I_3130 (I55777,I56018,I56153);
nor I_3131 (I55765,I55888,I56153);
not I_3132 (I56321,I3042);
DFFARX1 I_3133 (I740075,I3035,I56321,I56347,);
not I_3134 (I56355,I56347);
nand I_3135 (I56372,I740069,I740090);
and I_3136 (I56389,I56372,I740066);
DFFARX1 I_3137 (I56389,I3035,I56321,I56415,);
DFFARX1 I_3138 (I740087,I3035,I56321,I56432,);
and I_3139 (I56440,I56432,I740084);
nor I_3140 (I56457,I56415,I56440);
DFFARX1 I_3141 (I56457,I3035,I56321,I56289,);
nand I_3142 (I56488,I56432,I740084);
nand I_3143 (I56505,I56355,I56488);
not I_3144 (I56301,I56505);
DFFARX1 I_3145 (I740072,I3035,I56321,I56545,);
DFFARX1 I_3146 (I56545,I3035,I56321,I56310,);
nand I_3147 (I56567,I740081,I740078);
and I_3148 (I56584,I56567,I740063);
DFFARX1 I_3149 (I56584,I3035,I56321,I56610,);
DFFARX1 I_3150 (I56610,I3035,I56321,I56627,);
not I_3151 (I56313,I56627);
not I_3152 (I56649,I56610);
nand I_3153 (I56298,I56649,I56488);
nor I_3154 (I56680,I740063,I740078);
not I_3155 (I56697,I56680);
nor I_3156 (I56714,I56649,I56697);
nor I_3157 (I56731,I56355,I56714);
DFFARX1 I_3158 (I56731,I3035,I56321,I56307,);
nor I_3159 (I56762,I56415,I56697);
nor I_3160 (I56295,I56610,I56762);
nor I_3161 (I56304,I56545,I56680);
nor I_3162 (I56292,I56415,I56680);
not I_3163 (I56848,I3042);
DFFARX1 I_3164 (I211458,I3035,I56848,I56874,);
not I_3165 (I56882,I56874);
nand I_3166 (I56899,I211440,I211455);
and I_3167 (I56916,I56899,I211431);
DFFARX1 I_3168 (I56916,I3035,I56848,I56942,);
DFFARX1 I_3169 (I211434,I3035,I56848,I56959,);
and I_3170 (I56967,I56959,I211449);
nor I_3171 (I56984,I56942,I56967);
DFFARX1 I_3172 (I56984,I3035,I56848,I56816,);
nand I_3173 (I57015,I56959,I211449);
nand I_3174 (I57032,I56882,I57015);
not I_3175 (I56828,I57032);
DFFARX1 I_3176 (I211452,I3035,I56848,I57072,);
DFFARX1 I_3177 (I57072,I3035,I56848,I56837,);
nand I_3178 (I57094,I211431,I211443);
and I_3179 (I57111,I57094,I211437);
DFFARX1 I_3180 (I57111,I3035,I56848,I57137,);
DFFARX1 I_3181 (I57137,I3035,I56848,I57154,);
not I_3182 (I56840,I57154);
not I_3183 (I57176,I57137);
nand I_3184 (I56825,I57176,I57015);
nor I_3185 (I57207,I211446,I211443);
not I_3186 (I57224,I57207);
nor I_3187 (I57241,I57176,I57224);
nor I_3188 (I57258,I56882,I57241);
DFFARX1 I_3189 (I57258,I3035,I56848,I56834,);
nor I_3190 (I57289,I56942,I57224);
nor I_3191 (I56822,I57137,I57289);
nor I_3192 (I56831,I57072,I57207);
nor I_3193 (I56819,I56942,I57207);
not I_3194 (I57375,I3042);
DFFARX1 I_3195 (I297199,I3035,I57375,I57401,);
not I_3196 (I57409,I57401);
nand I_3197 (I57426,I297220,I297214);
and I_3198 (I57443,I57426,I297196);
DFFARX1 I_3199 (I57443,I3035,I57375,I57469,);
DFFARX1 I_3200 (I297199,I3035,I57375,I57486,);
and I_3201 (I57494,I57486,I297208);
nor I_3202 (I57511,I57469,I57494);
DFFARX1 I_3203 (I57511,I3035,I57375,I57343,);
nand I_3204 (I57542,I57486,I297208);
nand I_3205 (I57559,I57409,I57542);
not I_3206 (I57355,I57559);
DFFARX1 I_3207 (I297205,I3035,I57375,I57599,);
DFFARX1 I_3208 (I57599,I3035,I57375,I57364,);
nand I_3209 (I57621,I297211,I297202);
and I_3210 (I57638,I57621,I297196);
DFFARX1 I_3211 (I57638,I3035,I57375,I57664,);
DFFARX1 I_3212 (I57664,I3035,I57375,I57681,);
not I_3213 (I57367,I57681);
not I_3214 (I57703,I57664);
nand I_3215 (I57352,I57703,I57542);
nor I_3216 (I57734,I297217,I297202);
not I_3217 (I57751,I57734);
nor I_3218 (I57768,I57703,I57751);
nor I_3219 (I57785,I57409,I57768);
DFFARX1 I_3220 (I57785,I3035,I57375,I57361,);
nor I_3221 (I57816,I57469,I57751);
nor I_3222 (I57349,I57664,I57816);
nor I_3223 (I57358,I57599,I57734);
nor I_3224 (I57346,I57469,I57734);
not I_3225 (I57902,I3042);
DFFARX1 I_3226 (I134246,I3035,I57902,I57928,);
not I_3227 (I57936,I57928);
nand I_3228 (I57953,I134240,I134234);
and I_3229 (I57970,I57953,I134255);
DFFARX1 I_3230 (I57970,I3035,I57902,I57996,);
DFFARX1 I_3231 (I134252,I3035,I57902,I58013,);
and I_3232 (I58021,I58013,I134249);
nor I_3233 (I58038,I57996,I58021);
DFFARX1 I_3234 (I58038,I3035,I57902,I57870,);
nand I_3235 (I58069,I58013,I134249);
nand I_3236 (I58086,I57936,I58069);
not I_3237 (I57882,I58086);
DFFARX1 I_3238 (I134234,I3035,I57902,I58126,);
DFFARX1 I_3239 (I58126,I3035,I57902,I57891,);
nand I_3240 (I58148,I134237,I134237);
and I_3241 (I58165,I58148,I134258);
DFFARX1 I_3242 (I58165,I3035,I57902,I58191,);
DFFARX1 I_3243 (I58191,I3035,I57902,I58208,);
not I_3244 (I57894,I58208);
not I_3245 (I58230,I58191);
nand I_3246 (I57879,I58230,I58069);
nor I_3247 (I58261,I134243,I134237);
not I_3248 (I58278,I58261);
nor I_3249 (I58295,I58230,I58278);
nor I_3250 (I58312,I57936,I58295);
DFFARX1 I_3251 (I58312,I3035,I57902,I57888,);
nor I_3252 (I58343,I57996,I58278);
nor I_3253 (I57876,I58191,I58343);
nor I_3254 (I57885,I58126,I58261);
nor I_3255 (I57873,I57996,I58261);
not I_3256 (I58429,I3042);
DFFARX1 I_3257 (I438254,I3035,I58429,I58455,);
not I_3258 (I58463,I58455);
nand I_3259 (I58480,I438251,I438266);
and I_3260 (I58497,I58480,I438248);
DFFARX1 I_3261 (I58497,I3035,I58429,I58523,);
DFFARX1 I_3262 (I438245,I3035,I58429,I58540,);
and I_3263 (I58548,I58540,I438245);
nor I_3264 (I58565,I58523,I58548);
DFFARX1 I_3265 (I58565,I3035,I58429,I58397,);
nand I_3266 (I58596,I58540,I438245);
nand I_3267 (I58613,I58463,I58596);
not I_3268 (I58409,I58613);
DFFARX1 I_3269 (I438248,I3035,I58429,I58653,);
DFFARX1 I_3270 (I58653,I3035,I58429,I58418,);
nand I_3271 (I58675,I438260,I438251);
and I_3272 (I58692,I58675,I438263);
DFFARX1 I_3273 (I58692,I3035,I58429,I58718,);
DFFARX1 I_3274 (I58718,I3035,I58429,I58735,);
not I_3275 (I58421,I58735);
not I_3276 (I58757,I58718);
nand I_3277 (I58406,I58757,I58596);
nor I_3278 (I58788,I438257,I438251);
not I_3279 (I58805,I58788);
nor I_3280 (I58822,I58757,I58805);
nor I_3281 (I58839,I58463,I58822);
DFFARX1 I_3282 (I58839,I3035,I58429,I58415,);
nor I_3283 (I58870,I58523,I58805);
nor I_3284 (I58403,I58718,I58870);
nor I_3285 (I58412,I58653,I58788);
nor I_3286 (I58400,I58523,I58788);
not I_3287 (I58956,I3042);
DFFARX1 I_3288 (I729960,I3035,I58956,I58982,);
not I_3289 (I58990,I58982);
nand I_3290 (I59007,I729954,I729975);
and I_3291 (I59024,I59007,I729951);
DFFARX1 I_3292 (I59024,I3035,I58956,I59050,);
DFFARX1 I_3293 (I729972,I3035,I58956,I59067,);
and I_3294 (I59075,I59067,I729969);
nor I_3295 (I59092,I59050,I59075);
DFFARX1 I_3296 (I59092,I3035,I58956,I58924,);
nand I_3297 (I59123,I59067,I729969);
nand I_3298 (I59140,I58990,I59123);
not I_3299 (I58936,I59140);
DFFARX1 I_3300 (I729957,I3035,I58956,I59180,);
DFFARX1 I_3301 (I59180,I3035,I58956,I58945,);
nand I_3302 (I59202,I729966,I729963);
and I_3303 (I59219,I59202,I729948);
DFFARX1 I_3304 (I59219,I3035,I58956,I59245,);
DFFARX1 I_3305 (I59245,I3035,I58956,I59262,);
not I_3306 (I58948,I59262);
not I_3307 (I59284,I59245);
nand I_3308 (I58933,I59284,I59123);
nor I_3309 (I59315,I729948,I729963);
not I_3310 (I59332,I59315);
nor I_3311 (I59349,I59284,I59332);
nor I_3312 (I59366,I58990,I59349);
DFFARX1 I_3313 (I59366,I3035,I58956,I58942,);
nor I_3314 (I59397,I59050,I59332);
nor I_3315 (I58930,I59245,I59397);
nor I_3316 (I58939,I59180,I59315);
nor I_3317 (I58927,I59050,I59315);
not I_3318 (I59483,I3042);
DFFARX1 I_3319 (I399004,I3035,I59483,I59509,);
not I_3320 (I59517,I59509);
nand I_3321 (I59534,I398995,I399013);
and I_3322 (I59551,I59534,I398992);
DFFARX1 I_3323 (I59551,I3035,I59483,I59577,);
DFFARX1 I_3324 (I398995,I3035,I59483,I59594,);
and I_3325 (I59602,I59594,I398998);
nor I_3326 (I59619,I59577,I59602);
DFFARX1 I_3327 (I59619,I3035,I59483,I59451,);
nand I_3328 (I59650,I59594,I398998);
nand I_3329 (I59667,I59517,I59650);
not I_3330 (I59463,I59667);
DFFARX1 I_3331 (I398992,I3035,I59483,I59707,);
DFFARX1 I_3332 (I59707,I3035,I59483,I59472,);
nand I_3333 (I59729,I399010,I399001);
and I_3334 (I59746,I59729,I399016);
DFFARX1 I_3335 (I59746,I3035,I59483,I59772,);
DFFARX1 I_3336 (I59772,I3035,I59483,I59789,);
not I_3337 (I59475,I59789);
not I_3338 (I59811,I59772);
nand I_3339 (I59460,I59811,I59650);
nor I_3340 (I59842,I399007,I399001);
not I_3341 (I59859,I59842);
nor I_3342 (I59876,I59811,I59859);
nor I_3343 (I59893,I59517,I59876);
DFFARX1 I_3344 (I59893,I3035,I59483,I59469,);
nor I_3345 (I59924,I59577,I59859);
nor I_3346 (I59457,I59772,I59924);
nor I_3347 (I59466,I59707,I59842);
nor I_3348 (I59454,I59577,I59842);
not I_3349 (I60010,I3042);
DFFARX1 I_3350 (I109851,I3035,I60010,I60036,);
not I_3351 (I60044,I60036);
nand I_3352 (I60061,I109845,I109839);
and I_3353 (I60078,I60061,I109860);
DFFARX1 I_3354 (I60078,I3035,I60010,I60104,);
DFFARX1 I_3355 (I109857,I3035,I60010,I60121,);
and I_3356 (I60129,I60121,I109854);
nor I_3357 (I60146,I60104,I60129);
DFFARX1 I_3358 (I60146,I3035,I60010,I59978,);
nand I_3359 (I60177,I60121,I109854);
nand I_3360 (I60194,I60044,I60177);
not I_3361 (I59990,I60194);
DFFARX1 I_3362 (I109839,I3035,I60010,I60234,);
DFFARX1 I_3363 (I60234,I3035,I60010,I59999,);
nand I_3364 (I60256,I109842,I109842);
and I_3365 (I60273,I60256,I109863);
DFFARX1 I_3366 (I60273,I3035,I60010,I60299,);
DFFARX1 I_3367 (I60299,I3035,I60010,I60316,);
not I_3368 (I60002,I60316);
not I_3369 (I60338,I60299);
nand I_3370 (I59987,I60338,I60177);
nor I_3371 (I60369,I109848,I109842);
not I_3372 (I60386,I60369);
nor I_3373 (I60403,I60338,I60386);
nor I_3374 (I60420,I60044,I60403);
DFFARX1 I_3375 (I60420,I3035,I60010,I59996,);
nor I_3376 (I60451,I60104,I60386);
nor I_3377 (I59984,I60299,I60451);
nor I_3378 (I59993,I60234,I60369);
nor I_3379 (I59981,I60104,I60369);
not I_3380 (I60537,I3042);
DFFARX1 I_3381 (I269079,I3035,I60537,I60563,);
not I_3382 (I60571,I60563);
nand I_3383 (I60588,I269073,I269064);
and I_3384 (I60605,I60588,I269085);
DFFARX1 I_3385 (I60605,I3035,I60537,I60631,);
DFFARX1 I_3386 (I269067,I3035,I60537,I60648,);
and I_3387 (I60656,I60648,I269061);
nor I_3388 (I60673,I60631,I60656);
DFFARX1 I_3389 (I60673,I3035,I60537,I60505,);
nand I_3390 (I60704,I60648,I269061);
nand I_3391 (I60721,I60571,I60704);
not I_3392 (I60517,I60721);
DFFARX1 I_3393 (I269061,I3035,I60537,I60761,);
DFFARX1 I_3394 (I60761,I3035,I60537,I60526,);
nand I_3395 (I60783,I269088,I269070);
and I_3396 (I60800,I60783,I269076);
DFFARX1 I_3397 (I60800,I3035,I60537,I60826,);
DFFARX1 I_3398 (I60826,I3035,I60537,I60843,);
not I_3399 (I60529,I60843);
not I_3400 (I60865,I60826);
nand I_3401 (I60514,I60865,I60704);
nor I_3402 (I60896,I269082,I269070);
not I_3403 (I60913,I60896);
nor I_3404 (I60930,I60865,I60913);
nor I_3405 (I60947,I60571,I60930);
DFFARX1 I_3406 (I60947,I3035,I60537,I60523,);
nor I_3407 (I60978,I60631,I60913);
nor I_3408 (I60511,I60826,I60978);
nor I_3409 (I60520,I60761,I60896);
nor I_3410 (I60508,I60631,I60896);
not I_3411 (I61064,I3042);
DFFARX1 I_3412 (I356232,I3035,I61064,I61090,);
not I_3413 (I61098,I61090);
nand I_3414 (I61115,I356223,I356241);
and I_3415 (I61132,I61115,I356220);
DFFARX1 I_3416 (I61132,I3035,I61064,I61158,);
DFFARX1 I_3417 (I356223,I3035,I61064,I61175,);
and I_3418 (I61183,I61175,I356226);
nor I_3419 (I61200,I61158,I61183);
DFFARX1 I_3420 (I61200,I3035,I61064,I61032,);
nand I_3421 (I61231,I61175,I356226);
nand I_3422 (I61248,I61098,I61231);
not I_3423 (I61044,I61248);
DFFARX1 I_3424 (I356220,I3035,I61064,I61288,);
DFFARX1 I_3425 (I61288,I3035,I61064,I61053,);
nand I_3426 (I61310,I356238,I356229);
and I_3427 (I61327,I61310,I356244);
DFFARX1 I_3428 (I61327,I3035,I61064,I61353,);
DFFARX1 I_3429 (I61353,I3035,I61064,I61370,);
not I_3430 (I61056,I61370);
not I_3431 (I61392,I61353);
nand I_3432 (I61041,I61392,I61231);
nor I_3433 (I61423,I356235,I356229);
not I_3434 (I61440,I61423);
nor I_3435 (I61457,I61392,I61440);
nor I_3436 (I61474,I61098,I61457);
DFFARX1 I_3437 (I61474,I3035,I61064,I61050,);
nor I_3438 (I61505,I61158,I61440);
nor I_3439 (I61038,I61353,I61505);
nor I_3440 (I61047,I61288,I61423);
nor I_3441 (I61035,I61158,I61423);
not I_3442 (I61591,I3042);
DFFARX1 I_3443 (I180892,I3035,I61591,I61617,);
not I_3444 (I61625,I61617);
nand I_3445 (I61642,I180874,I180889);
and I_3446 (I61659,I61642,I180865);
DFFARX1 I_3447 (I61659,I3035,I61591,I61685,);
DFFARX1 I_3448 (I180868,I3035,I61591,I61702,);
and I_3449 (I61710,I61702,I180883);
nor I_3450 (I61727,I61685,I61710);
DFFARX1 I_3451 (I61727,I3035,I61591,I61559,);
nand I_3452 (I61758,I61702,I180883);
nand I_3453 (I61775,I61625,I61758);
not I_3454 (I61571,I61775);
DFFARX1 I_3455 (I180886,I3035,I61591,I61815,);
DFFARX1 I_3456 (I61815,I3035,I61591,I61580,);
nand I_3457 (I61837,I180865,I180877);
and I_3458 (I61854,I61837,I180871);
DFFARX1 I_3459 (I61854,I3035,I61591,I61880,);
DFFARX1 I_3460 (I61880,I3035,I61591,I61897,);
not I_3461 (I61583,I61897);
not I_3462 (I61919,I61880);
nand I_3463 (I61568,I61919,I61758);
nor I_3464 (I61950,I180880,I180877);
not I_3465 (I61967,I61950);
nor I_3466 (I61984,I61919,I61967);
nor I_3467 (I62001,I61625,I61984);
DFFARX1 I_3468 (I62001,I3035,I61591,I61577,);
nor I_3469 (I62032,I61685,I61967);
nor I_3470 (I61565,I61880,I62032);
nor I_3471 (I61574,I61815,I61950);
nor I_3472 (I61562,I61685,I61950);
not I_3473 (I62118,I3042);
DFFARX1 I_3474 (I180365,I3035,I62118,I62144,);
not I_3475 (I62152,I62144);
nand I_3476 (I62169,I180347,I180362);
and I_3477 (I62186,I62169,I180338);
DFFARX1 I_3478 (I62186,I3035,I62118,I62212,);
DFFARX1 I_3479 (I180341,I3035,I62118,I62229,);
and I_3480 (I62237,I62229,I180356);
nor I_3481 (I62254,I62212,I62237);
DFFARX1 I_3482 (I62254,I3035,I62118,I62086,);
nand I_3483 (I62285,I62229,I180356);
nand I_3484 (I62302,I62152,I62285);
not I_3485 (I62098,I62302);
DFFARX1 I_3486 (I180359,I3035,I62118,I62342,);
DFFARX1 I_3487 (I62342,I3035,I62118,I62107,);
nand I_3488 (I62364,I180338,I180350);
and I_3489 (I62381,I62364,I180344);
DFFARX1 I_3490 (I62381,I3035,I62118,I62407,);
DFFARX1 I_3491 (I62407,I3035,I62118,I62424,);
not I_3492 (I62110,I62424);
not I_3493 (I62446,I62407);
nand I_3494 (I62095,I62446,I62285);
nor I_3495 (I62477,I180353,I180350);
not I_3496 (I62494,I62477);
nor I_3497 (I62511,I62446,I62494);
nor I_3498 (I62528,I62152,I62511);
DFFARX1 I_3499 (I62528,I3035,I62118,I62104,);
nor I_3500 (I62559,I62212,I62494);
nor I_3501 (I62092,I62407,I62559);
nor I_3502 (I62101,I62342,I62477);
nor I_3503 (I62089,I62212,I62477);
not I_3504 (I62645,I3042);
DFFARX1 I_3505 (I175095,I3035,I62645,I62671,);
not I_3506 (I62679,I62671);
nand I_3507 (I62696,I175077,I175092);
and I_3508 (I62713,I62696,I175068);
DFFARX1 I_3509 (I62713,I3035,I62645,I62739,);
DFFARX1 I_3510 (I175071,I3035,I62645,I62756,);
and I_3511 (I62764,I62756,I175086);
nor I_3512 (I62781,I62739,I62764);
DFFARX1 I_3513 (I62781,I3035,I62645,I62613,);
nand I_3514 (I62812,I62756,I175086);
nand I_3515 (I62829,I62679,I62812);
not I_3516 (I62625,I62829);
DFFARX1 I_3517 (I175089,I3035,I62645,I62869,);
DFFARX1 I_3518 (I62869,I3035,I62645,I62634,);
nand I_3519 (I62891,I175068,I175080);
and I_3520 (I62908,I62891,I175074);
DFFARX1 I_3521 (I62908,I3035,I62645,I62934,);
DFFARX1 I_3522 (I62934,I3035,I62645,I62951,);
not I_3523 (I62637,I62951);
not I_3524 (I62973,I62934);
nand I_3525 (I62622,I62973,I62812);
nor I_3526 (I63004,I175083,I175080);
not I_3527 (I63021,I63004);
nor I_3528 (I63038,I62973,I63021);
nor I_3529 (I63055,I62679,I63038);
DFFARX1 I_3530 (I63055,I3035,I62645,I62631,);
nor I_3531 (I63086,I62739,I63021);
nor I_3532 (I62619,I62934,I63086);
nor I_3533 (I62628,I62869,I63004);
nor I_3534 (I62616,I62739,I63004);
not I_3535 (I63172,I3042);
DFFARX1 I_3536 (I529697,I3035,I63172,I63198,);
not I_3537 (I63206,I63198);
nand I_3538 (I63223,I529715,I529709);
and I_3539 (I63240,I63223,I529688);
DFFARX1 I_3540 (I63240,I3035,I63172,I63266,);
DFFARX1 I_3541 (I529706,I3035,I63172,I63283,);
and I_3542 (I63291,I63283,I529691);
nor I_3543 (I63308,I63266,I63291);
DFFARX1 I_3544 (I63308,I3035,I63172,I63140,);
nand I_3545 (I63339,I63283,I529691);
nand I_3546 (I63356,I63206,I63339);
not I_3547 (I63152,I63356);
DFFARX1 I_3548 (I529703,I3035,I63172,I63396,);
DFFARX1 I_3549 (I63396,I3035,I63172,I63161,);
nand I_3550 (I63418,I529712,I529700);
and I_3551 (I63435,I63418,I529694);
DFFARX1 I_3552 (I63435,I3035,I63172,I63461,);
DFFARX1 I_3553 (I63461,I3035,I63172,I63478,);
not I_3554 (I63164,I63478);
not I_3555 (I63500,I63461);
nand I_3556 (I63149,I63500,I63339);
nor I_3557 (I63531,I529688,I529700);
not I_3558 (I63548,I63531);
nor I_3559 (I63565,I63500,I63548);
nor I_3560 (I63582,I63206,I63565);
DFFARX1 I_3561 (I63582,I3035,I63172,I63158,);
nor I_3562 (I63613,I63266,I63548);
nor I_3563 (I63146,I63461,I63613);
nor I_3564 (I63155,I63396,I63531);
nor I_3565 (I63143,I63266,I63531);
not I_3566 (I63699,I3042);
DFFARX1 I_3567 (I516777,I3035,I63699,I63725,);
not I_3568 (I63733,I63725);
nand I_3569 (I63750,I516795,I516789);
and I_3570 (I63767,I63750,I516768);
DFFARX1 I_3571 (I63767,I3035,I63699,I63793,);
DFFARX1 I_3572 (I516786,I3035,I63699,I63810,);
and I_3573 (I63818,I63810,I516771);
nor I_3574 (I63835,I63793,I63818);
DFFARX1 I_3575 (I63835,I3035,I63699,I63667,);
nand I_3576 (I63866,I63810,I516771);
nand I_3577 (I63883,I63733,I63866);
not I_3578 (I63679,I63883);
DFFARX1 I_3579 (I516783,I3035,I63699,I63923,);
DFFARX1 I_3580 (I63923,I3035,I63699,I63688,);
nand I_3581 (I63945,I516792,I516780);
and I_3582 (I63962,I63945,I516774);
DFFARX1 I_3583 (I63962,I3035,I63699,I63988,);
DFFARX1 I_3584 (I63988,I3035,I63699,I64005,);
not I_3585 (I63691,I64005);
not I_3586 (I64027,I63988);
nand I_3587 (I63676,I64027,I63866);
nor I_3588 (I64058,I516768,I516780);
not I_3589 (I64075,I64058);
nor I_3590 (I64092,I64027,I64075);
nor I_3591 (I64109,I63733,I64092);
DFFARX1 I_3592 (I64109,I3035,I63699,I63685,);
nor I_3593 (I64140,I63793,I64075);
nor I_3594 (I63673,I63988,I64140);
nor I_3595 (I63682,I63923,I64058);
nor I_3596 (I63670,I63793,I64058);
not I_3597 (I64226,I3042);
DFFARX1 I_3598 (I738885,I3035,I64226,I64252,);
not I_3599 (I64260,I64252);
nand I_3600 (I64277,I738879,I738900);
and I_3601 (I64294,I64277,I738876);
DFFARX1 I_3602 (I64294,I3035,I64226,I64320,);
DFFARX1 I_3603 (I738897,I3035,I64226,I64337,);
and I_3604 (I64345,I64337,I738894);
nor I_3605 (I64362,I64320,I64345);
DFFARX1 I_3606 (I64362,I3035,I64226,I64194,);
nand I_3607 (I64393,I64337,I738894);
nand I_3608 (I64410,I64260,I64393);
not I_3609 (I64206,I64410);
DFFARX1 I_3610 (I738882,I3035,I64226,I64450,);
DFFARX1 I_3611 (I64450,I3035,I64226,I64215,);
nand I_3612 (I64472,I738891,I738888);
and I_3613 (I64489,I64472,I738873);
DFFARX1 I_3614 (I64489,I3035,I64226,I64515,);
DFFARX1 I_3615 (I64515,I3035,I64226,I64532,);
not I_3616 (I64218,I64532);
not I_3617 (I64554,I64515);
nand I_3618 (I64203,I64554,I64393);
nor I_3619 (I64585,I738873,I738888);
not I_3620 (I64602,I64585);
nor I_3621 (I64619,I64554,I64602);
nor I_3622 (I64636,I64260,I64619);
DFFARX1 I_3623 (I64636,I3035,I64226,I64212,);
nor I_3624 (I64667,I64320,I64602);
nor I_3625 (I64200,I64515,I64667);
nor I_3626 (I64209,I64450,I64585);
nor I_3627 (I64197,I64320,I64585);
not I_3628 (I64753,I3042);
DFFARX1 I_3629 (I382820,I3035,I64753,I64779,);
not I_3630 (I64787,I64779);
nand I_3631 (I64804,I382811,I382829);
and I_3632 (I64821,I64804,I382808);
DFFARX1 I_3633 (I64821,I3035,I64753,I64847,);
DFFARX1 I_3634 (I382811,I3035,I64753,I64864,);
and I_3635 (I64872,I64864,I382814);
nor I_3636 (I64889,I64847,I64872);
DFFARX1 I_3637 (I64889,I3035,I64753,I64721,);
nand I_3638 (I64920,I64864,I382814);
nand I_3639 (I64937,I64787,I64920);
not I_3640 (I64733,I64937);
DFFARX1 I_3641 (I382808,I3035,I64753,I64977,);
DFFARX1 I_3642 (I64977,I3035,I64753,I64742,);
nand I_3643 (I64999,I382826,I382817);
and I_3644 (I65016,I64999,I382832);
DFFARX1 I_3645 (I65016,I3035,I64753,I65042,);
DFFARX1 I_3646 (I65042,I3035,I64753,I65059,);
not I_3647 (I64745,I65059);
not I_3648 (I65081,I65042);
nand I_3649 (I64730,I65081,I64920);
nor I_3650 (I65112,I382823,I382817);
not I_3651 (I65129,I65112);
nor I_3652 (I65146,I65081,I65129);
nor I_3653 (I65163,I64787,I65146);
DFFARX1 I_3654 (I65163,I3035,I64753,I64739,);
nor I_3655 (I65194,I64847,I65129);
nor I_3656 (I64727,I65042,I65194);
nor I_3657 (I64736,I64977,I65112);
nor I_3658 (I64724,I64847,I65112);
not I_3659 (I65280,I3042);
DFFARX1 I_3660 (I300163,I3035,I65280,I65306,);
not I_3661 (I65314,I65306);
nand I_3662 (I65331,I300175,I300160);
and I_3663 (I65348,I65331,I300154);
DFFARX1 I_3664 (I65348,I3035,I65280,I65374,);
DFFARX1 I_3665 (I300169,I3035,I65280,I65391,);
and I_3666 (I65399,I65391,I300157);
nor I_3667 (I65416,I65374,I65399);
DFFARX1 I_3668 (I65416,I3035,I65280,I65248,);
nand I_3669 (I65447,I65391,I300157);
nand I_3670 (I65464,I65314,I65447);
not I_3671 (I65260,I65464);
DFFARX1 I_3672 (I300166,I3035,I65280,I65504,);
DFFARX1 I_3673 (I65504,I3035,I65280,I65269,);
nand I_3674 (I65526,I300172,I300178);
and I_3675 (I65543,I65526,I300154);
DFFARX1 I_3676 (I65543,I3035,I65280,I65569,);
DFFARX1 I_3677 (I65569,I3035,I65280,I65586,);
not I_3678 (I65272,I65586);
not I_3679 (I65608,I65569);
nand I_3680 (I65257,I65608,I65447);
nor I_3681 (I65639,I300157,I300178);
not I_3682 (I65656,I65639);
nor I_3683 (I65673,I65608,I65656);
nor I_3684 (I65690,I65314,I65673);
DFFARX1 I_3685 (I65690,I3035,I65280,I65266,);
nor I_3686 (I65721,I65374,I65656);
nor I_3687 (I65254,I65569,I65721);
nor I_3688 (I65263,I65504,I65639);
nor I_3689 (I65251,I65374,I65639);
not I_3690 (I65807,I3042);
DFFARX1 I_3691 (I378774,I3035,I65807,I65833,);
not I_3692 (I65841,I65833);
nand I_3693 (I65858,I378765,I378783);
and I_3694 (I65875,I65858,I378762);
DFFARX1 I_3695 (I65875,I3035,I65807,I65901,);
DFFARX1 I_3696 (I378765,I3035,I65807,I65918,);
and I_3697 (I65926,I65918,I378768);
nor I_3698 (I65943,I65901,I65926);
DFFARX1 I_3699 (I65943,I3035,I65807,I65775,);
nand I_3700 (I65974,I65918,I378768);
nand I_3701 (I65991,I65841,I65974);
not I_3702 (I65787,I65991);
DFFARX1 I_3703 (I378762,I3035,I65807,I66031,);
DFFARX1 I_3704 (I66031,I3035,I65807,I65796,);
nand I_3705 (I66053,I378780,I378771);
and I_3706 (I66070,I66053,I378786);
DFFARX1 I_3707 (I66070,I3035,I65807,I66096,);
DFFARX1 I_3708 (I66096,I3035,I65807,I66113,);
not I_3709 (I65799,I66113);
not I_3710 (I66135,I66096);
nand I_3711 (I65784,I66135,I65974);
nor I_3712 (I66166,I378777,I378771);
not I_3713 (I66183,I66166);
nor I_3714 (I66200,I66135,I66183);
nor I_3715 (I66217,I65841,I66200);
DFFARX1 I_3716 (I66217,I3035,I65807,I65793,);
nor I_3717 (I66248,I65901,I66183);
nor I_3718 (I65781,I66096,I66248);
nor I_3719 (I65790,I66031,I66166);
nor I_3720 (I65778,I65901,I66166);
not I_3721 (I66334,I3042);
DFFARX1 I_3722 (I613334,I3035,I66334,I66360,);
not I_3723 (I66368,I66360);
nand I_3724 (I66385,I613349,I613328);
and I_3725 (I66402,I66385,I613331);
DFFARX1 I_3726 (I66402,I3035,I66334,I66428,);
DFFARX1 I_3727 (I613352,I3035,I66334,I66445,);
and I_3728 (I66453,I66445,I613331);
nor I_3729 (I66470,I66428,I66453);
DFFARX1 I_3730 (I66470,I3035,I66334,I66302,);
nand I_3731 (I66501,I66445,I613331);
nand I_3732 (I66518,I66368,I66501);
not I_3733 (I66314,I66518);
DFFARX1 I_3734 (I613328,I3035,I66334,I66558,);
DFFARX1 I_3735 (I66558,I3035,I66334,I66323,);
nand I_3736 (I66580,I613340,I613337);
and I_3737 (I66597,I66580,I613343);
DFFARX1 I_3738 (I66597,I3035,I66334,I66623,);
DFFARX1 I_3739 (I66623,I3035,I66334,I66640,);
not I_3740 (I66326,I66640);
not I_3741 (I66662,I66623);
nand I_3742 (I66311,I66662,I66501);
nor I_3743 (I66693,I613346,I613337);
not I_3744 (I66710,I66693);
nor I_3745 (I66727,I66662,I66710);
nor I_3746 (I66744,I66368,I66727);
DFFARX1 I_3747 (I66744,I3035,I66334,I66320,);
nor I_3748 (I66775,I66428,I66710);
nor I_3749 (I66308,I66623,I66775);
nor I_3750 (I66317,I66558,I66693);
nor I_3751 (I66305,I66428,I66693);
not I_3752 (I66861,I3042);
DFFARX1 I_3753 (I117586,I3035,I66861,I66887,);
not I_3754 (I66895,I66887);
nand I_3755 (I66912,I117580,I117574);
and I_3756 (I66929,I66912,I117595);
DFFARX1 I_3757 (I66929,I3035,I66861,I66955,);
DFFARX1 I_3758 (I117592,I3035,I66861,I66972,);
and I_3759 (I66980,I66972,I117589);
nor I_3760 (I66997,I66955,I66980);
DFFARX1 I_3761 (I66997,I3035,I66861,I66829,);
nand I_3762 (I67028,I66972,I117589);
nand I_3763 (I67045,I66895,I67028);
not I_3764 (I66841,I67045);
DFFARX1 I_3765 (I117574,I3035,I66861,I67085,);
DFFARX1 I_3766 (I67085,I3035,I66861,I66850,);
nand I_3767 (I67107,I117577,I117577);
and I_3768 (I67124,I67107,I117598);
DFFARX1 I_3769 (I67124,I3035,I66861,I67150,);
DFFARX1 I_3770 (I67150,I3035,I66861,I67167,);
not I_3771 (I66853,I67167);
not I_3772 (I67189,I67150);
nand I_3773 (I66838,I67189,I67028);
nor I_3774 (I67220,I117583,I117577);
not I_3775 (I67237,I67220);
nor I_3776 (I67254,I67189,I67237);
nor I_3777 (I67271,I66895,I67254);
DFFARX1 I_3778 (I67271,I3035,I66861,I66847,);
nor I_3779 (I67302,I66955,I67237);
nor I_3780 (I66835,I67150,I67302);
nor I_3781 (I66844,I67085,I67220);
nor I_3782 (I66832,I66955,I67220);
not I_3783 (I67388,I3042);
DFFARX1 I_3784 (I368370,I3035,I67388,I67414,);
not I_3785 (I67422,I67414);
nand I_3786 (I67439,I368361,I368379);
and I_3787 (I67456,I67439,I368358);
DFFARX1 I_3788 (I67456,I3035,I67388,I67482,);
DFFARX1 I_3789 (I368361,I3035,I67388,I67499,);
and I_3790 (I67507,I67499,I368364);
nor I_3791 (I67524,I67482,I67507);
DFFARX1 I_3792 (I67524,I3035,I67388,I67356,);
nand I_3793 (I67555,I67499,I368364);
nand I_3794 (I67572,I67422,I67555);
not I_3795 (I67368,I67572);
DFFARX1 I_3796 (I368358,I3035,I67388,I67612,);
DFFARX1 I_3797 (I67612,I3035,I67388,I67377,);
nand I_3798 (I67634,I368376,I368367);
and I_3799 (I67651,I67634,I368382);
DFFARX1 I_3800 (I67651,I3035,I67388,I67677,);
DFFARX1 I_3801 (I67677,I3035,I67388,I67694,);
not I_3802 (I67380,I67694);
not I_3803 (I67716,I67677);
nand I_3804 (I67365,I67716,I67555);
nor I_3805 (I67747,I368373,I368367);
not I_3806 (I67764,I67747);
nor I_3807 (I67781,I67716,I67764);
nor I_3808 (I67798,I67422,I67781);
DFFARX1 I_3809 (I67798,I3035,I67388,I67374,);
nor I_3810 (I67829,I67482,I67764);
nor I_3811 (I67362,I67677,I67829);
nor I_3812 (I67371,I67612,I67747);
nor I_3813 (I67359,I67482,I67747);
not I_3814 (I67915,I3042);
DFFARX1 I_3815 (I694979,I3035,I67915,I67941,);
not I_3816 (I67949,I67941);
nand I_3817 (I67966,I694985,I695003);
and I_3818 (I67983,I67966,I695000);
DFFARX1 I_3819 (I67983,I3035,I67915,I68009,);
DFFARX1 I_3820 (I694997,I3035,I67915,I68026,);
and I_3821 (I68034,I68026,I694991);
nor I_3822 (I68051,I68009,I68034);
DFFARX1 I_3823 (I68051,I3035,I67915,I67883,);
nand I_3824 (I68082,I68026,I694991);
nand I_3825 (I68099,I67949,I68082);
not I_3826 (I67895,I68099);
DFFARX1 I_3827 (I694979,I3035,I67915,I68139,);
DFFARX1 I_3828 (I68139,I3035,I67915,I67904,);
nand I_3829 (I68161,I694994,I694982);
and I_3830 (I68178,I68161,I695006);
DFFARX1 I_3831 (I68178,I3035,I67915,I68204,);
DFFARX1 I_3832 (I68204,I3035,I67915,I68221,);
not I_3833 (I67907,I68221);
not I_3834 (I68243,I68204);
nand I_3835 (I67892,I68243,I68082);
nor I_3836 (I68274,I694988,I694982);
not I_3837 (I68291,I68274);
nor I_3838 (I68308,I68243,I68291);
nor I_3839 (I68325,I67949,I68308);
DFFARX1 I_3840 (I68325,I3035,I67915,I67901,);
nor I_3841 (I68356,I68009,I68291);
nor I_3842 (I67889,I68204,I68356);
nor I_3843 (I67898,I68139,I68274);
nor I_3844 (I67886,I68009,I68274);
not I_3845 (I68442,I3042);
DFFARX1 I_3846 (I177730,I3035,I68442,I68468,);
not I_3847 (I68476,I68468);
nand I_3848 (I68493,I177712,I177727);
and I_3849 (I68510,I68493,I177703);
DFFARX1 I_3850 (I68510,I3035,I68442,I68536,);
DFFARX1 I_3851 (I177706,I3035,I68442,I68553,);
and I_3852 (I68561,I68553,I177721);
nor I_3853 (I68578,I68536,I68561);
DFFARX1 I_3854 (I68578,I3035,I68442,I68410,);
nand I_3855 (I68609,I68553,I177721);
nand I_3856 (I68626,I68476,I68609);
not I_3857 (I68422,I68626);
DFFARX1 I_3858 (I177724,I3035,I68442,I68666,);
DFFARX1 I_3859 (I68666,I3035,I68442,I68431,);
nand I_3860 (I68688,I177703,I177715);
and I_3861 (I68705,I68688,I177709);
DFFARX1 I_3862 (I68705,I3035,I68442,I68731,);
DFFARX1 I_3863 (I68731,I3035,I68442,I68748,);
not I_3864 (I68434,I68748);
not I_3865 (I68770,I68731);
nand I_3866 (I68419,I68770,I68609);
nor I_3867 (I68801,I177718,I177715);
not I_3868 (I68818,I68801);
nor I_3869 (I68835,I68770,I68818);
nor I_3870 (I68852,I68476,I68835);
DFFARX1 I_3871 (I68852,I3035,I68442,I68428,);
nor I_3872 (I68883,I68536,I68818);
nor I_3873 (I68416,I68731,I68883);
nor I_3874 (I68425,I68666,I68801);
nor I_3875 (I68413,I68536,I68801);
not I_3876 (I68969,I3042);
DFFARX1 I_3877 (I574608,I3035,I68969,I68995,);
not I_3878 (I69003,I68995);
nand I_3879 (I69020,I574623,I574602);
and I_3880 (I69037,I69020,I574605);
DFFARX1 I_3881 (I69037,I3035,I68969,I69063,);
DFFARX1 I_3882 (I574626,I3035,I68969,I69080,);
and I_3883 (I69088,I69080,I574605);
nor I_3884 (I69105,I69063,I69088);
DFFARX1 I_3885 (I69105,I3035,I68969,I68937,);
nand I_3886 (I69136,I69080,I574605);
nand I_3887 (I69153,I69003,I69136);
not I_3888 (I68949,I69153);
DFFARX1 I_3889 (I574602,I3035,I68969,I69193,);
DFFARX1 I_3890 (I69193,I3035,I68969,I68958,);
nand I_3891 (I69215,I574614,I574611);
and I_3892 (I69232,I69215,I574617);
DFFARX1 I_3893 (I69232,I3035,I68969,I69258,);
DFFARX1 I_3894 (I69258,I3035,I68969,I69275,);
not I_3895 (I68961,I69275);
not I_3896 (I69297,I69258);
nand I_3897 (I68946,I69297,I69136);
nor I_3898 (I69328,I574620,I574611);
not I_3899 (I69345,I69328);
nor I_3900 (I69362,I69297,I69345);
nor I_3901 (I69379,I69003,I69362);
DFFARX1 I_3902 (I69379,I3035,I68969,I68955,);
nor I_3903 (I69410,I69063,I69345);
nor I_3904 (I68943,I69258,I69410);
nor I_3905 (I68952,I69193,I69328);
nor I_3906 (I68940,I69063,I69328);
not I_3907 (I69496,I3042);
DFFARX1 I_3908 (I193540,I3035,I69496,I69522,);
not I_3909 (I69530,I69522);
nand I_3910 (I69547,I193522,I193537);
and I_3911 (I69564,I69547,I193513);
DFFARX1 I_3912 (I69564,I3035,I69496,I69590,);
DFFARX1 I_3913 (I193516,I3035,I69496,I69607,);
and I_3914 (I69615,I69607,I193531);
nor I_3915 (I69632,I69590,I69615);
DFFARX1 I_3916 (I69632,I3035,I69496,I69464,);
nand I_3917 (I69663,I69607,I193531);
nand I_3918 (I69680,I69530,I69663);
not I_3919 (I69476,I69680);
DFFARX1 I_3920 (I193534,I3035,I69496,I69720,);
DFFARX1 I_3921 (I69720,I3035,I69496,I69485,);
nand I_3922 (I69742,I193513,I193525);
and I_3923 (I69759,I69742,I193519);
DFFARX1 I_3924 (I69759,I3035,I69496,I69785,);
DFFARX1 I_3925 (I69785,I3035,I69496,I69802,);
not I_3926 (I69488,I69802);
not I_3927 (I69824,I69785);
nand I_3928 (I69473,I69824,I69663);
nor I_3929 (I69855,I193528,I193525);
not I_3930 (I69872,I69855);
nor I_3931 (I69889,I69824,I69872);
nor I_3932 (I69906,I69530,I69889);
DFFARX1 I_3933 (I69906,I3035,I69496,I69482,);
nor I_3934 (I69937,I69590,I69872);
nor I_3935 (I69470,I69785,I69937);
nor I_3936 (I69479,I69720,I69855);
nor I_3937 (I69467,I69590,I69855);
not I_3938 (I70023,I3042);
DFFARX1 I_3939 (I131271,I3035,I70023,I70049,);
not I_3940 (I70057,I70049);
nand I_3941 (I70074,I131265,I131259);
and I_3942 (I70091,I70074,I131280);
DFFARX1 I_3943 (I70091,I3035,I70023,I70117,);
DFFARX1 I_3944 (I131277,I3035,I70023,I70134,);
and I_3945 (I70142,I70134,I131274);
nor I_3946 (I70159,I70117,I70142);
DFFARX1 I_3947 (I70159,I3035,I70023,I69991,);
nand I_3948 (I70190,I70134,I131274);
nand I_3949 (I70207,I70057,I70190);
not I_3950 (I70003,I70207);
DFFARX1 I_3951 (I131259,I3035,I70023,I70247,);
DFFARX1 I_3952 (I70247,I3035,I70023,I70012,);
nand I_3953 (I70269,I131262,I131262);
and I_3954 (I70286,I70269,I131283);
DFFARX1 I_3955 (I70286,I3035,I70023,I70312,);
DFFARX1 I_3956 (I70312,I3035,I70023,I70329,);
not I_3957 (I70015,I70329);
not I_3958 (I70351,I70312);
nand I_3959 (I70000,I70351,I70190);
nor I_3960 (I70382,I131268,I131262);
not I_3961 (I70399,I70382);
nor I_3962 (I70416,I70351,I70399);
nor I_3963 (I70433,I70057,I70416);
DFFARX1 I_3964 (I70433,I3035,I70023,I70009,);
nor I_3965 (I70464,I70117,I70399);
nor I_3966 (I69997,I70312,I70464);
nor I_3967 (I70006,I70247,I70382);
nor I_3968 (I69994,I70117,I70382);
not I_3969 (I70550,I3042);
DFFARX1 I_3970 (I652332,I3035,I70550,I70576,);
not I_3971 (I70584,I70576);
nand I_3972 (I70601,I652326,I652347);
and I_3973 (I70618,I70601,I652338);
DFFARX1 I_3974 (I70618,I3035,I70550,I70644,);
DFFARX1 I_3975 (I652329,I3035,I70550,I70661,);
and I_3976 (I70669,I70661,I652341);
nor I_3977 (I70686,I70644,I70669);
DFFARX1 I_3978 (I70686,I3035,I70550,I70518,);
nand I_3979 (I70717,I70661,I652341);
nand I_3980 (I70734,I70584,I70717);
not I_3981 (I70530,I70734);
DFFARX1 I_3982 (I652329,I3035,I70550,I70774,);
DFFARX1 I_3983 (I70774,I3035,I70550,I70539,);
nand I_3984 (I70796,I652350,I652335);
and I_3985 (I70813,I70796,I652326);
DFFARX1 I_3986 (I70813,I3035,I70550,I70839,);
DFFARX1 I_3987 (I70839,I3035,I70550,I70856,);
not I_3988 (I70542,I70856);
not I_3989 (I70878,I70839);
nand I_3990 (I70527,I70878,I70717);
nor I_3991 (I70909,I652344,I652335);
not I_3992 (I70926,I70909);
nor I_3993 (I70943,I70878,I70926);
nor I_3994 (I70960,I70584,I70943);
DFFARX1 I_3995 (I70960,I3035,I70550,I70536,);
nor I_3996 (I70991,I70644,I70926);
nor I_3997 (I70524,I70839,I70991);
nor I_3998 (I70533,I70774,I70909);
nor I_3999 (I70521,I70644,I70909);
not I_4000 (I71077,I3042);
DFFARX1 I_4001 (I592526,I3035,I71077,I71103,);
not I_4002 (I71111,I71103);
nand I_4003 (I71128,I592541,I592520);
and I_4004 (I71145,I71128,I592523);
DFFARX1 I_4005 (I71145,I3035,I71077,I71171,);
DFFARX1 I_4006 (I592544,I3035,I71077,I71188,);
and I_4007 (I71196,I71188,I592523);
nor I_4008 (I71213,I71171,I71196);
DFFARX1 I_4009 (I71213,I3035,I71077,I71045,);
nand I_4010 (I71244,I71188,I592523);
nand I_4011 (I71261,I71111,I71244);
not I_4012 (I71057,I71261);
DFFARX1 I_4013 (I592520,I3035,I71077,I71301,);
DFFARX1 I_4014 (I71301,I3035,I71077,I71066,);
nand I_4015 (I71323,I592532,I592529);
and I_4016 (I71340,I71323,I592535);
DFFARX1 I_4017 (I71340,I3035,I71077,I71366,);
DFFARX1 I_4018 (I71366,I3035,I71077,I71383,);
not I_4019 (I71069,I71383);
not I_4020 (I71405,I71366);
nand I_4021 (I71054,I71405,I71244);
nor I_4022 (I71436,I592538,I592529);
not I_4023 (I71453,I71436);
nor I_4024 (I71470,I71405,I71453);
nor I_4025 (I71487,I71111,I71470);
DFFARX1 I_4026 (I71487,I3035,I71077,I71063,);
nor I_4027 (I71518,I71171,I71453);
nor I_4028 (I71051,I71366,I71518);
nor I_4029 (I71060,I71301,I71436);
nor I_4030 (I71048,I71171,I71436);
not I_4031 (I71604,I3042);
DFFARX1 I_4032 (I199337,I3035,I71604,I71630,);
not I_4033 (I71638,I71630);
nand I_4034 (I71655,I199319,I199334);
and I_4035 (I71672,I71655,I199310);
DFFARX1 I_4036 (I71672,I3035,I71604,I71698,);
DFFARX1 I_4037 (I199313,I3035,I71604,I71715,);
and I_4038 (I71723,I71715,I199328);
nor I_4039 (I71740,I71698,I71723);
DFFARX1 I_4040 (I71740,I3035,I71604,I71572,);
nand I_4041 (I71771,I71715,I199328);
nand I_4042 (I71788,I71638,I71771);
not I_4043 (I71584,I71788);
DFFARX1 I_4044 (I199331,I3035,I71604,I71828,);
DFFARX1 I_4045 (I71828,I3035,I71604,I71593,);
nand I_4046 (I71850,I199310,I199322);
and I_4047 (I71867,I71850,I199316);
DFFARX1 I_4048 (I71867,I3035,I71604,I71893,);
DFFARX1 I_4049 (I71893,I3035,I71604,I71910,);
not I_4050 (I71596,I71910);
not I_4051 (I71932,I71893);
nand I_4052 (I71581,I71932,I71771);
nor I_4053 (I71963,I199325,I199322);
not I_4054 (I71980,I71963);
nor I_4055 (I71997,I71932,I71980);
nor I_4056 (I72014,I71638,I71997);
DFFARX1 I_4057 (I72014,I3035,I71604,I71590,);
nor I_4058 (I72045,I71698,I71980);
nor I_4059 (I71578,I71893,I72045);
nor I_4060 (I71587,I71828,I71963);
nor I_4061 (I71575,I71698,I71963);
not I_4062 (I72131,I3042);
DFFARX1 I_4063 (I348718,I3035,I72131,I72157,);
not I_4064 (I72165,I72157);
nand I_4065 (I72182,I348709,I348727);
and I_4066 (I72199,I72182,I348706);
DFFARX1 I_4067 (I72199,I3035,I72131,I72225,);
DFFARX1 I_4068 (I348709,I3035,I72131,I72242,);
and I_4069 (I72250,I72242,I348712);
nor I_4070 (I72267,I72225,I72250);
DFFARX1 I_4071 (I72267,I3035,I72131,I72099,);
nand I_4072 (I72298,I72242,I348712);
nand I_4073 (I72315,I72165,I72298);
not I_4074 (I72111,I72315);
DFFARX1 I_4075 (I348706,I3035,I72131,I72355,);
DFFARX1 I_4076 (I72355,I3035,I72131,I72120,);
nand I_4077 (I72377,I348724,I348715);
and I_4078 (I72394,I72377,I348730);
DFFARX1 I_4079 (I72394,I3035,I72131,I72420,);
DFFARX1 I_4080 (I72420,I3035,I72131,I72437,);
not I_4081 (I72123,I72437);
not I_4082 (I72459,I72420);
nand I_4083 (I72108,I72459,I72298);
nor I_4084 (I72490,I348721,I348715);
not I_4085 (I72507,I72490);
nor I_4086 (I72524,I72459,I72507);
nor I_4087 (I72541,I72165,I72524);
DFFARX1 I_4088 (I72541,I3035,I72131,I72117,);
nor I_4089 (I72572,I72225,I72507);
nor I_4090 (I72105,I72420,I72572);
nor I_4091 (I72114,I72355,I72490);
nor I_4092 (I72102,I72225,I72490);
not I_4093 (I72658,I3042);
DFFARX1 I_4094 (I533573,I3035,I72658,I72684,);
not I_4095 (I72692,I72684);
nand I_4096 (I72709,I533591,I533585);
and I_4097 (I72726,I72709,I533564);
DFFARX1 I_4098 (I72726,I3035,I72658,I72752,);
DFFARX1 I_4099 (I533582,I3035,I72658,I72769,);
and I_4100 (I72777,I72769,I533567);
nor I_4101 (I72794,I72752,I72777);
DFFARX1 I_4102 (I72794,I3035,I72658,I72626,);
nand I_4103 (I72825,I72769,I533567);
nand I_4104 (I72842,I72692,I72825);
not I_4105 (I72638,I72842);
DFFARX1 I_4106 (I533579,I3035,I72658,I72882,);
DFFARX1 I_4107 (I72882,I3035,I72658,I72647,);
nand I_4108 (I72904,I533588,I533576);
and I_4109 (I72921,I72904,I533570);
DFFARX1 I_4110 (I72921,I3035,I72658,I72947,);
DFFARX1 I_4111 (I72947,I3035,I72658,I72964,);
not I_4112 (I72650,I72964);
not I_4113 (I72986,I72947);
nand I_4114 (I72635,I72986,I72825);
nor I_4115 (I73017,I533564,I533576);
not I_4116 (I73034,I73017);
nor I_4117 (I73051,I72986,I73034);
nor I_4118 (I73068,I72692,I73051);
DFFARX1 I_4119 (I73068,I3035,I72658,I72644,);
nor I_4120 (I73099,I72752,I73034);
nor I_4121 (I72632,I72947,I73099);
nor I_4122 (I72641,I72882,I73017);
nor I_4123 (I72629,I72752,I73017);
not I_4124 (I73185,I3042);
DFFARX1 I_4125 (I152434,I3035,I73185,I73211,);
not I_4126 (I73219,I73211);
nand I_4127 (I73236,I152416,I152431);
and I_4128 (I73253,I73236,I152407);
DFFARX1 I_4129 (I73253,I3035,I73185,I73279,);
DFFARX1 I_4130 (I152410,I3035,I73185,I73296,);
and I_4131 (I73304,I73296,I152425);
nor I_4132 (I73321,I73279,I73304);
DFFARX1 I_4133 (I73321,I3035,I73185,I73153,);
nand I_4134 (I73352,I73296,I152425);
nand I_4135 (I73369,I73219,I73352);
not I_4136 (I73165,I73369);
DFFARX1 I_4137 (I152428,I3035,I73185,I73409,);
DFFARX1 I_4138 (I73409,I3035,I73185,I73174,);
nand I_4139 (I73431,I152407,I152419);
and I_4140 (I73448,I73431,I152413);
DFFARX1 I_4141 (I73448,I3035,I73185,I73474,);
DFFARX1 I_4142 (I73474,I3035,I73185,I73491,);
not I_4143 (I73177,I73491);
not I_4144 (I73513,I73474);
nand I_4145 (I73162,I73513,I73352);
nor I_4146 (I73544,I152422,I152419);
not I_4147 (I73561,I73544);
nor I_4148 (I73578,I73513,I73561);
nor I_4149 (I73595,I73219,I73578);
DFFARX1 I_4150 (I73595,I3035,I73185,I73171,);
nor I_4151 (I73626,I73279,I73561);
nor I_4152 (I73159,I73474,I73626);
nor I_4153 (I73168,I73409,I73544);
nor I_4154 (I73156,I73279,I73544);
not I_4155 (I73712,I3042);
DFFARX1 I_4156 (I248407,I3035,I73712,I73738,);
not I_4157 (I73746,I73738);
nand I_4158 (I73763,I248401,I248392);
and I_4159 (I73780,I73763,I248413);
DFFARX1 I_4160 (I73780,I3035,I73712,I73806,);
DFFARX1 I_4161 (I248395,I3035,I73712,I73823,);
and I_4162 (I73831,I73823,I248389);
nor I_4163 (I73848,I73806,I73831);
DFFARX1 I_4164 (I73848,I3035,I73712,I73680,);
nand I_4165 (I73879,I73823,I248389);
nand I_4166 (I73896,I73746,I73879);
not I_4167 (I73692,I73896);
DFFARX1 I_4168 (I248389,I3035,I73712,I73936,);
DFFARX1 I_4169 (I73936,I3035,I73712,I73701,);
nand I_4170 (I73958,I248416,I248398);
and I_4171 (I73975,I73958,I248404);
DFFARX1 I_4172 (I73975,I3035,I73712,I74001,);
DFFARX1 I_4173 (I74001,I3035,I73712,I74018,);
not I_4174 (I73704,I74018);
not I_4175 (I74040,I74001);
nand I_4176 (I73689,I74040,I73879);
nor I_4177 (I74071,I248410,I248398);
not I_4178 (I74088,I74071);
nor I_4179 (I74105,I74040,I74088);
nor I_4180 (I74122,I73746,I74105);
DFFARX1 I_4181 (I74122,I3035,I73712,I73698,);
nor I_4182 (I74153,I73806,I74088);
nor I_4183 (I73686,I74001,I74153);
nor I_4184 (I73695,I73936,I74071);
nor I_4185 (I73683,I73806,I74071);
not I_4186 (I74239,I3042);
DFFARX1 I_4187 (I441416,I3035,I74239,I74265,);
not I_4188 (I74273,I74265);
nand I_4189 (I74290,I441413,I441428);
and I_4190 (I74307,I74290,I441410);
DFFARX1 I_4191 (I74307,I3035,I74239,I74333,);
DFFARX1 I_4192 (I441407,I3035,I74239,I74350,);
and I_4193 (I74358,I74350,I441407);
nor I_4194 (I74375,I74333,I74358);
DFFARX1 I_4195 (I74375,I3035,I74239,I74207,);
nand I_4196 (I74406,I74350,I441407);
nand I_4197 (I74423,I74273,I74406);
not I_4198 (I74219,I74423);
DFFARX1 I_4199 (I441410,I3035,I74239,I74463,);
DFFARX1 I_4200 (I74463,I3035,I74239,I74228,);
nand I_4201 (I74485,I441422,I441413);
and I_4202 (I74502,I74485,I441425);
DFFARX1 I_4203 (I74502,I3035,I74239,I74528,);
DFFARX1 I_4204 (I74528,I3035,I74239,I74545,);
not I_4205 (I74231,I74545);
not I_4206 (I74567,I74528);
nand I_4207 (I74216,I74567,I74406);
nor I_4208 (I74598,I441419,I441413);
not I_4209 (I74615,I74598);
nor I_4210 (I74632,I74567,I74615);
nor I_4211 (I74649,I74273,I74632);
DFFARX1 I_4212 (I74649,I3035,I74239,I74225,);
nor I_4213 (I74680,I74333,I74615);
nor I_4214 (I74213,I74528,I74680);
nor I_4215 (I74222,I74463,I74598);
nor I_4216 (I74210,I74333,I74598);
not I_4217 (I74769,I3042);
DFFARX1 I_4218 (I287688,I3035,I74769,I74795,);
not I_4219 (I74803,I74795);
DFFARX1 I_4220 (I287694,I3035,I74769,I74829,);
not I_4221 (I74837,I287676);
or I_4222 (I74854,I287700,I287676);
nor I_4223 (I74871,I74829,I287700);
nand I_4224 (I74746,I74837,I74871);
nor I_4225 (I74902,I287691,I287700);
nand I_4226 (I74740,I74902,I74837);
not I_4227 (I74933,I287682);
nand I_4228 (I74950,I74837,I74933);
nor I_4229 (I74967,I287685,I287679);
not I_4230 (I74984,I74967);
nor I_4231 (I75001,I74984,I74950);
nor I_4232 (I75018,I74902,I75001);
DFFARX1 I_4233 (I75018,I3035,I74769,I74755,);
nor I_4234 (I74752,I74967,I74854);
DFFARX1 I_4235 (I74967,I3035,I74769,I74758,);
nor I_4236 (I75077,I74933,I287685);
nor I_4237 (I75094,I75077,I287676);
nor I_4238 (I75111,I287697,I287676);
DFFARX1 I_4239 (I75111,I3035,I74769,I75137,);
nor I_4240 (I74737,I75137,I75094);
DFFARX1 I_4241 (I75137,I3035,I74769,I75168,);
nand I_4242 (I75176,I75168,I287679);
nor I_4243 (I74761,I74803,I75176);
not I_4244 (I75207,I75137);
nand I_4245 (I75224,I75207,I287679);
nor I_4246 (I75241,I74803,I75224);
nor I_4247 (I74743,I74829,I75241);
nor I_4248 (I75272,I287697,I287691);
nor I_4249 (I75289,I74829,I75272);
DFFARX1 I_4250 (I75289,I3035,I74769,I74734,);
and I_4251 (I74749,I74902,I287697);
not I_4252 (I75364,I3042);
DFFARX1 I_4253 (I130688,I3035,I75364,I75390,);
not I_4254 (I75398,I75390);
DFFARX1 I_4255 (I130682,I3035,I75364,I75424,);
not I_4256 (I75432,I130667);
or I_4257 (I75449,I130676,I130667);
nor I_4258 (I75466,I75424,I130676);
nand I_4259 (I75341,I75432,I75466);
nor I_4260 (I75497,I130664,I130676);
nand I_4261 (I75335,I75497,I75432);
not I_4262 (I75528,I130670);
nand I_4263 (I75545,I75432,I75528);
nor I_4264 (I75562,I130673,I130685);
not I_4265 (I75579,I75562);
nor I_4266 (I75596,I75579,I75545);
nor I_4267 (I75613,I75497,I75596);
DFFARX1 I_4268 (I75613,I3035,I75364,I75350,);
nor I_4269 (I75347,I75562,I75449);
DFFARX1 I_4270 (I75562,I3035,I75364,I75353,);
nor I_4271 (I75672,I75528,I130673);
nor I_4272 (I75689,I75672,I130667);
nor I_4273 (I75706,I130679,I130667);
DFFARX1 I_4274 (I75706,I3035,I75364,I75732,);
nor I_4275 (I75332,I75732,I75689);
DFFARX1 I_4276 (I75732,I3035,I75364,I75763,);
nand I_4277 (I75771,I75763,I130664);
nor I_4278 (I75356,I75398,I75771);
not I_4279 (I75802,I75732);
nand I_4280 (I75819,I75802,I130664);
nor I_4281 (I75836,I75398,I75819);
nor I_4282 (I75338,I75424,I75836);
nor I_4283 (I75867,I130679,I130664);
nor I_4284 (I75884,I75424,I75867);
DFFARX1 I_4285 (I75884,I3035,I75364,I75329,);
and I_4286 (I75344,I75497,I130679);
not I_4287 (I75959,I3042);
DFFARX1 I_4288 (I107483,I3035,I75959,I75985,);
not I_4289 (I75993,I75985);
DFFARX1 I_4290 (I107477,I3035,I75959,I76019,);
not I_4291 (I76027,I107462);
or I_4292 (I76044,I107471,I107462);
nor I_4293 (I76061,I76019,I107471);
nand I_4294 (I75936,I76027,I76061);
nor I_4295 (I76092,I107459,I107471);
nand I_4296 (I75930,I76092,I76027);
not I_4297 (I76123,I107465);
nand I_4298 (I76140,I76027,I76123);
nor I_4299 (I76157,I107468,I107480);
not I_4300 (I76174,I76157);
nor I_4301 (I76191,I76174,I76140);
nor I_4302 (I76208,I76092,I76191);
DFFARX1 I_4303 (I76208,I3035,I75959,I75945,);
nor I_4304 (I75942,I76157,I76044);
DFFARX1 I_4305 (I76157,I3035,I75959,I75948,);
nor I_4306 (I76267,I76123,I107468);
nor I_4307 (I76284,I76267,I107462);
nor I_4308 (I76301,I107474,I107462);
DFFARX1 I_4309 (I76301,I3035,I75959,I76327,);
nor I_4310 (I75927,I76327,I76284);
DFFARX1 I_4311 (I76327,I3035,I75959,I76358,);
nand I_4312 (I76366,I76358,I107459);
nor I_4313 (I75951,I75993,I76366);
not I_4314 (I76397,I76327);
nand I_4315 (I76414,I76397,I107459);
nor I_4316 (I76431,I75993,I76414);
nor I_4317 (I75933,I76019,I76431);
nor I_4318 (I76462,I107474,I107459);
nor I_4319 (I76479,I76019,I76462);
DFFARX1 I_4320 (I76479,I3035,I75959,I75924,);
and I_4321 (I75939,I76092,I107474);
not I_4322 (I76554,I3042);
DFFARX1 I_4323 (I249501,I3035,I76554,I76580,);
not I_4324 (I76588,I76580);
DFFARX1 I_4325 (I249495,I3035,I76554,I76614,);
not I_4326 (I76622,I249492);
or I_4327 (I76639,I249483,I249492);
nor I_4328 (I76656,I76614,I249483);
nand I_4329 (I76531,I76622,I76656);
nor I_4330 (I76687,I249486,I249483);
nand I_4331 (I76525,I76687,I76622);
not I_4332 (I76718,I249489);
nand I_4333 (I76735,I76622,I76718);
nor I_4334 (I76752,I249477,I249504);
not I_4335 (I76769,I76752);
nor I_4336 (I76786,I76769,I76735);
nor I_4337 (I76803,I76687,I76786);
DFFARX1 I_4338 (I76803,I3035,I76554,I76540,);
nor I_4339 (I76537,I76752,I76639);
DFFARX1 I_4340 (I76752,I3035,I76554,I76543,);
nor I_4341 (I76862,I76718,I249477);
nor I_4342 (I76879,I76862,I249492);
nor I_4343 (I76896,I249480,I249477);
DFFARX1 I_4344 (I76896,I3035,I76554,I76922,);
nor I_4345 (I76522,I76922,I76879);
DFFARX1 I_4346 (I76922,I3035,I76554,I76953,);
nand I_4347 (I76961,I76953,I249498);
nor I_4348 (I76546,I76588,I76961);
not I_4349 (I76992,I76922);
nand I_4350 (I77009,I76992,I249498);
nor I_4351 (I77026,I76588,I77009);
nor I_4352 (I76528,I76614,I77026);
nor I_4353 (I77057,I249480,I249486);
nor I_4354 (I77074,I76614,I77057);
DFFARX1 I_4355 (I77074,I3035,I76554,I76519,);
and I_4356 (I76534,I76687,I249480);
not I_4357 (I77149,I3042);
DFFARX1 I_4358 (I494164,I3035,I77149,I77175,);
not I_4359 (I77183,I77175);
DFFARX1 I_4360 (I494185,I3035,I77149,I77209,);
not I_4361 (I77217,I494167);
or I_4362 (I77234,I494158,I494167);
nor I_4363 (I77251,I77209,I494158);
nand I_4364 (I77126,I77217,I77251);
nor I_4365 (I77282,I494170,I494158);
nand I_4366 (I77120,I77282,I77217);
not I_4367 (I77313,I494161);
nand I_4368 (I77330,I77217,I77313);
nor I_4369 (I77347,I494179,I494182);
not I_4370 (I77364,I77347);
nor I_4371 (I77381,I77364,I77330);
nor I_4372 (I77398,I77282,I77381);
DFFARX1 I_4373 (I77398,I3035,I77149,I77135,);
nor I_4374 (I77132,I77347,I77234);
DFFARX1 I_4375 (I77347,I3035,I77149,I77138,);
nor I_4376 (I77457,I77313,I494179);
nor I_4377 (I77474,I77457,I494167);
nor I_4378 (I77491,I494173,I494176);
DFFARX1 I_4379 (I77491,I3035,I77149,I77517,);
nor I_4380 (I77117,I77517,I77474);
DFFARX1 I_4381 (I77517,I3035,I77149,I77548,);
nand I_4382 (I77556,I77548,I494158);
nor I_4383 (I77141,I77183,I77556);
not I_4384 (I77587,I77517);
nand I_4385 (I77604,I77587,I494158);
nor I_4386 (I77621,I77183,I77604);
nor I_4387 (I77123,I77209,I77621);
nor I_4388 (I77652,I494173,I494170);
nor I_4389 (I77669,I77209,I77652);
DFFARX1 I_4390 (I77669,I3035,I77149,I77114,);
and I_4391 (I77129,I77282,I494173);
not I_4392 (I77744,I3042);
DFFARX1 I_4393 (I374138,I3035,I77744,I77770,);
not I_4394 (I77778,I77770);
DFFARX1 I_4395 (I374159,I3035,I77744,I77804,);
not I_4396 (I77812,I374138);
or I_4397 (I77829,I374150,I374138);
nor I_4398 (I77846,I77804,I374150);
nand I_4399 (I77721,I77812,I77846);
nor I_4400 (I77877,I374147,I374150);
nand I_4401 (I77715,I77877,I77812);
not I_4402 (I77908,I374156);
nand I_4403 (I77925,I77812,I77908);
nor I_4404 (I77942,I374141,I374141);
not I_4405 (I77959,I77942);
nor I_4406 (I77976,I77959,I77925);
nor I_4407 (I77993,I77877,I77976);
DFFARX1 I_4408 (I77993,I3035,I77744,I77730,);
nor I_4409 (I77727,I77942,I77829);
DFFARX1 I_4410 (I77942,I3035,I77744,I77733,);
nor I_4411 (I78052,I77908,I374141);
nor I_4412 (I78069,I78052,I374138);
nor I_4413 (I78086,I374162,I374144);
DFFARX1 I_4414 (I78086,I3035,I77744,I78112,);
nor I_4415 (I77712,I78112,I78069);
DFFARX1 I_4416 (I78112,I3035,I77744,I78143,);
nand I_4417 (I78151,I78143,I374153);
nor I_4418 (I77736,I77778,I78151);
not I_4419 (I78182,I78112);
nand I_4420 (I78199,I78182,I374153);
nor I_4421 (I78216,I77778,I78199);
nor I_4422 (I77718,I77804,I78216);
nor I_4423 (I78247,I374162,I374147);
nor I_4424 (I78264,I77804,I78247);
DFFARX1 I_4425 (I78264,I3035,I77744,I77709,);
and I_4426 (I77724,I77877,I374162);
not I_4427 (I78339,I3042);
DFFARX1 I_4428 (I342926,I3035,I78339,I78365,);
not I_4429 (I78373,I78365);
DFFARX1 I_4430 (I342947,I3035,I78339,I78399,);
not I_4431 (I78407,I342926);
or I_4432 (I78424,I342938,I342926);
nor I_4433 (I78441,I78399,I342938);
nand I_4434 (I78316,I78407,I78441);
nor I_4435 (I78472,I342935,I342938);
nand I_4436 (I78310,I78472,I78407);
not I_4437 (I78503,I342944);
nand I_4438 (I78520,I78407,I78503);
nor I_4439 (I78537,I342929,I342929);
not I_4440 (I78554,I78537);
nor I_4441 (I78571,I78554,I78520);
nor I_4442 (I78588,I78472,I78571);
DFFARX1 I_4443 (I78588,I3035,I78339,I78325,);
nor I_4444 (I78322,I78537,I78424);
DFFARX1 I_4445 (I78537,I3035,I78339,I78328,);
nor I_4446 (I78647,I78503,I342929);
nor I_4447 (I78664,I78647,I342926);
nor I_4448 (I78681,I342950,I342932);
DFFARX1 I_4449 (I78681,I3035,I78339,I78707,);
nor I_4450 (I78307,I78707,I78664);
DFFARX1 I_4451 (I78707,I3035,I78339,I78738,);
nand I_4452 (I78746,I78738,I342941);
nor I_4453 (I78331,I78373,I78746);
not I_4454 (I78777,I78707);
nand I_4455 (I78794,I78777,I342941);
nor I_4456 (I78811,I78373,I78794);
nor I_4457 (I78313,I78399,I78811);
nor I_4458 (I78842,I342950,I342935);
nor I_4459 (I78859,I78399,I78842);
DFFARX1 I_4460 (I78859,I3035,I78339,I78304,);
and I_4461 (I78319,I78472,I342950);
not I_4462 (I78931,I3042);
DFFARX1 I_4463 (I698434,I3035,I78931,I78957,);
DFFARX1 I_4464 (I78957,I3035,I78931,I78974,);
not I_4465 (I78923,I78974);
not I_4466 (I78996,I78957);
DFFARX1 I_4467 (I698425,I3035,I78931,I79022,);
not I_4468 (I79030,I79022);
and I_4469 (I79047,I78996,I698419);
not I_4470 (I79064,I698413);
nand I_4471 (I79081,I79064,I698419);
not I_4472 (I79098,I698440);
nor I_4473 (I79115,I79098,I698413);
nand I_4474 (I79132,I79115,I698437);
nor I_4475 (I79149,I79132,I79081);
DFFARX1 I_4476 (I79149,I3035,I78931,I78899,);
not I_4477 (I79180,I79132);
not I_4478 (I79197,I698413);
nand I_4479 (I79214,I79197,I698419);
nor I_4480 (I79231,I698413,I698413);
nand I_4481 (I78911,I79047,I79231);
nand I_4482 (I78905,I78996,I698413);
nand I_4483 (I79276,I79098,I698422);
DFFARX1 I_4484 (I79276,I3035,I78931,I78920,);
DFFARX1 I_4485 (I79276,I3035,I78931,I78914,);
not I_4486 (I79321,I698422);
nor I_4487 (I79338,I79321,I698428);
and I_4488 (I79355,I79338,I698431);
or I_4489 (I79372,I79355,I698416);
DFFARX1 I_4490 (I79372,I3035,I78931,I79398,);
nand I_4491 (I79406,I79398,I79064);
nor I_4492 (I78908,I79406,I79214);
nor I_4493 (I78902,I79398,I79030);
DFFARX1 I_4494 (I79398,I3035,I78931,I79460,);
not I_4495 (I79468,I79460);
nor I_4496 (I78917,I79468,I79180);
not I_4497 (I79526,I3042);
DFFARX1 I_4498 (I576914,I3035,I79526,I79552,);
DFFARX1 I_4499 (I79552,I3035,I79526,I79569,);
not I_4500 (I79518,I79569);
not I_4501 (I79591,I79552);
DFFARX1 I_4502 (I576914,I3035,I79526,I79617,);
not I_4503 (I79625,I79617);
and I_4504 (I79642,I79591,I576917);
not I_4505 (I79659,I576929);
nand I_4506 (I79676,I79659,I576917);
not I_4507 (I79693,I576935);
nor I_4508 (I79710,I79693,I576926);
nand I_4509 (I79727,I79710,I576932);
nor I_4510 (I79744,I79727,I79676);
DFFARX1 I_4511 (I79744,I3035,I79526,I79494,);
not I_4512 (I79775,I79727);
not I_4513 (I79792,I576926);
nand I_4514 (I79809,I79792,I576917);
nor I_4515 (I79826,I576926,I576929);
nand I_4516 (I79506,I79642,I79826);
nand I_4517 (I79500,I79591,I576926);
nand I_4518 (I79871,I79693,I576923);
DFFARX1 I_4519 (I79871,I3035,I79526,I79515,);
DFFARX1 I_4520 (I79871,I3035,I79526,I79509,);
not I_4521 (I79916,I576923);
nor I_4522 (I79933,I79916,I576920);
and I_4523 (I79950,I79933,I576938);
or I_4524 (I79967,I79950,I576917);
DFFARX1 I_4525 (I79967,I3035,I79526,I79993,);
nand I_4526 (I80001,I79993,I79659);
nor I_4527 (I79503,I80001,I79809);
nor I_4528 (I79497,I79993,I79625);
DFFARX1 I_4529 (I79993,I3035,I79526,I80055,);
not I_4530 (I80063,I80055);
nor I_4531 (I79512,I80063,I79775);
not I_4532 (I80121,I3042);
DFFARX1 I_4533 (I509677,I3035,I80121,I80147,);
DFFARX1 I_4534 (I80147,I3035,I80121,I80164,);
not I_4535 (I80113,I80164);
not I_4536 (I80186,I80147);
DFFARX1 I_4537 (I509686,I3035,I80121,I80212,);
not I_4538 (I80220,I80212);
and I_4539 (I80237,I80186,I509674);
not I_4540 (I80254,I509665);
nand I_4541 (I80271,I80254,I509674);
not I_4542 (I80288,I509671);
nor I_4543 (I80305,I80288,I509689);
nand I_4544 (I80322,I80305,I509662);
nor I_4545 (I80339,I80322,I80271);
DFFARX1 I_4546 (I80339,I3035,I80121,I80089,);
not I_4547 (I80370,I80322);
not I_4548 (I80387,I509689);
nand I_4549 (I80404,I80387,I509674);
nor I_4550 (I80421,I509689,I509665);
nand I_4551 (I80101,I80237,I80421);
nand I_4552 (I80095,I80186,I509689);
nand I_4553 (I80466,I80288,I509668);
DFFARX1 I_4554 (I80466,I3035,I80121,I80110,);
DFFARX1 I_4555 (I80466,I3035,I80121,I80104,);
not I_4556 (I80511,I509668);
nor I_4557 (I80528,I80511,I509680);
and I_4558 (I80545,I80528,I509662);
or I_4559 (I80562,I80545,I509683);
DFFARX1 I_4560 (I80562,I3035,I80121,I80588,);
nand I_4561 (I80596,I80588,I80254);
nor I_4562 (I80098,I80596,I80404);
nor I_4563 (I80092,I80588,I80220);
DFFARX1 I_4564 (I80588,I3035,I80121,I80650,);
not I_4565 (I80658,I80650);
nor I_4566 (I80107,I80658,I80370);
not I_4567 (I80716,I3042);
DFFARX1 I_4568 (I673647,I3035,I80716,I80742,);
DFFARX1 I_4569 (I80742,I3035,I80716,I80759,);
not I_4570 (I80708,I80759);
not I_4571 (I80781,I80742);
DFFARX1 I_4572 (I673659,I3035,I80716,I80807,);
not I_4573 (I80815,I80807);
and I_4574 (I80832,I80781,I673653);
not I_4575 (I80849,I673665);
nand I_4576 (I80866,I80849,I673653);
not I_4577 (I80883,I673650);
nor I_4578 (I80900,I80883,I673662);
nand I_4579 (I80917,I80900,I673644);
nor I_4580 (I80934,I80917,I80866);
DFFARX1 I_4581 (I80934,I3035,I80716,I80684,);
not I_4582 (I80965,I80917);
not I_4583 (I80982,I673662);
nand I_4584 (I80999,I80982,I673653);
nor I_4585 (I81016,I673662,I673665);
nand I_4586 (I80696,I80832,I81016);
nand I_4587 (I80690,I80781,I673662);
nand I_4588 (I81061,I80883,I673656);
DFFARX1 I_4589 (I81061,I3035,I80716,I80705,);
DFFARX1 I_4590 (I81061,I3035,I80716,I80699,);
not I_4591 (I81106,I673656);
nor I_4592 (I81123,I81106,I673647);
and I_4593 (I81140,I81123,I673644);
or I_4594 (I81157,I81140,I673668);
DFFARX1 I_4595 (I81157,I3035,I80716,I81183,);
nand I_4596 (I81191,I81183,I80849);
nor I_4597 (I80693,I81191,I80999);
nor I_4598 (I80687,I81183,I80815);
DFFARX1 I_4599 (I81183,I3035,I80716,I81245,);
not I_4600 (I81253,I81245);
nor I_4601 (I80702,I81253,I80965);
not I_4602 (I81311,I3042);
DFFARX1 I_4603 (I235901,I3035,I81311,I81337,);
DFFARX1 I_4604 (I81337,I3035,I81311,I81354,);
not I_4605 (I81303,I81354);
not I_4606 (I81376,I81337);
DFFARX1 I_4607 (I235889,I3035,I81311,I81402,);
not I_4608 (I81410,I81402);
and I_4609 (I81427,I81376,I235898);
not I_4610 (I81444,I235895);
nand I_4611 (I81461,I81444,I235898);
not I_4612 (I81478,I235886);
nor I_4613 (I81495,I81478,I235892);
nand I_4614 (I81512,I81495,I235877);
nor I_4615 (I81529,I81512,I81461);
DFFARX1 I_4616 (I81529,I3035,I81311,I81279,);
not I_4617 (I81560,I81512);
not I_4618 (I81577,I235892);
nand I_4619 (I81594,I81577,I235898);
nor I_4620 (I81611,I235892,I235895);
nand I_4621 (I81291,I81427,I81611);
nand I_4622 (I81285,I81376,I235892);
nand I_4623 (I81656,I81478,I235877);
DFFARX1 I_4624 (I81656,I3035,I81311,I81300,);
DFFARX1 I_4625 (I81656,I3035,I81311,I81294,);
not I_4626 (I81701,I235877);
nor I_4627 (I81718,I81701,I235883);
and I_4628 (I81735,I81718,I235880);
or I_4629 (I81752,I81735,I235904);
DFFARX1 I_4630 (I81752,I3035,I81311,I81778,);
nand I_4631 (I81786,I81778,I81444);
nor I_4632 (I81288,I81786,I81594);
nor I_4633 (I81282,I81778,I81410);
DFFARX1 I_4634 (I81778,I3035,I81311,I81840,);
not I_4635 (I81848,I81840);
nor I_4636 (I81297,I81848,I81560);
not I_4637 (I81906,I3042);
DFFARX1 I_4638 (I188243,I3035,I81906,I81932,);
DFFARX1 I_4639 (I81932,I3035,I81906,I81949,);
not I_4640 (I81898,I81949);
not I_4641 (I81971,I81932);
DFFARX1 I_4642 (I188258,I3035,I81906,I81997,);
not I_4643 (I82005,I81997);
and I_4644 (I82022,I81971,I188255);
not I_4645 (I82039,I188243);
nand I_4646 (I82056,I82039,I188255);
not I_4647 (I82073,I188252);
nor I_4648 (I82090,I82073,I188267);
nand I_4649 (I82107,I82090,I188264);
nor I_4650 (I82124,I82107,I82056);
DFFARX1 I_4651 (I82124,I3035,I81906,I81874,);
not I_4652 (I82155,I82107);
not I_4653 (I82172,I188267);
nand I_4654 (I82189,I82172,I188255);
nor I_4655 (I82206,I188267,I188243);
nand I_4656 (I81886,I82022,I82206);
nand I_4657 (I81880,I81971,I188267);
nand I_4658 (I82251,I82073,I188261);
DFFARX1 I_4659 (I82251,I3035,I81906,I81895,);
DFFARX1 I_4660 (I82251,I3035,I81906,I81889,);
not I_4661 (I82296,I188261);
nor I_4662 (I82313,I82296,I188249);
and I_4663 (I82330,I82313,I188270);
or I_4664 (I82347,I82330,I188246);
DFFARX1 I_4665 (I82347,I3035,I81906,I82373,);
nand I_4666 (I82381,I82373,I82039);
nor I_4667 (I81883,I82381,I82189);
nor I_4668 (I81877,I82373,I82005);
DFFARX1 I_4669 (I82373,I3035,I81906,I82435,);
not I_4670 (I82443,I82435);
nor I_4671 (I81892,I82443,I82155);
not I_4672 (I82501,I3042);
DFFARX1 I_4673 (I424022,I3035,I82501,I82527,);
DFFARX1 I_4674 (I82527,I3035,I82501,I82544,);
not I_4675 (I82493,I82544);
not I_4676 (I82566,I82527);
DFFARX1 I_4677 (I424016,I3035,I82501,I82592,);
not I_4678 (I82600,I82592);
and I_4679 (I82617,I82566,I424034);
not I_4680 (I82634,I424022);
nand I_4681 (I82651,I82634,I424034);
not I_4682 (I82668,I424016);
nor I_4683 (I82685,I82668,I424028);
nand I_4684 (I82702,I82685,I424019);
nor I_4685 (I82719,I82702,I82651);
DFFARX1 I_4686 (I82719,I3035,I82501,I82469,);
not I_4687 (I82750,I82702);
not I_4688 (I82767,I424028);
nand I_4689 (I82784,I82767,I424034);
nor I_4690 (I82801,I424028,I424022);
nand I_4691 (I82481,I82617,I82801);
nand I_4692 (I82475,I82566,I424028);
nand I_4693 (I82846,I82668,I424031);
DFFARX1 I_4694 (I82846,I3035,I82501,I82490,);
DFFARX1 I_4695 (I82846,I3035,I82501,I82484,);
not I_4696 (I82891,I424031);
nor I_4697 (I82908,I82891,I424037);
and I_4698 (I82925,I82908,I424019);
or I_4699 (I82942,I82925,I424025);
DFFARX1 I_4700 (I82942,I3035,I82501,I82968,);
nand I_4701 (I82976,I82968,I82634);
nor I_4702 (I82478,I82976,I82784);
nor I_4703 (I82472,I82968,I82600);
DFFARX1 I_4704 (I82968,I3035,I82501,I83030,);
not I_4705 (I83038,I83030);
nor I_4706 (I82487,I83038,I82750);
not I_4707 (I83096,I3042);
DFFARX1 I_4708 (I363168,I3035,I83096,I83122,);
DFFARX1 I_4709 (I83122,I3035,I83096,I83139,);
not I_4710 (I83088,I83139);
not I_4711 (I83161,I83122);
DFFARX1 I_4712 (I363165,I3035,I83096,I83187,);
not I_4713 (I83195,I83187);
and I_4714 (I83212,I83161,I363171);
not I_4715 (I83229,I363156);
nand I_4716 (I83246,I83229,I363171);
not I_4717 (I83263,I363159);
nor I_4718 (I83280,I83263,I363180);
nand I_4719 (I83297,I83280,I363177);
nor I_4720 (I83314,I83297,I83246);
DFFARX1 I_4721 (I83314,I3035,I83096,I83064,);
not I_4722 (I83345,I83297);
not I_4723 (I83362,I363180);
nand I_4724 (I83379,I83362,I363171);
nor I_4725 (I83396,I363180,I363156);
nand I_4726 (I83076,I83212,I83396);
nand I_4727 (I83070,I83161,I363180);
nand I_4728 (I83441,I83263,I363156);
DFFARX1 I_4729 (I83441,I3035,I83096,I83085,);
DFFARX1 I_4730 (I83441,I3035,I83096,I83079,);
not I_4731 (I83486,I363156);
nor I_4732 (I83503,I83486,I363162);
and I_4733 (I83520,I83503,I363174);
or I_4734 (I83537,I83520,I363159);
DFFARX1 I_4735 (I83537,I3035,I83096,I83563,);
nand I_4736 (I83571,I83563,I83229);
nor I_4737 (I83073,I83571,I83379);
nor I_4738 (I83067,I83563,I83195);
DFFARX1 I_4739 (I83563,I3035,I83096,I83625,);
not I_4740 (I83633,I83625);
nor I_4741 (I83082,I83633,I83345);
not I_4742 (I83691,I3042);
DFFARX1 I_4743 (I54190,I3035,I83691,I83717,);
DFFARX1 I_4744 (I83717,I3035,I83691,I83734,);
not I_4745 (I83683,I83734);
not I_4746 (I83756,I83717);
DFFARX1 I_4747 (I54184,I3035,I83691,I83782,);
not I_4748 (I83790,I83782);
and I_4749 (I83807,I83756,I54181);
not I_4750 (I83824,I54202);
nand I_4751 (I83841,I83824,I54181);
not I_4752 (I83858,I54196);
nor I_4753 (I83875,I83858,I54187);
nand I_4754 (I83892,I83875,I54193);
nor I_4755 (I83909,I83892,I83841);
DFFARX1 I_4756 (I83909,I3035,I83691,I83659,);
not I_4757 (I83940,I83892);
not I_4758 (I83957,I54187);
nand I_4759 (I83974,I83957,I54181);
nor I_4760 (I83991,I54187,I54202);
nand I_4761 (I83671,I83807,I83991);
nand I_4762 (I83665,I83756,I54187);
nand I_4763 (I84036,I83858,I54181);
DFFARX1 I_4764 (I84036,I3035,I83691,I83680,);
DFFARX1 I_4765 (I84036,I3035,I83691,I83674,);
not I_4766 (I84081,I54181);
nor I_4767 (I84098,I84081,I54199);
and I_4768 (I84115,I84098,I54205);
or I_4769 (I84132,I84115,I54184);
DFFARX1 I_4770 (I84132,I3035,I83691,I84158,);
nand I_4771 (I84166,I84158,I83824);
nor I_4772 (I83668,I84166,I83974);
nor I_4773 (I83662,I84158,I83790);
DFFARX1 I_4774 (I84158,I3035,I83691,I84220,);
not I_4775 (I84228,I84220);
nor I_4776 (I83677,I84228,I83940);
not I_4777 (I84286,I3042);
DFFARX1 I_4778 (I693323,I3035,I84286,I84312,);
DFFARX1 I_4779 (I84312,I3035,I84286,I84329,);
not I_4780 (I84278,I84329);
not I_4781 (I84351,I84312);
DFFARX1 I_4782 (I693296,I3035,I84286,I84377,);
not I_4783 (I84385,I84377);
and I_4784 (I84402,I84351,I693320);
not I_4785 (I84419,I693317);
nand I_4786 (I84436,I84419,I693320);
not I_4787 (I84453,I693296);
nor I_4788 (I84470,I84453,I693314);
nand I_4789 (I84487,I84470,I693302);
nor I_4790 (I84504,I84487,I84436);
DFFARX1 I_4791 (I84504,I3035,I84286,I84254,);
not I_4792 (I84535,I84487);
not I_4793 (I84552,I693314);
nand I_4794 (I84569,I84552,I693320);
nor I_4795 (I84586,I693314,I693317);
nand I_4796 (I84266,I84402,I84586);
nand I_4797 (I84260,I84351,I693314);
nand I_4798 (I84631,I84453,I693308);
DFFARX1 I_4799 (I84631,I3035,I84286,I84275,);
DFFARX1 I_4800 (I84631,I3035,I84286,I84269,);
not I_4801 (I84676,I693308);
nor I_4802 (I84693,I84676,I693311);
and I_4803 (I84710,I84693,I693299);
or I_4804 (I84727,I84710,I693305);
DFFARX1 I_4805 (I84727,I3035,I84286,I84753,);
nand I_4806 (I84761,I84753,I84419);
nor I_4807 (I84263,I84761,I84569);
nor I_4808 (I84257,I84753,I84385);
DFFARX1 I_4809 (I84753,I3035,I84286,I84815,);
not I_4810 (I84823,I84815);
nor I_4811 (I84272,I84823,I84535);
not I_4812 (I84881,I3042);
DFFARX1 I_4813 (I530995,I3035,I84881,I84907,);
DFFARX1 I_4814 (I84907,I3035,I84881,I84924,);
not I_4815 (I84873,I84924);
not I_4816 (I84946,I84907);
DFFARX1 I_4817 (I531004,I3035,I84881,I84972,);
not I_4818 (I84980,I84972);
and I_4819 (I84997,I84946,I530992);
not I_4820 (I85014,I530983);
nand I_4821 (I85031,I85014,I530992);
not I_4822 (I85048,I530989);
nor I_4823 (I85065,I85048,I531007);
nand I_4824 (I85082,I85065,I530980);
nor I_4825 (I85099,I85082,I85031);
DFFARX1 I_4826 (I85099,I3035,I84881,I84849,);
not I_4827 (I85130,I85082);
not I_4828 (I85147,I531007);
nand I_4829 (I85164,I85147,I530992);
nor I_4830 (I85181,I531007,I530983);
nand I_4831 (I84861,I84997,I85181);
nand I_4832 (I84855,I84946,I531007);
nand I_4833 (I85226,I85048,I530986);
DFFARX1 I_4834 (I85226,I3035,I84881,I84870,);
DFFARX1 I_4835 (I85226,I3035,I84881,I84864,);
not I_4836 (I85271,I530986);
nor I_4837 (I85288,I85271,I530998);
and I_4838 (I85305,I85288,I530980);
or I_4839 (I85322,I85305,I531001);
DFFARX1 I_4840 (I85322,I3035,I84881,I85348,);
nand I_4841 (I85356,I85348,I85014);
nor I_4842 (I84858,I85356,I85164);
nor I_4843 (I84852,I85348,I84980);
DFFARX1 I_4844 (I85348,I3035,I84881,I85410,);
not I_4845 (I85418,I85410);
nor I_4846 (I84867,I85418,I85130);
not I_4847 (I85476,I3042);
DFFARX1 I_4848 (I503217,I3035,I85476,I85502,);
DFFARX1 I_4849 (I85502,I3035,I85476,I85519,);
not I_4850 (I85468,I85519);
not I_4851 (I85541,I85502);
DFFARX1 I_4852 (I503226,I3035,I85476,I85567,);
not I_4853 (I85575,I85567);
and I_4854 (I85592,I85541,I503214);
not I_4855 (I85609,I503205);
nand I_4856 (I85626,I85609,I503214);
not I_4857 (I85643,I503211);
nor I_4858 (I85660,I85643,I503229);
nand I_4859 (I85677,I85660,I503202);
nor I_4860 (I85694,I85677,I85626);
DFFARX1 I_4861 (I85694,I3035,I85476,I85444,);
not I_4862 (I85725,I85677);
not I_4863 (I85742,I503229);
nand I_4864 (I85759,I85742,I503214);
nor I_4865 (I85776,I503229,I503205);
nand I_4866 (I85456,I85592,I85776);
nand I_4867 (I85450,I85541,I503229);
nand I_4868 (I85821,I85643,I503208);
DFFARX1 I_4869 (I85821,I3035,I85476,I85465,);
DFFARX1 I_4870 (I85821,I3035,I85476,I85459,);
not I_4871 (I85866,I503208);
nor I_4872 (I85883,I85866,I503220);
and I_4873 (I85900,I85883,I503202);
or I_4874 (I85917,I85900,I503223);
DFFARX1 I_4875 (I85917,I3035,I85476,I85943,);
nand I_4876 (I85951,I85943,I85609);
nor I_4877 (I85453,I85951,I85759);
nor I_4878 (I85447,I85943,I85575);
DFFARX1 I_4879 (I85943,I3035,I85476,I86005,);
not I_4880 (I86013,I86005);
nor I_4881 (I85462,I86013,I85725);
not I_4882 (I86071,I3042);
DFFARX1 I_4883 (I325023,I3035,I86071,I86097,);
DFFARX1 I_4884 (I86097,I3035,I86071,I86114,);
not I_4885 (I86063,I86114);
not I_4886 (I86136,I86097);
DFFARX1 I_4887 (I325014,I3035,I86071,I86162,);
not I_4888 (I86170,I86162);
and I_4889 (I86187,I86136,I325032);
not I_4890 (I86204,I325029);
nand I_4891 (I86221,I86204,I325032);
not I_4892 (I86238,I325008);
nor I_4893 (I86255,I86238,I325011);
nand I_4894 (I86272,I86255,I325020);
nor I_4895 (I86289,I86272,I86221);
DFFARX1 I_4896 (I86289,I3035,I86071,I86039,);
not I_4897 (I86320,I86272);
not I_4898 (I86337,I325011);
nand I_4899 (I86354,I86337,I325032);
nor I_4900 (I86371,I325011,I325029);
nand I_4901 (I86051,I86187,I86371);
nand I_4902 (I86045,I86136,I325011);
nand I_4903 (I86416,I86238,I325026);
DFFARX1 I_4904 (I86416,I3035,I86071,I86060,);
DFFARX1 I_4905 (I86416,I3035,I86071,I86054,);
not I_4906 (I86461,I325026);
nor I_4907 (I86478,I86461,I325008);
and I_4908 (I86495,I86478,I325017);
or I_4909 (I86512,I86495,I325011);
DFFARX1 I_4910 (I86512,I3035,I86071,I86538,);
nand I_4911 (I86546,I86538,I86204);
nor I_4912 (I86048,I86546,I86354);
nor I_4913 (I86042,I86538,I86170);
DFFARX1 I_4914 (I86538,I3035,I86071,I86600,);
not I_4915 (I86608,I86600);
nor I_4916 (I86057,I86608,I86320);
not I_4917 (I86666,I3042);
DFFARX1 I_4918 (I632402,I3035,I86666,I86692,);
DFFARX1 I_4919 (I86692,I3035,I86666,I86709,);
not I_4920 (I86658,I86709);
not I_4921 (I86731,I86692);
DFFARX1 I_4922 (I632402,I3035,I86666,I86757,);
not I_4923 (I86765,I86757);
and I_4924 (I86782,I86731,I632405);
not I_4925 (I86799,I632417);
nand I_4926 (I86816,I86799,I632405);
not I_4927 (I86833,I632423);
nor I_4928 (I86850,I86833,I632414);
nand I_4929 (I86867,I86850,I632420);
nor I_4930 (I86884,I86867,I86816);
DFFARX1 I_4931 (I86884,I3035,I86666,I86634,);
not I_4932 (I86915,I86867);
not I_4933 (I86932,I632414);
nand I_4934 (I86949,I86932,I632405);
nor I_4935 (I86966,I632414,I632417);
nand I_4936 (I86646,I86782,I86966);
nand I_4937 (I86640,I86731,I632414);
nand I_4938 (I87011,I86833,I632411);
DFFARX1 I_4939 (I87011,I3035,I86666,I86655,);
DFFARX1 I_4940 (I87011,I3035,I86666,I86649,);
not I_4941 (I87056,I632411);
nor I_4942 (I87073,I87056,I632408);
and I_4943 (I87090,I87073,I632426);
or I_4944 (I87107,I87090,I632405);
DFFARX1 I_4945 (I87107,I3035,I86666,I87133,);
nand I_4946 (I87141,I87133,I86799);
nor I_4947 (I86643,I87141,I86949);
nor I_4948 (I86637,I87133,I86765);
DFFARX1 I_4949 (I87133,I3035,I86666,I87195,);
not I_4950 (I87203,I87195);
nor I_4951 (I86652,I87203,I86915);
not I_4952 (I87261,I3042);
DFFARX1 I_4953 (I155042,I3035,I87261,I87287,);
DFFARX1 I_4954 (I87287,I3035,I87261,I87304,);
not I_4955 (I87253,I87304);
not I_4956 (I87326,I87287);
DFFARX1 I_4957 (I155057,I3035,I87261,I87352,);
not I_4958 (I87360,I87352);
and I_4959 (I87377,I87326,I155054);
not I_4960 (I87394,I155042);
nand I_4961 (I87411,I87394,I155054);
not I_4962 (I87428,I155051);
nor I_4963 (I87445,I87428,I155066);
nand I_4964 (I87462,I87445,I155063);
nor I_4965 (I87479,I87462,I87411);
DFFARX1 I_4966 (I87479,I3035,I87261,I87229,);
not I_4967 (I87510,I87462);
not I_4968 (I87527,I155066);
nand I_4969 (I87544,I87527,I155054);
nor I_4970 (I87561,I155066,I155042);
nand I_4971 (I87241,I87377,I87561);
nand I_4972 (I87235,I87326,I155066);
nand I_4973 (I87606,I87428,I155060);
DFFARX1 I_4974 (I87606,I3035,I87261,I87250,);
DFFARX1 I_4975 (I87606,I3035,I87261,I87244,);
not I_4976 (I87651,I155060);
nor I_4977 (I87668,I87651,I155048);
and I_4978 (I87685,I87668,I155069);
or I_4979 (I87702,I87685,I155045);
DFFARX1 I_4980 (I87702,I3035,I87261,I87728,);
nand I_4981 (I87736,I87728,I87394);
nor I_4982 (I87238,I87736,I87544);
nor I_4983 (I87232,I87728,I87360);
DFFARX1 I_4984 (I87728,I3035,I87261,I87790,);
not I_4985 (I87798,I87790);
nor I_4986 (I87247,I87798,I87510);
not I_4987 (I87856,I3042);
DFFARX1 I_4988 (I728184,I3035,I87856,I87882,);
DFFARX1 I_4989 (I87882,I3035,I87856,I87899,);
not I_4990 (I87848,I87899);
not I_4991 (I87921,I87882);
DFFARX1 I_4992 (I728175,I3035,I87856,I87947,);
not I_4993 (I87955,I87947);
and I_4994 (I87972,I87921,I728169);
not I_4995 (I87989,I728163);
nand I_4996 (I88006,I87989,I728169);
not I_4997 (I88023,I728190);
nor I_4998 (I88040,I88023,I728163);
nand I_4999 (I88057,I88040,I728187);
nor I_5000 (I88074,I88057,I88006);
DFFARX1 I_5001 (I88074,I3035,I87856,I87824,);
not I_5002 (I88105,I88057);
not I_5003 (I88122,I728163);
nand I_5004 (I88139,I88122,I728169);
nor I_5005 (I88156,I728163,I728163);
nand I_5006 (I87836,I87972,I88156);
nand I_5007 (I87830,I87921,I728163);
nand I_5008 (I88201,I88023,I728172);
DFFARX1 I_5009 (I88201,I3035,I87856,I87845,);
DFFARX1 I_5010 (I88201,I3035,I87856,I87839,);
not I_5011 (I88246,I728172);
nor I_5012 (I88263,I88246,I728178);
and I_5013 (I88280,I88263,I728181);
or I_5014 (I88297,I88280,I728166);
DFFARX1 I_5015 (I88297,I3035,I87856,I88323,);
nand I_5016 (I88331,I88323,I87989);
nor I_5017 (I87833,I88331,I88139);
nor I_5018 (I87827,I88323,I87955);
DFFARX1 I_5019 (I88323,I3035,I87856,I88385,);
not I_5020 (I88393,I88385);
nor I_5021 (I87842,I88393,I88105);
not I_5022 (I88451,I3042);
DFFARX1 I_5023 (I2220,I3035,I88451,I88477,);
DFFARX1 I_5024 (I88477,I3035,I88451,I88494,);
not I_5025 (I88443,I88494);
not I_5026 (I88516,I88477);
DFFARX1 I_5027 (I1732,I3035,I88451,I88542,);
not I_5028 (I88550,I88542);
and I_5029 (I88567,I88516,I2420);
not I_5030 (I88584,I2148);
nand I_5031 (I88601,I88584,I2420);
not I_5032 (I88618,I3028);
nor I_5033 (I88635,I88618,I2596);
nand I_5034 (I88652,I88635,I2084);
nor I_5035 (I88669,I88652,I88601);
DFFARX1 I_5036 (I88669,I3035,I88451,I88419,);
not I_5037 (I88700,I88652);
not I_5038 (I88717,I2596);
nand I_5039 (I88734,I88717,I2420);
nor I_5040 (I88751,I2596,I2148);
nand I_5041 (I88431,I88567,I88751);
nand I_5042 (I88425,I88516,I2596);
nand I_5043 (I88796,I88618,I2732);
DFFARX1 I_5044 (I88796,I3035,I88451,I88440,);
DFFARX1 I_5045 (I88796,I3035,I88451,I88434,);
not I_5046 (I88841,I2732);
nor I_5047 (I88858,I88841,I2780);
and I_5048 (I88875,I88858,I2364);
or I_5049 (I88892,I88875,I1492);
DFFARX1 I_5050 (I88892,I3035,I88451,I88918,);
nand I_5051 (I88926,I88918,I88584);
nor I_5052 (I88428,I88926,I88734);
nor I_5053 (I88422,I88918,I88550);
DFFARX1 I_5054 (I88918,I3035,I88451,I88980,);
not I_5055 (I88988,I88980);
nor I_5056 (I88437,I88988,I88700);
not I_5057 (I89046,I3042);
DFFARX1 I_5058 (I49447,I3035,I89046,I89072,);
DFFARX1 I_5059 (I89072,I3035,I89046,I89089,);
not I_5060 (I89038,I89089);
not I_5061 (I89111,I89072);
DFFARX1 I_5062 (I49441,I3035,I89046,I89137,);
not I_5063 (I89145,I89137);
and I_5064 (I89162,I89111,I49438);
not I_5065 (I89179,I49459);
nand I_5066 (I89196,I89179,I49438);
not I_5067 (I89213,I49453);
nor I_5068 (I89230,I89213,I49444);
nand I_5069 (I89247,I89230,I49450);
nor I_5070 (I89264,I89247,I89196);
DFFARX1 I_5071 (I89264,I3035,I89046,I89014,);
not I_5072 (I89295,I89247);
not I_5073 (I89312,I49444);
nand I_5074 (I89329,I89312,I49438);
nor I_5075 (I89346,I49444,I49459);
nand I_5076 (I89026,I89162,I89346);
nand I_5077 (I89020,I89111,I49444);
nand I_5078 (I89391,I89213,I49438);
DFFARX1 I_5079 (I89391,I3035,I89046,I89035,);
DFFARX1 I_5080 (I89391,I3035,I89046,I89029,);
not I_5081 (I89436,I49438);
nor I_5082 (I89453,I89436,I49456);
and I_5083 (I89470,I89453,I49462);
or I_5084 (I89487,I89470,I49441);
DFFARX1 I_5085 (I89487,I3035,I89046,I89513,);
nand I_5086 (I89521,I89513,I89179);
nor I_5087 (I89023,I89521,I89329);
nor I_5088 (I89017,I89513,I89145);
DFFARX1 I_5089 (I89513,I3035,I89046,I89575,);
not I_5090 (I89583,I89575);
nor I_5091 (I89032,I89583,I89295);
not I_5092 (I89641,I3042);
DFFARX1 I_5093 (I709739,I3035,I89641,I89667,);
DFFARX1 I_5094 (I89667,I3035,I89641,I89684,);
not I_5095 (I89633,I89684);
not I_5096 (I89706,I89667);
DFFARX1 I_5097 (I709730,I3035,I89641,I89732,);
not I_5098 (I89740,I89732);
and I_5099 (I89757,I89706,I709724);
not I_5100 (I89774,I709718);
nand I_5101 (I89791,I89774,I709724);
not I_5102 (I89808,I709745);
nor I_5103 (I89825,I89808,I709718);
nand I_5104 (I89842,I89825,I709742);
nor I_5105 (I89859,I89842,I89791);
DFFARX1 I_5106 (I89859,I3035,I89641,I89609,);
not I_5107 (I89890,I89842);
not I_5108 (I89907,I709718);
nand I_5109 (I89924,I89907,I709724);
nor I_5110 (I89941,I709718,I709718);
nand I_5111 (I89621,I89757,I89941);
nand I_5112 (I89615,I89706,I709718);
nand I_5113 (I89986,I89808,I709727);
DFFARX1 I_5114 (I89986,I3035,I89641,I89630,);
DFFARX1 I_5115 (I89986,I3035,I89641,I89624,);
not I_5116 (I90031,I709727);
nor I_5117 (I90048,I90031,I709733);
and I_5118 (I90065,I90048,I709736);
or I_5119 (I90082,I90065,I709721);
DFFARX1 I_5120 (I90082,I3035,I89641,I90108,);
nand I_5121 (I90116,I90108,I89774);
nor I_5122 (I89618,I90116,I89924);
nor I_5123 (I89612,I90108,I89740);
DFFARX1 I_5124 (I90108,I3035,I89641,I90170,);
not I_5125 (I90178,I90170);
nor I_5126 (I89627,I90178,I89890);
not I_5127 (I90236,I3042);
DFFARX1 I_5128 (I744249,I3035,I90236,I90262,);
DFFARX1 I_5129 (I90262,I3035,I90236,I90279,);
not I_5130 (I90228,I90279);
not I_5131 (I90301,I90262);
DFFARX1 I_5132 (I744240,I3035,I90236,I90327,);
not I_5133 (I90335,I90327);
and I_5134 (I90352,I90301,I744234);
not I_5135 (I90369,I744228);
nand I_5136 (I90386,I90369,I744234);
not I_5137 (I90403,I744255);
nor I_5138 (I90420,I90403,I744228);
nand I_5139 (I90437,I90420,I744252);
nor I_5140 (I90454,I90437,I90386);
DFFARX1 I_5141 (I90454,I3035,I90236,I90204,);
not I_5142 (I90485,I90437);
not I_5143 (I90502,I744228);
nand I_5144 (I90519,I90502,I744234);
nor I_5145 (I90536,I744228,I744228);
nand I_5146 (I90216,I90352,I90536);
nand I_5147 (I90210,I90301,I744228);
nand I_5148 (I90581,I90403,I744237);
DFFARX1 I_5149 (I90581,I3035,I90236,I90225,);
DFFARX1 I_5150 (I90581,I3035,I90236,I90219,);
not I_5151 (I90626,I744237);
nor I_5152 (I90643,I90626,I744243);
and I_5153 (I90660,I90643,I744246);
or I_5154 (I90677,I90660,I744231);
DFFARX1 I_5155 (I90677,I3035,I90236,I90703,);
nand I_5156 (I90711,I90703,I90369);
nor I_5157 (I90213,I90711,I90519);
nor I_5158 (I90207,I90703,I90335);
DFFARX1 I_5159 (I90703,I3035,I90236,I90765,);
not I_5160 (I90773,I90765);
nor I_5161 (I90222,I90773,I90485);
not I_5162 (I90831,I3042);
DFFARX1 I_5163 (I499987,I3035,I90831,I90857,);
DFFARX1 I_5164 (I90857,I3035,I90831,I90874,);
not I_5165 (I90823,I90874);
not I_5166 (I90896,I90857);
DFFARX1 I_5167 (I499996,I3035,I90831,I90922,);
not I_5168 (I90930,I90922);
and I_5169 (I90947,I90896,I499984);
not I_5170 (I90964,I499975);
nand I_5171 (I90981,I90964,I499984);
not I_5172 (I90998,I499981);
nor I_5173 (I91015,I90998,I499999);
nand I_5174 (I91032,I91015,I499972);
nor I_5175 (I91049,I91032,I90981);
DFFARX1 I_5176 (I91049,I3035,I90831,I90799,);
not I_5177 (I91080,I91032);
not I_5178 (I91097,I499999);
nand I_5179 (I91114,I91097,I499984);
nor I_5180 (I91131,I499999,I499975);
nand I_5181 (I90811,I90947,I91131);
nand I_5182 (I90805,I90896,I499999);
nand I_5183 (I91176,I90998,I499978);
DFFARX1 I_5184 (I91176,I3035,I90831,I90820,);
DFFARX1 I_5185 (I91176,I3035,I90831,I90814,);
not I_5186 (I91221,I499978);
nor I_5187 (I91238,I91221,I499990);
and I_5188 (I91255,I91238,I499972);
or I_5189 (I91272,I91255,I499993);
DFFARX1 I_5190 (I91272,I3035,I90831,I91298,);
nand I_5191 (I91306,I91298,I90964);
nor I_5192 (I90808,I91306,I91114);
nor I_5193 (I90802,I91298,I90930);
DFFARX1 I_5194 (I91298,I3035,I90831,I91360,);
not I_5195 (I91368,I91360);
nor I_5196 (I90817,I91368,I91080);
not I_5197 (I91426,I3042);
DFFARX1 I_5198 (I675959,I3035,I91426,I91452,);
DFFARX1 I_5199 (I91452,I3035,I91426,I91469,);
not I_5200 (I91418,I91469);
not I_5201 (I91491,I91452);
DFFARX1 I_5202 (I675971,I3035,I91426,I91517,);
not I_5203 (I91525,I91517);
and I_5204 (I91542,I91491,I675965);
not I_5205 (I91559,I675977);
nand I_5206 (I91576,I91559,I675965);
not I_5207 (I91593,I675962);
nor I_5208 (I91610,I91593,I675974);
nand I_5209 (I91627,I91610,I675956);
nor I_5210 (I91644,I91627,I91576);
DFFARX1 I_5211 (I91644,I3035,I91426,I91394,);
not I_5212 (I91675,I91627);
not I_5213 (I91692,I675974);
nand I_5214 (I91709,I91692,I675965);
nor I_5215 (I91726,I675974,I675977);
nand I_5216 (I91406,I91542,I91726);
nand I_5217 (I91400,I91491,I675974);
nand I_5218 (I91771,I91593,I675968);
DFFARX1 I_5219 (I91771,I3035,I91426,I91415,);
DFFARX1 I_5220 (I91771,I3035,I91426,I91409,);
not I_5221 (I91816,I675968);
nor I_5222 (I91833,I91816,I675959);
and I_5223 (I91850,I91833,I675956);
or I_5224 (I91867,I91850,I675980);
DFFARX1 I_5225 (I91867,I3035,I91426,I91893,);
nand I_5226 (I91901,I91893,I91559);
nor I_5227 (I91403,I91901,I91709);
nor I_5228 (I91397,I91893,I91525);
DFFARX1 I_5229 (I91893,I3035,I91426,I91955,);
not I_5230 (I91963,I91955);
nor I_5231 (I91412,I91963,I91675);
not I_5232 (I92021,I3042);
DFFARX1 I_5233 (I30475,I3035,I92021,I92047,);
DFFARX1 I_5234 (I92047,I3035,I92021,I92064,);
not I_5235 (I92013,I92064);
not I_5236 (I92086,I92047);
DFFARX1 I_5237 (I30469,I3035,I92021,I92112,);
not I_5238 (I92120,I92112);
and I_5239 (I92137,I92086,I30466);
not I_5240 (I92154,I30487);
nand I_5241 (I92171,I92154,I30466);
not I_5242 (I92188,I30481);
nor I_5243 (I92205,I92188,I30472);
nand I_5244 (I92222,I92205,I30478);
nor I_5245 (I92239,I92222,I92171);
DFFARX1 I_5246 (I92239,I3035,I92021,I91989,);
not I_5247 (I92270,I92222);
not I_5248 (I92287,I30472);
nand I_5249 (I92304,I92287,I30466);
nor I_5250 (I92321,I30472,I30487);
nand I_5251 (I92001,I92137,I92321);
nand I_5252 (I91995,I92086,I30472);
nand I_5253 (I92366,I92188,I30466);
DFFARX1 I_5254 (I92366,I3035,I92021,I92010,);
DFFARX1 I_5255 (I92366,I3035,I92021,I92004,);
not I_5256 (I92411,I30466);
nor I_5257 (I92428,I92411,I30484);
and I_5258 (I92445,I92428,I30490);
or I_5259 (I92462,I92445,I30469);
DFFARX1 I_5260 (I92462,I3035,I92021,I92488,);
nand I_5261 (I92496,I92488,I92154);
nor I_5262 (I91998,I92496,I92304);
nor I_5263 (I91992,I92488,I92120);
DFFARX1 I_5264 (I92488,I3035,I92021,I92550,);
not I_5265 (I92558,I92550);
nor I_5266 (I92007,I92558,I92270);
not I_5267 (I92616,I3042);
DFFARX1 I_5268 (I479961,I3035,I92616,I92642,);
DFFARX1 I_5269 (I92642,I3035,I92616,I92659,);
not I_5270 (I92608,I92659);
not I_5271 (I92681,I92642);
DFFARX1 I_5272 (I479970,I3035,I92616,I92707,);
not I_5273 (I92715,I92707);
and I_5274 (I92732,I92681,I479958);
not I_5275 (I92749,I479949);
nand I_5276 (I92766,I92749,I479958);
not I_5277 (I92783,I479955);
nor I_5278 (I92800,I92783,I479973);
nand I_5279 (I92817,I92800,I479946);
nor I_5280 (I92834,I92817,I92766);
DFFARX1 I_5281 (I92834,I3035,I92616,I92584,);
not I_5282 (I92865,I92817);
not I_5283 (I92882,I479973);
nand I_5284 (I92899,I92882,I479958);
nor I_5285 (I92916,I479973,I479949);
nand I_5286 (I92596,I92732,I92916);
nand I_5287 (I92590,I92681,I479973);
nand I_5288 (I92961,I92783,I479952);
DFFARX1 I_5289 (I92961,I3035,I92616,I92605,);
DFFARX1 I_5290 (I92961,I3035,I92616,I92599,);
not I_5291 (I93006,I479952);
nor I_5292 (I93023,I93006,I479964);
and I_5293 (I93040,I93023,I479946);
or I_5294 (I93057,I93040,I479967);
DFFARX1 I_5295 (I93057,I3035,I92616,I93083,);
nand I_5296 (I93091,I93083,I92749);
nor I_5297 (I92593,I93091,I92899);
nor I_5298 (I92587,I93083,I92715);
DFFARX1 I_5299 (I93083,I3035,I92616,I93145,);
not I_5300 (I93153,I93145);
nor I_5301 (I92602,I93153,I92865);
not I_5302 (I93211,I3042);
DFFARX1 I_5303 (I547609,I3035,I93211,I93237,);
DFFARX1 I_5304 (I93237,I3035,I93211,I93254,);
not I_5305 (I93203,I93254);
not I_5306 (I93276,I93237);
DFFARX1 I_5307 (I547618,I3035,I93211,I93302,);
not I_5308 (I93310,I93302);
and I_5309 (I93327,I93276,I547612);
not I_5310 (I93344,I547606);
nand I_5311 (I93361,I93344,I547612);
not I_5312 (I93378,I547621);
nor I_5313 (I93395,I93378,I547609);
nand I_5314 (I93412,I93395,I547615);
nor I_5315 (I93429,I93412,I93361);
DFFARX1 I_5316 (I93429,I3035,I93211,I93179,);
not I_5317 (I93460,I93412);
not I_5318 (I93477,I547609);
nand I_5319 (I93494,I93477,I547612);
nor I_5320 (I93511,I547609,I547606);
nand I_5321 (I93191,I93327,I93511);
nand I_5322 (I93185,I93276,I547609);
nand I_5323 (I93556,I93378,I547612);
DFFARX1 I_5324 (I93556,I3035,I93211,I93200,);
DFFARX1 I_5325 (I93556,I3035,I93211,I93194,);
not I_5326 (I93601,I547612);
nor I_5327 (I93618,I93601,I547627);
and I_5328 (I93635,I93618,I547624);
or I_5329 (I93652,I93635,I547606);
DFFARX1 I_5330 (I93652,I3035,I93211,I93678,);
nand I_5331 (I93686,I93678,I93344);
nor I_5332 (I93188,I93686,I93494);
nor I_5333 (I93182,I93678,I93310);
DFFARX1 I_5334 (I93678,I3035,I93211,I93740,);
not I_5335 (I93748,I93740);
nor I_5336 (I93197,I93748,I93460);
not I_5337 (I93806,I3042);
DFFARX1 I_5338 (I334849,I3035,I93806,I93832,);
DFFARX1 I_5339 (I93832,I3035,I93806,I93849,);
not I_5340 (I93798,I93849);
not I_5341 (I93871,I93832);
DFFARX1 I_5342 (I334840,I3035,I93806,I93897,);
not I_5343 (I93905,I93897);
and I_5344 (I93922,I93871,I334858);
not I_5345 (I93939,I334855);
nand I_5346 (I93956,I93939,I334858);
not I_5347 (I93973,I334834);
nor I_5348 (I93990,I93973,I334837);
nand I_5349 (I94007,I93990,I334846);
nor I_5350 (I94024,I94007,I93956);
DFFARX1 I_5351 (I94024,I3035,I93806,I93774,);
not I_5352 (I94055,I94007);
not I_5353 (I94072,I334837);
nand I_5354 (I94089,I94072,I334858);
nor I_5355 (I94106,I334837,I334855);
nand I_5356 (I93786,I93922,I94106);
nand I_5357 (I93780,I93871,I334837);
nand I_5358 (I94151,I93973,I334852);
DFFARX1 I_5359 (I94151,I3035,I93806,I93795,);
DFFARX1 I_5360 (I94151,I3035,I93806,I93789,);
not I_5361 (I94196,I334852);
nor I_5362 (I94213,I94196,I334834);
and I_5363 (I94230,I94213,I334843);
or I_5364 (I94247,I94230,I334837);
DFFARX1 I_5365 (I94247,I3035,I93806,I94273,);
nand I_5366 (I94281,I94273,I93939);
nor I_5367 (I93783,I94281,I94089);
nor I_5368 (I93777,I94273,I93905);
DFFARX1 I_5369 (I94273,I3035,I93806,I94335,);
not I_5370 (I94343,I94335);
nor I_5371 (I93792,I94343,I94055);
not I_5372 (I94401,I3042);
DFFARX1 I_5373 (I357966,I3035,I94401,I94427,);
DFFARX1 I_5374 (I94427,I3035,I94401,I94444,);
not I_5375 (I94393,I94444);
not I_5376 (I94466,I94427);
DFFARX1 I_5377 (I357963,I3035,I94401,I94492,);
not I_5378 (I94500,I94492);
and I_5379 (I94517,I94466,I357969);
not I_5380 (I94534,I357954);
nand I_5381 (I94551,I94534,I357969);
not I_5382 (I94568,I357957);
nor I_5383 (I94585,I94568,I357978);
nand I_5384 (I94602,I94585,I357975);
nor I_5385 (I94619,I94602,I94551);
DFFARX1 I_5386 (I94619,I3035,I94401,I94369,);
not I_5387 (I94650,I94602);
not I_5388 (I94667,I357978);
nand I_5389 (I94684,I94667,I357969);
nor I_5390 (I94701,I357978,I357954);
nand I_5391 (I94381,I94517,I94701);
nand I_5392 (I94375,I94466,I357978);
nand I_5393 (I94746,I94568,I357954);
DFFARX1 I_5394 (I94746,I3035,I94401,I94390,);
DFFARX1 I_5395 (I94746,I3035,I94401,I94384,);
not I_5396 (I94791,I357954);
nor I_5397 (I94808,I94791,I357960);
and I_5398 (I94825,I94808,I357972);
or I_5399 (I94842,I94825,I357957);
DFFARX1 I_5400 (I94842,I3035,I94401,I94868,);
nand I_5401 (I94876,I94868,I94534);
nor I_5402 (I94378,I94876,I94684);
nor I_5403 (I94372,I94868,I94500);
DFFARX1 I_5404 (I94868,I3035,I94401,I94930,);
not I_5405 (I94938,I94930);
nor I_5406 (I94387,I94938,I94650);
not I_5407 (I94996,I3042);
DFFARX1 I_5408 (I219336,I3035,I94996,I95022,);
DFFARX1 I_5409 (I95022,I3035,I94996,I95039,);
not I_5410 (I94988,I95039);
not I_5411 (I95061,I95022);
DFFARX1 I_5412 (I219351,I3035,I94996,I95087,);
not I_5413 (I95095,I95087);
and I_5414 (I95112,I95061,I219348);
not I_5415 (I95129,I219336);
nand I_5416 (I95146,I95129,I219348);
not I_5417 (I95163,I219345);
nor I_5418 (I95180,I95163,I219360);
nand I_5419 (I95197,I95180,I219357);
nor I_5420 (I95214,I95197,I95146);
DFFARX1 I_5421 (I95214,I3035,I94996,I94964,);
not I_5422 (I95245,I95197);
not I_5423 (I95262,I219360);
nand I_5424 (I95279,I95262,I219348);
nor I_5425 (I95296,I219360,I219336);
nand I_5426 (I94976,I95112,I95296);
nand I_5427 (I94970,I95061,I219360);
nand I_5428 (I95341,I95163,I219354);
DFFARX1 I_5429 (I95341,I3035,I94996,I94985,);
DFFARX1 I_5430 (I95341,I3035,I94996,I94979,);
not I_5431 (I95386,I219354);
nor I_5432 (I95403,I95386,I219342);
and I_5433 (I95420,I95403,I219363);
or I_5434 (I95437,I95420,I219339);
DFFARX1 I_5435 (I95437,I3035,I94996,I95463,);
nand I_5436 (I95471,I95463,I95129);
nor I_5437 (I94973,I95471,I95279);
nor I_5438 (I94967,I95463,I95095);
DFFARX1 I_5439 (I95463,I3035,I94996,I95525,);
not I_5440 (I95533,I95525);
nor I_5441 (I94982,I95533,I95245);
not I_5442 (I95591,I3042);
DFFARX1 I_5443 (I722234,I3035,I95591,I95617,);
DFFARX1 I_5444 (I95617,I3035,I95591,I95634,);
not I_5445 (I95583,I95634);
not I_5446 (I95656,I95617);
DFFARX1 I_5447 (I722225,I3035,I95591,I95682,);
not I_5448 (I95690,I95682);
and I_5449 (I95707,I95656,I722219);
not I_5450 (I95724,I722213);
nand I_5451 (I95741,I95724,I722219);
not I_5452 (I95758,I722240);
nor I_5453 (I95775,I95758,I722213);
nand I_5454 (I95792,I95775,I722237);
nor I_5455 (I95809,I95792,I95741);
DFFARX1 I_5456 (I95809,I3035,I95591,I95559,);
not I_5457 (I95840,I95792);
not I_5458 (I95857,I722213);
nand I_5459 (I95874,I95857,I722219);
nor I_5460 (I95891,I722213,I722213);
nand I_5461 (I95571,I95707,I95891);
nand I_5462 (I95565,I95656,I722213);
nand I_5463 (I95936,I95758,I722222);
DFFARX1 I_5464 (I95936,I3035,I95591,I95580,);
DFFARX1 I_5465 (I95936,I3035,I95591,I95574,);
not I_5466 (I95981,I722222);
nor I_5467 (I95998,I95981,I722228);
and I_5468 (I96015,I95998,I722231);
or I_5469 (I96032,I96015,I722216);
DFFARX1 I_5470 (I96032,I3035,I95591,I96058,);
nand I_5471 (I96066,I96058,I95724);
nor I_5472 (I95568,I96066,I95874);
nor I_5473 (I95562,I96058,I95690);
DFFARX1 I_5474 (I96058,I3035,I95591,I96120,);
not I_5475 (I96128,I96120);
nor I_5476 (I95577,I96128,I95840);
not I_5477 (I96186,I3042);
DFFARX1 I_5478 (I161893,I3035,I96186,I96212,);
DFFARX1 I_5479 (I96212,I3035,I96186,I96229,);
not I_5480 (I96178,I96229);
not I_5481 (I96251,I96212);
DFFARX1 I_5482 (I161908,I3035,I96186,I96277,);
not I_5483 (I96285,I96277);
and I_5484 (I96302,I96251,I161905);
not I_5485 (I96319,I161893);
nand I_5486 (I96336,I96319,I161905);
not I_5487 (I96353,I161902);
nor I_5488 (I96370,I96353,I161917);
nand I_5489 (I96387,I96370,I161914);
nor I_5490 (I96404,I96387,I96336);
DFFARX1 I_5491 (I96404,I3035,I96186,I96154,);
not I_5492 (I96435,I96387);
not I_5493 (I96452,I161917);
nand I_5494 (I96469,I96452,I161905);
nor I_5495 (I96486,I161917,I161893);
nand I_5496 (I96166,I96302,I96486);
nand I_5497 (I96160,I96251,I161917);
nand I_5498 (I96531,I96353,I161911);
DFFARX1 I_5499 (I96531,I3035,I96186,I96175,);
DFFARX1 I_5500 (I96531,I3035,I96186,I96169,);
not I_5501 (I96576,I161911);
nor I_5502 (I96593,I96576,I161899);
and I_5503 (I96610,I96593,I161920);
or I_5504 (I96627,I96610,I161896);
DFFARX1 I_5505 (I96627,I3035,I96186,I96653,);
nand I_5506 (I96661,I96653,I96319);
nor I_5507 (I96163,I96661,I96469);
nor I_5508 (I96157,I96653,I96285);
DFFARX1 I_5509 (I96653,I3035,I96186,I96715,);
not I_5510 (I96723,I96715);
nor I_5511 (I96172,I96723,I96435);
not I_5512 (I96781,I3042);
DFFARX1 I_5513 (I162947,I3035,I96781,I96807,);
DFFARX1 I_5514 (I96807,I3035,I96781,I96824,);
not I_5515 (I96773,I96824);
not I_5516 (I96846,I96807);
DFFARX1 I_5517 (I162962,I3035,I96781,I96872,);
not I_5518 (I96880,I96872);
and I_5519 (I96897,I96846,I162959);
not I_5520 (I96914,I162947);
nand I_5521 (I96931,I96914,I162959);
not I_5522 (I96948,I162956);
nor I_5523 (I96965,I96948,I162971);
nand I_5524 (I96982,I96965,I162968);
nor I_5525 (I96999,I96982,I96931);
DFFARX1 I_5526 (I96999,I3035,I96781,I96749,);
not I_5527 (I97030,I96982);
not I_5528 (I97047,I162971);
nand I_5529 (I97064,I97047,I162959);
nor I_5530 (I97081,I162971,I162947);
nand I_5531 (I96761,I96897,I97081);
nand I_5532 (I96755,I96846,I162971);
nand I_5533 (I97126,I96948,I162965);
DFFARX1 I_5534 (I97126,I3035,I96781,I96770,);
DFFARX1 I_5535 (I97126,I3035,I96781,I96764,);
not I_5536 (I97171,I162965);
nor I_5537 (I97188,I97171,I162953);
and I_5538 (I97205,I97188,I162974);
or I_5539 (I97222,I97205,I162950);
DFFARX1 I_5540 (I97222,I3035,I96781,I97248,);
nand I_5541 (I97256,I97248,I96914);
nor I_5542 (I96758,I97256,I97064);
nor I_5543 (I96752,I97248,I96880);
DFFARX1 I_5544 (I97248,I3035,I96781,I97310,);
not I_5545 (I97318,I97310);
nor I_5546 (I96767,I97318,I97030);
not I_5547 (I97376,I3042);
DFFARX1 I_5548 (I666488,I3035,I97376,I97402,);
DFFARX1 I_5549 (I97402,I3035,I97376,I97419,);
not I_5550 (I97368,I97419);
not I_5551 (I97441,I97402);
DFFARX1 I_5552 (I666473,I3035,I97376,I97467,);
not I_5553 (I97475,I97467);
and I_5554 (I97492,I97441,I666491);
not I_5555 (I97509,I666473);
nand I_5556 (I97526,I97509,I666491);
not I_5557 (I97543,I666494);
nor I_5558 (I97560,I97543,I666485);
nand I_5559 (I97577,I97560,I666482);
nor I_5560 (I97594,I97577,I97526);
DFFARX1 I_5561 (I97594,I3035,I97376,I97344,);
not I_5562 (I97625,I97577);
not I_5563 (I97642,I666485);
nand I_5564 (I97659,I97642,I666491);
nor I_5565 (I97676,I666485,I666473);
nand I_5566 (I97356,I97492,I97676);
nand I_5567 (I97350,I97441,I666485);
nand I_5568 (I97721,I97543,I666479);
DFFARX1 I_5569 (I97721,I3035,I97376,I97365,);
DFFARX1 I_5570 (I97721,I3035,I97376,I97359,);
not I_5571 (I97766,I666479);
nor I_5572 (I97783,I97766,I666470);
and I_5573 (I97800,I97783,I666476);
or I_5574 (I97817,I97800,I666470);
DFFARX1 I_5575 (I97817,I3035,I97376,I97843,);
nand I_5576 (I97851,I97843,I97509);
nor I_5577 (I97353,I97851,I97659);
nor I_5578 (I97347,I97843,I97475);
DFFARX1 I_5579 (I97843,I3035,I97376,I97905,);
not I_5580 (I97913,I97905);
nor I_5581 (I97362,I97913,I97625);
not I_5582 (I97971,I3042);
DFFARX1 I_5583 (I633558,I3035,I97971,I97997,);
DFFARX1 I_5584 (I97997,I3035,I97971,I98014,);
not I_5585 (I97963,I98014);
not I_5586 (I98036,I97997);
DFFARX1 I_5587 (I633558,I3035,I97971,I98062,);
not I_5588 (I98070,I98062);
and I_5589 (I98087,I98036,I633561);
not I_5590 (I98104,I633573);
nand I_5591 (I98121,I98104,I633561);
not I_5592 (I98138,I633579);
nor I_5593 (I98155,I98138,I633570);
nand I_5594 (I98172,I98155,I633576);
nor I_5595 (I98189,I98172,I98121);
DFFARX1 I_5596 (I98189,I3035,I97971,I97939,);
not I_5597 (I98220,I98172);
not I_5598 (I98237,I633570);
nand I_5599 (I98254,I98237,I633561);
nor I_5600 (I98271,I633570,I633573);
nand I_5601 (I97951,I98087,I98271);
nand I_5602 (I97945,I98036,I633570);
nand I_5603 (I98316,I98138,I633567);
DFFARX1 I_5604 (I98316,I3035,I97971,I97960,);
DFFARX1 I_5605 (I98316,I3035,I97971,I97954,);
not I_5606 (I98361,I633567);
nor I_5607 (I98378,I98361,I633564);
and I_5608 (I98395,I98378,I633582);
or I_5609 (I98412,I98395,I633561);
DFFARX1 I_5610 (I98412,I3035,I97971,I98438,);
nand I_5611 (I98446,I98438,I98104);
nor I_5612 (I97948,I98446,I98254);
nor I_5613 (I97942,I98438,I98070);
DFFARX1 I_5614 (I98438,I3035,I97971,I98500,);
not I_5615 (I98508,I98500);
nor I_5616 (I97957,I98508,I98220);
not I_5617 (I98566,I3042);
DFFARX1 I_5618 (I617374,I3035,I98566,I98592,);
DFFARX1 I_5619 (I98592,I3035,I98566,I98609,);
not I_5620 (I98558,I98609);
not I_5621 (I98631,I98592);
DFFARX1 I_5622 (I617374,I3035,I98566,I98657,);
not I_5623 (I98665,I98657);
and I_5624 (I98682,I98631,I617377);
not I_5625 (I98699,I617389);
nand I_5626 (I98716,I98699,I617377);
not I_5627 (I98733,I617395);
nor I_5628 (I98750,I98733,I617386);
nand I_5629 (I98767,I98750,I617392);
nor I_5630 (I98784,I98767,I98716);
DFFARX1 I_5631 (I98784,I3035,I98566,I98534,);
not I_5632 (I98815,I98767);
not I_5633 (I98832,I617386);
nand I_5634 (I98849,I98832,I617377);
nor I_5635 (I98866,I617386,I617389);
nand I_5636 (I98546,I98682,I98866);
nand I_5637 (I98540,I98631,I617386);
nand I_5638 (I98911,I98733,I617383);
DFFARX1 I_5639 (I98911,I3035,I98566,I98555,);
DFFARX1 I_5640 (I98911,I3035,I98566,I98549,);
not I_5641 (I98956,I617383);
nor I_5642 (I98973,I98956,I617380);
and I_5643 (I98990,I98973,I617398);
or I_5644 (I99007,I98990,I617377);
DFFARX1 I_5645 (I99007,I3035,I98566,I99033,);
nand I_5646 (I99041,I99033,I98699);
nor I_5647 (I98543,I99041,I98849);
nor I_5648 (I98537,I99033,I98665);
DFFARX1 I_5649 (I99033,I3035,I98566,I99095,);
not I_5650 (I99103,I99095);
nor I_5651 (I98552,I99103,I98815);
not I_5652 (I99161,I3042);
DFFARX1 I_5653 (I531641,I3035,I99161,I99187,);
DFFARX1 I_5654 (I99187,I3035,I99161,I99204,);
not I_5655 (I99153,I99204);
not I_5656 (I99226,I99187);
DFFARX1 I_5657 (I531650,I3035,I99161,I99252,);
not I_5658 (I99260,I99252);
and I_5659 (I99277,I99226,I531638);
not I_5660 (I99294,I531629);
nand I_5661 (I99311,I99294,I531638);
not I_5662 (I99328,I531635);
nor I_5663 (I99345,I99328,I531653);
nand I_5664 (I99362,I99345,I531626);
nor I_5665 (I99379,I99362,I99311);
DFFARX1 I_5666 (I99379,I3035,I99161,I99129,);
not I_5667 (I99410,I99362);
not I_5668 (I99427,I531653);
nand I_5669 (I99444,I99427,I531638);
nor I_5670 (I99461,I531653,I531629);
nand I_5671 (I99141,I99277,I99461);
nand I_5672 (I99135,I99226,I531653);
nand I_5673 (I99506,I99328,I531632);
DFFARX1 I_5674 (I99506,I3035,I99161,I99150,);
DFFARX1 I_5675 (I99506,I3035,I99161,I99144,);
not I_5676 (I99551,I531632);
nor I_5677 (I99568,I99551,I531644);
and I_5678 (I99585,I99568,I531626);
or I_5679 (I99602,I99585,I531647);
DFFARX1 I_5680 (I99602,I3035,I99161,I99628,);
nand I_5681 (I99636,I99628,I99294);
nor I_5682 (I99138,I99636,I99444);
nor I_5683 (I99132,I99628,I99260);
DFFARX1 I_5684 (I99628,I3035,I99161,I99690,);
not I_5685 (I99698,I99690);
nor I_5686 (I99147,I99698,I99410);
not I_5687 (I99756,I3042);
DFFARX1 I_5688 (I593676,I3035,I99756,I99782,);
DFFARX1 I_5689 (I99782,I3035,I99756,I99799,);
not I_5690 (I99748,I99799);
not I_5691 (I99821,I99782);
DFFARX1 I_5692 (I593676,I3035,I99756,I99847,);
not I_5693 (I99855,I99847);
and I_5694 (I99872,I99821,I593679);
not I_5695 (I99889,I593691);
nand I_5696 (I99906,I99889,I593679);
not I_5697 (I99923,I593697);
nor I_5698 (I99940,I99923,I593688);
nand I_5699 (I99957,I99940,I593694);
nor I_5700 (I99974,I99957,I99906);
DFFARX1 I_5701 (I99974,I3035,I99756,I99724,);
not I_5702 (I100005,I99957);
not I_5703 (I100022,I593688);
nand I_5704 (I100039,I100022,I593679);
nor I_5705 (I100056,I593688,I593691);
nand I_5706 (I99736,I99872,I100056);
nand I_5707 (I99730,I99821,I593688);
nand I_5708 (I100101,I99923,I593685);
DFFARX1 I_5709 (I100101,I3035,I99756,I99745,);
DFFARX1 I_5710 (I100101,I3035,I99756,I99739,);
not I_5711 (I100146,I593685);
nor I_5712 (I100163,I100146,I593682);
and I_5713 (I100180,I100163,I593700);
or I_5714 (I100197,I100180,I593679);
DFFARX1 I_5715 (I100197,I3035,I99756,I100223,);
nand I_5716 (I100231,I100223,I99889);
nor I_5717 (I99733,I100231,I100039);
nor I_5718 (I99727,I100223,I99855);
DFFARX1 I_5719 (I100223,I3035,I99756,I100285,);
not I_5720 (I100293,I100285);
nor I_5721 (I99742,I100293,I100005);
not I_5722 (I100351,I3042);
DFFARX1 I_5723 (I17842,I3035,I100351,I100377,);
DFFARX1 I_5724 (I100377,I3035,I100351,I100394,);
not I_5725 (I100343,I100394);
not I_5726 (I100416,I100377);
DFFARX1 I_5727 (I17818,I3035,I100351,I100442,);
not I_5728 (I100450,I100442);
and I_5729 (I100467,I100416,I17833);
not I_5730 (I100484,I17821);
nand I_5731 (I100501,I100484,I17833);
not I_5732 (I100518,I17824);
nor I_5733 (I100535,I100518,I17836);
nand I_5734 (I100552,I100535,I17827);
nor I_5735 (I100569,I100552,I100501);
DFFARX1 I_5736 (I100569,I3035,I100351,I100319,);
not I_5737 (I100600,I100552);
not I_5738 (I100617,I17836);
nand I_5739 (I100634,I100617,I17833);
nor I_5740 (I100651,I17836,I17821);
nand I_5741 (I100331,I100467,I100651);
nand I_5742 (I100325,I100416,I17836);
nand I_5743 (I100696,I100518,I17830);
DFFARX1 I_5744 (I100696,I3035,I100351,I100340,);
DFFARX1 I_5745 (I100696,I3035,I100351,I100334,);
not I_5746 (I100741,I17830);
nor I_5747 (I100758,I100741,I17821);
and I_5748 (I100775,I100758,I17818);
or I_5749 (I100792,I100775,I17839);
DFFARX1 I_5750 (I100792,I3035,I100351,I100818,);
nand I_5751 (I100826,I100818,I100484);
nor I_5752 (I100328,I100826,I100634);
nor I_5753 (I100322,I100818,I100450);
DFFARX1 I_5754 (I100818,I3035,I100351,I100880,);
not I_5755 (I100888,I100880);
nor I_5756 (I100337,I100888,I100600);
not I_5757 (I100946,I3042);
DFFARX1 I_5758 (I409986,I3035,I100946,I100972,);
DFFARX1 I_5759 (I100972,I3035,I100946,I100989,);
not I_5760 (I100938,I100989);
not I_5761 (I101011,I100972);
DFFARX1 I_5762 (I409983,I3035,I100946,I101037,);
not I_5763 (I101045,I101037);
and I_5764 (I101062,I101011,I409989);
not I_5765 (I101079,I409974);
nand I_5766 (I101096,I101079,I409989);
not I_5767 (I101113,I409977);
nor I_5768 (I101130,I101113,I409998);
nand I_5769 (I101147,I101130,I409995);
nor I_5770 (I101164,I101147,I101096);
DFFARX1 I_5771 (I101164,I3035,I100946,I100914,);
not I_5772 (I101195,I101147);
not I_5773 (I101212,I409998);
nand I_5774 (I101229,I101212,I409989);
nor I_5775 (I101246,I409998,I409974);
nand I_5776 (I100926,I101062,I101246);
nand I_5777 (I100920,I101011,I409998);
nand I_5778 (I101291,I101113,I409974);
DFFARX1 I_5779 (I101291,I3035,I100946,I100935,);
DFFARX1 I_5780 (I101291,I3035,I100946,I100929,);
not I_5781 (I101336,I409974);
nor I_5782 (I101353,I101336,I409980);
and I_5783 (I101370,I101353,I409992);
or I_5784 (I101387,I101370,I409977);
DFFARX1 I_5785 (I101387,I3035,I100946,I101413,);
nand I_5786 (I101421,I101413,I101079);
nor I_5787 (I100923,I101421,I101229);
nor I_5788 (I100917,I101413,I101045);
DFFARX1 I_5789 (I101413,I3035,I100946,I101475,);
not I_5790 (I101483,I101475);
nor I_5791 (I100932,I101483,I101195);
not I_5792 (I101541,I3042);
DFFARX1 I_5793 (I351608,I3035,I101541,I101567,);
DFFARX1 I_5794 (I101567,I3035,I101541,I101584,);
not I_5795 (I101533,I101584);
not I_5796 (I101606,I101567);
DFFARX1 I_5797 (I351605,I3035,I101541,I101632,);
not I_5798 (I101640,I101632);
and I_5799 (I101657,I101606,I351611);
not I_5800 (I101674,I351596);
nand I_5801 (I101691,I101674,I351611);
not I_5802 (I101708,I351599);
nor I_5803 (I101725,I101708,I351620);
nand I_5804 (I101742,I101725,I351617);
nor I_5805 (I101759,I101742,I101691);
DFFARX1 I_5806 (I101759,I3035,I101541,I101509,);
not I_5807 (I101790,I101742);
not I_5808 (I101807,I351620);
nand I_5809 (I101824,I101807,I351611);
nor I_5810 (I101841,I351620,I351596);
nand I_5811 (I101521,I101657,I101841);
nand I_5812 (I101515,I101606,I351620);
nand I_5813 (I101886,I101708,I351596);
DFFARX1 I_5814 (I101886,I3035,I101541,I101530,);
DFFARX1 I_5815 (I101886,I3035,I101541,I101524,);
not I_5816 (I101931,I351596);
nor I_5817 (I101948,I101931,I351602);
and I_5818 (I101965,I101948,I351614);
or I_5819 (I101982,I101965,I351599);
DFFARX1 I_5820 (I101982,I3035,I101541,I102008,);
nand I_5821 (I102016,I102008,I101674);
nor I_5822 (I101518,I102016,I101824);
nor I_5823 (I101512,I102008,I101640);
DFFARX1 I_5824 (I102008,I3035,I101541,I102070,);
not I_5825 (I102078,I102070);
nor I_5826 (I101527,I102078,I101790);
not I_5827 (I102136,I3042);
DFFARX1 I_5828 (I396114,I3035,I102136,I102162,);
DFFARX1 I_5829 (I102162,I3035,I102136,I102179,);
not I_5830 (I102128,I102179);
not I_5831 (I102201,I102162);
DFFARX1 I_5832 (I396111,I3035,I102136,I102227,);
not I_5833 (I102235,I102227);
and I_5834 (I102252,I102201,I396117);
not I_5835 (I102269,I396102);
nand I_5836 (I102286,I102269,I396117);
not I_5837 (I102303,I396105);
nor I_5838 (I102320,I102303,I396126);
nand I_5839 (I102337,I102320,I396123);
nor I_5840 (I102354,I102337,I102286);
DFFARX1 I_5841 (I102354,I3035,I102136,I102104,);
not I_5842 (I102385,I102337);
not I_5843 (I102402,I396126);
nand I_5844 (I102419,I102402,I396117);
nor I_5845 (I102436,I396126,I396102);
nand I_5846 (I102116,I102252,I102436);
nand I_5847 (I102110,I102201,I396126);
nand I_5848 (I102481,I102303,I396102);
DFFARX1 I_5849 (I102481,I3035,I102136,I102125,);
DFFARX1 I_5850 (I102481,I3035,I102136,I102119,);
not I_5851 (I102526,I396102);
nor I_5852 (I102543,I102526,I396108);
and I_5853 (I102560,I102543,I396120);
or I_5854 (I102577,I102560,I396105);
DFFARX1 I_5855 (I102577,I3035,I102136,I102603,);
nand I_5856 (I102611,I102603,I102269);
nor I_5857 (I102113,I102611,I102419);
nor I_5858 (I102107,I102603,I102235);
DFFARX1 I_5859 (I102603,I3035,I102136,I102665,);
not I_5860 (I102673,I102665);
nor I_5861 (I102122,I102673,I102385);
not I_5862 (I102731,I3042);
DFFARX1 I_5863 (I445629,I3035,I102731,I102757,);
DFFARX1 I_5864 (I102757,I3035,I102731,I102774,);
not I_5865 (I102723,I102774);
not I_5866 (I102796,I102757);
DFFARX1 I_5867 (I445623,I3035,I102731,I102822,);
not I_5868 (I102830,I102822);
and I_5869 (I102847,I102796,I445641);
not I_5870 (I102864,I445629);
nand I_5871 (I102881,I102864,I445641);
not I_5872 (I102898,I445623);
nor I_5873 (I102915,I102898,I445635);
nand I_5874 (I102932,I102915,I445626);
nor I_5875 (I102949,I102932,I102881);
DFFARX1 I_5876 (I102949,I3035,I102731,I102699,);
not I_5877 (I102980,I102932);
not I_5878 (I102997,I445635);
nand I_5879 (I103014,I102997,I445641);
nor I_5880 (I103031,I445635,I445629);
nand I_5881 (I102711,I102847,I103031);
nand I_5882 (I102705,I102796,I445635);
nand I_5883 (I103076,I102898,I445638);
DFFARX1 I_5884 (I103076,I3035,I102731,I102720,);
DFFARX1 I_5885 (I103076,I3035,I102731,I102714,);
not I_5886 (I103121,I445638);
nor I_5887 (I103138,I103121,I445644);
and I_5888 (I103155,I103138,I445626);
or I_5889 (I103172,I103155,I445632);
DFFARX1 I_5890 (I103172,I3035,I102731,I103198,);
nand I_5891 (I103206,I103198,I102864);
nor I_5892 (I102708,I103206,I103014);
nor I_5893 (I102702,I103198,I102830);
DFFARX1 I_5894 (I103198,I3035,I102731,I103260,);
not I_5895 (I103268,I103260);
nor I_5896 (I102717,I103268,I102980);
not I_5897 (I103326,I3042);
DFFARX1 I_5898 (I36272,I3035,I103326,I103352,);
DFFARX1 I_5899 (I103352,I3035,I103326,I103369,);
not I_5900 (I103318,I103369);
not I_5901 (I103391,I103352);
DFFARX1 I_5902 (I36266,I3035,I103326,I103417,);
not I_5903 (I103425,I103417);
and I_5904 (I103442,I103391,I36263);
not I_5905 (I103459,I36284);
nand I_5906 (I103476,I103459,I36263);
not I_5907 (I103493,I36278);
nor I_5908 (I103510,I103493,I36269);
nand I_5909 (I103527,I103510,I36275);
nor I_5910 (I103544,I103527,I103476);
DFFARX1 I_5911 (I103544,I3035,I103326,I103294,);
not I_5912 (I103575,I103527);
not I_5913 (I103592,I36269);
nand I_5914 (I103609,I103592,I36263);
nor I_5915 (I103626,I36269,I36284);
nand I_5916 (I103306,I103442,I103626);
nand I_5917 (I103300,I103391,I36269);
nand I_5918 (I103671,I103493,I36263);
DFFARX1 I_5919 (I103671,I3035,I103326,I103315,);
DFFARX1 I_5920 (I103671,I3035,I103326,I103309,);
not I_5921 (I103716,I36263);
nor I_5922 (I103733,I103716,I36281);
and I_5923 (I103750,I103733,I36287);
or I_5924 (I103767,I103750,I36266);
DFFARX1 I_5925 (I103767,I3035,I103326,I103793,);
nand I_5926 (I103801,I103793,I103459);
nor I_5927 (I103303,I103801,I103609);
nor I_5928 (I103297,I103793,I103425);
DFFARX1 I_5929 (I103793,I3035,I103326,I103855,);
not I_5930 (I103863,I103855);
nor I_5931 (I103312,I103863,I103575);
not I_5932 (I103921,I3042);
DFFARX1 I_5933 (I261469,I3035,I103921,I103947,);
DFFARX1 I_5934 (I103947,I3035,I103921,I103964,);
not I_5935 (I103913,I103964);
not I_5936 (I103986,I103947);
DFFARX1 I_5937 (I261457,I3035,I103921,I104012,);
not I_5938 (I104020,I104012);
and I_5939 (I104037,I103986,I261466);
not I_5940 (I104054,I261463);
nand I_5941 (I104071,I104054,I261466);
not I_5942 (I104088,I261454);
nor I_5943 (I104105,I104088,I261460);
nand I_5944 (I104122,I104105,I261445);
nor I_5945 (I104139,I104122,I104071);
DFFARX1 I_5946 (I104139,I3035,I103921,I103889,);
not I_5947 (I104170,I104122);
not I_5948 (I104187,I261460);
nand I_5949 (I104204,I104187,I261466);
nor I_5950 (I104221,I261460,I261463);
nand I_5951 (I103901,I104037,I104221);
nand I_5952 (I103895,I103986,I261460);
nand I_5953 (I104266,I104088,I261445);
DFFARX1 I_5954 (I104266,I3035,I103921,I103910,);
DFFARX1 I_5955 (I104266,I3035,I103921,I103904,);
not I_5956 (I104311,I261445);
nor I_5957 (I104328,I104311,I261451);
and I_5958 (I104345,I104328,I261448);
or I_5959 (I104362,I104345,I261472);
DFFARX1 I_5960 (I104362,I3035,I103921,I104388,);
nand I_5961 (I104396,I104388,I104054);
nor I_5962 (I103898,I104396,I104204);
nor I_5963 (I103892,I104388,I104020);
DFFARX1 I_5964 (I104388,I3035,I103921,I104450,);
not I_5965 (I104458,I104450);
nor I_5966 (I103907,I104458,I104170);
not I_5967 (I104516,I3042);
DFFARX1 I_5968 (I68946,I3035,I104516,I104542,);
DFFARX1 I_5969 (I104542,I3035,I104516,I104559,);
not I_5970 (I104508,I104559);
not I_5971 (I104581,I104542);
DFFARX1 I_5972 (I68940,I3035,I104516,I104607,);
not I_5973 (I104615,I104607);
and I_5974 (I104632,I104581,I68937);
not I_5975 (I104649,I68958);
nand I_5976 (I104666,I104649,I68937);
not I_5977 (I104683,I68952);
nor I_5978 (I104700,I104683,I68943);
nand I_5979 (I104717,I104700,I68949);
nor I_5980 (I104734,I104717,I104666);
DFFARX1 I_5981 (I104734,I3035,I104516,I104484,);
not I_5982 (I104765,I104717);
not I_5983 (I104782,I68943);
nand I_5984 (I104799,I104782,I68937);
nor I_5985 (I104816,I68943,I68958);
nand I_5986 (I104496,I104632,I104816);
nand I_5987 (I104490,I104581,I68943);
nand I_5988 (I104861,I104683,I68937);
DFFARX1 I_5989 (I104861,I3035,I104516,I104505,);
DFFARX1 I_5990 (I104861,I3035,I104516,I104499,);
not I_5991 (I104906,I68937);
nor I_5992 (I104923,I104906,I68955);
and I_5993 (I104940,I104923,I68961);
or I_5994 (I104957,I104940,I68940);
DFFARX1 I_5995 (I104957,I3035,I104516,I104983,);
nand I_5996 (I104991,I104983,I104649);
nor I_5997 (I104493,I104991,I104799);
nor I_5998 (I104487,I104983,I104615);
DFFARX1 I_5999 (I104983,I3035,I104516,I105045,);
not I_6000 (I105053,I105045);
nor I_6001 (I104502,I105053,I104765);
not I_6002 (I105111,I3042);
DFFARX1 I_6003 (I245693,I3035,I105111,I105137,);
DFFARX1 I_6004 (I105137,I3035,I105111,I105154,);
not I_6005 (I105103,I105154);
not I_6006 (I105176,I105137);
DFFARX1 I_6007 (I245681,I3035,I105111,I105202,);
not I_6008 (I105210,I105202);
and I_6009 (I105227,I105176,I245690);
not I_6010 (I105244,I245687);
nand I_6011 (I105261,I105244,I245690);
not I_6012 (I105278,I245678);
nor I_6013 (I105295,I105278,I245684);
nand I_6014 (I105312,I105295,I245669);
nor I_6015 (I105329,I105312,I105261);
DFFARX1 I_6016 (I105329,I3035,I105111,I105079,);
not I_6017 (I105360,I105312);
not I_6018 (I105377,I245684);
nand I_6019 (I105394,I105377,I245690);
nor I_6020 (I105411,I245684,I245687);
nand I_6021 (I105091,I105227,I105411);
nand I_6022 (I105085,I105176,I245684);
nand I_6023 (I105456,I105278,I245669);
DFFARX1 I_6024 (I105456,I3035,I105111,I105100,);
DFFARX1 I_6025 (I105456,I3035,I105111,I105094,);
not I_6026 (I105501,I245669);
nor I_6027 (I105518,I105501,I245675);
and I_6028 (I105535,I105518,I245672);
or I_6029 (I105552,I105535,I245696);
DFFARX1 I_6030 (I105552,I3035,I105111,I105578,);
nand I_6031 (I105586,I105578,I105244);
nor I_6032 (I105088,I105586,I105394);
nor I_6033 (I105082,I105578,I105210);
DFFARX1 I_6034 (I105578,I3035,I105111,I105640,);
not I_6035 (I105648,I105640);
nor I_6036 (I105097,I105648,I105360);
not I_6037 (I105706,I3042);
DFFARX1 I_6038 (I77132,I3035,I105706,I105732,);
DFFARX1 I_6039 (I105732,I3035,I105706,I105749,);
not I_6040 (I105698,I105749);
not I_6041 (I105771,I105732);
DFFARX1 I_6042 (I77117,I3035,I105706,I105797,);
not I_6043 (I105805,I105797);
and I_6044 (I105822,I105771,I77138);
not I_6045 (I105839,I77129);
nand I_6046 (I105856,I105839,I77138);
not I_6047 (I105873,I77114);
nor I_6048 (I105890,I105873,I77126);
nand I_6049 (I105907,I105890,I77141);
nor I_6050 (I105924,I105907,I105856);
DFFARX1 I_6051 (I105924,I3035,I105706,I105674,);
not I_6052 (I105955,I105907);
not I_6053 (I105972,I77126);
nand I_6054 (I105989,I105972,I77138);
nor I_6055 (I106006,I77126,I77129);
nand I_6056 (I105686,I105822,I106006);
nand I_6057 (I105680,I105771,I77126);
nand I_6058 (I106051,I105873,I77120);
DFFARX1 I_6059 (I106051,I3035,I105706,I105695,);
DFFARX1 I_6060 (I106051,I3035,I105706,I105689,);
not I_6061 (I106096,I77120);
nor I_6062 (I106113,I106096,I77123);
and I_6063 (I106130,I106113,I77114);
or I_6064 (I106147,I106130,I77135);
DFFARX1 I_6065 (I106147,I3035,I105706,I106173,);
nand I_6066 (I106181,I106173,I105839);
nor I_6067 (I105683,I106181,I105989);
nor I_6068 (I105677,I106173,I105805);
DFFARX1 I_6069 (I106173,I3035,I105706,I106235,);
not I_6070 (I106243,I106235);
nor I_6071 (I105692,I106243,I105955);
not I_6072 (I106301,I3042);
DFFARX1 I_6073 (I15207,I3035,I106301,I106327,);
DFFARX1 I_6074 (I106327,I3035,I106301,I106344,);
not I_6075 (I106293,I106344);
not I_6076 (I106366,I106327);
DFFARX1 I_6077 (I15183,I3035,I106301,I106392,);
not I_6078 (I106400,I106392);
and I_6079 (I106417,I106366,I15198);
not I_6080 (I106434,I15186);
nand I_6081 (I106451,I106434,I15198);
not I_6082 (I106468,I15189);
nor I_6083 (I106485,I106468,I15201);
nand I_6084 (I106502,I106485,I15192);
nor I_6085 (I106519,I106502,I106451);
DFFARX1 I_6086 (I106519,I3035,I106301,I106269,);
not I_6087 (I106550,I106502);
not I_6088 (I106567,I15201);
nand I_6089 (I106584,I106567,I15198);
nor I_6090 (I106601,I15201,I15186);
nand I_6091 (I106281,I106417,I106601);
nand I_6092 (I106275,I106366,I15201);
nand I_6093 (I106646,I106468,I15195);
DFFARX1 I_6094 (I106646,I3035,I106301,I106290,);
DFFARX1 I_6095 (I106646,I3035,I106301,I106284,);
not I_6096 (I106691,I15195);
nor I_6097 (I106708,I106691,I15186);
and I_6098 (I106725,I106708,I15183);
or I_6099 (I106742,I106725,I15204);
DFFARX1 I_6100 (I106742,I3035,I106301,I106768,);
nand I_6101 (I106776,I106768,I106434);
nor I_6102 (I106278,I106776,I106584);
nor I_6103 (I106272,I106768,I106400);
DFFARX1 I_6104 (I106768,I3035,I106301,I106830,);
not I_6105 (I106838,I106830);
nor I_6106 (I106287,I106838,I106550);
not I_6107 (I106896,I3042);
DFFARX1 I_6108 (I567805,I3035,I106896,I106922,);
DFFARX1 I_6109 (I106922,I3035,I106896,I106939,);
not I_6110 (I106888,I106939);
not I_6111 (I106961,I106922);
DFFARX1 I_6112 (I567814,I3035,I106896,I106987,);
not I_6113 (I106995,I106987);
and I_6114 (I107012,I106961,I567808);
not I_6115 (I107029,I567802);
nand I_6116 (I107046,I107029,I567808);
not I_6117 (I107063,I567817);
nor I_6118 (I107080,I107063,I567805);
nand I_6119 (I107097,I107080,I567811);
nor I_6120 (I107114,I107097,I107046);
DFFARX1 I_6121 (I107114,I3035,I106896,I106864,);
not I_6122 (I107145,I107097);
not I_6123 (I107162,I567805);
nand I_6124 (I107179,I107162,I567808);
nor I_6125 (I107196,I567805,I567802);
nand I_6126 (I106876,I107012,I107196);
nand I_6127 (I106870,I106961,I567805);
nand I_6128 (I107241,I107063,I567808);
DFFARX1 I_6129 (I107241,I3035,I106896,I106885,);
DFFARX1 I_6130 (I107241,I3035,I106896,I106879,);
not I_6131 (I107286,I567808);
nor I_6132 (I107303,I107286,I567823);
and I_6133 (I107320,I107303,I567820);
or I_6134 (I107337,I107320,I567802);
DFFARX1 I_6135 (I107337,I3035,I106896,I107363,);
nand I_6136 (I107371,I107363,I107029);
nor I_6137 (I106873,I107371,I107179);
nor I_6138 (I106867,I107363,I106995);
DFFARX1 I_6139 (I107363,I3035,I106896,I107425,);
not I_6140 (I107433,I107425);
nor I_6141 (I106882,I107433,I107145);
not I_6142 (I107491,I3042);
DFFARX1 I_6143 (I415188,I3035,I107491,I107517,);
DFFARX1 I_6144 (I107517,I3035,I107491,I107534,);
not I_6145 (I107483,I107534);
not I_6146 (I107556,I107517);
DFFARX1 I_6147 (I415185,I3035,I107491,I107582,);
not I_6148 (I107590,I107582);
and I_6149 (I107607,I107556,I415191);
not I_6150 (I107624,I415176);
nand I_6151 (I107641,I107624,I415191);
not I_6152 (I107658,I415179);
nor I_6153 (I107675,I107658,I415200);
nand I_6154 (I107692,I107675,I415197);
nor I_6155 (I107709,I107692,I107641);
DFFARX1 I_6156 (I107709,I3035,I107491,I107459,);
not I_6157 (I107740,I107692);
not I_6158 (I107757,I415200);
nand I_6159 (I107774,I107757,I415191);
nor I_6160 (I107791,I415200,I415176);
nand I_6161 (I107471,I107607,I107791);
nand I_6162 (I107465,I107556,I415200);
nand I_6163 (I107836,I107658,I415176);
DFFARX1 I_6164 (I107836,I3035,I107491,I107480,);
DFFARX1 I_6165 (I107836,I3035,I107491,I107474,);
not I_6166 (I107881,I415176);
nor I_6167 (I107898,I107881,I415182);
and I_6168 (I107915,I107898,I415194);
or I_6169 (I107932,I107915,I415179);
DFFARX1 I_6170 (I107932,I3035,I107491,I107958,);
nand I_6171 (I107966,I107958,I107624);
nor I_6172 (I107468,I107966,I107774);
nor I_6173 (I107462,I107958,I107590);
DFFARX1 I_6174 (I107958,I3035,I107491,I108020,);
not I_6175 (I108028,I108020);
nor I_6176 (I107477,I108028,I107740);
not I_6177 (I108086,I3042);
DFFARX1 I_6178 (I411720,I3035,I108086,I108112,);
DFFARX1 I_6179 (I108112,I3035,I108086,I108129,);
not I_6180 (I108078,I108129);
not I_6181 (I108151,I108112);
DFFARX1 I_6182 (I411717,I3035,I108086,I108177,);
not I_6183 (I108185,I108177);
and I_6184 (I108202,I108151,I411723);
not I_6185 (I108219,I411708);
nand I_6186 (I108236,I108219,I411723);
not I_6187 (I108253,I411711);
nor I_6188 (I108270,I108253,I411732);
nand I_6189 (I108287,I108270,I411729);
nor I_6190 (I108304,I108287,I108236);
DFFARX1 I_6191 (I108304,I3035,I108086,I108054,);
not I_6192 (I108335,I108287);
not I_6193 (I108352,I411732);
nand I_6194 (I108369,I108352,I411723);
nor I_6195 (I108386,I411732,I411708);
nand I_6196 (I108066,I108202,I108386);
nand I_6197 (I108060,I108151,I411732);
nand I_6198 (I108431,I108253,I411708);
DFFARX1 I_6199 (I108431,I3035,I108086,I108075,);
DFFARX1 I_6200 (I108431,I3035,I108086,I108069,);
not I_6201 (I108476,I411708);
nor I_6202 (I108493,I108476,I411714);
and I_6203 (I108510,I108493,I411726);
or I_6204 (I108527,I108510,I411711);
DFFARX1 I_6205 (I108527,I3035,I108086,I108553,);
nand I_6206 (I108561,I108553,I108219);
nor I_6207 (I108063,I108561,I108369);
nor I_6208 (I108057,I108553,I108185);
DFFARX1 I_6209 (I108553,I3035,I108086,I108615,);
not I_6210 (I108623,I108615);
nor I_6211 (I108072,I108623,I108335);
not I_6212 (I108681,I3042);
DFFARX1 I_6213 (I271805,I3035,I108681,I108707,);
DFFARX1 I_6214 (I108707,I3035,I108681,I108724,);
not I_6215 (I108673,I108724);
not I_6216 (I108746,I108707);
DFFARX1 I_6217 (I271793,I3035,I108681,I108772,);
not I_6218 (I108780,I108772);
and I_6219 (I108797,I108746,I271802);
not I_6220 (I108814,I271799);
nand I_6221 (I108831,I108814,I271802);
not I_6222 (I108848,I271790);
nor I_6223 (I108865,I108848,I271796);
nand I_6224 (I108882,I108865,I271781);
nor I_6225 (I108899,I108882,I108831);
DFFARX1 I_6226 (I108899,I3035,I108681,I108649,);
not I_6227 (I108930,I108882);
not I_6228 (I108947,I271796);
nand I_6229 (I108964,I108947,I271802);
nor I_6230 (I108981,I271796,I271799);
nand I_6231 (I108661,I108797,I108981);
nand I_6232 (I108655,I108746,I271796);
nand I_6233 (I109026,I108848,I271781);
DFFARX1 I_6234 (I109026,I3035,I108681,I108670,);
DFFARX1 I_6235 (I109026,I3035,I108681,I108664,);
not I_6236 (I109071,I271781);
nor I_6237 (I109088,I109071,I271787);
and I_6238 (I109105,I109088,I271784);
or I_6239 (I109122,I109105,I271808);
DFFARX1 I_6240 (I109122,I3035,I108681,I109148,);
nand I_6241 (I109156,I109148,I108814);
nor I_6242 (I108658,I109156,I108964);
nor I_6243 (I108652,I109148,I108780);
DFFARX1 I_6244 (I109148,I3035,I108681,I109210,);
not I_6245 (I109218,I109210);
nor I_6246 (I108667,I109218,I108930);
not I_6247 (I109276,I3042);
DFFARX1 I_6248 (I680005,I3035,I109276,I109302,);
DFFARX1 I_6249 (I109302,I3035,I109276,I109319,);
not I_6250 (I109268,I109319);
not I_6251 (I109341,I109302);
DFFARX1 I_6252 (I680017,I3035,I109276,I109367,);
not I_6253 (I109375,I109367);
and I_6254 (I109392,I109341,I680011);
not I_6255 (I109409,I680023);
nand I_6256 (I109426,I109409,I680011);
not I_6257 (I109443,I680008);
nor I_6258 (I109460,I109443,I680020);
nand I_6259 (I109477,I109460,I680002);
nor I_6260 (I109494,I109477,I109426);
DFFARX1 I_6261 (I109494,I3035,I109276,I109244,);
not I_6262 (I109525,I109477);
not I_6263 (I109542,I680020);
nand I_6264 (I109559,I109542,I680011);
nor I_6265 (I109576,I680020,I680023);
nand I_6266 (I109256,I109392,I109576);
nand I_6267 (I109250,I109341,I680020);
nand I_6268 (I109621,I109443,I680014);
DFFARX1 I_6269 (I109621,I3035,I109276,I109265,);
DFFARX1 I_6270 (I109621,I3035,I109276,I109259,);
not I_6271 (I109666,I680014);
nor I_6272 (I109683,I109666,I680005);
and I_6273 (I109700,I109683,I680002);
or I_6274 (I109717,I109700,I680026);
DFFARX1 I_6275 (I109717,I3035,I109276,I109743,);
nand I_6276 (I109751,I109743,I109409);
nor I_6277 (I109253,I109751,I109559);
nor I_6278 (I109247,I109743,I109375);
DFFARX1 I_6279 (I109743,I3035,I109276,I109805,);
not I_6280 (I109813,I109805);
nor I_6281 (I109262,I109813,I109525);
not I_6282 (I109871,I3042);
DFFARX1 I_6283 (I231005,I3035,I109871,I109897,);
DFFARX1 I_6284 (I109897,I3035,I109871,I109914,);
not I_6285 (I109863,I109914);
not I_6286 (I109936,I109897);
DFFARX1 I_6287 (I230993,I3035,I109871,I109962,);
not I_6288 (I109970,I109962);
and I_6289 (I109987,I109936,I231002);
not I_6290 (I110004,I230999);
nand I_6291 (I110021,I110004,I231002);
not I_6292 (I110038,I230990);
nor I_6293 (I110055,I110038,I230996);
nand I_6294 (I110072,I110055,I230981);
nor I_6295 (I110089,I110072,I110021);
DFFARX1 I_6296 (I110089,I3035,I109871,I109839,);
not I_6297 (I110120,I110072);
not I_6298 (I110137,I230996);
nand I_6299 (I110154,I110137,I231002);
nor I_6300 (I110171,I230996,I230999);
nand I_6301 (I109851,I109987,I110171);
nand I_6302 (I109845,I109936,I230996);
nand I_6303 (I110216,I110038,I230981);
DFFARX1 I_6304 (I110216,I3035,I109871,I109860,);
DFFARX1 I_6305 (I110216,I3035,I109871,I109854,);
not I_6306 (I110261,I230981);
nor I_6307 (I110278,I110261,I230987);
and I_6308 (I110295,I110278,I230984);
or I_6309 (I110312,I110295,I231008);
DFFARX1 I_6310 (I110312,I3035,I109871,I110338,);
nand I_6311 (I110346,I110338,I110004);
nor I_6312 (I109848,I110346,I110154);
nor I_6313 (I109842,I110338,I109970);
DFFARX1 I_6314 (I110338,I3035,I109871,I110400,);
not I_6315 (I110408,I110400);
nor I_6316 (I109857,I110408,I110120);
not I_6317 (I110466,I3042);
DFFARX1 I_6318 (I662680,I3035,I110466,I110492,);
DFFARX1 I_6319 (I110492,I3035,I110466,I110509,);
not I_6320 (I110458,I110509);
not I_6321 (I110531,I110492);
DFFARX1 I_6322 (I662665,I3035,I110466,I110557,);
not I_6323 (I110565,I110557);
and I_6324 (I110582,I110531,I662683);
not I_6325 (I110599,I662665);
nand I_6326 (I110616,I110599,I662683);
not I_6327 (I110633,I662686);
nor I_6328 (I110650,I110633,I662677);
nand I_6329 (I110667,I110650,I662674);
nor I_6330 (I110684,I110667,I110616);
DFFARX1 I_6331 (I110684,I3035,I110466,I110434,);
not I_6332 (I110715,I110667);
not I_6333 (I110732,I662677);
nand I_6334 (I110749,I110732,I662683);
nor I_6335 (I110766,I662677,I662665);
nand I_6336 (I110446,I110582,I110766);
nand I_6337 (I110440,I110531,I662677);
nand I_6338 (I110811,I110633,I662671);
DFFARX1 I_6339 (I110811,I3035,I110466,I110455,);
DFFARX1 I_6340 (I110811,I3035,I110466,I110449,);
not I_6341 (I110856,I662671);
nor I_6342 (I110873,I110856,I662662);
and I_6343 (I110890,I110873,I662668);
or I_6344 (I110907,I110890,I662662);
DFFARX1 I_6345 (I110907,I3035,I110466,I110933,);
nand I_6346 (I110941,I110933,I110599);
nor I_6347 (I110443,I110941,I110749);
nor I_6348 (I110437,I110933,I110565);
DFFARX1 I_6349 (I110933,I3035,I110466,I110995,);
not I_6350 (I111003,I110995);
nor I_6351 (I110452,I111003,I110715);
not I_6352 (I111061,I3042);
DFFARX1 I_6353 (I597722,I3035,I111061,I111087,);
DFFARX1 I_6354 (I111087,I3035,I111061,I111104,);
not I_6355 (I111053,I111104);
not I_6356 (I111126,I111087);
DFFARX1 I_6357 (I597722,I3035,I111061,I111152,);
not I_6358 (I111160,I111152);
and I_6359 (I111177,I111126,I597725);
not I_6360 (I111194,I597737);
nand I_6361 (I111211,I111194,I597725);
not I_6362 (I111228,I597743);
nor I_6363 (I111245,I111228,I597734);
nand I_6364 (I111262,I111245,I597740);
nor I_6365 (I111279,I111262,I111211);
DFFARX1 I_6366 (I111279,I3035,I111061,I111029,);
not I_6367 (I111310,I111262);
not I_6368 (I111327,I597734);
nand I_6369 (I111344,I111327,I597725);
nor I_6370 (I111361,I597734,I597737);
nand I_6371 (I111041,I111177,I111361);
nand I_6372 (I111035,I111126,I597734);
nand I_6373 (I111406,I111228,I597731);
DFFARX1 I_6374 (I111406,I3035,I111061,I111050,);
DFFARX1 I_6375 (I111406,I3035,I111061,I111044,);
not I_6376 (I111451,I597731);
nor I_6377 (I111468,I111451,I597728);
and I_6378 (I111485,I111468,I597746);
or I_6379 (I111502,I111485,I597725);
DFFARX1 I_6380 (I111502,I3035,I111061,I111528,);
nand I_6381 (I111536,I111528,I111194);
nor I_6382 (I111038,I111536,I111344);
nor I_6383 (I111032,I111528,I111160);
DFFARX1 I_6384 (I111528,I3035,I111061,I111590,);
not I_6385 (I111598,I111590);
nor I_6386 (I111047,I111598,I111310);
not I_6387 (I111656,I3042);
DFFARX1 I_6388 (I546487,I3035,I111656,I111682,);
DFFARX1 I_6389 (I111682,I3035,I111656,I111699,);
not I_6390 (I111648,I111699);
not I_6391 (I111721,I111682);
DFFARX1 I_6392 (I546496,I3035,I111656,I111747,);
not I_6393 (I111755,I111747);
and I_6394 (I111772,I111721,I546490);
not I_6395 (I111789,I546484);
nand I_6396 (I111806,I111789,I546490);
not I_6397 (I111823,I546499);
nor I_6398 (I111840,I111823,I546487);
nand I_6399 (I111857,I111840,I546493);
nor I_6400 (I111874,I111857,I111806);
DFFARX1 I_6401 (I111874,I3035,I111656,I111624,);
not I_6402 (I111905,I111857);
not I_6403 (I111922,I546487);
nand I_6404 (I111939,I111922,I546490);
nor I_6405 (I111956,I546487,I546484);
nand I_6406 (I111636,I111772,I111956);
nand I_6407 (I111630,I111721,I546487);
nand I_6408 (I112001,I111823,I546490);
DFFARX1 I_6409 (I112001,I3035,I111656,I111645,);
DFFARX1 I_6410 (I112001,I3035,I111656,I111639,);
not I_6411 (I112046,I546490);
nor I_6412 (I112063,I112046,I546505);
and I_6413 (I112080,I112063,I546502);
or I_6414 (I112097,I112080,I546484);
DFFARX1 I_6415 (I112097,I3035,I111656,I112123,);
nand I_6416 (I112131,I112123,I111789);
nor I_6417 (I111633,I112131,I111939);
nor I_6418 (I111627,I112123,I111755);
DFFARX1 I_6419 (I112123,I3035,I111656,I112185,);
not I_6420 (I112193,I112185);
nor I_6421 (I111642,I112193,I111905);
not I_6422 (I112251,I3042);
DFFARX1 I_6423 (I562756,I3035,I112251,I112277,);
DFFARX1 I_6424 (I112277,I3035,I112251,I112294,);
not I_6425 (I112243,I112294);
not I_6426 (I112316,I112277);
DFFARX1 I_6427 (I562765,I3035,I112251,I112342,);
not I_6428 (I112350,I112342);
and I_6429 (I112367,I112316,I562759);
not I_6430 (I112384,I562753);
nand I_6431 (I112401,I112384,I562759);
not I_6432 (I112418,I562768);
nor I_6433 (I112435,I112418,I562756);
nand I_6434 (I112452,I112435,I562762);
nor I_6435 (I112469,I112452,I112401);
DFFARX1 I_6436 (I112469,I3035,I112251,I112219,);
not I_6437 (I112500,I112452);
not I_6438 (I112517,I562756);
nand I_6439 (I112534,I112517,I562759);
nor I_6440 (I112551,I562756,I562753);
nand I_6441 (I112231,I112367,I112551);
nand I_6442 (I112225,I112316,I562756);
nand I_6443 (I112596,I112418,I562759);
DFFARX1 I_6444 (I112596,I3035,I112251,I112240,);
DFFARX1 I_6445 (I112596,I3035,I112251,I112234,);
not I_6446 (I112641,I562759);
nor I_6447 (I112658,I112641,I562774);
and I_6448 (I112675,I112658,I562771);
or I_6449 (I112692,I112675,I562753);
DFFARX1 I_6450 (I112692,I3035,I112251,I112718,);
nand I_6451 (I112726,I112718,I112384);
nor I_6452 (I112228,I112726,I112534);
nor I_6453 (I112222,I112718,I112350);
DFFARX1 I_6454 (I112718,I3035,I112251,I112780,);
not I_6455 (I112788,I112780);
nor I_6456 (I112237,I112788,I112500);
not I_6457 (I112846,I3042);
DFFARX1 I_6458 (I520013,I3035,I112846,I112872,);
DFFARX1 I_6459 (I112872,I3035,I112846,I112889,);
not I_6460 (I112838,I112889);
not I_6461 (I112911,I112872);
DFFARX1 I_6462 (I520022,I3035,I112846,I112937,);
not I_6463 (I112945,I112937);
and I_6464 (I112962,I112911,I520010);
not I_6465 (I112979,I520001);
nand I_6466 (I112996,I112979,I520010);
not I_6467 (I113013,I520007);
nor I_6468 (I113030,I113013,I520025);
nand I_6469 (I113047,I113030,I519998);
nor I_6470 (I113064,I113047,I112996);
DFFARX1 I_6471 (I113064,I3035,I112846,I112814,);
not I_6472 (I113095,I113047);
not I_6473 (I113112,I520025);
nand I_6474 (I113129,I113112,I520010);
nor I_6475 (I113146,I520025,I520001);
nand I_6476 (I112826,I112962,I113146);
nand I_6477 (I112820,I112911,I520025);
nand I_6478 (I113191,I113013,I520004);
DFFARX1 I_6479 (I113191,I3035,I112846,I112835,);
DFFARX1 I_6480 (I113191,I3035,I112846,I112829,);
not I_6481 (I113236,I520004);
nor I_6482 (I113253,I113236,I520016);
and I_6483 (I113270,I113253,I519998);
or I_6484 (I113287,I113270,I520019);
DFFARX1 I_6485 (I113287,I3035,I112846,I113313,);
nand I_6486 (I113321,I113313,I112979);
nor I_6487 (I112823,I113321,I113129);
nor I_6488 (I112817,I113313,I112945);
DFFARX1 I_6489 (I113313,I3035,I112846,I113375,);
not I_6490 (I113383,I113375);
nor I_6491 (I112832,I113383,I113095);
not I_6492 (I113441,I3042);
DFFARX1 I_6493 (I558829,I3035,I113441,I113467,);
DFFARX1 I_6494 (I113467,I3035,I113441,I113484,);
not I_6495 (I113433,I113484);
not I_6496 (I113506,I113467);
DFFARX1 I_6497 (I558838,I3035,I113441,I113532,);
not I_6498 (I113540,I113532);
and I_6499 (I113557,I113506,I558832);
not I_6500 (I113574,I558826);
nand I_6501 (I113591,I113574,I558832);
not I_6502 (I113608,I558841);
nor I_6503 (I113625,I113608,I558829);
nand I_6504 (I113642,I113625,I558835);
nor I_6505 (I113659,I113642,I113591);
DFFARX1 I_6506 (I113659,I3035,I113441,I113409,);
not I_6507 (I113690,I113642);
not I_6508 (I113707,I558829);
nand I_6509 (I113724,I113707,I558832);
nor I_6510 (I113741,I558829,I558826);
nand I_6511 (I113421,I113557,I113741);
nand I_6512 (I113415,I113506,I558829);
nand I_6513 (I113786,I113608,I558832);
DFFARX1 I_6514 (I113786,I3035,I113441,I113430,);
DFFARX1 I_6515 (I113786,I3035,I113441,I113424,);
not I_6516 (I113831,I558832);
nor I_6517 (I113848,I113831,I558847);
and I_6518 (I113865,I113848,I558844);
or I_6519 (I113882,I113865,I558826);
DFFARX1 I_6520 (I113882,I3035,I113441,I113908,);
nand I_6521 (I113916,I113908,I113574);
nor I_6522 (I113418,I113916,I113724);
nor I_6523 (I113412,I113908,I113540);
DFFARX1 I_6524 (I113908,I3035,I113441,I113970,);
not I_6525 (I113978,I113970);
nor I_6526 (I113427,I113978,I113690);
not I_6527 (I114036,I3042);
DFFARX1 I_6528 (I50501,I3035,I114036,I114062,);
DFFARX1 I_6529 (I114062,I3035,I114036,I114079,);
not I_6530 (I114028,I114079);
not I_6531 (I114101,I114062);
DFFARX1 I_6532 (I50495,I3035,I114036,I114127,);
not I_6533 (I114135,I114127);
and I_6534 (I114152,I114101,I50492);
not I_6535 (I114169,I50513);
nand I_6536 (I114186,I114169,I50492);
not I_6537 (I114203,I50507);
nor I_6538 (I114220,I114203,I50498);
nand I_6539 (I114237,I114220,I50504);
nor I_6540 (I114254,I114237,I114186);
DFFARX1 I_6541 (I114254,I3035,I114036,I114004,);
not I_6542 (I114285,I114237);
not I_6543 (I114302,I50498);
nand I_6544 (I114319,I114302,I50492);
nor I_6545 (I114336,I50498,I50513);
nand I_6546 (I114016,I114152,I114336);
nand I_6547 (I114010,I114101,I50498);
nand I_6548 (I114381,I114203,I50492);
DFFARX1 I_6549 (I114381,I3035,I114036,I114025,);
DFFARX1 I_6550 (I114381,I3035,I114036,I114019,);
not I_6551 (I114426,I50492);
nor I_6552 (I114443,I114426,I50510);
and I_6553 (I114460,I114443,I50516);
or I_6554 (I114477,I114460,I50495);
DFFARX1 I_6555 (I114477,I3035,I114036,I114503,);
nand I_6556 (I114511,I114503,I114169);
nor I_6557 (I114013,I114511,I114319);
nor I_6558 (I114007,I114503,I114135);
DFFARX1 I_6559 (I114503,I3035,I114036,I114565,);
not I_6560 (I114573,I114565);
nor I_6561 (I114022,I114573,I114285);
not I_6562 (I114631,I3042);
DFFARX1 I_6563 (I635292,I3035,I114631,I114657,);
DFFARX1 I_6564 (I114657,I3035,I114631,I114674,);
not I_6565 (I114623,I114674);
not I_6566 (I114696,I114657);
DFFARX1 I_6567 (I635292,I3035,I114631,I114722,);
not I_6568 (I114730,I114722);
and I_6569 (I114747,I114696,I635295);
not I_6570 (I114764,I635307);
nand I_6571 (I114781,I114764,I635295);
not I_6572 (I114798,I635313);
nor I_6573 (I114815,I114798,I635304);
nand I_6574 (I114832,I114815,I635310);
nor I_6575 (I114849,I114832,I114781);
DFFARX1 I_6576 (I114849,I3035,I114631,I114599,);
not I_6577 (I114880,I114832);
not I_6578 (I114897,I635304);
nand I_6579 (I114914,I114897,I635295);
nor I_6580 (I114931,I635304,I635307);
nand I_6581 (I114611,I114747,I114931);
nand I_6582 (I114605,I114696,I635304);
nand I_6583 (I114976,I114798,I635301);
DFFARX1 I_6584 (I114976,I3035,I114631,I114620,);
DFFARX1 I_6585 (I114976,I3035,I114631,I114614,);
not I_6586 (I115021,I635301);
nor I_6587 (I115038,I115021,I635298);
and I_6588 (I115055,I115038,I635316);
or I_6589 (I115072,I115055,I635295);
DFFARX1 I_6590 (I115072,I3035,I114631,I115098,);
nand I_6591 (I115106,I115098,I114764);
nor I_6592 (I114608,I115106,I114914);
nor I_6593 (I114602,I115098,I114730);
DFFARX1 I_6594 (I115098,I3035,I114631,I115160,);
not I_6595 (I115168,I115160);
nor I_6596 (I114617,I115168,I114880);
not I_6597 (I115226,I3042);
DFFARX1 I_6598 (I623732,I3035,I115226,I115252,);
DFFARX1 I_6599 (I115252,I3035,I115226,I115269,);
not I_6600 (I115218,I115269);
not I_6601 (I115291,I115252);
DFFARX1 I_6602 (I623732,I3035,I115226,I115317,);
not I_6603 (I115325,I115317);
and I_6604 (I115342,I115291,I623735);
not I_6605 (I115359,I623747);
nand I_6606 (I115376,I115359,I623735);
not I_6607 (I115393,I623753);
nor I_6608 (I115410,I115393,I623744);
nand I_6609 (I115427,I115410,I623750);
nor I_6610 (I115444,I115427,I115376);
DFFARX1 I_6611 (I115444,I3035,I115226,I115194,);
not I_6612 (I115475,I115427);
not I_6613 (I115492,I623744);
nand I_6614 (I115509,I115492,I623735);
nor I_6615 (I115526,I623744,I623747);
nand I_6616 (I115206,I115342,I115526);
nand I_6617 (I115200,I115291,I623744);
nand I_6618 (I115571,I115393,I623741);
DFFARX1 I_6619 (I115571,I3035,I115226,I115215,);
DFFARX1 I_6620 (I115571,I3035,I115226,I115209,);
not I_6621 (I115616,I623741);
nor I_6622 (I115633,I115616,I623738);
and I_6623 (I115650,I115633,I623756);
or I_6624 (I115667,I115650,I623735);
DFFARX1 I_6625 (I115667,I3035,I115226,I115693,);
nand I_6626 (I115701,I115693,I115359);
nor I_6627 (I115203,I115701,I115509);
nor I_6628 (I115197,I115693,I115325);
DFFARX1 I_6629 (I115693,I3035,I115226,I115755,);
not I_6630 (I115763,I115755);
nor I_6631 (I115212,I115763,I115475);
not I_6632 (I115821,I3042);
DFFARX1 I_6633 (I426657,I3035,I115821,I115847,);
DFFARX1 I_6634 (I115847,I3035,I115821,I115864,);
not I_6635 (I115813,I115864);
not I_6636 (I115886,I115847);
DFFARX1 I_6637 (I426651,I3035,I115821,I115912,);
not I_6638 (I115920,I115912);
and I_6639 (I115937,I115886,I426669);
not I_6640 (I115954,I426657);
nand I_6641 (I115971,I115954,I426669);
not I_6642 (I115988,I426651);
nor I_6643 (I116005,I115988,I426663);
nand I_6644 (I116022,I116005,I426654);
nor I_6645 (I116039,I116022,I115971);
DFFARX1 I_6646 (I116039,I3035,I115821,I115789,);
not I_6647 (I116070,I116022);
not I_6648 (I116087,I426663);
nand I_6649 (I116104,I116087,I426669);
nor I_6650 (I116121,I426663,I426657);
nand I_6651 (I115801,I115937,I116121);
nand I_6652 (I115795,I115886,I426663);
nand I_6653 (I116166,I115988,I426666);
DFFARX1 I_6654 (I116166,I3035,I115821,I115810,);
DFFARX1 I_6655 (I116166,I3035,I115821,I115804,);
not I_6656 (I116211,I426666);
nor I_6657 (I116228,I116211,I426672);
and I_6658 (I116245,I116228,I426654);
or I_6659 (I116262,I116245,I426660);
DFFARX1 I_6660 (I116262,I3035,I115821,I116288,);
nand I_6661 (I116296,I116288,I115954);
nor I_6662 (I115798,I116296,I116104);
nor I_6663 (I115792,I116288,I115920);
DFFARX1 I_6664 (I116288,I3035,I115821,I116350,);
not I_6665 (I116358,I116350);
nor I_6666 (I115807,I116358,I116070);
not I_6667 (I116416,I3042);
DFFARX1 I_6668 (I327913,I3035,I116416,I116442,);
DFFARX1 I_6669 (I116442,I3035,I116416,I116459,);
not I_6670 (I116408,I116459);
not I_6671 (I116481,I116442);
DFFARX1 I_6672 (I327904,I3035,I116416,I116507,);
not I_6673 (I116515,I116507);
and I_6674 (I116532,I116481,I327922);
not I_6675 (I116549,I327919);
nand I_6676 (I116566,I116549,I327922);
not I_6677 (I116583,I327898);
nor I_6678 (I116600,I116583,I327901);
nand I_6679 (I116617,I116600,I327910);
nor I_6680 (I116634,I116617,I116566);
DFFARX1 I_6681 (I116634,I3035,I116416,I116384,);
not I_6682 (I116665,I116617);
not I_6683 (I116682,I327901);
nand I_6684 (I116699,I116682,I327922);
nor I_6685 (I116716,I327901,I327919);
nand I_6686 (I116396,I116532,I116716);
nand I_6687 (I116390,I116481,I327901);
nand I_6688 (I116761,I116583,I327916);
DFFARX1 I_6689 (I116761,I3035,I116416,I116405,);
DFFARX1 I_6690 (I116761,I3035,I116416,I116399,);
not I_6691 (I116806,I327916);
nor I_6692 (I116823,I116806,I327898);
and I_6693 (I116840,I116823,I327907);
or I_6694 (I116857,I116840,I327901);
DFFARX1 I_6695 (I116857,I3035,I116416,I116883,);
nand I_6696 (I116891,I116883,I116549);
nor I_6697 (I116393,I116891,I116699);
nor I_6698 (I116387,I116883,I116515);
DFFARX1 I_6699 (I116883,I3035,I116416,I116945,);
not I_6700 (I116953,I116945);
nor I_6701 (I116402,I116953,I116665);
not I_6702 (I117011,I3042);
DFFARX1 I_6703 (I396692,I3035,I117011,I117037,);
DFFARX1 I_6704 (I117037,I3035,I117011,I117054,);
not I_6705 (I117003,I117054);
not I_6706 (I117076,I117037);
DFFARX1 I_6707 (I396689,I3035,I117011,I117102,);
not I_6708 (I117110,I117102);
and I_6709 (I117127,I117076,I396695);
not I_6710 (I117144,I396680);
nand I_6711 (I117161,I117144,I396695);
not I_6712 (I117178,I396683);
nor I_6713 (I117195,I117178,I396704);
nand I_6714 (I117212,I117195,I396701);
nor I_6715 (I117229,I117212,I117161);
DFFARX1 I_6716 (I117229,I3035,I117011,I116979,);
not I_6717 (I117260,I117212);
not I_6718 (I117277,I396704);
nand I_6719 (I117294,I117277,I396695);
nor I_6720 (I117311,I396704,I396680);
nand I_6721 (I116991,I117127,I117311);
nand I_6722 (I116985,I117076,I396704);
nand I_6723 (I117356,I117178,I396680);
DFFARX1 I_6724 (I117356,I3035,I117011,I117000,);
DFFARX1 I_6725 (I117356,I3035,I117011,I116994,);
not I_6726 (I117401,I396680);
nor I_6727 (I117418,I117401,I396686);
and I_6728 (I117435,I117418,I396698);
or I_6729 (I117452,I117435,I396683);
DFFARX1 I_6730 (I117452,I3035,I117011,I117478,);
nand I_6731 (I117486,I117478,I117144);
nor I_6732 (I116988,I117486,I117294);
nor I_6733 (I116982,I117478,I117110);
DFFARX1 I_6734 (I117478,I3035,I117011,I117540,);
not I_6735 (I117548,I117540);
nor I_6736 (I116997,I117548,I117260);
not I_6737 (I117606,I3042);
DFFARX1 I_6738 (I366636,I3035,I117606,I117632,);
DFFARX1 I_6739 (I117632,I3035,I117606,I117649,);
not I_6740 (I117598,I117649);
not I_6741 (I117671,I117632);
DFFARX1 I_6742 (I366633,I3035,I117606,I117697,);
not I_6743 (I117705,I117697);
and I_6744 (I117722,I117671,I366639);
not I_6745 (I117739,I366624);
nand I_6746 (I117756,I117739,I366639);
not I_6747 (I117773,I366627);
nor I_6748 (I117790,I117773,I366648);
nand I_6749 (I117807,I117790,I366645);
nor I_6750 (I117824,I117807,I117756);
DFFARX1 I_6751 (I117824,I3035,I117606,I117574,);
not I_6752 (I117855,I117807);
not I_6753 (I117872,I366648);
nand I_6754 (I117889,I117872,I366639);
nor I_6755 (I117906,I366648,I366624);
nand I_6756 (I117586,I117722,I117906);
nand I_6757 (I117580,I117671,I366648);
nand I_6758 (I117951,I117773,I366624);
DFFARX1 I_6759 (I117951,I3035,I117606,I117595,);
DFFARX1 I_6760 (I117951,I3035,I117606,I117589,);
not I_6761 (I117996,I366624);
nor I_6762 (I118013,I117996,I366630);
and I_6763 (I118030,I118013,I366642);
or I_6764 (I118047,I118030,I366627);
DFFARX1 I_6765 (I118047,I3035,I117606,I118073,);
nand I_6766 (I118081,I118073,I117739);
nor I_6767 (I117583,I118081,I117889);
nor I_6768 (I117577,I118073,I117705);
DFFARX1 I_6769 (I118073,I3035,I117606,I118135,);
not I_6770 (I118143,I118135);
nor I_6771 (I117592,I118143,I117855);
not I_6772 (I118201,I3042);
DFFARX1 I_6773 (I564439,I3035,I118201,I118227,);
DFFARX1 I_6774 (I118227,I3035,I118201,I118244,);
not I_6775 (I118193,I118244);
not I_6776 (I118266,I118227);
DFFARX1 I_6777 (I564448,I3035,I118201,I118292,);
not I_6778 (I118300,I118292);
and I_6779 (I118317,I118266,I564442);
not I_6780 (I118334,I564436);
nand I_6781 (I118351,I118334,I564442);
not I_6782 (I118368,I564451);
nor I_6783 (I118385,I118368,I564439);
nand I_6784 (I118402,I118385,I564445);
nor I_6785 (I118419,I118402,I118351);
DFFARX1 I_6786 (I118419,I3035,I118201,I118169,);
not I_6787 (I118450,I118402);
not I_6788 (I118467,I564439);
nand I_6789 (I118484,I118467,I564442);
nor I_6790 (I118501,I564439,I564436);
nand I_6791 (I118181,I118317,I118501);
nand I_6792 (I118175,I118266,I564439);
nand I_6793 (I118546,I118368,I564442);
DFFARX1 I_6794 (I118546,I3035,I118201,I118190,);
DFFARX1 I_6795 (I118546,I3035,I118201,I118184,);
not I_6796 (I118591,I564442);
nor I_6797 (I118608,I118591,I564457);
and I_6798 (I118625,I118608,I564454);
or I_6799 (I118642,I118625,I564436);
DFFARX1 I_6800 (I118642,I3035,I118201,I118668,);
nand I_6801 (I118676,I118668,I118334);
nor I_6802 (I118178,I118676,I118484);
nor I_6803 (I118172,I118668,I118300);
DFFARX1 I_6804 (I118668,I3035,I118201,I118730,);
not I_6805 (I118738,I118730);
nor I_6806 (I118187,I118738,I118450);
not I_6807 (I118796,I3042);
DFFARX1 I_6808 (I236445,I3035,I118796,I118822,);
DFFARX1 I_6809 (I118822,I3035,I118796,I118839,);
not I_6810 (I118788,I118839);
not I_6811 (I118861,I118822);
DFFARX1 I_6812 (I236433,I3035,I118796,I118887,);
not I_6813 (I118895,I118887);
and I_6814 (I118912,I118861,I236442);
not I_6815 (I118929,I236439);
nand I_6816 (I118946,I118929,I236442);
not I_6817 (I118963,I236430);
nor I_6818 (I118980,I118963,I236436);
nand I_6819 (I118997,I118980,I236421);
nor I_6820 (I119014,I118997,I118946);
DFFARX1 I_6821 (I119014,I3035,I118796,I118764,);
not I_6822 (I119045,I118997);
not I_6823 (I119062,I236436);
nand I_6824 (I119079,I119062,I236442);
nor I_6825 (I119096,I236436,I236439);
nand I_6826 (I118776,I118912,I119096);
nand I_6827 (I118770,I118861,I236436);
nand I_6828 (I119141,I118963,I236421);
DFFARX1 I_6829 (I119141,I3035,I118796,I118785,);
DFFARX1 I_6830 (I119141,I3035,I118796,I118779,);
not I_6831 (I119186,I236421);
nor I_6832 (I119203,I119186,I236427);
and I_6833 (I119220,I119203,I236424);
or I_6834 (I119237,I119220,I236448);
DFFARX1 I_6835 (I119237,I3035,I118796,I119263,);
nand I_6836 (I119271,I119263,I118929);
nor I_6837 (I118773,I119271,I119079);
nor I_6838 (I118767,I119263,I118895);
DFFARX1 I_6839 (I119263,I3035,I118796,I119325,);
not I_6840 (I119333,I119325);
nor I_6841 (I118782,I119333,I119045);
not I_6842 (I119391,I3042);
DFFARX1 I_6843 (I583272,I3035,I119391,I119417,);
DFFARX1 I_6844 (I119417,I3035,I119391,I119434,);
not I_6845 (I119383,I119434);
not I_6846 (I119456,I119417);
DFFARX1 I_6847 (I583272,I3035,I119391,I119482,);
not I_6848 (I119490,I119482);
and I_6849 (I119507,I119456,I583275);
not I_6850 (I119524,I583287);
nand I_6851 (I119541,I119524,I583275);
not I_6852 (I119558,I583293);
nor I_6853 (I119575,I119558,I583284);
nand I_6854 (I119592,I119575,I583290);
nor I_6855 (I119609,I119592,I119541);
DFFARX1 I_6856 (I119609,I3035,I119391,I119359,);
not I_6857 (I119640,I119592);
not I_6858 (I119657,I583284);
nand I_6859 (I119674,I119657,I583275);
nor I_6860 (I119691,I583284,I583287);
nand I_6861 (I119371,I119507,I119691);
nand I_6862 (I119365,I119456,I583284);
nand I_6863 (I119736,I119558,I583281);
DFFARX1 I_6864 (I119736,I3035,I119391,I119380,);
DFFARX1 I_6865 (I119736,I3035,I119391,I119374,);
not I_6866 (I119781,I583281);
nor I_6867 (I119798,I119781,I583278);
and I_6868 (I119815,I119798,I583296);
or I_6869 (I119832,I119815,I583275);
DFFARX1 I_6870 (I119832,I3035,I119391,I119858,);
nand I_6871 (I119866,I119858,I119524);
nor I_6872 (I119368,I119866,I119674);
nor I_6873 (I119362,I119858,I119490);
DFFARX1 I_6874 (I119858,I3035,I119391,I119920,);
not I_6875 (I119928,I119920);
nor I_6876 (I119377,I119928,I119640);
not I_6877 (I119986,I3042);
DFFARX1 I_6878 (I384554,I3035,I119986,I120012,);
DFFARX1 I_6879 (I120012,I3035,I119986,I120029,);
not I_6880 (I119978,I120029);
not I_6881 (I120051,I120012);
DFFARX1 I_6882 (I384551,I3035,I119986,I120077,);
not I_6883 (I120085,I120077);
and I_6884 (I120102,I120051,I384557);
not I_6885 (I120119,I384542);
nand I_6886 (I120136,I120119,I384557);
not I_6887 (I120153,I384545);
nor I_6888 (I120170,I120153,I384566);
nand I_6889 (I120187,I120170,I384563);
nor I_6890 (I120204,I120187,I120136);
DFFARX1 I_6891 (I120204,I3035,I119986,I119954,);
not I_6892 (I120235,I120187);
not I_6893 (I120252,I384566);
nand I_6894 (I120269,I120252,I384557);
nor I_6895 (I120286,I384566,I384542);
nand I_6896 (I119966,I120102,I120286);
nand I_6897 (I119960,I120051,I384566);
nand I_6898 (I120331,I120153,I384542);
DFFARX1 I_6899 (I120331,I3035,I119986,I119975,);
DFFARX1 I_6900 (I120331,I3035,I119986,I119969,);
not I_6901 (I120376,I384542);
nor I_6902 (I120393,I120376,I384548);
and I_6903 (I120410,I120393,I384560);
or I_6904 (I120427,I120410,I384545);
DFFARX1 I_6905 (I120427,I3035,I119986,I120453,);
nand I_6906 (I120461,I120453,I120119);
nor I_6907 (I119963,I120461,I120269);
nor I_6908 (I119957,I120453,I120085);
DFFARX1 I_6909 (I120453,I3035,I119986,I120515,);
not I_6910 (I120523,I120515);
nor I_6911 (I119972,I120523,I120235);
not I_6912 (I120581,I3042);
DFFARX1 I_6913 (I629512,I3035,I120581,I120607,);
DFFARX1 I_6914 (I120607,I3035,I120581,I120624,);
not I_6915 (I120573,I120624);
not I_6916 (I120646,I120607);
DFFARX1 I_6917 (I629512,I3035,I120581,I120672,);
not I_6918 (I120680,I120672);
and I_6919 (I120697,I120646,I629515);
not I_6920 (I120714,I629527);
nand I_6921 (I120731,I120714,I629515);
not I_6922 (I120748,I629533);
nor I_6923 (I120765,I120748,I629524);
nand I_6924 (I120782,I120765,I629530);
nor I_6925 (I120799,I120782,I120731);
DFFARX1 I_6926 (I120799,I3035,I120581,I120549,);
not I_6927 (I120830,I120782);
not I_6928 (I120847,I629524);
nand I_6929 (I120864,I120847,I629515);
nor I_6930 (I120881,I629524,I629527);
nand I_6931 (I120561,I120697,I120881);
nand I_6932 (I120555,I120646,I629524);
nand I_6933 (I120926,I120748,I629521);
DFFARX1 I_6934 (I120926,I3035,I120581,I120570,);
DFFARX1 I_6935 (I120926,I3035,I120581,I120564,);
not I_6936 (I120971,I629521);
nor I_6937 (I120988,I120971,I629518);
and I_6938 (I121005,I120988,I629536);
or I_6939 (I121022,I121005,I629515);
DFFARX1 I_6940 (I121022,I3035,I120581,I121048,);
nand I_6941 (I121056,I121048,I120714);
nor I_6942 (I120558,I121056,I120864);
nor I_6943 (I120552,I121048,I120680);
DFFARX1 I_6944 (I121048,I3035,I120581,I121110,);
not I_6945 (I121118,I121110);
nor I_6946 (I120567,I121118,I120830);
not I_6947 (I121176,I3042);
DFFARX1 I_6948 (I45231,I3035,I121176,I121202,);
DFFARX1 I_6949 (I121202,I3035,I121176,I121219,);
not I_6950 (I121168,I121219);
not I_6951 (I121241,I121202);
DFFARX1 I_6952 (I45225,I3035,I121176,I121267,);
not I_6953 (I121275,I121267);
and I_6954 (I121292,I121241,I45222);
not I_6955 (I121309,I45243);
nand I_6956 (I121326,I121309,I45222);
not I_6957 (I121343,I45237);
nor I_6958 (I121360,I121343,I45228);
nand I_6959 (I121377,I121360,I45234);
nor I_6960 (I121394,I121377,I121326);
DFFARX1 I_6961 (I121394,I3035,I121176,I121144,);
not I_6962 (I121425,I121377);
not I_6963 (I121442,I45228);
nand I_6964 (I121459,I121442,I45222);
nor I_6965 (I121476,I45228,I45243);
nand I_6966 (I121156,I121292,I121476);
nand I_6967 (I121150,I121241,I45228);
nand I_6968 (I121521,I121343,I45222);
DFFARX1 I_6969 (I121521,I3035,I121176,I121165,);
DFFARX1 I_6970 (I121521,I3035,I121176,I121159,);
not I_6971 (I121566,I45222);
nor I_6972 (I121583,I121566,I45240);
and I_6973 (I121600,I121583,I45246);
or I_6974 (I121617,I121600,I45225);
DFFARX1 I_6975 (I121617,I3035,I121176,I121643,);
nand I_6976 (I121651,I121643,I121309);
nor I_6977 (I121153,I121651,I121459);
nor I_6978 (I121147,I121643,I121275);
DFFARX1 I_6979 (I121643,I3035,I121176,I121705,);
not I_6980 (I121713,I121705);
nor I_6981 (I121162,I121713,I121425);
not I_6982 (I121771,I3042);
DFFARX1 I_6983 (I726399,I3035,I121771,I121797,);
DFFARX1 I_6984 (I121797,I3035,I121771,I121814,);
not I_6985 (I121763,I121814);
not I_6986 (I121836,I121797);
DFFARX1 I_6987 (I726390,I3035,I121771,I121862,);
not I_6988 (I121870,I121862);
and I_6989 (I121887,I121836,I726384);
not I_6990 (I121904,I726378);
nand I_6991 (I121921,I121904,I726384);
not I_6992 (I121938,I726405);
nor I_6993 (I121955,I121938,I726378);
nand I_6994 (I121972,I121955,I726402);
nor I_6995 (I121989,I121972,I121921);
DFFARX1 I_6996 (I121989,I3035,I121771,I121739,);
not I_6997 (I122020,I121972);
not I_6998 (I122037,I726378);
nand I_6999 (I122054,I122037,I726384);
nor I_7000 (I122071,I726378,I726378);
nand I_7001 (I121751,I121887,I122071);
nand I_7002 (I121745,I121836,I726378);
nand I_7003 (I122116,I121938,I726387);
DFFARX1 I_7004 (I122116,I3035,I121771,I121760,);
DFFARX1 I_7005 (I122116,I3035,I121771,I121754,);
not I_7006 (I122161,I726387);
nor I_7007 (I122178,I122161,I726393);
and I_7008 (I122195,I122178,I726396);
or I_7009 (I122212,I122195,I726381);
DFFARX1 I_7010 (I122212,I3035,I121771,I122238,);
nand I_7011 (I122246,I122238,I121904);
nor I_7012 (I121748,I122246,I122054);
nor I_7013 (I121742,I122238,I121870);
DFFARX1 I_7014 (I122238,I3035,I121771,I122300,);
not I_7015 (I122308,I122300);
nor I_7016 (I121757,I122308,I122020);
not I_7017 (I122366,I3042);
DFFARX1 I_7018 (I12045,I3035,I122366,I122392,);
DFFARX1 I_7019 (I122392,I3035,I122366,I122409,);
not I_7020 (I122358,I122409);
not I_7021 (I122431,I122392);
DFFARX1 I_7022 (I12021,I3035,I122366,I122457,);
not I_7023 (I122465,I122457);
and I_7024 (I122482,I122431,I12036);
not I_7025 (I122499,I12024);
nand I_7026 (I122516,I122499,I12036);
not I_7027 (I122533,I12027);
nor I_7028 (I122550,I122533,I12039);
nand I_7029 (I122567,I122550,I12030);
nor I_7030 (I122584,I122567,I122516);
DFFARX1 I_7031 (I122584,I3035,I122366,I122334,);
not I_7032 (I122615,I122567);
not I_7033 (I122632,I12039);
nand I_7034 (I122649,I122632,I12036);
nor I_7035 (I122666,I12039,I12024);
nand I_7036 (I122346,I122482,I122666);
nand I_7037 (I122340,I122431,I12039);
nand I_7038 (I122711,I122533,I12033);
DFFARX1 I_7039 (I122711,I3035,I122366,I122355,);
DFFARX1 I_7040 (I122711,I3035,I122366,I122349,);
not I_7041 (I122756,I12033);
nor I_7042 (I122773,I122756,I12024);
and I_7043 (I122790,I122773,I12021);
or I_7044 (I122807,I122790,I12042);
DFFARX1 I_7045 (I122807,I3035,I122366,I122833,);
nand I_7046 (I122841,I122833,I122499);
nor I_7047 (I122343,I122841,I122649);
nor I_7048 (I122337,I122833,I122465);
DFFARX1 I_7049 (I122833,I3035,I122366,I122895,);
not I_7050 (I122903,I122895);
nor I_7051 (I122352,I122903,I122615);
not I_7052 (I122961,I3042);
DFFARX1 I_7053 (I2964,I3035,I122961,I122987,);
DFFARX1 I_7054 (I122987,I3035,I122961,I123004,);
not I_7055 (I122953,I123004);
not I_7056 (I123026,I122987);
DFFARX1 I_7057 (I2860,I3035,I122961,I123052,);
not I_7058 (I123060,I123052);
and I_7059 (I123077,I123026,I1756);
not I_7060 (I123094,I1596);
nand I_7061 (I123111,I123094,I1756);
not I_7062 (I123128,I1660);
nor I_7063 (I123145,I123128,I1388);
nand I_7064 (I123162,I123145,I1948);
nor I_7065 (I123179,I123162,I123111);
DFFARX1 I_7066 (I123179,I3035,I122961,I122929,);
not I_7067 (I123210,I123162);
not I_7068 (I123227,I1388);
nand I_7069 (I123244,I123227,I1756);
nor I_7070 (I123261,I1388,I1596);
nand I_7071 (I122941,I123077,I123261);
nand I_7072 (I122935,I123026,I1388);
nand I_7073 (I123306,I123128,I1980);
DFFARX1 I_7074 (I123306,I3035,I122961,I122950,);
DFFARX1 I_7075 (I123306,I3035,I122961,I122944,);
not I_7076 (I123351,I1980);
nor I_7077 (I123368,I123351,I2268);
and I_7078 (I123385,I123368,I1804);
or I_7079 (I123402,I123385,I2412);
DFFARX1 I_7080 (I123402,I3035,I122961,I123428,);
nand I_7081 (I123436,I123428,I123094);
nor I_7082 (I122938,I123436,I123244);
nor I_7083 (I122932,I123428,I123060);
DFFARX1 I_7084 (I123428,I3035,I122961,I123490,);
not I_7085 (I123498,I123490);
nor I_7086 (I122947,I123498,I123210);
not I_7087 (I123556,I3042);
DFFARX1 I_7088 (I548170,I3035,I123556,I123582,);
DFFARX1 I_7089 (I123582,I3035,I123556,I123599,);
not I_7090 (I123548,I123599);
not I_7091 (I123621,I123582);
DFFARX1 I_7092 (I548179,I3035,I123556,I123647,);
not I_7093 (I123655,I123647);
and I_7094 (I123672,I123621,I548173);
not I_7095 (I123689,I548167);
nand I_7096 (I123706,I123689,I548173);
not I_7097 (I123723,I548182);
nor I_7098 (I123740,I123723,I548170);
nand I_7099 (I123757,I123740,I548176);
nor I_7100 (I123774,I123757,I123706);
DFFARX1 I_7101 (I123774,I3035,I123556,I123524,);
not I_7102 (I123805,I123757);
not I_7103 (I123822,I548170);
nand I_7104 (I123839,I123822,I548173);
nor I_7105 (I123856,I548170,I548167);
nand I_7106 (I123536,I123672,I123856);
nand I_7107 (I123530,I123621,I548170);
nand I_7108 (I123901,I123723,I548173);
DFFARX1 I_7109 (I123901,I3035,I123556,I123545,);
DFFARX1 I_7110 (I123901,I3035,I123556,I123539,);
not I_7111 (I123946,I548173);
nor I_7112 (I123963,I123946,I548188);
and I_7113 (I123980,I123963,I548185);
or I_7114 (I123997,I123980,I548167);
DFFARX1 I_7115 (I123997,I3035,I123556,I124023,);
nand I_7116 (I124031,I124023,I123689);
nor I_7117 (I123533,I124031,I123839);
nor I_7118 (I123527,I124023,I123655);
DFFARX1 I_7119 (I124023,I3035,I123556,I124085,);
not I_7120 (I124093,I124085);
nor I_7121 (I123542,I124093,I123805);
not I_7122 (I124151,I3042);
DFFARX1 I_7123 (I317509,I3035,I124151,I124177,);
DFFARX1 I_7124 (I124177,I3035,I124151,I124194,);
not I_7125 (I124143,I124194);
not I_7126 (I124216,I124177);
DFFARX1 I_7127 (I317500,I3035,I124151,I124242,);
not I_7128 (I124250,I124242);
and I_7129 (I124267,I124216,I317518);
not I_7130 (I124284,I317515);
nand I_7131 (I124301,I124284,I317518);
not I_7132 (I124318,I317494);
nor I_7133 (I124335,I124318,I317497);
nand I_7134 (I124352,I124335,I317506);
nor I_7135 (I124369,I124352,I124301);
DFFARX1 I_7136 (I124369,I3035,I124151,I124119,);
not I_7137 (I124400,I124352);
not I_7138 (I124417,I317497);
nand I_7139 (I124434,I124417,I317518);
nor I_7140 (I124451,I317497,I317515);
nand I_7141 (I124131,I124267,I124451);
nand I_7142 (I124125,I124216,I317497);
nand I_7143 (I124496,I124318,I317512);
DFFARX1 I_7144 (I124496,I3035,I124151,I124140,);
DFFARX1 I_7145 (I124496,I3035,I124151,I124134,);
not I_7146 (I124541,I317512);
nor I_7147 (I124558,I124541,I317494);
and I_7148 (I124575,I124558,I317503);
or I_7149 (I124592,I124575,I317497);
DFFARX1 I_7150 (I124592,I3035,I124151,I124618,);
nand I_7151 (I124626,I124618,I124284);
nor I_7152 (I124128,I124626,I124434);
nor I_7153 (I124122,I124618,I124250);
DFFARX1 I_7154 (I124618,I3035,I124151,I124680,);
not I_7155 (I124688,I124680);
nor I_7156 (I124137,I124688,I124400);
not I_7157 (I124746,I3042);
DFFARX1 I_7158 (I618530,I3035,I124746,I124772,);
DFFARX1 I_7159 (I124772,I3035,I124746,I124789,);
not I_7160 (I124738,I124789);
not I_7161 (I124811,I124772);
DFFARX1 I_7162 (I618530,I3035,I124746,I124837,);
not I_7163 (I124845,I124837);
and I_7164 (I124862,I124811,I618533);
not I_7165 (I124879,I618545);
nand I_7166 (I124896,I124879,I618533);
not I_7167 (I124913,I618551);
nor I_7168 (I124930,I124913,I618542);
nand I_7169 (I124947,I124930,I618548);
nor I_7170 (I124964,I124947,I124896);
DFFARX1 I_7171 (I124964,I3035,I124746,I124714,);
not I_7172 (I124995,I124947);
not I_7173 (I125012,I618542);
nand I_7174 (I125029,I125012,I618533);
nor I_7175 (I125046,I618542,I618545);
nand I_7176 (I124726,I124862,I125046);
nand I_7177 (I124720,I124811,I618542);
nand I_7178 (I125091,I124913,I618539);
DFFARX1 I_7179 (I125091,I3035,I124746,I124735,);
DFFARX1 I_7180 (I125091,I3035,I124746,I124729,);
not I_7181 (I125136,I618539);
nor I_7182 (I125153,I125136,I618536);
and I_7183 (I125170,I125153,I618554);
or I_7184 (I125187,I125170,I618533);
DFFARX1 I_7185 (I125187,I3035,I124746,I125213,);
nand I_7186 (I125221,I125213,I124879);
nor I_7187 (I124723,I125221,I125029);
nor I_7188 (I124717,I125213,I124845);
DFFARX1 I_7189 (I125213,I3035,I124746,I125275,);
not I_7190 (I125283,I125275);
nor I_7191 (I124732,I125283,I124995);
not I_7192 (I125341,I3042);
DFFARX1 I_7193 (I349874,I3035,I125341,I125367,);
DFFARX1 I_7194 (I125367,I3035,I125341,I125384,);
not I_7195 (I125333,I125384);
not I_7196 (I125406,I125367);
DFFARX1 I_7197 (I349871,I3035,I125341,I125432,);
not I_7198 (I125440,I125432);
and I_7199 (I125457,I125406,I349877);
not I_7200 (I125474,I349862);
nand I_7201 (I125491,I125474,I349877);
not I_7202 (I125508,I349865);
nor I_7203 (I125525,I125508,I349886);
nand I_7204 (I125542,I125525,I349883);
nor I_7205 (I125559,I125542,I125491);
DFFARX1 I_7206 (I125559,I3035,I125341,I125309,);
not I_7207 (I125590,I125542);
not I_7208 (I125607,I349886);
nand I_7209 (I125624,I125607,I349877);
nor I_7210 (I125641,I349886,I349862);
nand I_7211 (I125321,I125457,I125641);
nand I_7212 (I125315,I125406,I349886);
nand I_7213 (I125686,I125508,I349862);
DFFARX1 I_7214 (I125686,I3035,I125341,I125330,);
DFFARX1 I_7215 (I125686,I3035,I125341,I125324,);
not I_7216 (I125731,I349862);
nor I_7217 (I125748,I125731,I349868);
and I_7218 (I125765,I125748,I349880);
or I_7219 (I125782,I125765,I349865);
DFFARX1 I_7220 (I125782,I3035,I125341,I125808,);
nand I_7221 (I125816,I125808,I125474);
nor I_7222 (I125318,I125816,I125624);
nor I_7223 (I125312,I125808,I125440);
DFFARX1 I_7224 (I125808,I3035,I125341,I125870,);
not I_7225 (I125878,I125870);
nor I_7226 (I125327,I125878,I125590);
not I_7227 (I125936,I3042);
DFFARX1 I_7228 (I35218,I3035,I125936,I125962,);
DFFARX1 I_7229 (I125962,I3035,I125936,I125979,);
not I_7230 (I125928,I125979);
not I_7231 (I126001,I125962);
DFFARX1 I_7232 (I35212,I3035,I125936,I126027,);
not I_7233 (I126035,I126027);
and I_7234 (I126052,I126001,I35209);
not I_7235 (I126069,I35230);
nand I_7236 (I126086,I126069,I35209);
not I_7237 (I126103,I35224);
nor I_7238 (I126120,I126103,I35215);
nand I_7239 (I126137,I126120,I35221);
nor I_7240 (I126154,I126137,I126086);
DFFARX1 I_7241 (I126154,I3035,I125936,I125904,);
not I_7242 (I126185,I126137);
not I_7243 (I126202,I35215);
nand I_7244 (I126219,I126202,I35209);
nor I_7245 (I126236,I35215,I35230);
nand I_7246 (I125916,I126052,I126236);
nand I_7247 (I125910,I126001,I35215);
nand I_7248 (I126281,I126103,I35209);
DFFARX1 I_7249 (I126281,I3035,I125936,I125925,);
DFFARX1 I_7250 (I126281,I3035,I125936,I125919,);
not I_7251 (I126326,I35209);
nor I_7252 (I126343,I126326,I35227);
and I_7253 (I126360,I126343,I35233);
or I_7254 (I126377,I126360,I35212);
DFFARX1 I_7255 (I126377,I3035,I125936,I126403,);
nand I_7256 (I126411,I126403,I126069);
nor I_7257 (I125913,I126411,I126219);
nor I_7258 (I125907,I126403,I126035);
DFFARX1 I_7259 (I126403,I3035,I125936,I126465,);
not I_7260 (I126473,I126465);
nor I_7261 (I125922,I126473,I126185);
not I_7262 (I126531,I3042);
DFFARX1 I_7263 (I402472,I3035,I126531,I126557,);
DFFARX1 I_7264 (I126557,I3035,I126531,I126574,);
not I_7265 (I126523,I126574);
not I_7266 (I126596,I126557);
DFFARX1 I_7267 (I402469,I3035,I126531,I126622,);
not I_7268 (I126630,I126622);
and I_7269 (I126647,I126596,I402475);
not I_7270 (I126664,I402460);
nand I_7271 (I126681,I126664,I402475);
not I_7272 (I126698,I402463);
nor I_7273 (I126715,I126698,I402484);
nand I_7274 (I126732,I126715,I402481);
nor I_7275 (I126749,I126732,I126681);
DFFARX1 I_7276 (I126749,I3035,I126531,I126499,);
not I_7277 (I126780,I126732);
not I_7278 (I126797,I402484);
nand I_7279 (I126814,I126797,I402475);
nor I_7280 (I126831,I402484,I402460);
nand I_7281 (I126511,I126647,I126831);
nand I_7282 (I126505,I126596,I402484);
nand I_7283 (I126876,I126698,I402460);
DFFARX1 I_7284 (I126876,I3035,I126531,I126520,);
DFFARX1 I_7285 (I126876,I3035,I126531,I126514,);
not I_7286 (I126921,I402460);
nor I_7287 (I126938,I126921,I402466);
and I_7288 (I126955,I126938,I402478);
or I_7289 (I126972,I126955,I402463);
DFFARX1 I_7290 (I126972,I3035,I126531,I126998,);
nand I_7291 (I127006,I126998,I126664);
nor I_7292 (I126508,I127006,I126814);
nor I_7293 (I126502,I126998,I126630);
DFFARX1 I_7294 (I126998,I3035,I126531,I127060,);
not I_7295 (I127068,I127060);
nor I_7296 (I126517,I127068,I126780);
not I_7297 (I127126,I3042);
DFFARX1 I_7298 (I367214,I3035,I127126,I127152,);
DFFARX1 I_7299 (I127152,I3035,I127126,I127169,);
not I_7300 (I127118,I127169);
not I_7301 (I127191,I127152);
DFFARX1 I_7302 (I367211,I3035,I127126,I127217,);
not I_7303 (I127225,I127217);
and I_7304 (I127242,I127191,I367217);
not I_7305 (I127259,I367202);
nand I_7306 (I127276,I127259,I367217);
not I_7307 (I127293,I367205);
nor I_7308 (I127310,I127293,I367226);
nand I_7309 (I127327,I127310,I367223);
nor I_7310 (I127344,I127327,I127276);
DFFARX1 I_7311 (I127344,I3035,I127126,I127094,);
not I_7312 (I127375,I127327);
not I_7313 (I127392,I367226);
nand I_7314 (I127409,I127392,I367217);
nor I_7315 (I127426,I367226,I367202);
nand I_7316 (I127106,I127242,I127426);
nand I_7317 (I127100,I127191,I367226);
nand I_7318 (I127471,I127293,I367202);
DFFARX1 I_7319 (I127471,I3035,I127126,I127115,);
DFFARX1 I_7320 (I127471,I3035,I127126,I127109,);
not I_7321 (I127516,I367202);
nor I_7322 (I127533,I127516,I367208);
and I_7323 (I127550,I127533,I367220);
or I_7324 (I127567,I127550,I367205);
DFFARX1 I_7325 (I127567,I3035,I127126,I127593,);
nand I_7326 (I127601,I127593,I127259);
nor I_7327 (I127103,I127601,I127409);
nor I_7328 (I127097,I127593,I127225);
DFFARX1 I_7329 (I127593,I3035,I127126,I127655,);
not I_7330 (I127663,I127655);
nor I_7331 (I127112,I127663,I127375);
not I_7332 (I127721,I3042);
DFFARX1 I_7333 (I227768,I3035,I127721,I127747,);
DFFARX1 I_7334 (I127747,I3035,I127721,I127764,);
not I_7335 (I127713,I127764);
not I_7336 (I127786,I127747);
DFFARX1 I_7337 (I227783,I3035,I127721,I127812,);
not I_7338 (I127820,I127812);
and I_7339 (I127837,I127786,I227780);
not I_7340 (I127854,I227768);
nand I_7341 (I127871,I127854,I227780);
not I_7342 (I127888,I227777);
nor I_7343 (I127905,I127888,I227792);
nand I_7344 (I127922,I127905,I227789);
nor I_7345 (I127939,I127922,I127871);
DFFARX1 I_7346 (I127939,I3035,I127721,I127689,);
not I_7347 (I127970,I127922);
not I_7348 (I127987,I227792);
nand I_7349 (I128004,I127987,I227780);
nor I_7350 (I128021,I227792,I227768);
nand I_7351 (I127701,I127837,I128021);
nand I_7352 (I127695,I127786,I227792);
nand I_7353 (I128066,I127888,I227786);
DFFARX1 I_7354 (I128066,I3035,I127721,I127710,);
DFFARX1 I_7355 (I128066,I3035,I127721,I127704,);
not I_7356 (I128111,I227786);
nor I_7357 (I128128,I128111,I227774);
and I_7358 (I128145,I128128,I227795);
or I_7359 (I128162,I128145,I227771);
DFFARX1 I_7360 (I128162,I3035,I127721,I128188,);
nand I_7361 (I128196,I128188,I127854);
nor I_7362 (I127698,I128196,I128004);
nor I_7363 (I127692,I128188,I127820);
DFFARX1 I_7364 (I128188,I3035,I127721,I128250,);
not I_7365 (I128258,I128250);
nor I_7366 (I127707,I128258,I127970);
not I_7367 (I128316,I3042);
DFFARX1 I_7368 (I13626,I3035,I128316,I128342,);
DFFARX1 I_7369 (I128342,I3035,I128316,I128359,);
not I_7370 (I128308,I128359);
not I_7371 (I128381,I128342);
DFFARX1 I_7372 (I13602,I3035,I128316,I128407,);
not I_7373 (I128415,I128407);
and I_7374 (I128432,I128381,I13617);
not I_7375 (I128449,I13605);
nand I_7376 (I128466,I128449,I13617);
not I_7377 (I128483,I13608);
nor I_7378 (I128500,I128483,I13620);
nand I_7379 (I128517,I128500,I13611);
nor I_7380 (I128534,I128517,I128466);
DFFARX1 I_7381 (I128534,I3035,I128316,I128284,);
not I_7382 (I128565,I128517);
not I_7383 (I128582,I13620);
nand I_7384 (I128599,I128582,I13617);
nor I_7385 (I128616,I13620,I13605);
nand I_7386 (I128296,I128432,I128616);
nand I_7387 (I128290,I128381,I13620);
nand I_7388 (I128661,I128483,I13614);
DFFARX1 I_7389 (I128661,I3035,I128316,I128305,);
DFFARX1 I_7390 (I128661,I3035,I128316,I128299,);
not I_7391 (I128706,I13614);
nor I_7392 (I128723,I128706,I13605);
and I_7393 (I128740,I128723,I13602);
or I_7394 (I128757,I128740,I13623);
DFFARX1 I_7395 (I128757,I3035,I128316,I128783,);
nand I_7396 (I128791,I128783,I128449);
nor I_7397 (I128293,I128791,I128599);
nor I_7398 (I128287,I128783,I128415);
DFFARX1 I_7399 (I128783,I3035,I128316,I128845,);
not I_7400 (I128853,I128845);
nor I_7401 (I128302,I128853,I128565);
not I_7402 (I128911,I3042);
DFFARX1 I_7403 (I469344,I3035,I128911,I128937,);
DFFARX1 I_7404 (I128937,I3035,I128911,I128954,);
not I_7405 (I128903,I128954);
not I_7406 (I128976,I128937);
DFFARX1 I_7407 (I469338,I3035,I128911,I129002,);
not I_7408 (I129010,I129002);
and I_7409 (I129027,I128976,I469356);
not I_7410 (I129044,I469344);
nand I_7411 (I129061,I129044,I469356);
not I_7412 (I129078,I469338);
nor I_7413 (I129095,I129078,I469350);
nand I_7414 (I129112,I129095,I469341);
nor I_7415 (I129129,I129112,I129061);
DFFARX1 I_7416 (I129129,I3035,I128911,I128879,);
not I_7417 (I129160,I129112);
not I_7418 (I129177,I469350);
nand I_7419 (I129194,I129177,I469356);
nor I_7420 (I129211,I469350,I469344);
nand I_7421 (I128891,I129027,I129211);
nand I_7422 (I128885,I128976,I469350);
nand I_7423 (I129256,I129078,I469353);
DFFARX1 I_7424 (I129256,I3035,I128911,I128900,);
DFFARX1 I_7425 (I129256,I3035,I128911,I128894,);
not I_7426 (I129301,I469353);
nor I_7427 (I129318,I129301,I469359);
and I_7428 (I129335,I129318,I469341);
or I_7429 (I129352,I129335,I469347);
DFFARX1 I_7430 (I129352,I3035,I128911,I129378,);
nand I_7431 (I129386,I129378,I129044);
nor I_7432 (I128888,I129386,I129194);
nor I_7433 (I128882,I129378,I129010);
DFFARX1 I_7434 (I129378,I3035,I128911,I129440,);
not I_7435 (I129448,I129440);
nor I_7436 (I128897,I129448,I129160);
not I_7437 (I129506,I3042);
DFFARX1 I_7438 (I418078,I3035,I129506,I129532,);
DFFARX1 I_7439 (I129532,I3035,I129506,I129549,);
not I_7440 (I129498,I129549);
not I_7441 (I129571,I129532);
DFFARX1 I_7442 (I418075,I3035,I129506,I129597,);
not I_7443 (I129605,I129597);
and I_7444 (I129622,I129571,I418081);
not I_7445 (I129639,I418066);
nand I_7446 (I129656,I129639,I418081);
not I_7447 (I129673,I418069);
nor I_7448 (I129690,I129673,I418090);
nand I_7449 (I129707,I129690,I418087);
nor I_7450 (I129724,I129707,I129656);
DFFARX1 I_7451 (I129724,I3035,I129506,I129474,);
not I_7452 (I129755,I129707);
not I_7453 (I129772,I418090);
nand I_7454 (I129789,I129772,I418081);
nor I_7455 (I129806,I418090,I418066);
nand I_7456 (I129486,I129622,I129806);
nand I_7457 (I129480,I129571,I418090);
nand I_7458 (I129851,I129673,I418066);
DFFARX1 I_7459 (I129851,I3035,I129506,I129495,);
DFFARX1 I_7460 (I129851,I3035,I129506,I129489,);
not I_7461 (I129896,I418066);
nor I_7462 (I129913,I129896,I418072);
and I_7463 (I129930,I129913,I418084);
or I_7464 (I129947,I129930,I418069);
DFFARX1 I_7465 (I129947,I3035,I129506,I129973,);
nand I_7466 (I129981,I129973,I129639);
nor I_7467 (I129483,I129981,I129789);
nor I_7468 (I129477,I129973,I129605);
DFFARX1 I_7469 (I129973,I3035,I129506,I130035,);
not I_7470 (I130043,I130035);
nor I_7471 (I129492,I130043,I129755);
not I_7472 (I130101,I3042);
DFFARX1 I_7473 (I517429,I3035,I130101,I130127,);
DFFARX1 I_7474 (I130127,I3035,I130101,I130144,);
not I_7475 (I130093,I130144);
not I_7476 (I130166,I130127);
DFFARX1 I_7477 (I517438,I3035,I130101,I130192,);
not I_7478 (I130200,I130192);
and I_7479 (I130217,I130166,I517426);
not I_7480 (I130234,I517417);
nand I_7481 (I130251,I130234,I517426);
not I_7482 (I130268,I517423);
nor I_7483 (I130285,I130268,I517441);
nand I_7484 (I130302,I130285,I517414);
nor I_7485 (I130319,I130302,I130251);
DFFARX1 I_7486 (I130319,I3035,I130101,I130069,);
not I_7487 (I130350,I130302);
not I_7488 (I130367,I517441);
nand I_7489 (I130384,I130367,I517426);
nor I_7490 (I130401,I517441,I517417);
nand I_7491 (I130081,I130217,I130401);
nand I_7492 (I130075,I130166,I517441);
nand I_7493 (I130446,I130268,I517420);
DFFARX1 I_7494 (I130446,I3035,I130101,I130090,);
DFFARX1 I_7495 (I130446,I3035,I130101,I130084,);
not I_7496 (I130491,I517420);
nor I_7497 (I130508,I130491,I517432);
and I_7498 (I130525,I130508,I517414);
or I_7499 (I130542,I130525,I517435);
DFFARX1 I_7500 (I130542,I3035,I130101,I130568,);
nand I_7501 (I130576,I130568,I130234);
nor I_7502 (I130078,I130576,I130384);
nor I_7503 (I130072,I130568,I130200);
DFFARX1 I_7504 (I130568,I3035,I130101,I130630,);
not I_7505 (I130638,I130630);
nor I_7506 (I130087,I130638,I130350);
not I_7507 (I130696,I3042);
DFFARX1 I_7508 (I230461,I3035,I130696,I130722,);
DFFARX1 I_7509 (I130722,I3035,I130696,I130739,);
not I_7510 (I130688,I130739);
not I_7511 (I130761,I130722);
DFFARX1 I_7512 (I230449,I3035,I130696,I130787,);
not I_7513 (I130795,I130787);
and I_7514 (I130812,I130761,I230458);
not I_7515 (I130829,I230455);
nand I_7516 (I130846,I130829,I230458);
not I_7517 (I130863,I230446);
nor I_7518 (I130880,I130863,I230452);
nand I_7519 (I130897,I130880,I230437);
nor I_7520 (I130914,I130897,I130846);
DFFARX1 I_7521 (I130914,I3035,I130696,I130664,);
not I_7522 (I130945,I130897);
not I_7523 (I130962,I230452);
nand I_7524 (I130979,I130962,I230458);
nor I_7525 (I130996,I230452,I230455);
nand I_7526 (I130676,I130812,I130996);
nand I_7527 (I130670,I130761,I230452);
nand I_7528 (I131041,I130863,I230437);
DFFARX1 I_7529 (I131041,I3035,I130696,I130685,);
DFFARX1 I_7530 (I131041,I3035,I130696,I130679,);
not I_7531 (I131086,I230437);
nor I_7532 (I131103,I131086,I230443);
and I_7533 (I131120,I131103,I230440);
or I_7534 (I131137,I131120,I230464);
DFFARX1 I_7535 (I131137,I3035,I130696,I131163,);
nand I_7536 (I131171,I131163,I130829);
nor I_7537 (I130673,I131171,I130979);
nor I_7538 (I130667,I131163,I130795);
DFFARX1 I_7539 (I131163,I3035,I130696,I131225,);
not I_7540 (I131233,I131225);
nor I_7541 (I130682,I131233,I130945);
not I_7542 (I131291,I3042);
DFFARX1 I_7543 (I435616,I3035,I131291,I131317,);
DFFARX1 I_7544 (I131317,I3035,I131291,I131334,);
not I_7545 (I131283,I131334);
not I_7546 (I131356,I131317);
DFFARX1 I_7547 (I435610,I3035,I131291,I131382,);
not I_7548 (I131390,I131382);
and I_7549 (I131407,I131356,I435628);
not I_7550 (I131424,I435616);
nand I_7551 (I131441,I131424,I435628);
not I_7552 (I131458,I435610);
nor I_7553 (I131475,I131458,I435622);
nand I_7554 (I131492,I131475,I435613);
nor I_7555 (I131509,I131492,I131441);
DFFARX1 I_7556 (I131509,I3035,I131291,I131259,);
not I_7557 (I131540,I131492);
not I_7558 (I131557,I435622);
nand I_7559 (I131574,I131557,I435628);
nor I_7560 (I131591,I435622,I435616);
nand I_7561 (I131271,I131407,I131591);
nand I_7562 (I131265,I131356,I435622);
nand I_7563 (I131636,I131458,I435625);
DFFARX1 I_7564 (I131636,I3035,I131291,I131280,);
DFFARX1 I_7565 (I131636,I3035,I131291,I131274,);
not I_7566 (I131681,I435625);
nor I_7567 (I131698,I131681,I435631);
and I_7568 (I131715,I131698,I435613);
or I_7569 (I131732,I131715,I435619);
DFFARX1 I_7570 (I131732,I3035,I131291,I131758,);
nand I_7571 (I131766,I131758,I131424);
nor I_7572 (I131268,I131766,I131574);
nor I_7573 (I131262,I131758,I131390);
DFFARX1 I_7574 (I131758,I3035,I131291,I131820,);
not I_7575 (I131828,I131820);
nor I_7576 (I131277,I131828,I131540);
not I_7577 (I131886,I3042);
DFFARX1 I_7578 (I52609,I3035,I131886,I131912,);
DFFARX1 I_7579 (I131912,I3035,I131886,I131929,);
not I_7580 (I131878,I131929);
not I_7581 (I131951,I131912);
DFFARX1 I_7582 (I52603,I3035,I131886,I131977,);
not I_7583 (I131985,I131977);
and I_7584 (I132002,I131951,I52600);
not I_7585 (I132019,I52621);
nand I_7586 (I132036,I132019,I52600);
not I_7587 (I132053,I52615);
nor I_7588 (I132070,I132053,I52606);
nand I_7589 (I132087,I132070,I52612);
nor I_7590 (I132104,I132087,I132036);
DFFARX1 I_7591 (I132104,I3035,I131886,I131854,);
not I_7592 (I132135,I132087);
not I_7593 (I132152,I52606);
nand I_7594 (I132169,I132152,I52600);
nor I_7595 (I132186,I52606,I52621);
nand I_7596 (I131866,I132002,I132186);
nand I_7597 (I131860,I131951,I52606);
nand I_7598 (I132231,I132053,I52600);
DFFARX1 I_7599 (I132231,I3035,I131886,I131875,);
DFFARX1 I_7600 (I132231,I3035,I131886,I131869,);
not I_7601 (I132276,I52600);
nor I_7602 (I132293,I132276,I52618);
and I_7603 (I132310,I132293,I52624);
or I_7604 (I132327,I132310,I52603);
DFFARX1 I_7605 (I132327,I3035,I131886,I132353,);
nand I_7606 (I132361,I132353,I132019);
nor I_7607 (I131863,I132361,I132169);
nor I_7608 (I131857,I132353,I131985);
DFFARX1 I_7609 (I132353,I3035,I131886,I132415,);
not I_7610 (I132423,I132415);
nor I_7611 (I131872,I132423,I132135);
not I_7612 (I132481,I3042);
DFFARX1 I_7613 (I632980,I3035,I132481,I132507,);
DFFARX1 I_7614 (I132507,I3035,I132481,I132524,);
not I_7615 (I132473,I132524);
not I_7616 (I132546,I132507);
DFFARX1 I_7617 (I632980,I3035,I132481,I132572,);
not I_7618 (I132580,I132572);
and I_7619 (I132597,I132546,I632983);
not I_7620 (I132614,I632995);
nand I_7621 (I132631,I132614,I632983);
not I_7622 (I132648,I633001);
nor I_7623 (I132665,I132648,I632992);
nand I_7624 (I132682,I132665,I632998);
nor I_7625 (I132699,I132682,I132631);
DFFARX1 I_7626 (I132699,I3035,I132481,I132449,);
not I_7627 (I132730,I132682);
not I_7628 (I132747,I632992);
nand I_7629 (I132764,I132747,I632983);
nor I_7630 (I132781,I632992,I632995);
nand I_7631 (I132461,I132597,I132781);
nand I_7632 (I132455,I132546,I632992);
nand I_7633 (I132826,I132648,I632989);
DFFARX1 I_7634 (I132826,I3035,I132481,I132470,);
DFFARX1 I_7635 (I132826,I3035,I132481,I132464,);
not I_7636 (I132871,I632989);
nor I_7637 (I132888,I132871,I632986);
and I_7638 (I132905,I132888,I633004);
or I_7639 (I132922,I132905,I632983);
DFFARX1 I_7640 (I132922,I3035,I132481,I132948,);
nand I_7641 (I132956,I132948,I132614);
nor I_7642 (I132458,I132956,I132764);
nor I_7643 (I132452,I132948,I132580);
DFFARX1 I_7644 (I132948,I3035,I132481,I133010,);
not I_7645 (I133018,I133010);
nor I_7646 (I132467,I133018,I132730);
not I_7647 (I133076,I3042);
DFFARX1 I_7648 (I290068,I3035,I133076,I133102,);
DFFARX1 I_7649 (I133102,I3035,I133076,I133119,);
not I_7650 (I133068,I133119);
not I_7651 (I133141,I133102);
DFFARX1 I_7652 (I290062,I3035,I133076,I133167,);
not I_7653 (I133175,I133167);
and I_7654 (I133192,I133141,I290077);
not I_7655 (I133209,I290074);
nand I_7656 (I133226,I133209,I290077);
not I_7657 (I133243,I290065);
nor I_7658 (I133260,I133243,I290056);
nand I_7659 (I133277,I133260,I290059);
nor I_7660 (I133294,I133277,I133226);
DFFARX1 I_7661 (I133294,I3035,I133076,I133044,);
not I_7662 (I133325,I133277);
not I_7663 (I133342,I290056);
nand I_7664 (I133359,I133342,I290077);
nor I_7665 (I133376,I290056,I290074);
nand I_7666 (I133056,I133192,I133376);
nand I_7667 (I133050,I133141,I290056);
nand I_7668 (I133421,I133243,I290080);
DFFARX1 I_7669 (I133421,I3035,I133076,I133065,);
DFFARX1 I_7670 (I133421,I3035,I133076,I133059,);
not I_7671 (I133466,I290080);
nor I_7672 (I133483,I133466,I290071);
and I_7673 (I133500,I133483,I290056);
or I_7674 (I133517,I133500,I290059);
DFFARX1 I_7675 (I133517,I3035,I133076,I133543,);
nand I_7676 (I133551,I133543,I133209);
nor I_7677 (I133053,I133551,I133359);
nor I_7678 (I133047,I133543,I133175);
DFFARX1 I_7679 (I133543,I3035,I133076,I133605,);
not I_7680 (I133613,I133605);
nor I_7681 (I133062,I133613,I133325);
not I_7682 (I133671,I3042);
DFFARX1 I_7683 (I527765,I3035,I133671,I133697,);
DFFARX1 I_7684 (I133697,I3035,I133671,I133714,);
not I_7685 (I133663,I133714);
not I_7686 (I133736,I133697);
DFFARX1 I_7687 (I527774,I3035,I133671,I133762,);
not I_7688 (I133770,I133762);
and I_7689 (I133787,I133736,I527762);
not I_7690 (I133804,I527753);
nand I_7691 (I133821,I133804,I527762);
not I_7692 (I133838,I527759);
nor I_7693 (I133855,I133838,I527777);
nand I_7694 (I133872,I133855,I527750);
nor I_7695 (I133889,I133872,I133821);
DFFARX1 I_7696 (I133889,I3035,I133671,I133639,);
not I_7697 (I133920,I133872);
not I_7698 (I133937,I527777);
nand I_7699 (I133954,I133937,I527762);
nor I_7700 (I133971,I527777,I527753);
nand I_7701 (I133651,I133787,I133971);
nand I_7702 (I133645,I133736,I527777);
nand I_7703 (I134016,I133838,I527756);
DFFARX1 I_7704 (I134016,I3035,I133671,I133660,);
DFFARX1 I_7705 (I134016,I3035,I133671,I133654,);
not I_7706 (I134061,I527756);
nor I_7707 (I134078,I134061,I527768);
and I_7708 (I134095,I134078,I527750);
or I_7709 (I134112,I134095,I527771);
DFFARX1 I_7710 (I134112,I3035,I133671,I134138,);
nand I_7711 (I134146,I134138,I133804);
nor I_7712 (I133648,I134146,I133954);
nor I_7713 (I133642,I134138,I133770);
DFFARX1 I_7714 (I134138,I3035,I133671,I134200,);
not I_7715 (I134208,I134200);
nor I_7716 (I133657,I134208,I133920);
not I_7717 (I134266,I3042);
DFFARX1 I_7718 (I161366,I3035,I134266,I134292,);
DFFARX1 I_7719 (I134292,I3035,I134266,I134309,);
not I_7720 (I134258,I134309);
not I_7721 (I134331,I134292);
DFFARX1 I_7722 (I161381,I3035,I134266,I134357,);
not I_7723 (I134365,I134357);
and I_7724 (I134382,I134331,I161378);
not I_7725 (I134399,I161366);
nand I_7726 (I134416,I134399,I161378);
not I_7727 (I134433,I161375);
nor I_7728 (I134450,I134433,I161390);
nand I_7729 (I134467,I134450,I161387);
nor I_7730 (I134484,I134467,I134416);
DFFARX1 I_7731 (I134484,I3035,I134266,I134234,);
not I_7732 (I134515,I134467);
not I_7733 (I134532,I161390);
nand I_7734 (I134549,I134532,I161378);
nor I_7735 (I134566,I161390,I161366);
nand I_7736 (I134246,I134382,I134566);
nand I_7737 (I134240,I134331,I161390);
nand I_7738 (I134611,I134433,I161384);
DFFARX1 I_7739 (I134611,I3035,I134266,I134255,);
DFFARX1 I_7740 (I134611,I3035,I134266,I134249,);
not I_7741 (I134656,I161384);
nor I_7742 (I134673,I134656,I161372);
and I_7743 (I134690,I134673,I161393);
or I_7744 (I134707,I134690,I161369);
DFFARX1 I_7745 (I134707,I3035,I134266,I134733,);
nand I_7746 (I134741,I134733,I134399);
nor I_7747 (I134243,I134741,I134549);
nor I_7748 (I134237,I134733,I134365);
DFFARX1 I_7749 (I134733,I3035,I134266,I134795,);
not I_7750 (I134803,I134795);
nor I_7751 (I134252,I134803,I134515);
not I_7752 (I134861,I3042);
DFFARX1 I_7753 (I187189,I3035,I134861,I134887,);
DFFARX1 I_7754 (I134887,I3035,I134861,I134904,);
not I_7755 (I134853,I134904);
not I_7756 (I134926,I134887);
DFFARX1 I_7757 (I187204,I3035,I134861,I134952,);
not I_7758 (I134960,I134952);
and I_7759 (I134977,I134926,I187201);
not I_7760 (I134994,I187189);
nand I_7761 (I135011,I134994,I187201);
not I_7762 (I135028,I187198);
nor I_7763 (I135045,I135028,I187213);
nand I_7764 (I135062,I135045,I187210);
nor I_7765 (I135079,I135062,I135011);
DFFARX1 I_7766 (I135079,I3035,I134861,I134829,);
not I_7767 (I135110,I135062);
not I_7768 (I135127,I187213);
nand I_7769 (I135144,I135127,I187201);
nor I_7770 (I135161,I187213,I187189);
nand I_7771 (I134841,I134977,I135161);
nand I_7772 (I134835,I134926,I187213);
nand I_7773 (I135206,I135028,I187207);
DFFARX1 I_7774 (I135206,I3035,I134861,I134850,);
DFFARX1 I_7775 (I135206,I3035,I134861,I134844,);
not I_7776 (I135251,I187207);
nor I_7777 (I135268,I135251,I187195);
and I_7778 (I135285,I135268,I187216);
or I_7779 (I135302,I135285,I187192);
DFFARX1 I_7780 (I135302,I3035,I134861,I135328,);
nand I_7781 (I135336,I135328,I134994);
nor I_7782 (I134838,I135336,I135144);
nor I_7783 (I134832,I135328,I134960);
DFFARX1 I_7784 (I135328,I3035,I134861,I135390,);
not I_7785 (I135398,I135390);
nor I_7786 (I134847,I135398,I135110);
not I_7787 (I135456,I3042);
DFFARX1 I_7788 (I501279,I3035,I135456,I135482,);
DFFARX1 I_7789 (I135482,I3035,I135456,I135499,);
not I_7790 (I135448,I135499);
not I_7791 (I135521,I135482);
DFFARX1 I_7792 (I501288,I3035,I135456,I135547,);
not I_7793 (I135555,I135547);
and I_7794 (I135572,I135521,I501276);
not I_7795 (I135589,I501267);
nand I_7796 (I135606,I135589,I501276);
not I_7797 (I135623,I501273);
nor I_7798 (I135640,I135623,I501291);
nand I_7799 (I135657,I135640,I501264);
nor I_7800 (I135674,I135657,I135606);
DFFARX1 I_7801 (I135674,I3035,I135456,I135424,);
not I_7802 (I135705,I135657);
not I_7803 (I135722,I501291);
nand I_7804 (I135739,I135722,I501276);
nor I_7805 (I135756,I501291,I501267);
nand I_7806 (I135436,I135572,I135756);
nand I_7807 (I135430,I135521,I501291);
nand I_7808 (I135801,I135623,I501270);
DFFARX1 I_7809 (I135801,I3035,I135456,I135445,);
DFFARX1 I_7810 (I135801,I3035,I135456,I135439,);
not I_7811 (I135846,I501270);
nor I_7812 (I135863,I135846,I501282);
and I_7813 (I135880,I135863,I501264);
or I_7814 (I135897,I135880,I501285);
DFFARX1 I_7815 (I135897,I3035,I135456,I135923,);
nand I_7816 (I135931,I135923,I135589);
nor I_7817 (I135433,I135931,I135739);
nor I_7818 (I135427,I135923,I135555);
DFFARX1 I_7819 (I135923,I3035,I135456,I135985,);
not I_7820 (I135993,I135985);
nor I_7821 (I135442,I135993,I135705);
not I_7822 (I136051,I3042);
DFFARX1 I_7823 (I156096,I3035,I136051,I136077,);
DFFARX1 I_7824 (I136077,I3035,I136051,I136094,);
not I_7825 (I136043,I136094);
not I_7826 (I136116,I136077);
DFFARX1 I_7827 (I156111,I3035,I136051,I136142,);
not I_7828 (I136150,I136142);
and I_7829 (I136167,I136116,I156108);
not I_7830 (I136184,I156096);
nand I_7831 (I136201,I136184,I156108);
not I_7832 (I136218,I156105);
nor I_7833 (I136235,I136218,I156120);
nand I_7834 (I136252,I136235,I156117);
nor I_7835 (I136269,I136252,I136201);
DFFARX1 I_7836 (I136269,I3035,I136051,I136019,);
not I_7837 (I136300,I136252);
not I_7838 (I136317,I156120);
nand I_7839 (I136334,I136317,I156108);
nor I_7840 (I136351,I156120,I156096);
nand I_7841 (I136031,I136167,I136351);
nand I_7842 (I136025,I136116,I156120);
nand I_7843 (I136396,I136218,I156114);
DFFARX1 I_7844 (I136396,I3035,I136051,I136040,);
DFFARX1 I_7845 (I136396,I3035,I136051,I136034,);
not I_7846 (I136441,I156114);
nor I_7847 (I136458,I136441,I156102);
and I_7848 (I136475,I136458,I156123);
or I_7849 (I136492,I136475,I156099);
DFFARX1 I_7850 (I136492,I3035,I136051,I136518,);
nand I_7851 (I136526,I136518,I136184);
nor I_7852 (I136028,I136526,I136334);
nor I_7853 (I136022,I136518,I136150);
DFFARX1 I_7854 (I136518,I3035,I136051,I136580,);
not I_7855 (I136588,I136580);
nor I_7856 (I136037,I136588,I136300);
not I_7857 (I136646,I3042);
DFFARX1 I_7858 (I194040,I3035,I136646,I136672,);
DFFARX1 I_7859 (I136672,I3035,I136646,I136689,);
not I_7860 (I136638,I136689);
not I_7861 (I136711,I136672);
DFFARX1 I_7862 (I194055,I3035,I136646,I136737,);
not I_7863 (I136745,I136737);
and I_7864 (I136762,I136711,I194052);
not I_7865 (I136779,I194040);
nand I_7866 (I136796,I136779,I194052);
not I_7867 (I136813,I194049);
nor I_7868 (I136830,I136813,I194064);
nand I_7869 (I136847,I136830,I194061);
nor I_7870 (I136864,I136847,I136796);
DFFARX1 I_7871 (I136864,I3035,I136646,I136614,);
not I_7872 (I136895,I136847);
not I_7873 (I136912,I194064);
nand I_7874 (I136929,I136912,I194052);
nor I_7875 (I136946,I194064,I194040);
nand I_7876 (I136626,I136762,I136946);
nand I_7877 (I136620,I136711,I194064);
nand I_7878 (I136991,I136813,I194058);
DFFARX1 I_7879 (I136991,I3035,I136646,I136635,);
DFFARX1 I_7880 (I136991,I3035,I136646,I136629,);
not I_7881 (I137036,I194058);
nor I_7882 (I137053,I137036,I194046);
and I_7883 (I137070,I137053,I194067);
or I_7884 (I137087,I137070,I194043);
DFFARX1 I_7885 (I137087,I3035,I136646,I137113,);
nand I_7886 (I137121,I137113,I136779);
nor I_7887 (I136623,I137121,I136929);
nor I_7888 (I136617,I137113,I136745);
DFFARX1 I_7889 (I137113,I3035,I136646,I137175,);
not I_7890 (I137183,I137175);
nor I_7891 (I136632,I137183,I136895);
not I_7892 (I137241,I3042);
DFFARX1 I_7893 (I266365,I3035,I137241,I137267,);
DFFARX1 I_7894 (I137267,I3035,I137241,I137284,);
not I_7895 (I137233,I137284);
not I_7896 (I137306,I137267);
DFFARX1 I_7897 (I266353,I3035,I137241,I137332,);
not I_7898 (I137340,I137332);
and I_7899 (I137357,I137306,I266362);
not I_7900 (I137374,I266359);
nand I_7901 (I137391,I137374,I266362);
not I_7902 (I137408,I266350);
nor I_7903 (I137425,I137408,I266356);
nand I_7904 (I137442,I137425,I266341);
nor I_7905 (I137459,I137442,I137391);
DFFARX1 I_7906 (I137459,I3035,I137241,I137209,);
not I_7907 (I137490,I137442);
not I_7908 (I137507,I266356);
nand I_7909 (I137524,I137507,I266362);
nor I_7910 (I137541,I266356,I266359);
nand I_7911 (I137221,I137357,I137541);
nand I_7912 (I137215,I137306,I266356);
nand I_7913 (I137586,I137408,I266341);
DFFARX1 I_7914 (I137586,I3035,I137241,I137230,);
DFFARX1 I_7915 (I137586,I3035,I137241,I137224,);
not I_7916 (I137631,I266341);
nor I_7917 (I137648,I137631,I266347);
and I_7918 (I137665,I137648,I266344);
or I_7919 (I137682,I137665,I266368);
DFFARX1 I_7920 (I137682,I3035,I137241,I137708,);
nand I_7921 (I137716,I137708,I137374);
nor I_7922 (I137218,I137716,I137524);
nor I_7923 (I137212,I137708,I137340);
DFFARX1 I_7924 (I137708,I3035,I137241,I137770,);
not I_7925 (I137778,I137770);
nor I_7926 (I137227,I137778,I137490);
not I_7927 (I137836,I3042);
DFFARX1 I_7928 (I178230,I3035,I137836,I137862,);
DFFARX1 I_7929 (I137862,I3035,I137836,I137879,);
not I_7930 (I137828,I137879);
not I_7931 (I137901,I137862);
DFFARX1 I_7932 (I178245,I3035,I137836,I137927,);
not I_7933 (I137935,I137927);
and I_7934 (I137952,I137901,I178242);
not I_7935 (I137969,I178230);
nand I_7936 (I137986,I137969,I178242);
not I_7937 (I138003,I178239);
nor I_7938 (I138020,I138003,I178254);
nand I_7939 (I138037,I138020,I178251);
nor I_7940 (I138054,I138037,I137986);
DFFARX1 I_7941 (I138054,I3035,I137836,I137804,);
not I_7942 (I138085,I138037);
not I_7943 (I138102,I178254);
nand I_7944 (I138119,I138102,I178242);
nor I_7945 (I138136,I178254,I178230);
nand I_7946 (I137816,I137952,I138136);
nand I_7947 (I137810,I137901,I178254);
nand I_7948 (I138181,I138003,I178248);
DFFARX1 I_7949 (I138181,I3035,I137836,I137825,);
DFFARX1 I_7950 (I138181,I3035,I137836,I137819,);
not I_7951 (I138226,I178248);
nor I_7952 (I138243,I138226,I178236);
and I_7953 (I138260,I138243,I178257);
or I_7954 (I138277,I138260,I178233);
DFFARX1 I_7955 (I138277,I3035,I137836,I138303,);
nand I_7956 (I138311,I138303,I137969);
nor I_7957 (I137813,I138311,I138119);
nor I_7958 (I137807,I138303,I137935);
DFFARX1 I_7959 (I138303,I3035,I137836,I138365,);
not I_7960 (I138373,I138365);
nor I_7961 (I137822,I138373,I138085);
not I_7962 (I138431,I3042);
DFFARX1 I_7963 (I589630,I3035,I138431,I138457,);
DFFARX1 I_7964 (I138457,I3035,I138431,I138474,);
not I_7965 (I138423,I138474);
not I_7966 (I138496,I138457);
DFFARX1 I_7967 (I589630,I3035,I138431,I138522,);
not I_7968 (I138530,I138522);
and I_7969 (I138547,I138496,I589633);
not I_7970 (I138564,I589645);
nand I_7971 (I138581,I138564,I589633);
not I_7972 (I138598,I589651);
nor I_7973 (I138615,I138598,I589642);
nand I_7974 (I138632,I138615,I589648);
nor I_7975 (I138649,I138632,I138581);
DFFARX1 I_7976 (I138649,I3035,I138431,I138399,);
not I_7977 (I138680,I138632);
not I_7978 (I138697,I589642);
nand I_7979 (I138714,I138697,I589633);
nor I_7980 (I138731,I589642,I589645);
nand I_7981 (I138411,I138547,I138731);
nand I_7982 (I138405,I138496,I589642);
nand I_7983 (I138776,I138598,I589639);
DFFARX1 I_7984 (I138776,I3035,I138431,I138420,);
DFFARX1 I_7985 (I138776,I3035,I138431,I138414,);
not I_7986 (I138821,I589639);
nor I_7987 (I138838,I138821,I589636);
and I_7988 (I138855,I138838,I589654);
or I_7989 (I138872,I138855,I589633);
DFFARX1 I_7990 (I138872,I3035,I138431,I138898,);
nand I_7991 (I138906,I138898,I138564);
nor I_7992 (I138408,I138906,I138714);
nor I_7993 (I138402,I138898,I138530);
DFFARX1 I_7994 (I138898,I3035,I138431,I138960,);
not I_7995 (I138968,I138960);
nor I_7996 (I138417,I138968,I138680);
not I_7997 (I139026,I3042);
DFFARX1 I_7998 (I664312,I3035,I139026,I139052,);
DFFARX1 I_7999 (I139052,I3035,I139026,I139069,);
not I_8000 (I139018,I139069);
not I_8001 (I139091,I139052);
DFFARX1 I_8002 (I664297,I3035,I139026,I139117,);
not I_8003 (I139125,I139117);
and I_8004 (I139142,I139091,I664315);
not I_8005 (I139159,I664297);
nand I_8006 (I139176,I139159,I664315);
not I_8007 (I139193,I664318);
nor I_8008 (I139210,I139193,I664309);
nand I_8009 (I139227,I139210,I664306);
nor I_8010 (I139244,I139227,I139176);
DFFARX1 I_8011 (I139244,I3035,I139026,I138994,);
not I_8012 (I139275,I139227);
not I_8013 (I139292,I664309);
nand I_8014 (I139309,I139292,I664315);
nor I_8015 (I139326,I664309,I664297);
nand I_8016 (I139006,I139142,I139326);
nand I_8017 (I139000,I139091,I664309);
nand I_8018 (I139371,I139193,I664303);
DFFARX1 I_8019 (I139371,I3035,I139026,I139015,);
DFFARX1 I_8020 (I139371,I3035,I139026,I139009,);
not I_8021 (I139416,I664303);
nor I_8022 (I139433,I139416,I664294);
and I_8023 (I139450,I139433,I664300);
or I_8024 (I139467,I139450,I664294);
DFFARX1 I_8025 (I139467,I3035,I139026,I139493,);
nand I_8026 (I139501,I139493,I139159);
nor I_8027 (I139003,I139501,I139309);
nor I_8028 (I138997,I139493,I139125);
DFFARX1 I_8029 (I139493,I3035,I139026,I139555,);
not I_8030 (I139563,I139555);
nor I_8031 (I139012,I139563,I139275);
not I_8032 (I139621,I3042);
DFFARX1 I_8033 (I648536,I3035,I139621,I139647,);
DFFARX1 I_8034 (I139647,I3035,I139621,I139664,);
not I_8035 (I139613,I139664);
not I_8036 (I139686,I139647);
DFFARX1 I_8037 (I648521,I3035,I139621,I139712,);
not I_8038 (I139720,I139712);
and I_8039 (I139737,I139686,I648539);
not I_8040 (I139754,I648521);
nand I_8041 (I139771,I139754,I648539);
not I_8042 (I139788,I648542);
nor I_8043 (I139805,I139788,I648533);
nand I_8044 (I139822,I139805,I648530);
nor I_8045 (I139839,I139822,I139771);
DFFARX1 I_8046 (I139839,I3035,I139621,I139589,);
not I_8047 (I139870,I139822);
not I_8048 (I139887,I648533);
nand I_8049 (I139904,I139887,I648539);
nor I_8050 (I139921,I648533,I648521);
nand I_8051 (I139601,I139737,I139921);
nand I_8052 (I139595,I139686,I648533);
nand I_8053 (I139966,I139788,I648527);
DFFARX1 I_8054 (I139966,I3035,I139621,I139610,);
DFFARX1 I_8055 (I139966,I3035,I139621,I139604,);
not I_8056 (I140011,I648527);
nor I_8057 (I140028,I140011,I648518);
and I_8058 (I140045,I140028,I648524);
or I_8059 (I140062,I140045,I648518);
DFFARX1 I_8060 (I140062,I3035,I139621,I140088,);
nand I_8061 (I140096,I140088,I139754);
nor I_8062 (I139598,I140096,I139904);
nor I_8063 (I139592,I140088,I139720);
DFFARX1 I_8064 (I140088,I3035,I139621,I140150,);
not I_8065 (I140158,I140150);
nor I_8066 (I139607,I140158,I139870);
not I_8067 (I140216,I3042);
DFFARX1 I_8068 (I155569,I3035,I140216,I140242,);
DFFARX1 I_8069 (I140242,I3035,I140216,I140259,);
not I_8070 (I140208,I140259);
not I_8071 (I140281,I140242);
DFFARX1 I_8072 (I155584,I3035,I140216,I140307,);
not I_8073 (I140315,I140307);
and I_8074 (I140332,I140281,I155581);
not I_8075 (I140349,I155569);
nand I_8076 (I140366,I140349,I155581);
not I_8077 (I140383,I155578);
nor I_8078 (I140400,I140383,I155593);
nand I_8079 (I140417,I140400,I155590);
nor I_8080 (I140434,I140417,I140366);
DFFARX1 I_8081 (I140434,I3035,I140216,I140184,);
not I_8082 (I140465,I140417);
not I_8083 (I140482,I155593);
nand I_8084 (I140499,I140482,I155581);
nor I_8085 (I140516,I155593,I155569);
nand I_8086 (I140196,I140332,I140516);
nand I_8087 (I140190,I140281,I155593);
nand I_8088 (I140561,I140383,I155587);
DFFARX1 I_8089 (I140561,I3035,I140216,I140205,);
DFFARX1 I_8090 (I140561,I3035,I140216,I140199,);
not I_8091 (I140606,I155587);
nor I_8092 (I140623,I140606,I155575);
and I_8093 (I140640,I140623,I155596);
or I_8094 (I140657,I140640,I155572);
DFFARX1 I_8095 (I140657,I3035,I140216,I140683,);
nand I_8096 (I140691,I140683,I140349);
nor I_8097 (I140193,I140691,I140499);
nor I_8098 (I140187,I140683,I140315);
DFFARX1 I_8099 (I140683,I3035,I140216,I140745,);
not I_8100 (I140753,I140745);
nor I_8101 (I140202,I140753,I140465);
not I_8102 (I140811,I3042);
DFFARX1 I_8103 (I463020,I3035,I140811,I140837,);
DFFARX1 I_8104 (I140837,I3035,I140811,I140854,);
not I_8105 (I140803,I140854);
not I_8106 (I140876,I140837);
DFFARX1 I_8107 (I463014,I3035,I140811,I140902,);
not I_8108 (I140910,I140902);
and I_8109 (I140927,I140876,I463032);
not I_8110 (I140944,I463020);
nand I_8111 (I140961,I140944,I463032);
not I_8112 (I140978,I463014);
nor I_8113 (I140995,I140978,I463026);
nand I_8114 (I141012,I140995,I463017);
nor I_8115 (I141029,I141012,I140961);
DFFARX1 I_8116 (I141029,I3035,I140811,I140779,);
not I_8117 (I141060,I141012);
not I_8118 (I141077,I463026);
nand I_8119 (I141094,I141077,I463032);
nor I_8120 (I141111,I463026,I463020);
nand I_8121 (I140791,I140927,I141111);
nand I_8122 (I140785,I140876,I463026);
nand I_8123 (I141156,I140978,I463029);
DFFARX1 I_8124 (I141156,I3035,I140811,I140800,);
DFFARX1 I_8125 (I141156,I3035,I140811,I140794,);
not I_8126 (I141201,I463029);
nor I_8127 (I141218,I141201,I463035);
and I_8128 (I141235,I141218,I463017);
or I_8129 (I141252,I141235,I463023);
DFFARX1 I_8130 (I141252,I3035,I140811,I141278,);
nand I_8131 (I141286,I141278,I140944);
nor I_8132 (I140788,I141286,I141094);
nor I_8133 (I140782,I141278,I140910);
DFFARX1 I_8134 (I141278,I3035,I140811,I141340,);
not I_8135 (I141348,I141340);
nor I_8136 (I140797,I141348,I141060);
not I_8137 (I141406,I3042);
DFFARX1 I_8138 (I667576,I3035,I141406,I141432,);
DFFARX1 I_8139 (I141432,I3035,I141406,I141449,);
not I_8140 (I141398,I141449);
not I_8141 (I141471,I141432);
DFFARX1 I_8142 (I667561,I3035,I141406,I141497,);
not I_8143 (I141505,I141497);
and I_8144 (I141522,I141471,I667579);
not I_8145 (I141539,I667561);
nand I_8146 (I141556,I141539,I667579);
not I_8147 (I141573,I667582);
nor I_8148 (I141590,I141573,I667573);
nand I_8149 (I141607,I141590,I667570);
nor I_8150 (I141624,I141607,I141556);
DFFARX1 I_8151 (I141624,I3035,I141406,I141374,);
not I_8152 (I141655,I141607);
not I_8153 (I141672,I667573);
nand I_8154 (I141689,I141672,I667579);
nor I_8155 (I141706,I667573,I667561);
nand I_8156 (I141386,I141522,I141706);
nand I_8157 (I141380,I141471,I667573);
nand I_8158 (I141751,I141573,I667567);
DFFARX1 I_8159 (I141751,I3035,I141406,I141395,);
DFFARX1 I_8160 (I141751,I3035,I141406,I141389,);
not I_8161 (I141796,I667567);
nor I_8162 (I141813,I141796,I667558);
and I_8163 (I141830,I141813,I667564);
or I_8164 (I141847,I141830,I667558);
DFFARX1 I_8165 (I141847,I3035,I141406,I141873,);
nand I_8166 (I141881,I141873,I141539);
nor I_8167 (I141383,I141881,I141689);
nor I_8168 (I141377,I141873,I141505);
DFFARX1 I_8169 (I141873,I3035,I141406,I141935,);
not I_8170 (I141943,I141935);
nor I_8171 (I141392,I141943,I141655);
not I_8172 (I142001,I3042);
DFFARX1 I_8173 (I590208,I3035,I142001,I142027,);
DFFARX1 I_8174 (I142027,I3035,I142001,I142044,);
not I_8175 (I141993,I142044);
not I_8176 (I142066,I142027);
DFFARX1 I_8177 (I590208,I3035,I142001,I142092,);
not I_8178 (I142100,I142092);
and I_8179 (I142117,I142066,I590211);
not I_8180 (I142134,I590223);
nand I_8181 (I142151,I142134,I590211);
not I_8182 (I142168,I590229);
nor I_8183 (I142185,I142168,I590220);
nand I_8184 (I142202,I142185,I590226);
nor I_8185 (I142219,I142202,I142151);
DFFARX1 I_8186 (I142219,I3035,I142001,I141969,);
not I_8187 (I142250,I142202);
not I_8188 (I142267,I590220);
nand I_8189 (I142284,I142267,I590211);
nor I_8190 (I142301,I590220,I590223);
nand I_8191 (I141981,I142117,I142301);
nand I_8192 (I141975,I142066,I590220);
nand I_8193 (I142346,I142168,I590217);
DFFARX1 I_8194 (I142346,I3035,I142001,I141990,);
DFFARX1 I_8195 (I142346,I3035,I142001,I141984,);
not I_8196 (I142391,I590217);
nor I_8197 (I142408,I142391,I590214);
and I_8198 (I142425,I142408,I590232);
or I_8199 (I142442,I142425,I590211);
DFFARX1 I_8200 (I142442,I3035,I142001,I142468,);
nand I_8201 (I142476,I142468,I142134);
nor I_8202 (I141978,I142476,I142284);
nor I_8203 (I141972,I142468,I142100);
DFFARX1 I_8204 (I142468,I3035,I142001,I142530,);
not I_8205 (I142538,I142530);
nor I_8206 (I141987,I142538,I142250);
not I_8207 (I142596,I3042);
DFFARX1 I_8208 (I296018,I3035,I142596,I142622,);
DFFARX1 I_8209 (I142622,I3035,I142596,I142639,);
not I_8210 (I142588,I142639);
not I_8211 (I142661,I142622);
DFFARX1 I_8212 (I296012,I3035,I142596,I142687,);
not I_8213 (I142695,I142687);
and I_8214 (I142712,I142661,I296027);
not I_8215 (I142729,I296024);
nand I_8216 (I142746,I142729,I296027);
not I_8217 (I142763,I296015);
nor I_8218 (I142780,I142763,I296006);
nand I_8219 (I142797,I142780,I296009);
nor I_8220 (I142814,I142797,I142746);
DFFARX1 I_8221 (I142814,I3035,I142596,I142564,);
not I_8222 (I142845,I142797);
not I_8223 (I142862,I296006);
nand I_8224 (I142879,I142862,I296027);
nor I_8225 (I142896,I296006,I296024);
nand I_8226 (I142576,I142712,I142896);
nand I_8227 (I142570,I142661,I296006);
nand I_8228 (I142941,I142763,I296030);
DFFARX1 I_8229 (I142941,I3035,I142596,I142585,);
DFFARX1 I_8230 (I142941,I3035,I142596,I142579,);
not I_8231 (I142986,I296030);
nor I_8232 (I143003,I142986,I296021);
and I_8233 (I143020,I143003,I296006);
or I_8234 (I143037,I143020,I296009);
DFFARX1 I_8235 (I143037,I3035,I142596,I143063,);
nand I_8236 (I143071,I143063,I142729);
nor I_8237 (I142573,I143071,I142879);
nor I_8238 (I142567,I143063,I142695);
DFFARX1 I_8239 (I143063,I3035,I142596,I143125,);
not I_8240 (I143133,I143125);
nor I_8241 (I142582,I143133,I142845);
not I_8242 (I143191,I3042);
DFFARX1 I_8243 (I74752,I3035,I143191,I143217,);
DFFARX1 I_8244 (I143217,I3035,I143191,I143234,);
not I_8245 (I143183,I143234);
not I_8246 (I143256,I143217);
DFFARX1 I_8247 (I74737,I3035,I143191,I143282,);
not I_8248 (I143290,I143282);
and I_8249 (I143307,I143256,I74758);
not I_8250 (I143324,I74749);
nand I_8251 (I143341,I143324,I74758);
not I_8252 (I143358,I74734);
nor I_8253 (I143375,I143358,I74746);
nand I_8254 (I143392,I143375,I74761);
nor I_8255 (I143409,I143392,I143341);
DFFARX1 I_8256 (I143409,I3035,I143191,I143159,);
not I_8257 (I143440,I143392);
not I_8258 (I143457,I74746);
nand I_8259 (I143474,I143457,I74758);
nor I_8260 (I143491,I74746,I74749);
nand I_8261 (I143171,I143307,I143491);
nand I_8262 (I143165,I143256,I74746);
nand I_8263 (I143536,I143358,I74740);
DFFARX1 I_8264 (I143536,I3035,I143191,I143180,);
DFFARX1 I_8265 (I143536,I3035,I143191,I143174,);
not I_8266 (I143581,I74740);
nor I_8267 (I143598,I143581,I74743);
and I_8268 (I143615,I143598,I74734);
or I_8269 (I143632,I143615,I74755);
DFFARX1 I_8270 (I143632,I3035,I143191,I143658,);
nand I_8271 (I143666,I143658,I143324);
nor I_8272 (I143168,I143666,I143474);
nor I_8273 (I143162,I143658,I143290);
DFFARX1 I_8274 (I143658,I3035,I143191,I143720,);
not I_8275 (I143728,I143720);
nor I_8276 (I143177,I143728,I143440);
not I_8277 (I143786,I3042);
DFFARX1 I_8278 (I57879,I3035,I143786,I143812,);
DFFARX1 I_8279 (I143812,I3035,I143786,I143829,);
not I_8280 (I143778,I143829);
not I_8281 (I143851,I143812);
DFFARX1 I_8282 (I57873,I3035,I143786,I143877,);
not I_8283 (I143885,I143877);
and I_8284 (I143902,I143851,I57870);
not I_8285 (I143919,I57891);
nand I_8286 (I143936,I143919,I57870);
not I_8287 (I143953,I57885);
nor I_8288 (I143970,I143953,I57876);
nand I_8289 (I143987,I143970,I57882);
nor I_8290 (I144004,I143987,I143936);
DFFARX1 I_8291 (I144004,I3035,I143786,I143754,);
not I_8292 (I144035,I143987);
not I_8293 (I144052,I57876);
nand I_8294 (I144069,I144052,I57870);
nor I_8295 (I144086,I57876,I57891);
nand I_8296 (I143766,I143902,I144086);
nand I_8297 (I143760,I143851,I57876);
nand I_8298 (I144131,I143953,I57870);
DFFARX1 I_8299 (I144131,I3035,I143786,I143775,);
DFFARX1 I_8300 (I144131,I3035,I143786,I143769,);
not I_8301 (I144176,I57870);
nor I_8302 (I144193,I144176,I57888);
and I_8303 (I144210,I144193,I57894);
or I_8304 (I144227,I144210,I57873);
DFFARX1 I_8305 (I144227,I3035,I143786,I144253,);
nand I_8306 (I144261,I144253,I143919);
nor I_8307 (I143763,I144261,I144069);
nor I_8308 (I143757,I144253,I143885);
DFFARX1 I_8309 (I144253,I3035,I143786,I144315,);
not I_8310 (I144323,I144315);
nor I_8311 (I143772,I144323,I144035);
not I_8312 (I144381,I3042);
DFFARX1 I_8313 (I401894,I3035,I144381,I144407,);
DFFARX1 I_8314 (I144407,I3035,I144381,I144424,);
not I_8315 (I144373,I144424);
not I_8316 (I144446,I144407);
DFFARX1 I_8317 (I401891,I3035,I144381,I144472,);
not I_8318 (I144480,I144472);
and I_8319 (I144497,I144446,I401897);
not I_8320 (I144514,I401882);
nand I_8321 (I144531,I144514,I401897);
not I_8322 (I144548,I401885);
nor I_8323 (I144565,I144548,I401906);
nand I_8324 (I144582,I144565,I401903);
nor I_8325 (I144599,I144582,I144531);
DFFARX1 I_8326 (I144599,I3035,I144381,I144349,);
not I_8327 (I144630,I144582);
not I_8328 (I144647,I401906);
nand I_8329 (I144664,I144647,I401897);
nor I_8330 (I144681,I401906,I401882);
nand I_8331 (I144361,I144497,I144681);
nand I_8332 (I144355,I144446,I401906);
nand I_8333 (I144726,I144548,I401882);
DFFARX1 I_8334 (I144726,I3035,I144381,I144370,);
DFFARX1 I_8335 (I144726,I3035,I144381,I144364,);
not I_8336 (I144771,I401882);
nor I_8337 (I144788,I144771,I401888);
and I_8338 (I144805,I144788,I401900);
or I_8339 (I144822,I144805,I401885);
DFFARX1 I_8340 (I144822,I3035,I144381,I144848,);
nand I_8341 (I144856,I144848,I144514);
nor I_8342 (I144358,I144856,I144664);
nor I_8343 (I144352,I144848,I144480);
DFFARX1 I_8344 (I144848,I3035,I144381,I144910,);
not I_8345 (I144918,I144910);
nor I_8346 (I144367,I144918,I144630);
not I_8347 (I144976,I3042);
DFFARX1 I_8348 (I409408,I3035,I144976,I145002,);
DFFARX1 I_8349 (I145002,I3035,I144976,I145019,);
not I_8350 (I144968,I145019);
not I_8351 (I145041,I145002);
DFFARX1 I_8352 (I409405,I3035,I144976,I145067,);
not I_8353 (I145075,I145067);
and I_8354 (I145092,I145041,I409411);
not I_8355 (I145109,I409396);
nand I_8356 (I145126,I145109,I409411);
not I_8357 (I145143,I409399);
nor I_8358 (I145160,I145143,I409420);
nand I_8359 (I145177,I145160,I409417);
nor I_8360 (I145194,I145177,I145126);
DFFARX1 I_8361 (I145194,I3035,I144976,I144944,);
not I_8362 (I145225,I145177);
not I_8363 (I145242,I409420);
nand I_8364 (I145259,I145242,I409411);
nor I_8365 (I145276,I409420,I409396);
nand I_8366 (I144956,I145092,I145276);
nand I_8367 (I144950,I145041,I409420);
nand I_8368 (I145321,I145143,I409396);
DFFARX1 I_8369 (I145321,I3035,I144976,I144965,);
DFFARX1 I_8370 (I145321,I3035,I144976,I144959,);
not I_8371 (I145366,I409396);
nor I_8372 (I145383,I145366,I409402);
and I_8373 (I145400,I145383,I409414);
or I_8374 (I145417,I145400,I409399);
DFFARX1 I_8375 (I145417,I3035,I144976,I145443,);
nand I_8376 (I145451,I145443,I145109);
nor I_8377 (I144953,I145451,I145259);
nor I_8378 (I144947,I145443,I145075);
DFFARX1 I_8379 (I145443,I3035,I144976,I145505,);
not I_8380 (I145513,I145505);
nor I_8381 (I144962,I145513,I145225);
not I_8382 (I145571,I3042);
DFFARX1 I_8383 (I375306,I3035,I145571,I145597,);
DFFARX1 I_8384 (I145597,I3035,I145571,I145614,);
not I_8385 (I145563,I145614);
not I_8386 (I145636,I145597);
DFFARX1 I_8387 (I375303,I3035,I145571,I145662,);
not I_8388 (I145670,I145662);
and I_8389 (I145687,I145636,I375309);
not I_8390 (I145704,I375294);
nand I_8391 (I145721,I145704,I375309);
not I_8392 (I145738,I375297);
nor I_8393 (I145755,I145738,I375318);
nand I_8394 (I145772,I145755,I375315);
nor I_8395 (I145789,I145772,I145721);
DFFARX1 I_8396 (I145789,I3035,I145571,I145539,);
not I_8397 (I145820,I145772);
not I_8398 (I145837,I375318);
nand I_8399 (I145854,I145837,I375309);
nor I_8400 (I145871,I375318,I375294);
nand I_8401 (I145551,I145687,I145871);
nand I_8402 (I145545,I145636,I375318);
nand I_8403 (I145916,I145738,I375294);
DFFARX1 I_8404 (I145916,I3035,I145571,I145560,);
DFFARX1 I_8405 (I145916,I3035,I145571,I145554,);
not I_8406 (I145961,I375294);
nor I_8407 (I145978,I145961,I375300);
and I_8408 (I145995,I145978,I375312);
or I_8409 (I146012,I145995,I375297);
DFFARX1 I_8410 (I146012,I3035,I145571,I146038,);
nand I_8411 (I146046,I146038,I145704);
nor I_8412 (I145548,I146046,I145854);
nor I_8413 (I145542,I146038,I145670);
DFFARX1 I_8414 (I146038,I3035,I145571,I146100,);
not I_8415 (I146108,I146100);
nor I_8416 (I145557,I146108,I145820);
not I_8417 (I146166,I3042);
DFFARX1 I_8418 (I474614,I3035,I146166,I146192,);
DFFARX1 I_8419 (I146192,I3035,I146166,I146209,);
not I_8420 (I146158,I146209);
not I_8421 (I146231,I146192);
DFFARX1 I_8422 (I474608,I3035,I146166,I146257,);
not I_8423 (I146265,I146257);
and I_8424 (I146282,I146231,I474626);
not I_8425 (I146299,I474614);
nand I_8426 (I146316,I146299,I474626);
not I_8427 (I146333,I474608);
nor I_8428 (I146350,I146333,I474620);
nand I_8429 (I146367,I146350,I474611);
nor I_8430 (I146384,I146367,I146316);
DFFARX1 I_8431 (I146384,I3035,I146166,I146134,);
not I_8432 (I146415,I146367);
not I_8433 (I146432,I474620);
nand I_8434 (I146449,I146432,I474626);
nor I_8435 (I146466,I474620,I474614);
nand I_8436 (I146146,I146282,I146466);
nand I_8437 (I146140,I146231,I474620);
nand I_8438 (I146511,I146333,I474623);
DFFARX1 I_8439 (I146511,I3035,I146166,I146155,);
DFFARX1 I_8440 (I146511,I3035,I146166,I146149,);
not I_8441 (I146556,I474623);
nor I_8442 (I146573,I146556,I474629);
and I_8443 (I146590,I146573,I474611);
or I_8444 (I146607,I146590,I474617);
DFFARX1 I_8445 (I146607,I3035,I146166,I146633,);
nand I_8446 (I146641,I146633,I146299);
nor I_8447 (I146143,I146641,I146449);
nor I_8448 (I146137,I146633,I146265);
DFFARX1 I_8449 (I146633,I3035,I146166,I146695,);
not I_8450 (I146703,I146695);
nor I_8451 (I146152,I146703,I146415);
not I_8452 (I146761,I3042);
DFFARX1 I_8453 (I75942,I3035,I146761,I146787,);
DFFARX1 I_8454 (I146787,I3035,I146761,I146804,);
not I_8455 (I146753,I146804);
not I_8456 (I146826,I146787);
DFFARX1 I_8457 (I75927,I3035,I146761,I146852,);
not I_8458 (I146860,I146852);
and I_8459 (I146877,I146826,I75948);
not I_8460 (I146894,I75939);
nand I_8461 (I146911,I146894,I75948);
not I_8462 (I146928,I75924);
nor I_8463 (I146945,I146928,I75936);
nand I_8464 (I146962,I146945,I75951);
nor I_8465 (I146979,I146962,I146911);
DFFARX1 I_8466 (I146979,I3035,I146761,I146729,);
not I_8467 (I147010,I146962);
not I_8468 (I147027,I75936);
nand I_8469 (I147044,I147027,I75948);
nor I_8470 (I147061,I75936,I75939);
nand I_8471 (I146741,I146877,I147061);
nand I_8472 (I146735,I146826,I75936);
nand I_8473 (I147106,I146928,I75930);
DFFARX1 I_8474 (I147106,I3035,I146761,I146750,);
DFFARX1 I_8475 (I147106,I3035,I146761,I146744,);
not I_8476 (I147151,I75930);
nor I_8477 (I147168,I147151,I75933);
and I_8478 (I147185,I147168,I75924);
or I_8479 (I147202,I147185,I75945);
DFFARX1 I_8480 (I147202,I3035,I146761,I147228,);
nand I_8481 (I147236,I147228,I146894);
nor I_8482 (I146738,I147236,I147044);
nor I_8483 (I146732,I147228,I146860);
DFFARX1 I_8484 (I147228,I3035,I146761,I147290,);
not I_8485 (I147298,I147290);
nor I_8486 (I146747,I147298,I147010);
not I_8487 (I147356,I3042);
DFFARX1 I_8488 (I693884,I3035,I147356,I147382,);
DFFARX1 I_8489 (I147382,I3035,I147356,I147399,);
not I_8490 (I147348,I147399);
not I_8491 (I147421,I147382);
DFFARX1 I_8492 (I693857,I3035,I147356,I147447,);
not I_8493 (I147455,I147447);
and I_8494 (I147472,I147421,I693881);
not I_8495 (I147489,I693878);
nand I_8496 (I147506,I147489,I693881);
not I_8497 (I147523,I693857);
nor I_8498 (I147540,I147523,I693875);
nand I_8499 (I147557,I147540,I693863);
nor I_8500 (I147574,I147557,I147506);
DFFARX1 I_8501 (I147574,I3035,I147356,I147324,);
not I_8502 (I147605,I147557);
not I_8503 (I147622,I693875);
nand I_8504 (I147639,I147622,I693881);
nor I_8505 (I147656,I693875,I693878);
nand I_8506 (I147336,I147472,I147656);
nand I_8507 (I147330,I147421,I693875);
nand I_8508 (I147701,I147523,I693869);
DFFARX1 I_8509 (I147701,I3035,I147356,I147345,);
DFFARX1 I_8510 (I147701,I3035,I147356,I147339,);
not I_8511 (I147746,I693869);
nor I_8512 (I147763,I147746,I693872);
and I_8513 (I147780,I147763,I693860);
or I_8514 (I147797,I147780,I693866);
DFFARX1 I_8515 (I147797,I3035,I147356,I147823,);
nand I_8516 (I147831,I147823,I147489);
nor I_8517 (I147333,I147831,I147639);
nor I_8518 (I147327,I147823,I147455);
DFFARX1 I_8519 (I147823,I3035,I147356,I147885,);
not I_8520 (I147893,I147885);
nor I_8521 (I147342,I147893,I147605);
not I_8522 (I147951,I3042);
DFFARX1 I_8523 (I630668,I3035,I147951,I147977,);
DFFARX1 I_8524 (I147977,I3035,I147951,I147994,);
not I_8525 (I147943,I147994);
not I_8526 (I148016,I147977);
DFFARX1 I_8527 (I630668,I3035,I147951,I148042,);
not I_8528 (I148050,I148042);
and I_8529 (I148067,I148016,I630671);
not I_8530 (I148084,I630683);
nand I_8531 (I148101,I148084,I630671);
not I_8532 (I148118,I630689);
nor I_8533 (I148135,I148118,I630680);
nand I_8534 (I148152,I148135,I630686);
nor I_8535 (I148169,I148152,I148101);
DFFARX1 I_8536 (I148169,I3035,I147951,I147919,);
not I_8537 (I148200,I148152);
not I_8538 (I148217,I630680);
nand I_8539 (I148234,I148217,I630671);
nor I_8540 (I148251,I630680,I630683);
nand I_8541 (I147931,I148067,I148251);
nand I_8542 (I147925,I148016,I630680);
nand I_8543 (I148296,I148118,I630677);
DFFARX1 I_8544 (I148296,I3035,I147951,I147940,);
DFFARX1 I_8545 (I148296,I3035,I147951,I147934,);
not I_8546 (I148341,I630677);
nor I_8547 (I148358,I148341,I630674);
and I_8548 (I148375,I148358,I630692);
or I_8549 (I148392,I148375,I630671);
DFFARX1 I_8550 (I148392,I3035,I147951,I148418,);
nand I_8551 (I148426,I148418,I148084);
nor I_8552 (I147928,I148426,I148234);
nor I_8553 (I147922,I148418,I148050);
DFFARX1 I_8554 (I148418,I3035,I147951,I148480,);
not I_8555 (I148488,I148480);
nor I_8556 (I147937,I148488,I148200);
not I_8557 (I148546,I3042);
DFFARX1 I_8558 (I510969,I3035,I148546,I148572,);
DFFARX1 I_8559 (I148572,I3035,I148546,I148589,);
not I_8560 (I148538,I148589);
not I_8561 (I148611,I148572);
DFFARX1 I_8562 (I510978,I3035,I148546,I148637,);
not I_8563 (I148645,I148637);
and I_8564 (I148662,I148611,I510966);
not I_8565 (I148679,I510957);
nand I_8566 (I148696,I148679,I510966);
not I_8567 (I148713,I510963);
nor I_8568 (I148730,I148713,I510981);
nand I_8569 (I148747,I148730,I510954);
nor I_8570 (I148764,I148747,I148696);
DFFARX1 I_8571 (I148764,I3035,I148546,I148514,);
not I_8572 (I148795,I148747);
not I_8573 (I148812,I510981);
nand I_8574 (I148829,I148812,I510966);
nor I_8575 (I148846,I510981,I510957);
nand I_8576 (I148526,I148662,I148846);
nand I_8577 (I148520,I148611,I510981);
nand I_8578 (I148891,I148713,I510960);
DFFARX1 I_8579 (I148891,I3035,I148546,I148535,);
DFFARX1 I_8580 (I148891,I3035,I148546,I148529,);
not I_8581 (I148936,I510960);
nor I_8582 (I148953,I148936,I510972);
and I_8583 (I148970,I148953,I510954);
or I_8584 (I148987,I148970,I510975);
DFFARX1 I_8585 (I148987,I3035,I148546,I149013,);
nand I_8586 (I149021,I149013,I148679);
nor I_8587 (I148523,I149021,I148829);
nor I_8588 (I148517,I149013,I148645);
DFFARX1 I_8589 (I149013,I3035,I148546,I149075,);
not I_8590 (I149083,I149075);
nor I_8591 (I148532,I149083,I148795);
not I_8592 (I149141,I3042);
DFFARX1 I_8593 (I538747,I3035,I149141,I149167,);
DFFARX1 I_8594 (I149167,I3035,I149141,I149184,);
not I_8595 (I149133,I149184);
not I_8596 (I149206,I149167);
DFFARX1 I_8597 (I538756,I3035,I149141,I149232,);
not I_8598 (I149240,I149232);
and I_8599 (I149257,I149206,I538744);
not I_8600 (I149274,I538735);
nand I_8601 (I149291,I149274,I538744);
not I_8602 (I149308,I538741);
nor I_8603 (I149325,I149308,I538759);
nand I_8604 (I149342,I149325,I538732);
nor I_8605 (I149359,I149342,I149291);
DFFARX1 I_8606 (I149359,I3035,I149141,I149109,);
not I_8607 (I149390,I149342);
not I_8608 (I149407,I538759);
nand I_8609 (I149424,I149407,I538744);
nor I_8610 (I149441,I538759,I538735);
nand I_8611 (I149121,I149257,I149441);
nand I_8612 (I149115,I149206,I538759);
nand I_8613 (I149486,I149308,I538738);
DFFARX1 I_8614 (I149486,I3035,I149141,I149130,);
DFFARX1 I_8615 (I149486,I3035,I149141,I149124,);
not I_8616 (I149531,I538738);
nor I_8617 (I149548,I149531,I538750);
and I_8618 (I149565,I149548,I538732);
or I_8619 (I149582,I149565,I538753);
DFFARX1 I_8620 (I149582,I3035,I149141,I149608,);
nand I_8621 (I149616,I149608,I149274);
nor I_8622 (I149118,I149616,I149424);
nor I_8623 (I149112,I149608,I149240);
DFFARX1 I_8624 (I149608,I3035,I149141,I149670,);
not I_8625 (I149678,I149670);
nor I_8626 (I149127,I149678,I149390);
not I_8627 (I149736,I3042);
DFFARX1 I_8628 (I205107,I3035,I149736,I149762,);
DFFARX1 I_8629 (I149762,I3035,I149736,I149779,);
not I_8630 (I149728,I149779);
not I_8631 (I149801,I149762);
DFFARX1 I_8632 (I205122,I3035,I149736,I149827,);
not I_8633 (I149835,I149827);
and I_8634 (I149852,I149801,I205119);
not I_8635 (I149869,I205107);
nand I_8636 (I149886,I149869,I205119);
not I_8637 (I149903,I205116);
nor I_8638 (I149920,I149903,I205131);
nand I_8639 (I149937,I149920,I205128);
nor I_8640 (I149954,I149937,I149886);
DFFARX1 I_8641 (I149954,I3035,I149736,I149704,);
not I_8642 (I149985,I149937);
not I_8643 (I150002,I205131);
nand I_8644 (I150019,I150002,I205119);
nor I_8645 (I150036,I205131,I205107);
nand I_8646 (I149716,I149852,I150036);
nand I_8647 (I149710,I149801,I205131);
nand I_8648 (I150081,I149903,I205125);
DFFARX1 I_8649 (I150081,I3035,I149736,I149725,);
DFFARX1 I_8650 (I150081,I3035,I149736,I149719,);
not I_8651 (I150126,I205125);
nor I_8652 (I150143,I150126,I205113);
and I_8653 (I150160,I150143,I205134);
or I_8654 (I150177,I150160,I205110);
DFFARX1 I_8655 (I150177,I3035,I149736,I150203,);
nand I_8656 (I150211,I150203,I149869);
nor I_8657 (I149713,I150211,I150019);
nor I_8658 (I149707,I150203,I149835);
DFFARX1 I_8659 (I150203,I3035,I149736,I150265,);
not I_8660 (I150273,I150265);
nor I_8661 (I149722,I150273,I149985);
not I_8662 (I150334,I3042);
DFFARX1 I_8663 (I542611,I3035,I150334,I150360,);
nand I_8664 (I150368,I542608,I542626);
and I_8665 (I150385,I150368,I542617);
DFFARX1 I_8666 (I150385,I3035,I150334,I150411,);
nor I_8667 (I150302,I150411,I150360);
not I_8668 (I150433,I150411);
DFFARX1 I_8669 (I542632,I3035,I150334,I150459,);
nand I_8670 (I150467,I150459,I542614);
not I_8671 (I150484,I150467);
DFFARX1 I_8672 (I150484,I3035,I150334,I150510,);
not I_8673 (I150326,I150510);
nor I_8674 (I150532,I150360,I150467);
nor I_8675 (I150308,I150411,I150532);
DFFARX1 I_8676 (I542620,I3035,I150334,I150572,);
DFFARX1 I_8677 (I150572,I3035,I150334,I150589,);
not I_8678 (I150597,I150589);
not I_8679 (I150614,I150572);
nand I_8680 (I150311,I150614,I150433);
nand I_8681 (I150645,I542608,I542635);
and I_8682 (I150662,I150645,I542623);
DFFARX1 I_8683 (I150662,I3035,I150334,I150688,);
nor I_8684 (I150696,I150688,I150360);
DFFARX1 I_8685 (I150696,I3035,I150334,I150299,);
DFFARX1 I_8686 (I150688,I3035,I150334,I150317,);
nor I_8687 (I150741,I542629,I542635);
not I_8688 (I150758,I150741);
nor I_8689 (I150320,I150597,I150758);
nand I_8690 (I150305,I150614,I150758);
nor I_8691 (I150314,I150360,I150741);
DFFARX1 I_8692 (I150741,I3035,I150334,I150323,);
not I_8693 (I150861,I3042);
DFFARX1 I_8694 (I445099,I3035,I150861,I150887,);
nand I_8695 (I150895,I445102,I445096);
and I_8696 (I150912,I150895,I445108);
DFFARX1 I_8697 (I150912,I3035,I150861,I150938,);
nor I_8698 (I150829,I150938,I150887);
not I_8699 (I150960,I150938);
DFFARX1 I_8700 (I445111,I3035,I150861,I150986,);
nand I_8701 (I150994,I150986,I445102);
not I_8702 (I151011,I150994);
DFFARX1 I_8703 (I151011,I3035,I150861,I151037,);
not I_8704 (I150853,I151037);
nor I_8705 (I151059,I150887,I150994);
nor I_8706 (I150835,I150938,I151059);
DFFARX1 I_8707 (I445114,I3035,I150861,I151099,);
DFFARX1 I_8708 (I151099,I3035,I150861,I151116,);
not I_8709 (I151124,I151116);
not I_8710 (I151141,I151099);
nand I_8711 (I150838,I151141,I150960);
nand I_8712 (I151172,I445096,I445105);
and I_8713 (I151189,I151172,I445099);
DFFARX1 I_8714 (I151189,I3035,I150861,I151215,);
nor I_8715 (I151223,I151215,I150887);
DFFARX1 I_8716 (I151223,I3035,I150861,I150826,);
DFFARX1 I_8717 (I151215,I3035,I150861,I150844,);
nor I_8718 (I151268,I445117,I445105);
not I_8719 (I151285,I151268);
nor I_8720 (I150847,I151124,I151285);
nand I_8721 (I150832,I151141,I151285);
nor I_8722 (I150841,I150887,I151268);
DFFARX1 I_8723 (I151268,I3035,I150861,I150850,);
not I_8724 (I151388,I3042);
DFFARX1 I_8725 (I291844,I3035,I151388,I151414,);
nand I_8726 (I151422,I291844,I291856);
and I_8727 (I151439,I151422,I291841);
DFFARX1 I_8728 (I151439,I3035,I151388,I151465,);
nor I_8729 (I151356,I151465,I151414);
not I_8730 (I151487,I151465);
DFFARX1 I_8731 (I291865,I3035,I151388,I151513,);
nand I_8732 (I151521,I151513,I291862);
not I_8733 (I151538,I151521);
DFFARX1 I_8734 (I151538,I3035,I151388,I151564,);
not I_8735 (I151380,I151564);
nor I_8736 (I151586,I151414,I151521);
nor I_8737 (I151362,I151465,I151586);
DFFARX1 I_8738 (I291853,I3035,I151388,I151626,);
DFFARX1 I_8739 (I151626,I3035,I151388,I151643,);
not I_8740 (I151651,I151643);
not I_8741 (I151668,I151626);
nand I_8742 (I151365,I151668,I151487);
nand I_8743 (I151699,I291841,I291850);
and I_8744 (I151716,I151699,I291859);
DFFARX1 I_8745 (I151716,I3035,I151388,I151742,);
nor I_8746 (I151750,I151742,I151414);
DFFARX1 I_8747 (I151750,I3035,I151388,I151353,);
DFFARX1 I_8748 (I151742,I3035,I151388,I151371,);
nor I_8749 (I151795,I291847,I291850);
not I_8750 (I151812,I151795);
nor I_8751 (I151374,I151651,I151812);
nand I_8752 (I151359,I151668,I151812);
nor I_8753 (I151368,I151414,I151795);
DFFARX1 I_8754 (I151795,I3035,I151388,I151377,);
not I_8755 (I151915,I3042);
DFFARX1 I_8756 (I471449,I3035,I151915,I151941,);
nand I_8757 (I151949,I471452,I471446);
and I_8758 (I151966,I151949,I471458);
DFFARX1 I_8759 (I151966,I3035,I151915,I151992,);
nor I_8760 (I151883,I151992,I151941);
not I_8761 (I152014,I151992);
DFFARX1 I_8762 (I471461,I3035,I151915,I152040,);
nand I_8763 (I152048,I152040,I471452);
not I_8764 (I152065,I152048);
DFFARX1 I_8765 (I152065,I3035,I151915,I152091,);
not I_8766 (I151907,I152091);
nor I_8767 (I152113,I151941,I152048);
nor I_8768 (I151889,I151992,I152113);
DFFARX1 I_8769 (I471464,I3035,I151915,I152153,);
DFFARX1 I_8770 (I152153,I3035,I151915,I152170,);
not I_8771 (I152178,I152170);
not I_8772 (I152195,I152153);
nand I_8773 (I151892,I152195,I152014);
nand I_8774 (I152226,I471446,I471455);
and I_8775 (I152243,I152226,I471449);
DFFARX1 I_8776 (I152243,I3035,I151915,I152269,);
nor I_8777 (I152277,I152269,I151941);
DFFARX1 I_8778 (I152277,I3035,I151915,I151880,);
DFFARX1 I_8779 (I152269,I3035,I151915,I151898,);
nor I_8780 (I152322,I471467,I471455);
not I_8781 (I152339,I152322);
nor I_8782 (I151901,I152178,I152339);
nand I_8783 (I151886,I152195,I152339);
nor I_8784 (I151895,I151941,I152322);
DFFARX1 I_8785 (I152322,I3035,I151915,I151904,);
not I_8786 (I152442,I3042);
DFFARX1 I_8787 (I291249,I3035,I152442,I152468,);
nand I_8788 (I152476,I291249,I291261);
and I_8789 (I152493,I152476,I291246);
DFFARX1 I_8790 (I152493,I3035,I152442,I152519,);
nor I_8791 (I152410,I152519,I152468);
not I_8792 (I152541,I152519);
DFFARX1 I_8793 (I291270,I3035,I152442,I152567,);
nand I_8794 (I152575,I152567,I291267);
not I_8795 (I152592,I152575);
DFFARX1 I_8796 (I152592,I3035,I152442,I152618,);
not I_8797 (I152434,I152618);
nor I_8798 (I152640,I152468,I152575);
nor I_8799 (I152416,I152519,I152640);
DFFARX1 I_8800 (I291258,I3035,I152442,I152680,);
DFFARX1 I_8801 (I152680,I3035,I152442,I152697,);
not I_8802 (I152705,I152697);
not I_8803 (I152722,I152680);
nand I_8804 (I152419,I152722,I152541);
nand I_8805 (I152753,I291246,I291255);
and I_8806 (I152770,I152753,I291264);
DFFARX1 I_8807 (I152770,I3035,I152442,I152796,);
nor I_8808 (I152804,I152796,I152468);
DFFARX1 I_8809 (I152804,I3035,I152442,I152407,);
DFFARX1 I_8810 (I152796,I3035,I152442,I152425,);
nor I_8811 (I152849,I291252,I291255);
not I_8812 (I152866,I152849);
nor I_8813 (I152428,I152705,I152866);
nand I_8814 (I152413,I152722,I152866);
nor I_8815 (I152422,I152468,I152849);
DFFARX1 I_8816 (I152849,I3035,I152442,I152431,);
not I_8817 (I152969,I3042);
DFFARX1 I_8818 (I690421,I3035,I152969,I152995,);
nand I_8819 (I153003,I690418,I690409);
and I_8820 (I153020,I153003,I690406);
DFFARX1 I_8821 (I153020,I3035,I152969,I153046,);
nor I_8822 (I152937,I153046,I152995);
not I_8823 (I153068,I153046);
DFFARX1 I_8824 (I690415,I3035,I152969,I153094,);
nand I_8825 (I153102,I153094,I690424);
not I_8826 (I153119,I153102);
DFFARX1 I_8827 (I153119,I3035,I152969,I153145,);
not I_8828 (I152961,I153145);
nor I_8829 (I153167,I152995,I153102);
nor I_8830 (I152943,I153046,I153167);
DFFARX1 I_8831 (I690427,I3035,I152969,I153207,);
DFFARX1 I_8832 (I153207,I3035,I152969,I153224,);
not I_8833 (I153232,I153224);
not I_8834 (I153249,I153207);
nand I_8835 (I152946,I153249,I153068);
nand I_8836 (I153280,I690406,I690412);
and I_8837 (I153297,I153280,I690430);
DFFARX1 I_8838 (I153297,I3035,I152969,I153323,);
nor I_8839 (I153331,I153323,I152995);
DFFARX1 I_8840 (I153331,I3035,I152969,I152934,);
DFFARX1 I_8841 (I153323,I3035,I152969,I152952,);
nor I_8842 (I153376,I690409,I690412);
not I_8843 (I153393,I153376);
nor I_8844 (I152955,I153232,I153393);
nand I_8845 (I152940,I153249,I153393);
nor I_8846 (I152949,I152995,I153376);
DFFARX1 I_8847 (I153376,I3035,I152969,I152958,);
not I_8848 (I153496,I3042);
DFFARX1 I_8849 (I458801,I3035,I153496,I153522,);
nand I_8850 (I153530,I458804,I458798);
and I_8851 (I153547,I153530,I458810);
DFFARX1 I_8852 (I153547,I3035,I153496,I153573,);
nor I_8853 (I153464,I153573,I153522);
not I_8854 (I153595,I153573);
DFFARX1 I_8855 (I458813,I3035,I153496,I153621,);
nand I_8856 (I153629,I153621,I458804);
not I_8857 (I153646,I153629);
DFFARX1 I_8858 (I153646,I3035,I153496,I153672,);
not I_8859 (I153488,I153672);
nor I_8860 (I153694,I153522,I153629);
nor I_8861 (I153470,I153573,I153694);
DFFARX1 I_8862 (I458816,I3035,I153496,I153734,);
DFFARX1 I_8863 (I153734,I3035,I153496,I153751,);
not I_8864 (I153759,I153751);
not I_8865 (I153776,I153734);
nand I_8866 (I153473,I153776,I153595);
nand I_8867 (I153807,I458798,I458807);
and I_8868 (I153824,I153807,I458801);
DFFARX1 I_8869 (I153824,I3035,I153496,I153850,);
nor I_8870 (I153858,I153850,I153522);
DFFARX1 I_8871 (I153858,I3035,I153496,I153461,);
DFFARX1 I_8872 (I153850,I3035,I153496,I153479,);
nor I_8873 (I153903,I458819,I458807);
not I_8874 (I153920,I153903);
nor I_8875 (I153482,I153759,I153920);
nand I_8876 (I153467,I153776,I153920);
nor I_8877 (I153476,I153522,I153903);
DFFARX1 I_8878 (I153903,I3035,I153496,I153485,);
not I_8879 (I154023,I3042);
DFFARX1 I_8880 (I737109,I3035,I154023,I154049,);
nand I_8881 (I154057,I737088,I737088);
and I_8882 (I154074,I154057,I737115);
DFFARX1 I_8883 (I154074,I3035,I154023,I154100,);
nor I_8884 (I153991,I154100,I154049);
not I_8885 (I154122,I154100);
DFFARX1 I_8886 (I737103,I3035,I154023,I154148,);
nand I_8887 (I154156,I154148,I737106);
not I_8888 (I154173,I154156);
DFFARX1 I_8889 (I154173,I3035,I154023,I154199,);
not I_8890 (I154015,I154199);
nor I_8891 (I154221,I154049,I154156);
nor I_8892 (I153997,I154100,I154221);
DFFARX1 I_8893 (I737097,I3035,I154023,I154261,);
DFFARX1 I_8894 (I154261,I3035,I154023,I154278,);
not I_8895 (I154286,I154278);
not I_8896 (I154303,I154261);
nand I_8897 (I154000,I154303,I154122);
nand I_8898 (I154334,I737094,I737091);
and I_8899 (I154351,I154334,I737112);
DFFARX1 I_8900 (I154351,I3035,I154023,I154377,);
nor I_8901 (I154385,I154377,I154049);
DFFARX1 I_8902 (I154385,I3035,I154023,I153988,);
DFFARX1 I_8903 (I154377,I3035,I154023,I154006,);
nor I_8904 (I154430,I737100,I737091);
not I_8905 (I154447,I154430);
nor I_8906 (I154009,I154286,I154447);
nand I_8907 (I153994,I154303,I154447);
nor I_8908 (I154003,I154049,I154430);
DFFARX1 I_8909 (I154430,I3035,I154023,I154012,);
not I_8910 (I154550,I3042);
DFFARX1 I_8911 (I658872,I3035,I154550,I154576,);
nand I_8912 (I154584,I658854,I658878);
and I_8913 (I154601,I154584,I658869);
DFFARX1 I_8914 (I154601,I3035,I154550,I154627,);
nor I_8915 (I154518,I154627,I154576);
not I_8916 (I154649,I154627);
DFFARX1 I_8917 (I658875,I3035,I154550,I154675,);
nand I_8918 (I154683,I154675,I658863);
not I_8919 (I154700,I154683);
DFFARX1 I_8920 (I154700,I3035,I154550,I154726,);
not I_8921 (I154542,I154726);
nor I_8922 (I154748,I154576,I154683);
nor I_8923 (I154524,I154627,I154748);
DFFARX1 I_8924 (I658854,I3035,I154550,I154788,);
DFFARX1 I_8925 (I154788,I3035,I154550,I154805,);
not I_8926 (I154813,I154805);
not I_8927 (I154830,I154788);
nand I_8928 (I154527,I154830,I154649);
nand I_8929 (I154861,I658860,I658857);
and I_8930 (I154878,I154861,I658866);
DFFARX1 I_8931 (I154878,I3035,I154550,I154904,);
nor I_8932 (I154912,I154904,I154576);
DFFARX1 I_8933 (I154912,I3035,I154550,I154515,);
DFFARX1 I_8934 (I154904,I3035,I154550,I154533,);
nor I_8935 (I154957,I658857,I658857);
not I_8936 (I154974,I154957);
nor I_8937 (I154536,I154813,I154974);
nand I_8938 (I154521,I154830,I154974);
nor I_8939 (I154530,I154576,I154957);
DFFARX1 I_8940 (I154957,I3035,I154550,I154539,);
not I_8941 (I155077,I3042);
DFFARX1 I_8942 (I14656,I3035,I155077,I155103,);
nand I_8943 (I155111,I14680,I14659);
and I_8944 (I155128,I155111,I14656);
DFFARX1 I_8945 (I155128,I3035,I155077,I155154,);
nor I_8946 (I155045,I155154,I155103);
not I_8947 (I155176,I155154);
DFFARX1 I_8948 (I14662,I3035,I155077,I155202,);
nand I_8949 (I155210,I155202,I14671);
not I_8950 (I155227,I155210);
DFFARX1 I_8951 (I155227,I3035,I155077,I155253,);
not I_8952 (I155069,I155253);
nor I_8953 (I155275,I155103,I155210);
nor I_8954 (I155051,I155154,I155275);
DFFARX1 I_8955 (I14665,I3035,I155077,I155315,);
DFFARX1 I_8956 (I155315,I3035,I155077,I155332,);
not I_8957 (I155340,I155332);
not I_8958 (I155357,I155315);
nand I_8959 (I155054,I155357,I155176);
nand I_8960 (I155388,I14677,I14659);
and I_8961 (I155405,I155388,I14668);
DFFARX1 I_8962 (I155405,I3035,I155077,I155431,);
nor I_8963 (I155439,I155431,I155103);
DFFARX1 I_8964 (I155439,I3035,I155077,I155042,);
DFFARX1 I_8965 (I155431,I3035,I155077,I155060,);
nor I_8966 (I155484,I14674,I14659);
not I_8967 (I155501,I155484);
nor I_8968 (I155063,I155340,I155501);
nand I_8969 (I155048,I155357,I155501);
nor I_8970 (I155057,I155103,I155484);
DFFARX1 I_8971 (I155484,I3035,I155077,I155066,);
not I_8972 (I155604,I3042);
DFFARX1 I_8973 (I619686,I3035,I155604,I155630,);
nand I_8974 (I155638,I619701,I619686);
and I_8975 (I155655,I155638,I619704);
DFFARX1 I_8976 (I155655,I3035,I155604,I155681,);
nor I_8977 (I155572,I155681,I155630);
not I_8978 (I155703,I155681);
DFFARX1 I_8979 (I619710,I3035,I155604,I155729,);
nand I_8980 (I155737,I155729,I619692);
not I_8981 (I155754,I155737);
DFFARX1 I_8982 (I155754,I3035,I155604,I155780,);
not I_8983 (I155596,I155780);
nor I_8984 (I155802,I155630,I155737);
nor I_8985 (I155578,I155681,I155802);
DFFARX1 I_8986 (I619689,I3035,I155604,I155842,);
DFFARX1 I_8987 (I155842,I3035,I155604,I155859,);
not I_8988 (I155867,I155859);
not I_8989 (I155884,I155842);
nand I_8990 (I155581,I155884,I155703);
nand I_8991 (I155915,I619689,I619695);
and I_8992 (I155932,I155915,I619707);
DFFARX1 I_8993 (I155932,I3035,I155604,I155958,);
nor I_8994 (I155966,I155958,I155630);
DFFARX1 I_8995 (I155966,I3035,I155604,I155569,);
DFFARX1 I_8996 (I155958,I3035,I155604,I155587,);
nor I_8997 (I156011,I619698,I619695);
not I_8998 (I156028,I156011);
nor I_8999 (I155590,I155867,I156028);
nand I_9000 (I155575,I155884,I156028);
nor I_9001 (I155584,I155630,I156011);
DFFARX1 I_9002 (I156011,I3035,I155604,I155593,);
not I_9003 (I156131,I3042);
DFFARX1 I_9004 (I1436,I3035,I156131,I156157,);
nand I_9005 (I156165,I1540,I1556);
and I_9006 (I156182,I156165,I1708);
DFFARX1 I_9007 (I156182,I3035,I156131,I156208,);
nor I_9008 (I156099,I156208,I156157);
not I_9009 (I156230,I156208);
DFFARX1 I_9010 (I2092,I3035,I156131,I156256,);
nand I_9011 (I156264,I156256,I1900);
not I_9012 (I156281,I156264);
DFFARX1 I_9013 (I156281,I3035,I156131,I156307,);
not I_9014 (I156123,I156307);
nor I_9015 (I156329,I156157,I156264);
nor I_9016 (I156105,I156208,I156329);
DFFARX1 I_9017 (I2476,I3035,I156131,I156369,);
DFFARX1 I_9018 (I156369,I3035,I156131,I156386,);
not I_9019 (I156394,I156386);
not I_9020 (I156411,I156369);
nand I_9021 (I156108,I156411,I156230);
nand I_9022 (I156442,I2772,I3020);
and I_9023 (I156459,I156442,I2196);
DFFARX1 I_9024 (I156459,I3035,I156131,I156485,);
nor I_9025 (I156493,I156485,I156157);
DFFARX1 I_9026 (I156493,I3035,I156131,I156096,);
DFFARX1 I_9027 (I156485,I3035,I156131,I156114,);
nor I_9028 (I156538,I1460,I3020);
not I_9029 (I156555,I156538);
nor I_9030 (I156117,I156394,I156555);
nand I_9031 (I156102,I156411,I156555);
nor I_9032 (I156111,I156157,I156538);
DFFARX1 I_9033 (I156538,I3035,I156131,I156120,);
not I_9034 (I156658,I3042);
DFFARX1 I_9035 (I93179,I3035,I156658,I156684,);
nand I_9036 (I156692,I93179,I93185);
and I_9037 (I156709,I156692,I93203);
DFFARX1 I_9038 (I156709,I3035,I156658,I156735,);
nor I_9039 (I156626,I156735,I156684);
not I_9040 (I156757,I156735);
DFFARX1 I_9041 (I93191,I3035,I156658,I156783,);
nand I_9042 (I156791,I156783,I93188);
not I_9043 (I156808,I156791);
DFFARX1 I_9044 (I156808,I3035,I156658,I156834,);
not I_9045 (I156650,I156834);
nor I_9046 (I156856,I156684,I156791);
nor I_9047 (I156632,I156735,I156856);
DFFARX1 I_9048 (I93197,I3035,I156658,I156896,);
DFFARX1 I_9049 (I156896,I3035,I156658,I156913,);
not I_9050 (I156921,I156913);
not I_9051 (I156938,I156896);
nand I_9052 (I156635,I156938,I156757);
nand I_9053 (I156969,I93182,I93182);
and I_9054 (I156986,I156969,I93194);
DFFARX1 I_9055 (I156986,I3035,I156658,I157012,);
nor I_9056 (I157020,I157012,I156684);
DFFARX1 I_9057 (I157020,I3035,I156658,I156623,);
DFFARX1 I_9058 (I157012,I3035,I156658,I156641,);
nor I_9059 (I157065,I93200,I93182);
not I_9060 (I157082,I157065);
nor I_9061 (I156644,I156921,I157082);
nand I_9062 (I156629,I156938,I157082);
nor I_9063 (I156638,I156684,I157065);
DFFARX1 I_9064 (I157065,I3035,I156658,I156647,);
not I_9065 (I157185,I3042);
DFFARX1 I_9066 (I725804,I3035,I157185,I157211,);
nand I_9067 (I157219,I725783,I725783);
and I_9068 (I157236,I157219,I725810);
DFFARX1 I_9069 (I157236,I3035,I157185,I157262,);
nor I_9070 (I157153,I157262,I157211);
not I_9071 (I157284,I157262);
DFFARX1 I_9072 (I725798,I3035,I157185,I157310,);
nand I_9073 (I157318,I157310,I725801);
not I_9074 (I157335,I157318);
DFFARX1 I_9075 (I157335,I3035,I157185,I157361,);
not I_9076 (I157177,I157361);
nor I_9077 (I157383,I157211,I157318);
nor I_9078 (I157159,I157262,I157383);
DFFARX1 I_9079 (I725792,I3035,I157185,I157423,);
DFFARX1 I_9080 (I157423,I3035,I157185,I157440,);
not I_9081 (I157448,I157440);
not I_9082 (I157465,I157423);
nand I_9083 (I157162,I157465,I157284);
nand I_9084 (I157496,I725789,I725786);
and I_9085 (I157513,I157496,I725807);
DFFARX1 I_9086 (I157513,I3035,I157185,I157539,);
nor I_9087 (I157547,I157539,I157211);
DFFARX1 I_9088 (I157547,I3035,I157185,I157150,);
DFFARX1 I_9089 (I157539,I3035,I157185,I157168,);
nor I_9090 (I157592,I725795,I725786);
not I_9091 (I157609,I157592);
nor I_9092 (I157171,I157448,I157609);
nand I_9093 (I157156,I157465,I157609);
nor I_9094 (I157165,I157211,I157592);
DFFARX1 I_9095 (I157592,I3035,I157185,I157174,);
not I_9096 (I157712,I3042);
DFFARX1 I_9097 (I234801,I3035,I157712,I157738,);
nand I_9098 (I157746,I234813,I234792);
and I_9099 (I157763,I157746,I234816);
DFFARX1 I_9100 (I157763,I3035,I157712,I157789,);
nor I_9101 (I157680,I157789,I157738);
not I_9102 (I157811,I157789);
DFFARX1 I_9103 (I234807,I3035,I157712,I157837,);
nand I_9104 (I157845,I157837,I234789);
not I_9105 (I157862,I157845);
DFFARX1 I_9106 (I157862,I3035,I157712,I157888,);
not I_9107 (I157704,I157888);
nor I_9108 (I157910,I157738,I157845);
nor I_9109 (I157686,I157789,I157910);
DFFARX1 I_9110 (I234804,I3035,I157712,I157950,);
DFFARX1 I_9111 (I157950,I3035,I157712,I157967,);
not I_9112 (I157975,I157967);
not I_9113 (I157992,I157950);
nand I_9114 (I157689,I157992,I157811);
nand I_9115 (I158023,I234789,I234795);
and I_9116 (I158040,I158023,I234798);
DFFARX1 I_9117 (I158040,I3035,I157712,I158066,);
nor I_9118 (I158074,I158066,I157738);
DFFARX1 I_9119 (I158074,I3035,I157712,I157677,);
DFFARX1 I_9120 (I158066,I3035,I157712,I157695,);
nor I_9121 (I158119,I234810,I234795);
not I_9122 (I158136,I158119);
nor I_9123 (I157698,I157975,I158136);
nand I_9124 (I157683,I157992,I158136);
nor I_9125 (I157692,I157738,I158119);
DFFARX1 I_9126 (I158119,I3035,I157712,I157701,);
not I_9127 (I158239,I3042);
DFFARX1 I_9128 (I361434,I3035,I158239,I158265,);
nand I_9129 (I158273,I361425,I361440);
and I_9130 (I158290,I158273,I361446);
DFFARX1 I_9131 (I158290,I3035,I158239,I158316,);
nor I_9132 (I158207,I158316,I158265);
not I_9133 (I158338,I158316);
DFFARX1 I_9134 (I361431,I3035,I158239,I158364,);
nand I_9135 (I158372,I158364,I361425);
not I_9136 (I158389,I158372);
DFFARX1 I_9137 (I158389,I3035,I158239,I158415,);
not I_9138 (I158231,I158415);
nor I_9139 (I158437,I158265,I158372);
nor I_9140 (I158213,I158316,I158437);
DFFARX1 I_9141 (I361428,I3035,I158239,I158477,);
DFFARX1 I_9142 (I158477,I3035,I158239,I158494,);
not I_9143 (I158502,I158494);
not I_9144 (I158519,I158477);
nand I_9145 (I158216,I158519,I158338);
nand I_9146 (I158550,I361422,I361437);
and I_9147 (I158567,I158550,I361422);
DFFARX1 I_9148 (I158567,I3035,I158239,I158593,);
nor I_9149 (I158601,I158593,I158265);
DFFARX1 I_9150 (I158601,I3035,I158239,I158204,);
DFFARX1 I_9151 (I158593,I3035,I158239,I158222,);
nor I_9152 (I158646,I361443,I361437);
not I_9153 (I158663,I158646);
nor I_9154 (I158225,I158502,I158663);
nand I_9155 (I158210,I158519,I158663);
nor I_9156 (I158219,I158265,I158646);
DFFARX1 I_9157 (I158646,I3035,I158239,I158228,);
not I_9158 (I158766,I3042);
DFFARX1 I_9159 (I720449,I3035,I158766,I158792,);
nand I_9160 (I158800,I720428,I720428);
and I_9161 (I158817,I158800,I720455);
DFFARX1 I_9162 (I158817,I3035,I158766,I158843,);
nor I_9163 (I158734,I158843,I158792);
not I_9164 (I158865,I158843);
DFFARX1 I_9165 (I720443,I3035,I158766,I158891,);
nand I_9166 (I158899,I158891,I720446);
not I_9167 (I158916,I158899);
DFFARX1 I_9168 (I158916,I3035,I158766,I158942,);
not I_9169 (I158758,I158942);
nor I_9170 (I158964,I158792,I158899);
nor I_9171 (I158740,I158843,I158964);
DFFARX1 I_9172 (I720437,I3035,I158766,I159004,);
DFFARX1 I_9173 (I159004,I3035,I158766,I159021,);
not I_9174 (I159029,I159021);
not I_9175 (I159046,I159004);
nand I_9176 (I158743,I159046,I158865);
nand I_9177 (I159077,I720434,I720431);
and I_9178 (I159094,I159077,I720452);
DFFARX1 I_9179 (I159094,I3035,I158766,I159120,);
nor I_9180 (I159128,I159120,I158792);
DFFARX1 I_9181 (I159128,I3035,I158766,I158731,);
DFFARX1 I_9182 (I159120,I3035,I158766,I158749,);
nor I_9183 (I159173,I720440,I720431);
not I_9184 (I159190,I159173);
nor I_9185 (I158752,I159029,I159190);
nand I_9186 (I158737,I159046,I159190);
nor I_9187 (I158746,I158792,I159173);
DFFARX1 I_9188 (I159173,I3035,I158766,I158755,);
not I_9189 (I159293,I3042);
DFFARX1 I_9190 (I373572,I3035,I159293,I159319,);
nand I_9191 (I159327,I373563,I373578);
and I_9192 (I159344,I159327,I373584);
DFFARX1 I_9193 (I159344,I3035,I159293,I159370,);
nor I_9194 (I159261,I159370,I159319);
not I_9195 (I159392,I159370);
DFFARX1 I_9196 (I373569,I3035,I159293,I159418,);
nand I_9197 (I159426,I159418,I373563);
not I_9198 (I159443,I159426);
DFFARX1 I_9199 (I159443,I3035,I159293,I159469,);
not I_9200 (I159285,I159469);
nor I_9201 (I159491,I159319,I159426);
nor I_9202 (I159267,I159370,I159491);
DFFARX1 I_9203 (I373566,I3035,I159293,I159531,);
DFFARX1 I_9204 (I159531,I3035,I159293,I159548,);
not I_9205 (I159556,I159548);
not I_9206 (I159573,I159531);
nand I_9207 (I159270,I159573,I159392);
nand I_9208 (I159604,I373560,I373575);
and I_9209 (I159621,I159604,I373560);
DFFARX1 I_9210 (I159621,I3035,I159293,I159647,);
nor I_9211 (I159655,I159647,I159319);
DFFARX1 I_9212 (I159655,I3035,I159293,I159258,);
DFFARX1 I_9213 (I159647,I3035,I159293,I159276,);
nor I_9214 (I159700,I373581,I373575);
not I_9215 (I159717,I159700);
nor I_9216 (I159279,I159556,I159717);
nand I_9217 (I159264,I159573,I159717);
nor I_9218 (I159273,I159319,I159700);
DFFARX1 I_9219 (I159700,I3035,I159293,I159282,);
not I_9220 (I159820,I3042);
DFFARX1 I_9221 (I78899,I3035,I159820,I159846,);
nand I_9222 (I159854,I78899,I78905);
and I_9223 (I159871,I159854,I78923);
DFFARX1 I_9224 (I159871,I3035,I159820,I159897,);
nor I_9225 (I159788,I159897,I159846);
not I_9226 (I159919,I159897);
DFFARX1 I_9227 (I78911,I3035,I159820,I159945,);
nand I_9228 (I159953,I159945,I78908);
not I_9229 (I159970,I159953);
DFFARX1 I_9230 (I159970,I3035,I159820,I159996,);
not I_9231 (I159812,I159996);
nor I_9232 (I160018,I159846,I159953);
nor I_9233 (I159794,I159897,I160018);
DFFARX1 I_9234 (I78917,I3035,I159820,I160058,);
DFFARX1 I_9235 (I160058,I3035,I159820,I160075,);
not I_9236 (I160083,I160075);
not I_9237 (I160100,I160058);
nand I_9238 (I159797,I160100,I159919);
nand I_9239 (I160131,I78902,I78902);
and I_9240 (I160148,I160131,I78914);
DFFARX1 I_9241 (I160148,I3035,I159820,I160174,);
nor I_9242 (I160182,I160174,I159846);
DFFARX1 I_9243 (I160182,I3035,I159820,I159785,);
DFFARX1 I_9244 (I160174,I3035,I159820,I159803,);
nor I_9245 (I160227,I78920,I78902);
not I_9246 (I160244,I160227);
nor I_9247 (I159806,I160083,I160244);
nand I_9248 (I159791,I160100,I160244);
nor I_9249 (I159800,I159846,I160227);
DFFARX1 I_9250 (I160227,I3035,I159820,I159809,);
not I_9251 (I160347,I3042);
DFFARX1 I_9252 (I383398,I3035,I160347,I160373,);
nand I_9253 (I160381,I383389,I383404);
and I_9254 (I160398,I160381,I383410);
DFFARX1 I_9255 (I160398,I3035,I160347,I160424,);
nor I_9256 (I160315,I160424,I160373);
not I_9257 (I160446,I160424);
DFFARX1 I_9258 (I383395,I3035,I160347,I160472,);
nand I_9259 (I160480,I160472,I383389);
not I_9260 (I160497,I160480);
DFFARX1 I_9261 (I160497,I3035,I160347,I160523,);
not I_9262 (I160339,I160523);
nor I_9263 (I160545,I160373,I160480);
nor I_9264 (I160321,I160424,I160545);
DFFARX1 I_9265 (I383392,I3035,I160347,I160585,);
DFFARX1 I_9266 (I160585,I3035,I160347,I160602,);
not I_9267 (I160610,I160602);
not I_9268 (I160627,I160585);
nand I_9269 (I160324,I160627,I160446);
nand I_9270 (I160658,I383386,I383401);
and I_9271 (I160675,I160658,I383386);
DFFARX1 I_9272 (I160675,I3035,I160347,I160701,);
nor I_9273 (I160709,I160701,I160373);
DFFARX1 I_9274 (I160709,I3035,I160347,I160312,);
DFFARX1 I_9275 (I160701,I3035,I160347,I160330,);
nor I_9276 (I160754,I383407,I383401);
not I_9277 (I160771,I160754);
nor I_9278 (I160333,I160610,I160771);
nand I_9279 (I160318,I160627,I160771);
nor I_9280 (I160327,I160373,I160754);
DFFARX1 I_9281 (I160754,I3035,I160347,I160336,);
not I_9282 (I160874,I3042);
DFFARX1 I_9283 (I707359,I3035,I160874,I160900,);
nand I_9284 (I160908,I707338,I707338);
and I_9285 (I160925,I160908,I707365);
DFFARX1 I_9286 (I160925,I3035,I160874,I160951,);
nor I_9287 (I160842,I160951,I160900);
not I_9288 (I160973,I160951);
DFFARX1 I_9289 (I707353,I3035,I160874,I160999,);
nand I_9290 (I161007,I160999,I707356);
not I_9291 (I161024,I161007);
DFFARX1 I_9292 (I161024,I3035,I160874,I161050,);
not I_9293 (I160866,I161050);
nor I_9294 (I161072,I160900,I161007);
nor I_9295 (I160848,I160951,I161072);
DFFARX1 I_9296 (I707347,I3035,I160874,I161112,);
DFFARX1 I_9297 (I161112,I3035,I160874,I161129,);
not I_9298 (I161137,I161129);
not I_9299 (I161154,I161112);
nand I_9300 (I160851,I161154,I160973);
nand I_9301 (I161185,I707344,I707341);
and I_9302 (I161202,I161185,I707362);
DFFARX1 I_9303 (I161202,I3035,I160874,I161228,);
nor I_9304 (I161236,I161228,I160900);
DFFARX1 I_9305 (I161236,I3035,I160874,I160839,);
DFFARX1 I_9306 (I161228,I3035,I160874,I160857,);
nor I_9307 (I161281,I707350,I707341);
not I_9308 (I161298,I161281);
nor I_9309 (I160860,I161137,I161298);
nand I_9310 (I160845,I161154,I161298);
nor I_9311 (I160854,I160900,I161281);
DFFARX1 I_9312 (I161281,I3035,I160874,I160863,);
not I_9313 (I161401,I3042);
DFFARX1 I_9314 (I53657,I3035,I161401,I161427,);
nand I_9315 (I161435,I53669,I53678);
and I_9316 (I161452,I161435,I53657);
DFFARX1 I_9317 (I161452,I3035,I161401,I161478,);
nor I_9318 (I161369,I161478,I161427);
not I_9319 (I161500,I161478);
DFFARX1 I_9320 (I53672,I3035,I161401,I161526,);
nand I_9321 (I161534,I161526,I53660);
not I_9322 (I161551,I161534);
DFFARX1 I_9323 (I161551,I3035,I161401,I161577,);
not I_9324 (I161393,I161577);
nor I_9325 (I161599,I161427,I161534);
nor I_9326 (I161375,I161478,I161599);
DFFARX1 I_9327 (I53663,I3035,I161401,I161639,);
DFFARX1 I_9328 (I161639,I3035,I161401,I161656,);
not I_9329 (I161664,I161656);
not I_9330 (I161681,I161639);
nand I_9331 (I161378,I161681,I161500);
nand I_9332 (I161712,I53654,I53654);
and I_9333 (I161729,I161712,I53666);
DFFARX1 I_9334 (I161729,I3035,I161401,I161755,);
nor I_9335 (I161763,I161755,I161427);
DFFARX1 I_9336 (I161763,I3035,I161401,I161366,);
DFFARX1 I_9337 (I161755,I3035,I161401,I161384,);
nor I_9338 (I161808,I53675,I53654);
not I_9339 (I161825,I161808);
nor I_9340 (I161387,I161664,I161825);
nand I_9341 (I161372,I161681,I161825);
nor I_9342 (I161381,I161427,I161808);
DFFARX1 I_9343 (I161808,I3035,I161401,I161390,);
not I_9344 (I161928,I3042);
DFFARX1 I_9345 (I476192,I3035,I161928,I161954,);
nand I_9346 (I161962,I476195,I476189);
and I_9347 (I161979,I161962,I476201);
DFFARX1 I_9348 (I161979,I3035,I161928,I162005,);
nor I_9349 (I161896,I162005,I161954);
not I_9350 (I162027,I162005);
DFFARX1 I_9351 (I476204,I3035,I161928,I162053,);
nand I_9352 (I162061,I162053,I476195);
not I_9353 (I162078,I162061);
DFFARX1 I_9354 (I162078,I3035,I161928,I162104,);
not I_9355 (I161920,I162104);
nor I_9356 (I162126,I161954,I162061);
nor I_9357 (I161902,I162005,I162126);
DFFARX1 I_9358 (I476207,I3035,I161928,I162166,);
DFFARX1 I_9359 (I162166,I3035,I161928,I162183,);
not I_9360 (I162191,I162183);
not I_9361 (I162208,I162166);
nand I_9362 (I161905,I162208,I162027);
nand I_9363 (I162239,I476189,I476198);
and I_9364 (I162256,I162239,I476192);
DFFARX1 I_9365 (I162256,I3035,I161928,I162282,);
nor I_9366 (I162290,I162282,I161954);
DFFARX1 I_9367 (I162290,I3035,I161928,I161893,);
DFFARX1 I_9368 (I162282,I3035,I161928,I161911,);
nor I_9369 (I162335,I476210,I476198);
not I_9370 (I162352,I162335);
nor I_9371 (I161914,I162191,I162352);
nand I_9372 (I161899,I162208,I162352);
nor I_9373 (I161908,I161954,I162335);
DFFARX1 I_9374 (I162335,I3035,I161928,I161917,);
not I_9375 (I162455,I3042);
DFFARX1 I_9376 (I695540,I3035,I162455,I162481,);
nand I_9377 (I162489,I695567,I695543);
and I_9378 (I162506,I162489,I695552);
DFFARX1 I_9379 (I162506,I3035,I162455,I162532,);
nor I_9380 (I162423,I162532,I162481);
not I_9381 (I162554,I162532);
DFFARX1 I_9382 (I695540,I3035,I162455,I162580,);
nand I_9383 (I162588,I162580,I695564);
not I_9384 (I162605,I162588);
DFFARX1 I_9385 (I162605,I3035,I162455,I162631,);
not I_9386 (I162447,I162631);
nor I_9387 (I162653,I162481,I162588);
nor I_9388 (I162429,I162532,I162653);
DFFARX1 I_9389 (I695546,I3035,I162455,I162693,);
DFFARX1 I_9390 (I162693,I3035,I162455,I162710,);
not I_9391 (I162718,I162710);
not I_9392 (I162735,I162693);
nand I_9393 (I162432,I162735,I162554);
nand I_9394 (I162766,I695561,I695549);
and I_9395 (I162783,I162766,I695555);
DFFARX1 I_9396 (I162783,I3035,I162455,I162809,);
nor I_9397 (I162817,I162809,I162481);
DFFARX1 I_9398 (I162817,I3035,I162455,I162420,);
DFFARX1 I_9399 (I162809,I3035,I162455,I162438,);
nor I_9400 (I162862,I695558,I695549);
not I_9401 (I162879,I162862);
nor I_9402 (I162441,I162718,I162879);
nand I_9403 (I162426,I162735,I162879);
nor I_9404 (I162435,I162481,I162862);
DFFARX1 I_9405 (I162862,I3035,I162455,I162444,);
not I_9406 (I162982,I3042);
DFFARX1 I_9407 (I128879,I3035,I162982,I163008,);
nand I_9408 (I163016,I128879,I128885);
and I_9409 (I163033,I163016,I128903);
DFFARX1 I_9410 (I163033,I3035,I162982,I163059,);
nor I_9411 (I162950,I163059,I163008);
not I_9412 (I163081,I163059);
DFFARX1 I_9413 (I128891,I3035,I162982,I163107,);
nand I_9414 (I163115,I163107,I128888);
not I_9415 (I163132,I163115);
DFFARX1 I_9416 (I163132,I3035,I162982,I163158,);
not I_9417 (I162974,I163158);
nor I_9418 (I163180,I163008,I163115);
nor I_9419 (I162956,I163059,I163180);
DFFARX1 I_9420 (I128897,I3035,I162982,I163220,);
DFFARX1 I_9421 (I163220,I3035,I162982,I163237,);
not I_9422 (I163245,I163237);
not I_9423 (I163262,I163220);
nand I_9424 (I162959,I163262,I163081);
nand I_9425 (I163293,I128882,I128882);
and I_9426 (I163310,I163293,I128894);
DFFARX1 I_9427 (I163310,I3035,I162982,I163336,);
nor I_9428 (I163344,I163336,I163008);
DFFARX1 I_9429 (I163344,I3035,I162982,I162947,);
DFFARX1 I_9430 (I163336,I3035,I162982,I162965,);
nor I_9431 (I163389,I128900,I128882);
not I_9432 (I163406,I163389);
nor I_9433 (I162968,I163245,I163406);
nand I_9434 (I162953,I163262,I163406);
nor I_9435 (I162962,I163008,I163389);
DFFARX1 I_9436 (I163389,I3035,I162982,I162971,);
not I_9437 (I163509,I3042);
DFFARX1 I_9438 (I368948,I3035,I163509,I163535,);
nand I_9439 (I163543,I368939,I368954);
and I_9440 (I163560,I163543,I368960);
DFFARX1 I_9441 (I163560,I3035,I163509,I163586,);
nor I_9442 (I163477,I163586,I163535);
not I_9443 (I163608,I163586);
DFFARX1 I_9444 (I368945,I3035,I163509,I163634,);
nand I_9445 (I163642,I163634,I368939);
not I_9446 (I163659,I163642);
DFFARX1 I_9447 (I163659,I3035,I163509,I163685,);
not I_9448 (I163501,I163685);
nor I_9449 (I163707,I163535,I163642);
nor I_9450 (I163483,I163586,I163707);
DFFARX1 I_9451 (I368942,I3035,I163509,I163747,);
DFFARX1 I_9452 (I163747,I3035,I163509,I163764,);
not I_9453 (I163772,I163764);
not I_9454 (I163789,I163747);
nand I_9455 (I163486,I163789,I163608);
nand I_9456 (I163820,I368936,I368951);
and I_9457 (I163837,I163820,I368936);
DFFARX1 I_9458 (I163837,I3035,I163509,I163863,);
nor I_9459 (I163871,I163863,I163535);
DFFARX1 I_9460 (I163871,I3035,I163509,I163474,);
DFFARX1 I_9461 (I163863,I3035,I163509,I163492,);
nor I_9462 (I163916,I368957,I368951);
not I_9463 (I163933,I163916);
nor I_9464 (I163495,I163772,I163933);
nand I_9465 (I163480,I163789,I163933);
nor I_9466 (I163489,I163535,I163916);
DFFARX1 I_9467 (I163916,I3035,I163509,I163498,);
not I_9468 (I164036,I3042);
DFFARX1 I_9469 (I559951,I3035,I164036,I164062,);
nand I_9470 (I164070,I559948,I559951);
and I_9471 (I164087,I164070,I559960);
DFFARX1 I_9472 (I164087,I3035,I164036,I164113,);
nor I_9473 (I164004,I164113,I164062);
not I_9474 (I164135,I164113);
DFFARX1 I_9475 (I559948,I3035,I164036,I164161,);
nand I_9476 (I164169,I164161,I559966);
not I_9477 (I164186,I164169);
DFFARX1 I_9478 (I164186,I3035,I164036,I164212,);
not I_9479 (I164028,I164212);
nor I_9480 (I164234,I164062,I164169);
nor I_9481 (I164010,I164113,I164234);
DFFARX1 I_9482 (I559954,I3035,I164036,I164274,);
DFFARX1 I_9483 (I164274,I3035,I164036,I164291,);
not I_9484 (I164299,I164291);
not I_9485 (I164316,I164274);
nand I_9486 (I164013,I164316,I164135);
nand I_9487 (I164347,I559963,I559969);
and I_9488 (I164364,I164347,I559954);
DFFARX1 I_9489 (I164364,I3035,I164036,I164390,);
nor I_9490 (I164398,I164390,I164062);
DFFARX1 I_9491 (I164398,I3035,I164036,I164001,);
DFFARX1 I_9492 (I164390,I3035,I164036,I164019,);
nor I_9493 (I164443,I559957,I559969);
not I_9494 (I164460,I164443);
nor I_9495 (I164022,I164299,I164460);
nand I_9496 (I164007,I164316,I164460);
nor I_9497 (I164016,I164062,I164443);
DFFARX1 I_9498 (I164443,I3035,I164036,I164025,);
not I_9499 (I164563,I3042);
DFFARX1 I_9500 (I550414,I3035,I164563,I164589,);
nand I_9501 (I164597,I550411,I550414);
and I_9502 (I164614,I164597,I550423);
DFFARX1 I_9503 (I164614,I3035,I164563,I164640,);
nor I_9504 (I164531,I164640,I164589);
not I_9505 (I164662,I164640);
DFFARX1 I_9506 (I550411,I3035,I164563,I164688,);
nand I_9507 (I164696,I164688,I550429);
not I_9508 (I164713,I164696);
DFFARX1 I_9509 (I164713,I3035,I164563,I164739,);
not I_9510 (I164555,I164739);
nor I_9511 (I164761,I164589,I164696);
nor I_9512 (I164537,I164640,I164761);
DFFARX1 I_9513 (I550417,I3035,I164563,I164801,);
DFFARX1 I_9514 (I164801,I3035,I164563,I164818,);
not I_9515 (I164826,I164818);
not I_9516 (I164843,I164801);
nand I_9517 (I164540,I164843,I164662);
nand I_9518 (I164874,I550426,I550432);
and I_9519 (I164891,I164874,I550417);
DFFARX1 I_9520 (I164891,I3035,I164563,I164917,);
nor I_9521 (I164925,I164917,I164589);
DFFARX1 I_9522 (I164925,I3035,I164563,I164528,);
DFFARX1 I_9523 (I164917,I3035,I164563,I164546,);
nor I_9524 (I164970,I550420,I550432);
not I_9525 (I164987,I164970);
nor I_9526 (I164549,I164826,I164987);
nand I_9527 (I164534,I164843,I164987);
nor I_9528 (I164543,I164589,I164970);
DFFARX1 I_9529 (I164970,I3035,I164563,I164552,);
not I_9530 (I165090,I3042);
DFFARX1 I_9531 (I133044,I3035,I165090,I165116,);
nand I_9532 (I165124,I133044,I133050);
and I_9533 (I165141,I165124,I133068);
DFFARX1 I_9534 (I165141,I3035,I165090,I165167,);
nor I_9535 (I165058,I165167,I165116);
not I_9536 (I165189,I165167);
DFFARX1 I_9537 (I133056,I3035,I165090,I165215,);
nand I_9538 (I165223,I165215,I133053);
not I_9539 (I165240,I165223);
DFFARX1 I_9540 (I165240,I3035,I165090,I165266,);
not I_9541 (I165082,I165266);
nor I_9542 (I165288,I165116,I165223);
nor I_9543 (I165064,I165167,I165288);
DFFARX1 I_9544 (I133062,I3035,I165090,I165328,);
DFFARX1 I_9545 (I165328,I3035,I165090,I165345,);
not I_9546 (I165353,I165345);
not I_9547 (I165370,I165328);
nand I_9548 (I165067,I165370,I165189);
nand I_9549 (I165401,I133047,I133047);
and I_9550 (I165418,I165401,I133059);
DFFARX1 I_9551 (I165418,I3035,I165090,I165444,);
nor I_9552 (I165452,I165444,I165116);
DFFARX1 I_9553 (I165452,I3035,I165090,I165055,);
DFFARX1 I_9554 (I165444,I3035,I165090,I165073,);
nor I_9555 (I165497,I133065,I133047);
not I_9556 (I165514,I165497);
nor I_9557 (I165076,I165353,I165514);
nand I_9558 (I165061,I165370,I165514);
nor I_9559 (I165070,I165116,I165497);
DFFARX1 I_9560 (I165497,I3035,I165090,I165079,);
not I_9561 (I165617,I3042);
DFFARX1 I_9562 (I87824,I3035,I165617,I165643,);
nand I_9563 (I165651,I87824,I87830);
and I_9564 (I165668,I165651,I87848);
DFFARX1 I_9565 (I165668,I3035,I165617,I165694,);
nor I_9566 (I165585,I165694,I165643);
not I_9567 (I165716,I165694);
DFFARX1 I_9568 (I87836,I3035,I165617,I165742,);
nand I_9569 (I165750,I165742,I87833);
not I_9570 (I165767,I165750);
DFFARX1 I_9571 (I165767,I3035,I165617,I165793,);
not I_9572 (I165609,I165793);
nor I_9573 (I165815,I165643,I165750);
nor I_9574 (I165591,I165694,I165815);
DFFARX1 I_9575 (I87842,I3035,I165617,I165855,);
DFFARX1 I_9576 (I165855,I3035,I165617,I165872,);
not I_9577 (I165880,I165872);
not I_9578 (I165897,I165855);
nand I_9579 (I165594,I165897,I165716);
nand I_9580 (I165928,I87827,I87827);
and I_9581 (I165945,I165928,I87839);
DFFARX1 I_9582 (I165945,I3035,I165617,I165971,);
nor I_9583 (I165979,I165971,I165643);
DFFARX1 I_9584 (I165979,I3035,I165617,I165582,);
DFFARX1 I_9585 (I165971,I3035,I165617,I165600,);
nor I_9586 (I166024,I87845,I87827);
not I_9587 (I166041,I166024);
nor I_9588 (I165603,I165880,I166041);
nand I_9589 (I165588,I165897,I166041);
nor I_9590 (I165597,I165643,I166024);
DFFARX1 I_9591 (I166024,I3035,I165617,I165606,);
not I_9592 (I166144,I3042);
DFFARX1 I_9593 (I2292,I3035,I166144,I166170,);
nand I_9594 (I166178,I2356,I2508);
and I_9595 (I166195,I166178,I2172);
DFFARX1 I_9596 (I166195,I3035,I166144,I166221,);
nor I_9597 (I166112,I166221,I166170);
not I_9598 (I166243,I166221);
DFFARX1 I_9599 (I2700,I3035,I166144,I166269,);
nand I_9600 (I166277,I166269,I1876);
not I_9601 (I166294,I166277);
DFFARX1 I_9602 (I166294,I3035,I166144,I166320,);
not I_9603 (I166136,I166320);
nor I_9604 (I166342,I166170,I166277);
nor I_9605 (I166118,I166221,I166342);
DFFARX1 I_9606 (I1892,I3035,I166144,I166382,);
DFFARX1 I_9607 (I166382,I3035,I166144,I166399,);
not I_9608 (I166407,I166399);
not I_9609 (I166424,I166382);
nand I_9610 (I166121,I166424,I166243);
nand I_9611 (I166455,I2956,I1916);
and I_9612 (I166472,I166455,I1612);
DFFARX1 I_9613 (I166472,I3035,I166144,I166498,);
nor I_9614 (I166506,I166498,I166170);
DFFARX1 I_9615 (I166506,I3035,I166144,I166109,);
DFFARX1 I_9616 (I166498,I3035,I166144,I166127,);
nor I_9617 (I166551,I2484,I1916);
not I_9618 (I166568,I166551);
nor I_9619 (I166130,I166407,I166568);
nand I_9620 (I166115,I166424,I166568);
nor I_9621 (I166124,I166170,I166551);
DFFARX1 I_9622 (I166551,I3035,I166144,I166133,);
not I_9623 (I166671,I3042);
DFFARX1 I_9624 (I136019,I3035,I166671,I166697,);
nand I_9625 (I166705,I136019,I136025);
and I_9626 (I166722,I166705,I136043);
DFFARX1 I_9627 (I166722,I3035,I166671,I166748,);
nor I_9628 (I166639,I166748,I166697);
not I_9629 (I166770,I166748);
DFFARX1 I_9630 (I136031,I3035,I166671,I166796,);
nand I_9631 (I166804,I166796,I136028);
not I_9632 (I166821,I166804);
DFFARX1 I_9633 (I166821,I3035,I166671,I166847,);
not I_9634 (I166663,I166847);
nor I_9635 (I166869,I166697,I166804);
nor I_9636 (I166645,I166748,I166869);
DFFARX1 I_9637 (I136037,I3035,I166671,I166909,);
DFFARX1 I_9638 (I166909,I3035,I166671,I166926,);
not I_9639 (I166934,I166926);
not I_9640 (I166951,I166909);
nand I_9641 (I166648,I166951,I166770);
nand I_9642 (I166982,I136022,I136022);
and I_9643 (I166999,I166982,I136034);
DFFARX1 I_9644 (I166999,I3035,I166671,I167025,);
nor I_9645 (I167033,I167025,I166697);
DFFARX1 I_9646 (I167033,I3035,I166671,I166636,);
DFFARX1 I_9647 (I167025,I3035,I166671,I166654,);
nor I_9648 (I167078,I136040,I136022);
not I_9649 (I167095,I167078);
nor I_9650 (I166657,I166934,I167095);
nand I_9651 (I166642,I166951,I167095);
nor I_9652 (I166651,I166697,I167078);
DFFARX1 I_9653 (I167078,I3035,I166671,I166660,);
not I_9654 (I167198,I3042);
DFFARX1 I_9655 (I449842,I3035,I167198,I167224,);
nand I_9656 (I167232,I449845,I449839);
and I_9657 (I167249,I167232,I449851);
DFFARX1 I_9658 (I167249,I3035,I167198,I167275,);
nor I_9659 (I167166,I167275,I167224);
not I_9660 (I167297,I167275);
DFFARX1 I_9661 (I449854,I3035,I167198,I167323,);
nand I_9662 (I167331,I167323,I449845);
not I_9663 (I167348,I167331);
DFFARX1 I_9664 (I167348,I3035,I167198,I167374,);
not I_9665 (I167190,I167374);
nor I_9666 (I167396,I167224,I167331);
nor I_9667 (I167172,I167275,I167396);
DFFARX1 I_9668 (I449857,I3035,I167198,I167436,);
DFFARX1 I_9669 (I167436,I3035,I167198,I167453,);
not I_9670 (I167461,I167453);
not I_9671 (I167478,I167436);
nand I_9672 (I167175,I167478,I167297);
nand I_9673 (I167509,I449839,I449848);
and I_9674 (I167526,I167509,I449842);
DFFARX1 I_9675 (I167526,I3035,I167198,I167552,);
nor I_9676 (I167560,I167552,I167224);
DFFARX1 I_9677 (I167560,I3035,I167198,I167163,);
DFFARX1 I_9678 (I167552,I3035,I167198,I167181,);
nor I_9679 (I167605,I449860,I449848);
not I_9680 (I167622,I167605);
nor I_9681 (I167184,I167461,I167622);
nand I_9682 (I167169,I167478,I167622);
nor I_9683 (I167178,I167224,I167605);
DFFARX1 I_9684 (I167605,I3035,I167198,I167187,);
not I_9685 (I167725,I3042);
DFFARX1 I_9686 (I530337,I3035,I167725,I167751,);
nand I_9687 (I167759,I530334,I530352);
and I_9688 (I167776,I167759,I530343);
DFFARX1 I_9689 (I167776,I3035,I167725,I167802,);
nor I_9690 (I167693,I167802,I167751);
not I_9691 (I167824,I167802);
DFFARX1 I_9692 (I530358,I3035,I167725,I167850,);
nand I_9693 (I167858,I167850,I530340);
not I_9694 (I167875,I167858);
DFFARX1 I_9695 (I167875,I3035,I167725,I167901,);
not I_9696 (I167717,I167901);
nor I_9697 (I167923,I167751,I167858);
nor I_9698 (I167699,I167802,I167923);
DFFARX1 I_9699 (I530346,I3035,I167725,I167963,);
DFFARX1 I_9700 (I167963,I3035,I167725,I167980,);
not I_9701 (I167988,I167980);
not I_9702 (I168005,I167963);
nand I_9703 (I167702,I168005,I167824);
nand I_9704 (I168036,I530334,I530361);
and I_9705 (I168053,I168036,I530349);
DFFARX1 I_9706 (I168053,I3035,I167725,I168079,);
nor I_9707 (I168087,I168079,I167751);
DFFARX1 I_9708 (I168087,I3035,I167725,I167690,);
DFFARX1 I_9709 (I168079,I3035,I167725,I167708,);
nor I_9710 (I168132,I530355,I530361);
not I_9711 (I168149,I168132);
nor I_9712 (I167711,I167988,I168149);
nand I_9713 (I167696,I168005,I168149);
nor I_9714 (I167705,I167751,I168132);
DFFARX1 I_9715 (I168132,I3035,I167725,I167714,);
not I_9716 (I168252,I3042);
DFFARX1 I_9717 (I405362,I3035,I168252,I168278,);
nand I_9718 (I168286,I405353,I405368);
and I_9719 (I168303,I168286,I405374);
DFFARX1 I_9720 (I168303,I3035,I168252,I168329,);
nor I_9721 (I168220,I168329,I168278);
not I_9722 (I168351,I168329);
DFFARX1 I_9723 (I405359,I3035,I168252,I168377,);
nand I_9724 (I168385,I168377,I405353);
not I_9725 (I168402,I168385);
DFFARX1 I_9726 (I168402,I3035,I168252,I168428,);
not I_9727 (I168244,I168428);
nor I_9728 (I168450,I168278,I168385);
nor I_9729 (I168226,I168329,I168450);
DFFARX1 I_9730 (I405356,I3035,I168252,I168490,);
DFFARX1 I_9731 (I168490,I3035,I168252,I168507,);
not I_9732 (I168515,I168507);
not I_9733 (I168532,I168490);
nand I_9734 (I168229,I168532,I168351);
nand I_9735 (I168563,I405350,I405365);
and I_9736 (I168580,I168563,I405350);
DFFARX1 I_9737 (I168580,I3035,I168252,I168606,);
nor I_9738 (I168614,I168606,I168278);
DFFARX1 I_9739 (I168614,I3035,I168252,I168217,);
DFFARX1 I_9740 (I168606,I3035,I168252,I168235,);
nor I_9741 (I168659,I405371,I405365);
not I_9742 (I168676,I168659);
nor I_9743 (I168238,I168515,I168676);
nand I_9744 (I168223,I168532,I168676);
nor I_9745 (I168232,I168278,I168659);
DFFARX1 I_9746 (I168659,I3035,I168252,I168241,);
not I_9747 (I168779,I3042);
DFFARX1 I_9748 (I133639,I3035,I168779,I168805,);
nand I_9749 (I168813,I133639,I133645);
and I_9750 (I168830,I168813,I133663);
DFFARX1 I_9751 (I168830,I3035,I168779,I168856,);
nor I_9752 (I168747,I168856,I168805);
not I_9753 (I168878,I168856);
DFFARX1 I_9754 (I133651,I3035,I168779,I168904,);
nand I_9755 (I168912,I168904,I133648);
not I_9756 (I168929,I168912);
DFFARX1 I_9757 (I168929,I3035,I168779,I168955,);
not I_9758 (I168771,I168955);
nor I_9759 (I168977,I168805,I168912);
nor I_9760 (I168753,I168856,I168977);
DFFARX1 I_9761 (I133657,I3035,I168779,I169017,);
DFFARX1 I_9762 (I169017,I3035,I168779,I169034,);
not I_9763 (I169042,I169034);
not I_9764 (I169059,I169017);
nand I_9765 (I168756,I169059,I168878);
nand I_9766 (I169090,I133642,I133642);
and I_9767 (I169107,I169090,I133654);
DFFARX1 I_9768 (I169107,I3035,I168779,I169133,);
nor I_9769 (I169141,I169133,I168805);
DFFARX1 I_9770 (I169141,I3035,I168779,I168744,);
DFFARX1 I_9771 (I169133,I3035,I168779,I168762,);
nor I_9772 (I169186,I133660,I133642);
not I_9773 (I169203,I169186);
nor I_9774 (I168765,I169042,I169203);
nand I_9775 (I168750,I169059,I169203);
nor I_9776 (I168759,I168805,I169186);
DFFARX1 I_9777 (I169186,I3035,I168779,I168768,);
not I_9778 (I169306,I3042);
DFFARX1 I_9779 (I302481,I3035,I169306,I169332,);
nand I_9780 (I169340,I302466,I302469);
and I_9781 (I169357,I169340,I302484);
DFFARX1 I_9782 (I169357,I3035,I169306,I169383,);
nor I_9783 (I169274,I169383,I169332);
not I_9784 (I169405,I169383);
DFFARX1 I_9785 (I302478,I3035,I169306,I169431,);
nand I_9786 (I169439,I169431,I302469);
not I_9787 (I169456,I169439);
DFFARX1 I_9788 (I169456,I3035,I169306,I169482,);
not I_9789 (I169298,I169482);
nor I_9790 (I169504,I169332,I169439);
nor I_9791 (I169280,I169383,I169504);
DFFARX1 I_9792 (I302475,I3035,I169306,I169544,);
DFFARX1 I_9793 (I169544,I3035,I169306,I169561,);
not I_9794 (I169569,I169561);
not I_9795 (I169586,I169544);
nand I_9796 (I169283,I169586,I169405);
nand I_9797 (I169617,I302490,I302466);
and I_9798 (I169634,I169617,I302487);
DFFARX1 I_9799 (I169634,I3035,I169306,I169660,);
nor I_9800 (I169668,I169660,I169332);
DFFARX1 I_9801 (I169668,I3035,I169306,I169271,);
DFFARX1 I_9802 (I169660,I3035,I169306,I169289,);
nor I_9803 (I169713,I302472,I302466);
not I_9804 (I169730,I169713);
nor I_9805 (I169292,I169569,I169730);
nand I_9806 (I169277,I169586,I169730);
nor I_9807 (I169286,I169332,I169713);
DFFARX1 I_9808 (I169713,I3035,I169306,I169295,);
not I_9809 (I169833,I3042);
DFFARX1 I_9810 (I576336,I3035,I169833,I169859,);
nand I_9811 (I169867,I576351,I576336);
and I_9812 (I169884,I169867,I576354);
DFFARX1 I_9813 (I169884,I3035,I169833,I169910,);
nor I_9814 (I169801,I169910,I169859);
not I_9815 (I169932,I169910);
DFFARX1 I_9816 (I576360,I3035,I169833,I169958,);
nand I_9817 (I169966,I169958,I576342);
not I_9818 (I169983,I169966);
DFFARX1 I_9819 (I169983,I3035,I169833,I170009,);
not I_9820 (I169825,I170009);
nor I_9821 (I170031,I169859,I169966);
nor I_9822 (I169807,I169910,I170031);
DFFARX1 I_9823 (I576339,I3035,I169833,I170071,);
DFFARX1 I_9824 (I170071,I3035,I169833,I170088,);
not I_9825 (I170096,I170088);
not I_9826 (I170113,I170071);
nand I_9827 (I169810,I170113,I169932);
nand I_9828 (I170144,I576339,I576345);
and I_9829 (I170161,I170144,I576357);
DFFARX1 I_9830 (I170161,I3035,I169833,I170187,);
nor I_9831 (I170195,I170187,I169859);
DFFARX1 I_9832 (I170195,I3035,I169833,I169798,);
DFFARX1 I_9833 (I170187,I3035,I169833,I169816,);
nor I_9834 (I170240,I576348,I576345);
not I_9835 (I170257,I170240);
nor I_9836 (I169819,I170096,I170257);
nand I_9837 (I169804,I170113,I170257);
nor I_9838 (I169813,I169859,I170240);
DFFARX1 I_9839 (I170240,I3035,I169833,I169822,);
not I_9840 (I170360,I3042);
DFFARX1 I_9841 (I1932,I3035,I170360,I170386,);
nand I_9842 (I170394,I2204,I1924);
and I_9843 (I170411,I170394,I1508);
DFFARX1 I_9844 (I170411,I3035,I170360,I170437,);
nor I_9845 (I170328,I170437,I170386);
not I_9846 (I170459,I170437);
DFFARX1 I_9847 (I1620,I3035,I170360,I170485,);
nand I_9848 (I170493,I170485,I2636);
not I_9849 (I170510,I170493);
DFFARX1 I_9850 (I170510,I3035,I170360,I170536,);
not I_9851 (I170352,I170536);
nor I_9852 (I170558,I170386,I170493);
nor I_9853 (I170334,I170437,I170558);
DFFARX1 I_9854 (I2380,I3035,I170360,I170598,);
DFFARX1 I_9855 (I170598,I3035,I170360,I170615,);
not I_9856 (I170623,I170615);
not I_9857 (I170640,I170598);
nand I_9858 (I170337,I170640,I170459);
nand I_9859 (I170671,I1476,I1572);
and I_9860 (I170688,I170671,I1484);
DFFARX1 I_9861 (I170688,I3035,I170360,I170714,);
nor I_9862 (I170722,I170714,I170386);
DFFARX1 I_9863 (I170722,I3035,I170360,I170325,);
DFFARX1 I_9864 (I170714,I3035,I170360,I170343,);
nor I_9865 (I170767,I2692,I1572);
not I_9866 (I170784,I170767);
nor I_9867 (I170346,I170623,I170784);
nand I_9868 (I170331,I170640,I170784);
nor I_9869 (I170340,I170386,I170767);
DFFARX1 I_9870 (I170767,I3035,I170360,I170349,);
not I_9871 (I170887,I3042);
DFFARX1 I_9872 (I439829,I3035,I170887,I170913,);
nand I_9873 (I170921,I439832,I439826);
and I_9874 (I170938,I170921,I439838);
DFFARX1 I_9875 (I170938,I3035,I170887,I170964,);
nor I_9876 (I170855,I170964,I170913);
not I_9877 (I170986,I170964);
DFFARX1 I_9878 (I439841,I3035,I170887,I171012,);
nand I_9879 (I171020,I171012,I439832);
not I_9880 (I171037,I171020);
DFFARX1 I_9881 (I171037,I3035,I170887,I171063,);
not I_9882 (I170879,I171063);
nor I_9883 (I171085,I170913,I171020);
nor I_9884 (I170861,I170964,I171085);
DFFARX1 I_9885 (I439844,I3035,I170887,I171125,);
DFFARX1 I_9886 (I171125,I3035,I170887,I171142,);
not I_9887 (I171150,I171142);
not I_9888 (I171167,I171125);
nand I_9889 (I170864,I171167,I170986);
nand I_9890 (I171198,I439826,I439835);
and I_9891 (I171215,I171198,I439829);
DFFARX1 I_9892 (I171215,I3035,I170887,I171241,);
nor I_9893 (I171249,I171241,I170913);
DFFARX1 I_9894 (I171249,I3035,I170887,I170852,);
DFFARX1 I_9895 (I171241,I3035,I170887,I170870,);
nor I_9896 (I171294,I439847,I439835);
not I_9897 (I171311,I171294);
nor I_9898 (I170873,I171150,I171311);
nand I_9899 (I170858,I171167,I171311);
nor I_9900 (I170867,I170913,I171294);
DFFARX1 I_9901 (I171294,I3035,I170887,I170876,);
not I_9902 (I171414,I3042);
DFFARX1 I_9903 (I61035,I3035,I171414,I171440,);
nand I_9904 (I171448,I61047,I61056);
and I_9905 (I171465,I171448,I61035);
DFFARX1 I_9906 (I171465,I3035,I171414,I171491,);
nor I_9907 (I171382,I171491,I171440);
not I_9908 (I171513,I171491);
DFFARX1 I_9909 (I61050,I3035,I171414,I171539,);
nand I_9910 (I171547,I171539,I61038);
not I_9911 (I171564,I171547);
DFFARX1 I_9912 (I171564,I3035,I171414,I171590,);
not I_9913 (I171406,I171590);
nor I_9914 (I171612,I171440,I171547);
nor I_9915 (I171388,I171491,I171612);
DFFARX1 I_9916 (I61041,I3035,I171414,I171652,);
DFFARX1 I_9917 (I171652,I3035,I171414,I171669,);
not I_9918 (I171677,I171669);
not I_9919 (I171694,I171652);
nand I_9920 (I171391,I171694,I171513);
nand I_9921 (I171725,I61032,I61032);
and I_9922 (I171742,I171725,I61044);
DFFARX1 I_9923 (I171742,I3035,I171414,I171768,);
nor I_9924 (I171776,I171768,I171440);
DFFARX1 I_9925 (I171776,I3035,I171414,I171379,);
DFFARX1 I_9926 (I171768,I3035,I171414,I171397,);
nor I_9927 (I171821,I61053,I61032);
not I_9928 (I171838,I171821);
nor I_9929 (I171400,I171677,I171838);
nand I_9930 (I171385,I171694,I171838);
nor I_9931 (I171394,I171440,I171821);
DFFARX1 I_9932 (I171821,I3035,I171414,I171403,);
not I_9933 (I171941,I3042);
DFFARX1 I_9934 (I670296,I3035,I171941,I171967,);
nand I_9935 (I171975,I670278,I670302);
and I_9936 (I171992,I171975,I670293);
DFFARX1 I_9937 (I171992,I3035,I171941,I172018,);
nor I_9938 (I171909,I172018,I171967);
not I_9939 (I172040,I172018);
DFFARX1 I_9940 (I670299,I3035,I171941,I172066,);
nand I_9941 (I172074,I172066,I670287);
not I_9942 (I172091,I172074);
DFFARX1 I_9943 (I172091,I3035,I171941,I172117,);
not I_9944 (I171933,I172117);
nor I_9945 (I172139,I171967,I172074);
nor I_9946 (I171915,I172018,I172139);
DFFARX1 I_9947 (I670278,I3035,I171941,I172179,);
DFFARX1 I_9948 (I172179,I3035,I171941,I172196,);
not I_9949 (I172204,I172196);
not I_9950 (I172221,I172179);
nand I_9951 (I171918,I172221,I172040);
nand I_9952 (I172252,I670284,I670281);
and I_9953 (I172269,I172252,I670290);
DFFARX1 I_9954 (I172269,I3035,I171941,I172295,);
nor I_9955 (I172303,I172295,I171967);
DFFARX1 I_9956 (I172303,I3035,I171941,I171906,);
DFFARX1 I_9957 (I172295,I3035,I171941,I171924,);
nor I_9958 (I172348,I670281,I670281);
not I_9959 (I172365,I172348);
nor I_9960 (I171927,I172204,I172365);
nand I_9961 (I171912,I172221,I172365);
nor I_9962 (I171921,I171967,I172348);
DFFARX1 I_9963 (I172348,I3035,I171941,I171930,);
not I_9964 (I172468,I3042);
DFFARX1 I_9965 (I473030,I3035,I172468,I172494,);
nand I_9966 (I172502,I473033,I473027);
and I_9967 (I172519,I172502,I473039);
DFFARX1 I_9968 (I172519,I3035,I172468,I172545,);
nor I_9969 (I172436,I172545,I172494);
not I_9970 (I172567,I172545);
DFFARX1 I_9971 (I473042,I3035,I172468,I172593,);
nand I_9972 (I172601,I172593,I473033);
not I_9973 (I172618,I172601);
DFFARX1 I_9974 (I172618,I3035,I172468,I172644,);
not I_9975 (I172460,I172644);
nor I_9976 (I172666,I172494,I172601);
nor I_9977 (I172442,I172545,I172666);
DFFARX1 I_9978 (I473045,I3035,I172468,I172706,);
DFFARX1 I_9979 (I172706,I3035,I172468,I172723,);
not I_9980 (I172731,I172723);
not I_9981 (I172748,I172706);
nand I_9982 (I172445,I172748,I172567);
nand I_9983 (I172779,I473027,I473036);
and I_9984 (I172796,I172779,I473030);
DFFARX1 I_9985 (I172796,I3035,I172468,I172822,);
nor I_9986 (I172830,I172822,I172494);
DFFARX1 I_9987 (I172830,I3035,I172468,I172433,);
DFFARX1 I_9988 (I172822,I3035,I172468,I172451,);
nor I_9989 (I172875,I473048,I473036);
not I_9990 (I172892,I172875);
nor I_9991 (I172454,I172731,I172892);
nand I_9992 (I172439,I172748,I172892);
nor I_9993 (I172448,I172494,I172875);
DFFARX1 I_9994 (I172875,I3035,I172468,I172457,);
not I_9995 (I172995,I3042);
DFFARX1 I_9996 (I460382,I3035,I172995,I173021,);
nand I_9997 (I173029,I460385,I460379);
and I_9998 (I173046,I173029,I460391);
DFFARX1 I_9999 (I173046,I3035,I172995,I173072,);
nor I_10000 (I172963,I173072,I173021);
not I_10001 (I173094,I173072);
DFFARX1 I_10002 (I460394,I3035,I172995,I173120,);
nand I_10003 (I173128,I173120,I460385);
not I_10004 (I173145,I173128);
DFFARX1 I_10005 (I173145,I3035,I172995,I173171,);
not I_10006 (I172987,I173171);
nor I_10007 (I173193,I173021,I173128);
nor I_10008 (I172969,I173072,I173193);
DFFARX1 I_10009 (I460397,I3035,I172995,I173233,);
DFFARX1 I_10010 (I173233,I3035,I172995,I173250,);
not I_10011 (I173258,I173250);
not I_10012 (I173275,I173233);
nand I_10013 (I172972,I173275,I173094);
nand I_10014 (I173306,I460379,I460388);
and I_10015 (I173323,I173306,I460382);
DFFARX1 I_10016 (I173323,I3035,I172995,I173349,);
nor I_10017 (I173357,I173349,I173021);
DFFARX1 I_10018 (I173357,I3035,I172995,I172960,);
DFFARX1 I_10019 (I173349,I3035,I172995,I172978,);
nor I_10020 (I173402,I460400,I460388);
not I_10021 (I173419,I173402);
nor I_10022 (I172981,I173258,I173419);
nand I_10023 (I172966,I173275,I173419);
nor I_10024 (I172975,I173021,I173402);
DFFARX1 I_10025 (I173402,I3035,I172995,I172984,);
not I_10026 (I173522,I3042);
DFFARX1 I_10027 (I616796,I3035,I173522,I173548,);
nand I_10028 (I173556,I616811,I616796);
and I_10029 (I173573,I173556,I616814);
DFFARX1 I_10030 (I173573,I3035,I173522,I173599,);
nor I_10031 (I173490,I173599,I173548);
not I_10032 (I173621,I173599);
DFFARX1 I_10033 (I616820,I3035,I173522,I173647,);
nand I_10034 (I173655,I173647,I616802);
not I_10035 (I173672,I173655);
DFFARX1 I_10036 (I173672,I3035,I173522,I173698,);
not I_10037 (I173514,I173698);
nor I_10038 (I173720,I173548,I173655);
nor I_10039 (I173496,I173599,I173720);
DFFARX1 I_10040 (I616799,I3035,I173522,I173760,);
DFFARX1 I_10041 (I173760,I3035,I173522,I173777,);
not I_10042 (I173785,I173777);
not I_10043 (I173802,I173760);
nand I_10044 (I173499,I173802,I173621);
nand I_10045 (I173833,I616799,I616805);
and I_10046 (I173850,I173833,I616817);
DFFARX1 I_10047 (I173850,I3035,I173522,I173876,);
nor I_10048 (I173884,I173876,I173548);
DFFARX1 I_10049 (I173884,I3035,I173522,I173487,);
DFFARX1 I_10050 (I173876,I3035,I173522,I173505,);
nor I_10051 (I173929,I616808,I616805);
not I_10052 (I173946,I173929);
nor I_10053 (I173508,I173785,I173946);
nand I_10054 (I173493,I173802,I173946);
nor I_10055 (I173502,I173548,I173929);
DFFARX1 I_10056 (I173929,I3035,I173522,I173511,);
not I_10057 (I174049,I3042);
DFFARX1 I_10058 (I661048,I3035,I174049,I174075,);
nand I_10059 (I174083,I661030,I661054);
and I_10060 (I174100,I174083,I661045);
DFFARX1 I_10061 (I174100,I3035,I174049,I174126,);
nor I_10062 (I174017,I174126,I174075);
not I_10063 (I174148,I174126);
DFFARX1 I_10064 (I661051,I3035,I174049,I174174,);
nand I_10065 (I174182,I174174,I661039);
not I_10066 (I174199,I174182);
DFFARX1 I_10067 (I174199,I3035,I174049,I174225,);
not I_10068 (I174041,I174225);
nor I_10069 (I174247,I174075,I174182);
nor I_10070 (I174023,I174126,I174247);
DFFARX1 I_10071 (I661030,I3035,I174049,I174287,);
DFFARX1 I_10072 (I174287,I3035,I174049,I174304,);
not I_10073 (I174312,I174304);
not I_10074 (I174329,I174287);
nand I_10075 (I174026,I174329,I174148);
nand I_10076 (I174360,I661036,I661033);
and I_10077 (I174377,I174360,I661042);
DFFARX1 I_10078 (I174377,I3035,I174049,I174403,);
nor I_10079 (I174411,I174403,I174075);
DFFARX1 I_10080 (I174411,I3035,I174049,I174014,);
DFFARX1 I_10081 (I174403,I3035,I174049,I174032,);
nor I_10082 (I174456,I661033,I661033);
not I_10083 (I174473,I174456);
nor I_10084 (I174035,I174312,I174473);
nand I_10085 (I174020,I174329,I174473);
nor I_10086 (I174029,I174075,I174456);
DFFARX1 I_10087 (I174456,I3035,I174049,I174038,);
not I_10088 (I174576,I3042);
DFFARX1 I_10089 (I518709,I3035,I174576,I174602,);
nand I_10090 (I174610,I518706,I518724);
and I_10091 (I174627,I174610,I518715);
DFFARX1 I_10092 (I174627,I3035,I174576,I174653,);
nor I_10093 (I174544,I174653,I174602);
not I_10094 (I174675,I174653);
DFFARX1 I_10095 (I518730,I3035,I174576,I174701,);
nand I_10096 (I174709,I174701,I518712);
not I_10097 (I174726,I174709);
DFFARX1 I_10098 (I174726,I3035,I174576,I174752,);
not I_10099 (I174568,I174752);
nor I_10100 (I174774,I174602,I174709);
nor I_10101 (I174550,I174653,I174774);
DFFARX1 I_10102 (I518718,I3035,I174576,I174814,);
DFFARX1 I_10103 (I174814,I3035,I174576,I174831,);
not I_10104 (I174839,I174831);
not I_10105 (I174856,I174814);
nand I_10106 (I174553,I174856,I174675);
nand I_10107 (I174887,I518706,I518733);
and I_10108 (I174904,I174887,I518721);
DFFARX1 I_10109 (I174904,I3035,I174576,I174930,);
nor I_10110 (I174938,I174930,I174602);
DFFARX1 I_10111 (I174938,I3035,I174576,I174541,);
DFFARX1 I_10112 (I174930,I3035,I174576,I174559,);
nor I_10113 (I174983,I518727,I518733);
not I_10114 (I175000,I174983);
nor I_10115 (I174562,I174839,I175000);
nand I_10116 (I174547,I174856,I175000);
nor I_10117 (I174556,I174602,I174983);
DFFARX1 I_10118 (I174983,I3035,I174576,I174565,);
not I_10119 (I175103,I3042);
DFFARX1 I_10120 (I665944,I3035,I175103,I175129,);
nand I_10121 (I175137,I665926,I665950);
and I_10122 (I175154,I175137,I665941);
DFFARX1 I_10123 (I175154,I3035,I175103,I175180,);
nor I_10124 (I175071,I175180,I175129);
not I_10125 (I175202,I175180);
DFFARX1 I_10126 (I665947,I3035,I175103,I175228,);
nand I_10127 (I175236,I175228,I665935);
not I_10128 (I175253,I175236);
DFFARX1 I_10129 (I175253,I3035,I175103,I175279,);
not I_10130 (I175095,I175279);
nor I_10131 (I175301,I175129,I175236);
nor I_10132 (I175077,I175180,I175301);
DFFARX1 I_10133 (I665926,I3035,I175103,I175341,);
DFFARX1 I_10134 (I175341,I3035,I175103,I175358,);
not I_10135 (I175366,I175358);
not I_10136 (I175383,I175341);
nand I_10137 (I175080,I175383,I175202);
nand I_10138 (I175414,I665932,I665929);
and I_10139 (I175431,I175414,I665938);
DFFARX1 I_10140 (I175431,I3035,I175103,I175457,);
nor I_10141 (I175465,I175457,I175129);
DFFARX1 I_10142 (I175465,I3035,I175103,I175068,);
DFFARX1 I_10143 (I175457,I3035,I175103,I175086,);
nor I_10144 (I175510,I665929,I665929);
not I_10145 (I175527,I175510);
nor I_10146 (I175089,I175366,I175527);
nand I_10147 (I175074,I175383,I175527);
nor I_10148 (I175083,I175129,I175510);
DFFARX1 I_10149 (I175510,I3035,I175103,I175092,);
not I_10150 (I175630,I3042);
DFFARX1 I_10151 (I371260,I3035,I175630,I175656,);
nand I_10152 (I175664,I371251,I371266);
and I_10153 (I175681,I175664,I371272);
DFFARX1 I_10154 (I175681,I3035,I175630,I175707,);
nor I_10155 (I175598,I175707,I175656);
not I_10156 (I175729,I175707);
DFFARX1 I_10157 (I371257,I3035,I175630,I175755,);
nand I_10158 (I175763,I175755,I371251);
not I_10159 (I175780,I175763);
DFFARX1 I_10160 (I175780,I3035,I175630,I175806,);
not I_10161 (I175622,I175806);
nor I_10162 (I175828,I175656,I175763);
nor I_10163 (I175604,I175707,I175828);
DFFARX1 I_10164 (I371254,I3035,I175630,I175868,);
DFFARX1 I_10165 (I175868,I3035,I175630,I175885,);
not I_10166 (I175893,I175885);
not I_10167 (I175910,I175868);
nand I_10168 (I175607,I175910,I175729);
nand I_10169 (I175941,I371248,I371263);
and I_10170 (I175958,I175941,I371248);
DFFARX1 I_10171 (I175958,I3035,I175630,I175984,);
nor I_10172 (I175992,I175984,I175656);
DFFARX1 I_10173 (I175992,I3035,I175630,I175595,);
DFFARX1 I_10174 (I175984,I3035,I175630,I175613,);
nor I_10175 (I176037,I371269,I371263);
not I_10176 (I176054,I176037);
nor I_10177 (I175616,I175893,I176054);
nand I_10178 (I175601,I175910,I176054);
nor I_10179 (I175610,I175656,I176037);
DFFARX1 I_10180 (I176037,I3035,I175630,I175619,);
not I_10181 (I176157,I3042);
DFFARX1 I_10182 (I525169,I3035,I176157,I176183,);
nand I_10183 (I176191,I525166,I525184);
and I_10184 (I176208,I176191,I525175);
DFFARX1 I_10185 (I176208,I3035,I176157,I176234,);
nor I_10186 (I176125,I176234,I176183);
not I_10187 (I176256,I176234);
DFFARX1 I_10188 (I525190,I3035,I176157,I176282,);
nand I_10189 (I176290,I176282,I525172);
not I_10190 (I176307,I176290);
DFFARX1 I_10191 (I176307,I3035,I176157,I176333,);
not I_10192 (I176149,I176333);
nor I_10193 (I176355,I176183,I176290);
nor I_10194 (I176131,I176234,I176355);
DFFARX1 I_10195 (I525178,I3035,I176157,I176395,);
DFFARX1 I_10196 (I176395,I3035,I176157,I176412,);
not I_10197 (I176420,I176412);
not I_10198 (I176437,I176395);
nand I_10199 (I176134,I176437,I176256);
nand I_10200 (I176468,I525166,I525193);
and I_10201 (I176485,I176468,I525181);
DFFARX1 I_10202 (I176485,I3035,I176157,I176511,);
nor I_10203 (I176519,I176511,I176183);
DFFARX1 I_10204 (I176519,I3035,I176157,I176122,);
DFFARX1 I_10205 (I176511,I3035,I176157,I176140,);
nor I_10206 (I176564,I525187,I525193);
not I_10207 (I176581,I176564);
nor I_10208 (I176143,I176420,I176581);
nand I_10209 (I176128,I176437,I176581);
nor I_10210 (I176137,I176183,I176564);
DFFARX1 I_10211 (I176564,I3035,I176157,I176146,);
not I_10212 (I176684,I3042);
DFFARX1 I_10213 (I552658,I3035,I176684,I176710,);
nand I_10214 (I176718,I552655,I552658);
and I_10215 (I176735,I176718,I552667);
DFFARX1 I_10216 (I176735,I3035,I176684,I176761,);
nor I_10217 (I176652,I176761,I176710);
not I_10218 (I176783,I176761);
DFFARX1 I_10219 (I552655,I3035,I176684,I176809,);
nand I_10220 (I176817,I176809,I552673);
not I_10221 (I176834,I176817);
DFFARX1 I_10222 (I176834,I3035,I176684,I176860,);
not I_10223 (I176676,I176860);
nor I_10224 (I176882,I176710,I176817);
nor I_10225 (I176658,I176761,I176882);
DFFARX1 I_10226 (I552661,I3035,I176684,I176922,);
DFFARX1 I_10227 (I176922,I3035,I176684,I176939,);
not I_10228 (I176947,I176939);
not I_10229 (I176964,I176922);
nand I_10230 (I176661,I176964,I176783);
nand I_10231 (I176995,I552670,I552676);
and I_10232 (I177012,I176995,I552661);
DFFARX1 I_10233 (I177012,I3035,I176684,I177038,);
nor I_10234 (I177046,I177038,I176710);
DFFARX1 I_10235 (I177046,I3035,I176684,I176649,);
DFFARX1 I_10236 (I177038,I3035,I176684,I176667,);
nor I_10237 (I177091,I552664,I552676);
not I_10238 (I177108,I177091);
nor I_10239 (I176670,I176947,I177108);
nand I_10240 (I176655,I176964,I177108);
nor I_10241 (I176664,I176710,I177091);
DFFARX1 I_10242 (I177091,I3035,I176684,I176673,);
not I_10243 (I177211,I3042);
DFFARX1 I_10244 (I412876,I3035,I177211,I177237,);
nand I_10245 (I177245,I412867,I412882);
and I_10246 (I177262,I177245,I412888);
DFFARX1 I_10247 (I177262,I3035,I177211,I177288,);
nor I_10248 (I177179,I177288,I177237);
not I_10249 (I177310,I177288);
DFFARX1 I_10250 (I412873,I3035,I177211,I177336,);
nand I_10251 (I177344,I177336,I412867);
not I_10252 (I177361,I177344);
DFFARX1 I_10253 (I177361,I3035,I177211,I177387,);
not I_10254 (I177203,I177387);
nor I_10255 (I177409,I177237,I177344);
nor I_10256 (I177185,I177288,I177409);
DFFARX1 I_10257 (I412870,I3035,I177211,I177449,);
DFFARX1 I_10258 (I177449,I3035,I177211,I177466,);
not I_10259 (I177474,I177466);
not I_10260 (I177491,I177449);
nand I_10261 (I177188,I177491,I177310);
nand I_10262 (I177522,I412864,I412879);
and I_10263 (I177539,I177522,I412864);
DFFARX1 I_10264 (I177539,I3035,I177211,I177565,);
nor I_10265 (I177573,I177565,I177237);
DFFARX1 I_10266 (I177573,I3035,I177211,I177176,);
DFFARX1 I_10267 (I177565,I3035,I177211,I177194,);
nor I_10268 (I177618,I412885,I412879);
not I_10269 (I177635,I177618);
nor I_10270 (I177197,I177474,I177635);
nand I_10271 (I177182,I177491,I177635);
nor I_10272 (I177191,I177237,I177618);
DFFARX1 I_10273 (I177618,I3035,I177211,I177200,);
not I_10274 (I177738,I3042);
DFFARX1 I_10275 (I420857,I3035,I177738,I177764,);
nand I_10276 (I177772,I420860,I420854);
and I_10277 (I177789,I177772,I420866);
DFFARX1 I_10278 (I177789,I3035,I177738,I177815,);
nor I_10279 (I177706,I177815,I177764);
not I_10280 (I177837,I177815);
DFFARX1 I_10281 (I420869,I3035,I177738,I177863,);
nand I_10282 (I177871,I177863,I420860);
not I_10283 (I177888,I177871);
DFFARX1 I_10284 (I177888,I3035,I177738,I177914,);
not I_10285 (I177730,I177914);
nor I_10286 (I177936,I177764,I177871);
nor I_10287 (I177712,I177815,I177936);
DFFARX1 I_10288 (I420872,I3035,I177738,I177976,);
DFFARX1 I_10289 (I177976,I3035,I177738,I177993,);
not I_10290 (I178001,I177993);
not I_10291 (I178018,I177976);
nand I_10292 (I177715,I178018,I177837);
nand I_10293 (I178049,I420854,I420863);
and I_10294 (I178066,I178049,I420857);
DFFARX1 I_10295 (I178066,I3035,I177738,I178092,);
nor I_10296 (I178100,I178092,I177764);
DFFARX1 I_10297 (I178100,I3035,I177738,I177703,);
DFFARX1 I_10298 (I178092,I3035,I177738,I177721,);
nor I_10299 (I178145,I420875,I420863);
not I_10300 (I178162,I178145);
nor I_10301 (I177724,I178001,I178162);
nand I_10302 (I177709,I178018,I178162);
nor I_10303 (I177718,I177764,I178145);
DFFARX1 I_10304 (I178145,I3035,I177738,I177727,);
not I_10305 (I178265,I3042);
DFFARX1 I_10306 (I699624,I3035,I178265,I178291,);
nand I_10307 (I178299,I699603,I699603);
and I_10308 (I178316,I178299,I699630);
DFFARX1 I_10309 (I178316,I3035,I178265,I178342,);
nor I_10310 (I178233,I178342,I178291);
not I_10311 (I178364,I178342);
DFFARX1 I_10312 (I699618,I3035,I178265,I178390,);
nand I_10313 (I178398,I178390,I699621);
not I_10314 (I178415,I178398);
DFFARX1 I_10315 (I178415,I3035,I178265,I178441,);
not I_10316 (I178257,I178441);
nor I_10317 (I178463,I178291,I178398);
nor I_10318 (I178239,I178342,I178463);
DFFARX1 I_10319 (I699612,I3035,I178265,I178503,);
DFFARX1 I_10320 (I178503,I3035,I178265,I178520,);
not I_10321 (I178528,I178520);
not I_10322 (I178545,I178503);
nand I_10323 (I178242,I178545,I178364);
nand I_10324 (I178576,I699609,I699606);
and I_10325 (I178593,I178576,I699627);
DFFARX1 I_10326 (I178593,I3035,I178265,I178619,);
nor I_10327 (I178627,I178619,I178291);
DFFARX1 I_10328 (I178627,I3035,I178265,I178230,);
DFFARX1 I_10329 (I178619,I3035,I178265,I178248,);
nor I_10330 (I178672,I699615,I699606);
not I_10331 (I178689,I178672);
nor I_10332 (I178251,I178528,I178689);
nand I_10333 (I178236,I178545,I178689);
nor I_10334 (I178245,I178291,I178672);
DFFARX1 I_10335 (I178672,I3035,I178265,I178254,);
not I_10336 (I178792,I3042);
DFFARX1 I_10337 (I405940,I3035,I178792,I178818,);
nand I_10338 (I178826,I405931,I405946);
and I_10339 (I178843,I178826,I405952);
DFFARX1 I_10340 (I178843,I3035,I178792,I178869,);
nor I_10341 (I178760,I178869,I178818);
not I_10342 (I178891,I178869);
DFFARX1 I_10343 (I405937,I3035,I178792,I178917,);
nand I_10344 (I178925,I178917,I405931);
not I_10345 (I178942,I178925);
DFFARX1 I_10346 (I178942,I3035,I178792,I178968,);
not I_10347 (I178784,I178968);
nor I_10348 (I178990,I178818,I178925);
nor I_10349 (I178766,I178869,I178990);
DFFARX1 I_10350 (I405934,I3035,I178792,I179030,);
DFFARX1 I_10351 (I179030,I3035,I178792,I179047,);
not I_10352 (I179055,I179047);
not I_10353 (I179072,I179030);
nand I_10354 (I178769,I179072,I178891);
nand I_10355 (I179103,I405928,I405943);
and I_10356 (I179120,I179103,I405928);
DFFARX1 I_10357 (I179120,I3035,I178792,I179146,);
nor I_10358 (I179154,I179146,I178818);
DFFARX1 I_10359 (I179154,I3035,I178792,I178757,);
DFFARX1 I_10360 (I179146,I3035,I178792,I178775,);
nor I_10361 (I179199,I405949,I405943);
not I_10362 (I179216,I179199);
nor I_10363 (I178778,I179055,I179216);
nand I_10364 (I178763,I179072,I179216);
nor I_10365 (I178772,I178818,I179199);
DFFARX1 I_10366 (I179199,I3035,I178792,I178781,);
not I_10367 (I179319,I3042);
DFFARX1 I_10368 (I367792,I3035,I179319,I179345,);
nand I_10369 (I179353,I367783,I367798);
and I_10370 (I179370,I179353,I367804);
DFFARX1 I_10371 (I179370,I3035,I179319,I179396,);
nor I_10372 (I179287,I179396,I179345);
not I_10373 (I179418,I179396);
DFFARX1 I_10374 (I367789,I3035,I179319,I179444,);
nand I_10375 (I179452,I179444,I367783);
not I_10376 (I179469,I179452);
DFFARX1 I_10377 (I179469,I3035,I179319,I179495,);
not I_10378 (I179311,I179495);
nor I_10379 (I179517,I179345,I179452);
nor I_10380 (I179293,I179396,I179517);
DFFARX1 I_10381 (I367786,I3035,I179319,I179557,);
DFFARX1 I_10382 (I179557,I3035,I179319,I179574,);
not I_10383 (I179582,I179574);
not I_10384 (I179599,I179557);
nand I_10385 (I179296,I179599,I179418);
nand I_10386 (I179630,I367780,I367795);
and I_10387 (I179647,I179630,I367780);
DFFARX1 I_10388 (I179647,I3035,I179319,I179673,);
nor I_10389 (I179681,I179673,I179345);
DFFARX1 I_10390 (I179681,I3035,I179319,I179284,);
DFFARX1 I_10391 (I179673,I3035,I179319,I179302,);
nor I_10392 (I179726,I367801,I367795);
not I_10393 (I179743,I179726);
nor I_10394 (I179305,I179582,I179743);
nand I_10395 (I179290,I179599,I179743);
nor I_10396 (I179299,I179345,I179726);
DFFARX1 I_10397 (I179726,I3035,I179319,I179308,);
not I_10398 (I179846,I3042);
DFFARX1 I_10399 (I381086,I3035,I179846,I179872,);
nand I_10400 (I179880,I381077,I381092);
and I_10401 (I179897,I179880,I381098);
DFFARX1 I_10402 (I179897,I3035,I179846,I179923,);
nor I_10403 (I179814,I179923,I179872);
not I_10404 (I179945,I179923);
DFFARX1 I_10405 (I381083,I3035,I179846,I179971,);
nand I_10406 (I179979,I179971,I381077);
not I_10407 (I179996,I179979);
DFFARX1 I_10408 (I179996,I3035,I179846,I180022,);
not I_10409 (I179838,I180022);
nor I_10410 (I180044,I179872,I179979);
nor I_10411 (I179820,I179923,I180044);
DFFARX1 I_10412 (I381080,I3035,I179846,I180084,);
DFFARX1 I_10413 (I180084,I3035,I179846,I180101,);
not I_10414 (I180109,I180101);
not I_10415 (I180126,I180084);
nand I_10416 (I179823,I180126,I179945);
nand I_10417 (I180157,I381074,I381089);
and I_10418 (I180174,I180157,I381074);
DFFARX1 I_10419 (I180174,I3035,I179846,I180200,);
nor I_10420 (I180208,I180200,I179872);
DFFARX1 I_10421 (I180208,I3035,I179846,I179811,);
DFFARX1 I_10422 (I180200,I3035,I179846,I179829,);
nor I_10423 (I180253,I381095,I381089);
not I_10424 (I180270,I180253);
nor I_10425 (I179832,I180109,I180270);
nand I_10426 (I179817,I180126,I180270);
nor I_10427 (I179826,I179872,I180253);
DFFARX1 I_10428 (I180253,I3035,I179846,I179835,);
not I_10429 (I180373,I3042);
DFFARX1 I_10430 (I449315,I3035,I180373,I180399,);
nand I_10431 (I180407,I449318,I449312);
and I_10432 (I180424,I180407,I449324);
DFFARX1 I_10433 (I180424,I3035,I180373,I180450,);
nor I_10434 (I180341,I180450,I180399);
not I_10435 (I180472,I180450);
DFFARX1 I_10436 (I449327,I3035,I180373,I180498,);
nand I_10437 (I180506,I180498,I449318);
not I_10438 (I180523,I180506);
DFFARX1 I_10439 (I180523,I3035,I180373,I180549,);
not I_10440 (I180365,I180549);
nor I_10441 (I180571,I180399,I180506);
nor I_10442 (I180347,I180450,I180571);
DFFARX1 I_10443 (I449330,I3035,I180373,I180611,);
DFFARX1 I_10444 (I180611,I3035,I180373,I180628,);
not I_10445 (I180636,I180628);
not I_10446 (I180653,I180611);
nand I_10447 (I180350,I180653,I180472);
nand I_10448 (I180684,I449312,I449321);
and I_10449 (I180701,I180684,I449315);
DFFARX1 I_10450 (I180701,I3035,I180373,I180727,);
nor I_10451 (I180735,I180727,I180399);
DFFARX1 I_10452 (I180735,I3035,I180373,I180338,);
DFFARX1 I_10453 (I180727,I3035,I180373,I180356,);
nor I_10454 (I180780,I449333,I449321);
not I_10455 (I180797,I180780);
nor I_10456 (I180359,I180636,I180797);
nand I_10457 (I180344,I180653,I180797);
nor I_10458 (I180353,I180399,I180780);
DFFARX1 I_10459 (I180780,I3035,I180373,I180362,);
not I_10460 (I180900,I3042);
DFFARX1 I_10461 (I613906,I3035,I180900,I180926,);
nand I_10462 (I180934,I613921,I613906);
and I_10463 (I180951,I180934,I613924);
DFFARX1 I_10464 (I180951,I3035,I180900,I180977,);
nor I_10465 (I180868,I180977,I180926);
not I_10466 (I180999,I180977);
DFFARX1 I_10467 (I613930,I3035,I180900,I181025,);
nand I_10468 (I181033,I181025,I613912);
not I_10469 (I181050,I181033);
DFFARX1 I_10470 (I181050,I3035,I180900,I181076,);
not I_10471 (I180892,I181076);
nor I_10472 (I181098,I180926,I181033);
nor I_10473 (I180874,I180977,I181098);
DFFARX1 I_10474 (I613909,I3035,I180900,I181138,);
DFFARX1 I_10475 (I181138,I3035,I180900,I181155,);
not I_10476 (I181163,I181155);
not I_10477 (I181180,I181138);
nand I_10478 (I180877,I181180,I180999);
nand I_10479 (I181211,I613909,I613915);
and I_10480 (I181228,I181211,I613927);
DFFARX1 I_10481 (I181228,I3035,I180900,I181254,);
nor I_10482 (I181262,I181254,I180926);
DFFARX1 I_10483 (I181262,I3035,I180900,I180865,);
DFFARX1 I_10484 (I181254,I3035,I180900,I180883,);
nor I_10485 (I181307,I613918,I613915);
not I_10486 (I181324,I181307);
nor I_10487 (I180886,I181163,I181324);
nand I_10488 (I180871,I181180,I181324);
nor I_10489 (I180880,I180926,I181307);
DFFARX1 I_10490 (I181307,I3035,I180900,I180889,);
not I_10491 (I181427,I3042);
DFFARX1 I_10492 (I595988,I3035,I181427,I181453,);
nand I_10493 (I181461,I596003,I595988);
and I_10494 (I181478,I181461,I596006);
DFFARX1 I_10495 (I181478,I3035,I181427,I181504,);
nor I_10496 (I181395,I181504,I181453);
not I_10497 (I181526,I181504);
DFFARX1 I_10498 (I596012,I3035,I181427,I181552,);
nand I_10499 (I181560,I181552,I595994);
not I_10500 (I181577,I181560);
DFFARX1 I_10501 (I181577,I3035,I181427,I181603,);
not I_10502 (I181419,I181603);
nor I_10503 (I181625,I181453,I181560);
nor I_10504 (I181401,I181504,I181625);
DFFARX1 I_10505 (I595991,I3035,I181427,I181665,);
DFFARX1 I_10506 (I181665,I3035,I181427,I181682,);
not I_10507 (I181690,I181682);
not I_10508 (I181707,I181665);
nand I_10509 (I181404,I181707,I181526);
nand I_10510 (I181738,I595991,I595997);
and I_10511 (I181755,I181738,I596009);
DFFARX1 I_10512 (I181755,I3035,I181427,I181781,);
nor I_10513 (I181789,I181781,I181453);
DFFARX1 I_10514 (I181789,I3035,I181427,I181392,);
DFFARX1 I_10515 (I181781,I3035,I181427,I181410,);
nor I_10516 (I181834,I596000,I595997);
not I_10517 (I181851,I181834);
nor I_10518 (I181413,I181690,I181851);
nand I_10519 (I181398,I181707,I181851);
nor I_10520 (I181407,I181453,I181834);
DFFARX1 I_10521 (I181834,I3035,I181427,I181416,);
not I_10522 (I181954,I3042);
DFFARX1 I_10523 (I408252,I3035,I181954,I181980,);
nand I_10524 (I181988,I408243,I408258);
and I_10525 (I182005,I181988,I408264);
DFFARX1 I_10526 (I182005,I3035,I181954,I182031,);
nor I_10527 (I181922,I182031,I181980);
not I_10528 (I182053,I182031);
DFFARX1 I_10529 (I408249,I3035,I181954,I182079,);
nand I_10530 (I182087,I182079,I408243);
not I_10531 (I182104,I182087);
DFFARX1 I_10532 (I182104,I3035,I181954,I182130,);
not I_10533 (I181946,I182130);
nor I_10534 (I182152,I181980,I182087);
nor I_10535 (I181928,I182031,I182152);
DFFARX1 I_10536 (I408246,I3035,I181954,I182192,);
DFFARX1 I_10537 (I182192,I3035,I181954,I182209,);
not I_10538 (I182217,I182209);
not I_10539 (I182234,I182192);
nand I_10540 (I181931,I182234,I182053);
nand I_10541 (I182265,I408240,I408255);
and I_10542 (I182282,I182265,I408240);
DFFARX1 I_10543 (I182282,I3035,I181954,I182308,);
nor I_10544 (I182316,I182308,I181980);
DFFARX1 I_10545 (I182316,I3035,I181954,I181919,);
DFFARX1 I_10546 (I182308,I3035,I181954,I181937,);
nor I_10547 (I182361,I408261,I408255);
not I_10548 (I182378,I182361);
nor I_10549 (I181940,I182217,I182378);
nand I_10550 (I181925,I182234,I182378);
nor I_10551 (I181934,I181980,I182361);
DFFARX1 I_10552 (I182361,I3035,I181954,I181943,);
not I_10553 (I182481,I3042);
DFFARX1 I_10554 (I259281,I3035,I182481,I182507,);
nand I_10555 (I182515,I259293,I259272);
and I_10556 (I182532,I182515,I259296);
DFFARX1 I_10557 (I182532,I3035,I182481,I182558,);
nor I_10558 (I182449,I182558,I182507);
not I_10559 (I182580,I182558);
DFFARX1 I_10560 (I259287,I3035,I182481,I182606,);
nand I_10561 (I182614,I182606,I259269);
not I_10562 (I182631,I182614);
DFFARX1 I_10563 (I182631,I3035,I182481,I182657,);
not I_10564 (I182473,I182657);
nor I_10565 (I182679,I182507,I182614);
nor I_10566 (I182455,I182558,I182679);
DFFARX1 I_10567 (I259284,I3035,I182481,I182719,);
DFFARX1 I_10568 (I182719,I3035,I182481,I182736,);
not I_10569 (I182744,I182736);
not I_10570 (I182761,I182719);
nand I_10571 (I182458,I182761,I182580);
nand I_10572 (I182792,I259269,I259275);
and I_10573 (I182809,I182792,I259278);
DFFARX1 I_10574 (I182809,I3035,I182481,I182835,);
nor I_10575 (I182843,I182835,I182507);
DFFARX1 I_10576 (I182843,I3035,I182481,I182446,);
DFFARX1 I_10577 (I182835,I3035,I182481,I182464,);
nor I_10578 (I182888,I259290,I259275);
not I_10579 (I182905,I182888);
nor I_10580 (I182467,I182744,I182905);
nand I_10581 (I182452,I182761,I182905);
nor I_10582 (I182461,I182507,I182888);
DFFARX1 I_10583 (I182888,I3035,I182481,I182470,);
not I_10584 (I183008,I3042);
DFFARX1 I_10585 (I90204,I3035,I183008,I183034,);
nand I_10586 (I183042,I90204,I90210);
and I_10587 (I183059,I183042,I90228);
DFFARX1 I_10588 (I183059,I3035,I183008,I183085,);
nor I_10589 (I182976,I183085,I183034);
not I_10590 (I183107,I183085);
DFFARX1 I_10591 (I90216,I3035,I183008,I183133,);
nand I_10592 (I183141,I183133,I90213);
not I_10593 (I183158,I183141);
DFFARX1 I_10594 (I183158,I3035,I183008,I183184,);
not I_10595 (I183000,I183184);
nor I_10596 (I183206,I183034,I183141);
nor I_10597 (I182982,I183085,I183206);
DFFARX1 I_10598 (I90222,I3035,I183008,I183246,);
DFFARX1 I_10599 (I183246,I3035,I183008,I183263,);
not I_10600 (I183271,I183263);
not I_10601 (I183288,I183246);
nand I_10602 (I182985,I183288,I183107);
nand I_10603 (I183319,I90207,I90207);
and I_10604 (I183336,I183319,I90219);
DFFARX1 I_10605 (I183336,I3035,I183008,I183362,);
nor I_10606 (I183370,I183362,I183034);
DFFARX1 I_10607 (I183370,I3035,I183008,I182973,);
DFFARX1 I_10608 (I183362,I3035,I183008,I182991,);
nor I_10609 (I183415,I90225,I90207);
not I_10610 (I183432,I183415);
nor I_10611 (I182994,I183271,I183432);
nand I_10612 (I182979,I183288,I183432);
nor I_10613 (I182988,I183034,I183415);
DFFARX1 I_10614 (I183415,I3035,I183008,I182997,);
not I_10615 (I183535,I3042);
DFFARX1 I_10616 (I46279,I3035,I183535,I183561,);
nand I_10617 (I183569,I46291,I46300);
and I_10618 (I183586,I183569,I46279);
DFFARX1 I_10619 (I183586,I3035,I183535,I183612,);
nor I_10620 (I183503,I183612,I183561);
not I_10621 (I183634,I183612);
DFFARX1 I_10622 (I46294,I3035,I183535,I183660,);
nand I_10623 (I183668,I183660,I46282);
not I_10624 (I183685,I183668);
DFFARX1 I_10625 (I183685,I3035,I183535,I183711,);
not I_10626 (I183527,I183711);
nor I_10627 (I183733,I183561,I183668);
nor I_10628 (I183509,I183612,I183733);
DFFARX1 I_10629 (I46285,I3035,I183535,I183773,);
DFFARX1 I_10630 (I183773,I3035,I183535,I183790,);
not I_10631 (I183798,I183790);
not I_10632 (I183815,I183773);
nand I_10633 (I183512,I183815,I183634);
nand I_10634 (I183846,I46276,I46276);
and I_10635 (I183863,I183846,I46288);
DFFARX1 I_10636 (I183863,I3035,I183535,I183889,);
nor I_10637 (I183897,I183889,I183561);
DFFARX1 I_10638 (I183897,I3035,I183535,I183500,);
DFFARX1 I_10639 (I183889,I3035,I183535,I183518,);
nor I_10640 (I183942,I46297,I46276);
not I_10641 (I183959,I183942);
nor I_10642 (I183521,I183798,I183959);
nand I_10643 (I183506,I183815,I183959);
nor I_10644 (I183515,I183561,I183942);
DFFARX1 I_10645 (I183942,I3035,I183535,I183524,);
not I_10646 (I184062,I3042);
DFFARX1 I_10647 (I674815,I3035,I184062,I184088,);
nand I_10648 (I184096,I674812,I674803);
and I_10649 (I184113,I184096,I674800);
DFFARX1 I_10650 (I184113,I3035,I184062,I184139,);
nor I_10651 (I184030,I184139,I184088);
not I_10652 (I184161,I184139);
DFFARX1 I_10653 (I674809,I3035,I184062,I184187,);
nand I_10654 (I184195,I184187,I674818);
not I_10655 (I184212,I184195);
DFFARX1 I_10656 (I184212,I3035,I184062,I184238,);
not I_10657 (I184054,I184238);
nor I_10658 (I184260,I184088,I184195);
nor I_10659 (I184036,I184139,I184260);
DFFARX1 I_10660 (I674821,I3035,I184062,I184300,);
DFFARX1 I_10661 (I184300,I3035,I184062,I184317,);
not I_10662 (I184325,I184317);
not I_10663 (I184342,I184300);
nand I_10664 (I184039,I184342,I184161);
nand I_10665 (I184373,I674800,I674806);
and I_10666 (I184390,I184373,I674824);
DFFARX1 I_10667 (I184390,I3035,I184062,I184416,);
nor I_10668 (I184424,I184416,I184088);
DFFARX1 I_10669 (I184424,I3035,I184062,I184027,);
DFFARX1 I_10670 (I184416,I3035,I184062,I184045,);
nor I_10671 (I184469,I674803,I674806);
not I_10672 (I184486,I184469);
nor I_10673 (I184048,I184325,I184486);
nand I_10674 (I184033,I184342,I184486);
nor I_10675 (I184042,I184088,I184469);
DFFARX1 I_10676 (I184469,I3035,I184062,I184051,);
not I_10677 (I184589,I3042);
DFFARX1 I_10678 (I669752,I3035,I184589,I184615,);
nand I_10679 (I184623,I669734,I669758);
and I_10680 (I184640,I184623,I669749);
DFFARX1 I_10681 (I184640,I3035,I184589,I184666,);
nor I_10682 (I184557,I184666,I184615);
not I_10683 (I184688,I184666);
DFFARX1 I_10684 (I669755,I3035,I184589,I184714,);
nand I_10685 (I184722,I184714,I669743);
not I_10686 (I184739,I184722);
DFFARX1 I_10687 (I184739,I3035,I184589,I184765,);
not I_10688 (I184581,I184765);
nor I_10689 (I184787,I184615,I184722);
nor I_10690 (I184563,I184666,I184787);
DFFARX1 I_10691 (I669734,I3035,I184589,I184827,);
DFFARX1 I_10692 (I184827,I3035,I184589,I184844,);
not I_10693 (I184852,I184844);
not I_10694 (I184869,I184827);
nand I_10695 (I184566,I184869,I184688);
nand I_10696 (I184900,I669740,I669737);
and I_10697 (I184917,I184900,I669746);
DFFARX1 I_10698 (I184917,I3035,I184589,I184943,);
nor I_10699 (I184951,I184943,I184615);
DFFARX1 I_10700 (I184951,I3035,I184589,I184554,);
DFFARX1 I_10701 (I184943,I3035,I184589,I184572,);
nor I_10702 (I184996,I669737,I669737);
not I_10703 (I185013,I184996);
nor I_10704 (I184575,I184852,I185013);
nand I_10705 (I184560,I184869,I185013);
nor I_10706 (I184569,I184615,I184996);
DFFARX1 I_10707 (I184996,I3035,I184589,I184578,);
not I_10708 (I185116,I3042);
DFFARX1 I_10709 (I143754,I3035,I185116,I185142,);
nand I_10710 (I185150,I143754,I143760);
and I_10711 (I185167,I185150,I143778);
DFFARX1 I_10712 (I185167,I3035,I185116,I185193,);
nor I_10713 (I185084,I185193,I185142);
not I_10714 (I185215,I185193);
DFFARX1 I_10715 (I143766,I3035,I185116,I185241,);
nand I_10716 (I185249,I185241,I143763);
not I_10717 (I185266,I185249);
DFFARX1 I_10718 (I185266,I3035,I185116,I185292,);
not I_10719 (I185108,I185292);
nor I_10720 (I185314,I185142,I185249);
nor I_10721 (I185090,I185193,I185314);
DFFARX1 I_10722 (I143772,I3035,I185116,I185354,);
DFFARX1 I_10723 (I185354,I3035,I185116,I185371,);
not I_10724 (I185379,I185371);
not I_10725 (I185396,I185354);
nand I_10726 (I185093,I185396,I185215);
nand I_10727 (I185427,I143757,I143757);
and I_10728 (I185444,I185427,I143769);
DFFARX1 I_10729 (I185444,I3035,I185116,I185470,);
nor I_10730 (I185478,I185470,I185142);
DFFARX1 I_10731 (I185478,I3035,I185116,I185081,);
DFFARX1 I_10732 (I185470,I3035,I185116,I185099,);
nor I_10733 (I185523,I143775,I143757);
not I_10734 (I185540,I185523);
nor I_10735 (I185102,I185379,I185540);
nand I_10736 (I185087,I185396,I185540);
nor I_10737 (I185096,I185142,I185523);
DFFARX1 I_10738 (I185523,I3035,I185116,I185105,);
not I_10739 (I185643,I3042);
DFFARX1 I_10740 (I570049,I3035,I185643,I185669,);
nand I_10741 (I185677,I570046,I570049);
and I_10742 (I185694,I185677,I570058);
DFFARX1 I_10743 (I185694,I3035,I185643,I185720,);
nor I_10744 (I185611,I185720,I185669);
not I_10745 (I185742,I185720);
DFFARX1 I_10746 (I570046,I3035,I185643,I185768,);
nand I_10747 (I185776,I185768,I570064);
not I_10748 (I185793,I185776);
DFFARX1 I_10749 (I185793,I3035,I185643,I185819,);
not I_10750 (I185635,I185819);
nor I_10751 (I185841,I185669,I185776);
nor I_10752 (I185617,I185720,I185841);
DFFARX1 I_10753 (I570052,I3035,I185643,I185881,);
DFFARX1 I_10754 (I185881,I3035,I185643,I185898,);
not I_10755 (I185906,I185898);
not I_10756 (I185923,I185881);
nand I_10757 (I185620,I185923,I185742);
nand I_10758 (I185954,I570061,I570067);
and I_10759 (I185971,I185954,I570052);
DFFARX1 I_10760 (I185971,I3035,I185643,I185997,);
nor I_10761 (I186005,I185997,I185669);
DFFARX1 I_10762 (I186005,I3035,I185643,I185608,);
DFFARX1 I_10763 (I185997,I3035,I185643,I185626,);
nor I_10764 (I186050,I570055,I570067);
not I_10765 (I186067,I186050);
nor I_10766 (I185629,I185906,I186067);
nand I_10767 (I185614,I185923,I186067);
nor I_10768 (I185623,I185669,I186050);
DFFARX1 I_10769 (I186050,I3035,I185643,I185632,);
not I_10770 (I186170,I3042);
DFFARX1 I_10771 (I79494,I3035,I186170,I186196,);
nand I_10772 (I186204,I79494,I79500);
and I_10773 (I186221,I186204,I79518);
DFFARX1 I_10774 (I186221,I3035,I186170,I186247,);
nor I_10775 (I186138,I186247,I186196);
not I_10776 (I186269,I186247);
DFFARX1 I_10777 (I79506,I3035,I186170,I186295,);
nand I_10778 (I186303,I186295,I79503);
not I_10779 (I186320,I186303);
DFFARX1 I_10780 (I186320,I3035,I186170,I186346,);
not I_10781 (I186162,I186346);
nor I_10782 (I186368,I186196,I186303);
nor I_10783 (I186144,I186247,I186368);
DFFARX1 I_10784 (I79512,I3035,I186170,I186408,);
DFFARX1 I_10785 (I186408,I3035,I186170,I186425,);
not I_10786 (I186433,I186425);
not I_10787 (I186450,I186408);
nand I_10788 (I186147,I186450,I186269);
nand I_10789 (I186481,I79497,I79497);
and I_10790 (I186498,I186481,I79509);
DFFARX1 I_10791 (I186498,I3035,I186170,I186524,);
nor I_10792 (I186532,I186524,I186196);
DFFARX1 I_10793 (I186532,I3035,I186170,I186135,);
DFFARX1 I_10794 (I186524,I3035,I186170,I186153,);
nor I_10795 (I186577,I79515,I79497);
not I_10796 (I186594,I186577);
nor I_10797 (I186156,I186433,I186594);
nand I_10798 (I186141,I186450,I186594);
nor I_10799 (I186150,I186196,I186577);
DFFARX1 I_10800 (I186577,I3035,I186170,I186159,);
not I_10801 (I186697,I3042);
DFFARX1 I_10802 (I284109,I3035,I186697,I186723,);
nand I_10803 (I186731,I284109,I284121);
and I_10804 (I186748,I186731,I284106);
DFFARX1 I_10805 (I186748,I3035,I186697,I186774,);
nor I_10806 (I186665,I186774,I186723);
not I_10807 (I186796,I186774);
DFFARX1 I_10808 (I284130,I3035,I186697,I186822,);
nand I_10809 (I186830,I186822,I284127);
not I_10810 (I186847,I186830);
DFFARX1 I_10811 (I186847,I3035,I186697,I186873,);
not I_10812 (I186689,I186873);
nor I_10813 (I186895,I186723,I186830);
nor I_10814 (I186671,I186774,I186895);
DFFARX1 I_10815 (I284118,I3035,I186697,I186935,);
DFFARX1 I_10816 (I186935,I3035,I186697,I186952,);
not I_10817 (I186960,I186952);
not I_10818 (I186977,I186935);
nand I_10819 (I186674,I186977,I186796);
nand I_10820 (I187008,I284106,I284115);
and I_10821 (I187025,I187008,I284124);
DFFARX1 I_10822 (I187025,I3035,I186697,I187051,);
nor I_10823 (I187059,I187051,I186723);
DFFARX1 I_10824 (I187059,I3035,I186697,I186662,);
DFFARX1 I_10825 (I187051,I3035,I186697,I186680,);
nor I_10826 (I187104,I284112,I284115);
not I_10827 (I187121,I187104);
nor I_10828 (I186683,I186960,I187121);
nand I_10829 (I186668,I186977,I187121);
nor I_10830 (I186677,I186723,I187104);
DFFARX1 I_10831 (I187104,I3035,I186697,I186686,);
not I_10832 (I187224,I3042);
DFFARX1 I_10833 (I146729,I3035,I187224,I187250,);
nand I_10834 (I187258,I146729,I146735);
and I_10835 (I187275,I187258,I146753);
DFFARX1 I_10836 (I187275,I3035,I187224,I187301,);
nor I_10837 (I187192,I187301,I187250);
not I_10838 (I187323,I187301);
DFFARX1 I_10839 (I146741,I3035,I187224,I187349,);
nand I_10840 (I187357,I187349,I146738);
not I_10841 (I187374,I187357);
DFFARX1 I_10842 (I187374,I3035,I187224,I187400,);
not I_10843 (I187216,I187400);
nor I_10844 (I187422,I187250,I187357);
nor I_10845 (I187198,I187301,I187422);
DFFARX1 I_10846 (I146747,I3035,I187224,I187462,);
DFFARX1 I_10847 (I187462,I3035,I187224,I187479,);
not I_10848 (I187487,I187479);
not I_10849 (I187504,I187462);
nand I_10850 (I187201,I187504,I187323);
nand I_10851 (I187535,I146732,I146732);
and I_10852 (I187552,I187535,I146744);
DFFARX1 I_10853 (I187552,I3035,I187224,I187578,);
nor I_10854 (I187586,I187578,I187250);
DFFARX1 I_10855 (I187586,I3035,I187224,I187189,);
DFFARX1 I_10856 (I187578,I3035,I187224,I187207,);
nor I_10857 (I187631,I146750,I146732);
not I_10858 (I187648,I187631);
nor I_10859 (I187210,I187487,I187648);
nand I_10860 (I187195,I187504,I187648);
nor I_10861 (I187204,I187250,I187631);
DFFARX1 I_10862 (I187631,I3035,I187224,I187213,);
not I_10863 (I187751,I3042);
DFFARX1 I_10864 (I742464,I3035,I187751,I187777,);
nand I_10865 (I187785,I742443,I742443);
and I_10866 (I187802,I187785,I742470);
DFFARX1 I_10867 (I187802,I3035,I187751,I187828,);
nor I_10868 (I187719,I187828,I187777);
not I_10869 (I187850,I187828);
DFFARX1 I_10870 (I742458,I3035,I187751,I187876,);
nand I_10871 (I187884,I187876,I742461);
not I_10872 (I187901,I187884);
DFFARX1 I_10873 (I187901,I3035,I187751,I187927,);
not I_10874 (I187743,I187927);
nor I_10875 (I187949,I187777,I187884);
nor I_10876 (I187725,I187828,I187949);
DFFARX1 I_10877 (I742452,I3035,I187751,I187989,);
DFFARX1 I_10878 (I187989,I3035,I187751,I188006,);
not I_10879 (I188014,I188006);
not I_10880 (I188031,I187989);
nand I_10881 (I187728,I188031,I187850);
nand I_10882 (I188062,I742449,I742446);
and I_10883 (I188079,I188062,I742467);
DFFARX1 I_10884 (I188079,I3035,I187751,I188105,);
nor I_10885 (I188113,I188105,I187777);
DFFARX1 I_10886 (I188113,I3035,I187751,I187716,);
DFFARX1 I_10887 (I188105,I3035,I187751,I187734,);
nor I_10888 (I188158,I742455,I742446);
not I_10889 (I188175,I188158);
nor I_10890 (I187737,I188014,I188175);
nand I_10891 (I187722,I188031,I188175);
nor I_10892 (I187731,I187777,I188158);
DFFARX1 I_10893 (I188158,I3035,I187751,I187740,);
not I_10894 (I188278,I3042);
DFFARX1 I_10895 (I481241,I3035,I188278,I188304,);
nand I_10896 (I188312,I481238,I481256);
and I_10897 (I188329,I188312,I481247);
DFFARX1 I_10898 (I188329,I3035,I188278,I188355,);
nor I_10899 (I188246,I188355,I188304);
not I_10900 (I188377,I188355);
DFFARX1 I_10901 (I481262,I3035,I188278,I188403,);
nand I_10902 (I188411,I188403,I481244);
not I_10903 (I188428,I188411);
DFFARX1 I_10904 (I188428,I3035,I188278,I188454,);
not I_10905 (I188270,I188454);
nor I_10906 (I188476,I188304,I188411);
nor I_10907 (I188252,I188355,I188476);
DFFARX1 I_10908 (I481250,I3035,I188278,I188516,);
DFFARX1 I_10909 (I188516,I3035,I188278,I188533,);
not I_10910 (I188541,I188533);
not I_10911 (I188558,I188516);
nand I_10912 (I188255,I188558,I188377);
nand I_10913 (I188589,I481238,I481265);
and I_10914 (I188606,I188589,I481253);
DFFARX1 I_10915 (I188606,I3035,I188278,I188632,);
nor I_10916 (I188640,I188632,I188304);
DFFARX1 I_10917 (I188640,I3035,I188278,I188243,);
DFFARX1 I_10918 (I188632,I3035,I188278,I188261,);
nor I_10919 (I188685,I481259,I481265);
not I_10920 (I188702,I188685);
nor I_10921 (I188264,I188541,I188702);
nand I_10922 (I188249,I188558,I188702);
nor I_10923 (I188258,I188304,I188685);
DFFARX1 I_10924 (I188685,I3035,I188278,I188267,);
not I_10925 (I188805,I3042);
DFFARX1 I_10926 (I711524,I3035,I188805,I188831,);
nand I_10927 (I188839,I711503,I711503);
and I_10928 (I188856,I188839,I711530);
DFFARX1 I_10929 (I188856,I3035,I188805,I188882,);
nor I_10930 (I188773,I188882,I188831);
not I_10931 (I188904,I188882);
DFFARX1 I_10932 (I711518,I3035,I188805,I188930,);
nand I_10933 (I188938,I188930,I711521);
not I_10934 (I188955,I188938);
DFFARX1 I_10935 (I188955,I3035,I188805,I188981,);
not I_10936 (I188797,I188981);
nor I_10937 (I189003,I188831,I188938);
nor I_10938 (I188779,I188882,I189003);
DFFARX1 I_10939 (I711512,I3035,I188805,I189043,);
DFFARX1 I_10940 (I189043,I3035,I188805,I189060,);
not I_10941 (I189068,I189060);
not I_10942 (I189085,I189043);
nand I_10943 (I188782,I189085,I188904);
nand I_10944 (I189116,I711509,I711506);
and I_10945 (I189133,I189116,I711527);
DFFARX1 I_10946 (I189133,I3035,I188805,I189159,);
nor I_10947 (I189167,I189159,I188831);
DFFARX1 I_10948 (I189167,I3035,I188805,I188770,);
DFFARX1 I_10949 (I189159,I3035,I188805,I188788,);
nor I_10950 (I189212,I711515,I711506);
not I_10951 (I189229,I189212);
nor I_10952 (I188791,I189068,I189229);
nand I_10953 (I188776,I189085,I189229);
nor I_10954 (I188785,I188831,I189212);
DFFARX1 I_10955 (I189212,I3035,I188805,I188794,);
not I_10956 (I189332,I3042);
DFFARX1 I_10957 (I323867,I3035,I189332,I189358,);
nand I_10958 (I189366,I323852,I323855);
and I_10959 (I189383,I189366,I323870);
DFFARX1 I_10960 (I189383,I3035,I189332,I189409,);
nor I_10961 (I189300,I189409,I189358);
not I_10962 (I189431,I189409);
DFFARX1 I_10963 (I323864,I3035,I189332,I189457,);
nand I_10964 (I189465,I189457,I323855);
not I_10965 (I189482,I189465);
DFFARX1 I_10966 (I189482,I3035,I189332,I189508,);
not I_10967 (I189324,I189508);
nor I_10968 (I189530,I189358,I189465);
nor I_10969 (I189306,I189409,I189530);
DFFARX1 I_10970 (I323861,I3035,I189332,I189570,);
DFFARX1 I_10971 (I189570,I3035,I189332,I189587,);
not I_10972 (I189595,I189587);
not I_10973 (I189612,I189570);
nand I_10974 (I189309,I189612,I189431);
nand I_10975 (I189643,I323876,I323852);
and I_10976 (I189660,I189643,I323873);
DFFARX1 I_10977 (I189660,I3035,I189332,I189686,);
nor I_10978 (I189694,I189686,I189358);
DFFARX1 I_10979 (I189694,I3035,I189332,I189297,);
DFFARX1 I_10980 (I189686,I3035,I189332,I189315,);
nor I_10981 (I189739,I323858,I323852);
not I_10982 (I189756,I189739);
nor I_10983 (I189318,I189595,I189756);
nand I_10984 (I189303,I189612,I189756);
nor I_10985 (I189312,I189358,I189739);
DFFARX1 I_10986 (I189739,I3035,I189332,I189321,);
not I_10987 (I189859,I3042);
DFFARX1 I_10988 (I372994,I3035,I189859,I189885,);
nand I_10989 (I189893,I372985,I373000);
and I_10990 (I189910,I189893,I373006);
DFFARX1 I_10991 (I189910,I3035,I189859,I189936,);
nor I_10992 (I189827,I189936,I189885);
not I_10993 (I189958,I189936);
DFFARX1 I_10994 (I372991,I3035,I189859,I189984,);
nand I_10995 (I189992,I189984,I372985);
not I_10996 (I190009,I189992);
DFFARX1 I_10997 (I190009,I3035,I189859,I190035,);
not I_10998 (I189851,I190035);
nor I_10999 (I190057,I189885,I189992);
nor I_11000 (I189833,I189936,I190057);
DFFARX1 I_11001 (I372988,I3035,I189859,I190097,);
DFFARX1 I_11002 (I190097,I3035,I189859,I190114,);
not I_11003 (I190122,I190114);
not I_11004 (I190139,I190097);
nand I_11005 (I189836,I190139,I189958);
nand I_11006 (I190170,I372982,I372997);
and I_11007 (I190187,I190170,I372982);
DFFARX1 I_11008 (I190187,I3035,I189859,I190213,);
nor I_11009 (I190221,I190213,I189885);
DFFARX1 I_11010 (I190221,I3035,I189859,I189824,);
DFFARX1 I_11011 (I190213,I3035,I189859,I189842,);
nor I_11012 (I190266,I373003,I372997);
not I_11013 (I190283,I190266);
nor I_11014 (I189845,I190122,I190283);
nand I_11015 (I189830,I190139,I190283);
nor I_11016 (I189839,I189885,I190266);
DFFARX1 I_11017 (I190266,I3035,I189859,I189848,);
not I_11018 (I190386,I3042);
DFFARX1 I_11019 (I628356,I3035,I190386,I190412,);
nand I_11020 (I190420,I628371,I628356);
and I_11021 (I190437,I190420,I628374);
DFFARX1 I_11022 (I190437,I3035,I190386,I190463,);
nor I_11023 (I190354,I190463,I190412);
not I_11024 (I190485,I190463);
DFFARX1 I_11025 (I628380,I3035,I190386,I190511,);
nand I_11026 (I190519,I190511,I628362);
not I_11027 (I190536,I190519);
DFFARX1 I_11028 (I190536,I3035,I190386,I190562,);
not I_11029 (I190378,I190562);
nor I_11030 (I190584,I190412,I190519);
nor I_11031 (I190360,I190463,I190584);
DFFARX1 I_11032 (I628359,I3035,I190386,I190624,);
DFFARX1 I_11033 (I190624,I3035,I190386,I190641,);
not I_11034 (I190649,I190641);
not I_11035 (I190666,I190624);
nand I_11036 (I190363,I190666,I190485);
nand I_11037 (I190697,I628359,I628365);
and I_11038 (I190714,I190697,I628377);
DFFARX1 I_11039 (I190714,I3035,I190386,I190740,);
nor I_11040 (I190748,I190740,I190412);
DFFARX1 I_11041 (I190748,I3035,I190386,I190351,);
DFFARX1 I_11042 (I190740,I3035,I190386,I190369,);
nor I_11043 (I190793,I628368,I628365);
not I_11044 (I190810,I190793);
nor I_11045 (I190372,I190649,I190810);
nand I_11046 (I190357,I190666,I190810);
nor I_11047 (I190366,I190412,I190793);
DFFARX1 I_11048 (I190793,I3035,I190386,I190375,);
not I_11049 (I190913,I3042);
DFFARX1 I_11050 (I38374,I3035,I190913,I190939,);
nand I_11051 (I190947,I38386,I38395);
and I_11052 (I190964,I190947,I38374);
DFFARX1 I_11053 (I190964,I3035,I190913,I190990,);
nor I_11054 (I190881,I190990,I190939);
not I_11055 (I191012,I190990);
DFFARX1 I_11056 (I38389,I3035,I190913,I191038,);
nand I_11057 (I191046,I191038,I38377);
not I_11058 (I191063,I191046);
DFFARX1 I_11059 (I191063,I3035,I190913,I191089,);
not I_11060 (I190905,I191089);
nor I_11061 (I191111,I190939,I191046);
nor I_11062 (I190887,I190990,I191111);
DFFARX1 I_11063 (I38380,I3035,I190913,I191151,);
DFFARX1 I_11064 (I191151,I3035,I190913,I191168,);
not I_11065 (I191176,I191168);
not I_11066 (I191193,I191151);
nand I_11067 (I190890,I191193,I191012);
nand I_11068 (I191224,I38371,I38371);
and I_11069 (I191241,I191224,I38383);
DFFARX1 I_11070 (I191241,I3035,I190913,I191267,);
nor I_11071 (I191275,I191267,I190939);
DFFARX1 I_11072 (I191275,I3035,I190913,I190878,);
DFFARX1 I_11073 (I191267,I3035,I190913,I190896,);
nor I_11074 (I191320,I38392,I38371);
not I_11075 (I191337,I191320);
nor I_11076 (I190899,I191176,I191337);
nand I_11077 (I190884,I191193,I191337);
nor I_11078 (I190893,I190939,I191320);
DFFARX1 I_11079 (I191320,I3035,I190913,I190902,);
not I_11080 (I191440,I3042);
DFFARX1 I_11081 (I97939,I3035,I191440,I191466,);
nand I_11082 (I191474,I97939,I97945);
and I_11083 (I191491,I191474,I97963);
DFFARX1 I_11084 (I191491,I3035,I191440,I191517,);
nor I_11085 (I191408,I191517,I191466);
not I_11086 (I191539,I191517);
DFFARX1 I_11087 (I97951,I3035,I191440,I191565,);
nand I_11088 (I191573,I191565,I97948);
not I_11089 (I191590,I191573);
DFFARX1 I_11090 (I191590,I3035,I191440,I191616,);
not I_11091 (I191432,I191616);
nor I_11092 (I191638,I191466,I191573);
nor I_11093 (I191414,I191517,I191638);
DFFARX1 I_11094 (I97957,I3035,I191440,I191678,);
DFFARX1 I_11095 (I191678,I3035,I191440,I191695,);
not I_11096 (I191703,I191695);
not I_11097 (I191720,I191678);
nand I_11098 (I191417,I191720,I191539);
nand I_11099 (I191751,I97942,I97942);
and I_11100 (I191768,I191751,I97954);
DFFARX1 I_11101 (I191768,I3035,I191440,I191794,);
nor I_11102 (I191802,I191794,I191466);
DFFARX1 I_11103 (I191802,I3035,I191440,I191405,);
DFFARX1 I_11104 (I191794,I3035,I191440,I191423,);
nor I_11105 (I191847,I97960,I97942);
not I_11106 (I191864,I191847);
nor I_11107 (I191426,I191703,I191864);
nand I_11108 (I191411,I191720,I191864);
nor I_11109 (I191420,I191466,I191847);
DFFARX1 I_11110 (I191847,I3035,I191440,I191429,);
not I_11111 (I191967,I3042);
DFFARX1 I_11112 (I47860,I3035,I191967,I191993,);
nand I_11113 (I192001,I47872,I47881);
and I_11114 (I192018,I192001,I47860);
DFFARX1 I_11115 (I192018,I3035,I191967,I192044,);
nor I_11116 (I191935,I192044,I191993);
not I_11117 (I192066,I192044);
DFFARX1 I_11118 (I47875,I3035,I191967,I192092,);
nand I_11119 (I192100,I192092,I47863);
not I_11120 (I192117,I192100);
DFFARX1 I_11121 (I192117,I3035,I191967,I192143,);
not I_11122 (I191959,I192143);
nor I_11123 (I192165,I191993,I192100);
nor I_11124 (I191941,I192044,I192165);
DFFARX1 I_11125 (I47866,I3035,I191967,I192205,);
DFFARX1 I_11126 (I192205,I3035,I191967,I192222,);
not I_11127 (I192230,I192222);
not I_11128 (I192247,I192205);
nand I_11129 (I191944,I192247,I192066);
nand I_11130 (I192278,I47857,I47857);
and I_11131 (I192295,I192278,I47869);
DFFARX1 I_11132 (I192295,I3035,I191967,I192321,);
nor I_11133 (I192329,I192321,I191993);
DFFARX1 I_11134 (I192329,I3035,I191967,I191932,);
DFFARX1 I_11135 (I192321,I3035,I191967,I191950,);
nor I_11136 (I192374,I47878,I47857);
not I_11137 (I192391,I192374);
nor I_11138 (I191953,I192230,I192391);
nand I_11139 (I191938,I192247,I192391);
nor I_11140 (I191947,I191993,I192374);
DFFARX1 I_11141 (I192374,I3035,I191967,I191956,);
not I_11142 (I192494,I3042);
DFFARX1 I_11143 (I444045,I3035,I192494,I192520,);
nand I_11144 (I192528,I444048,I444042);
and I_11145 (I192545,I192528,I444054);
DFFARX1 I_11146 (I192545,I3035,I192494,I192571,);
nor I_11147 (I192462,I192571,I192520);
not I_11148 (I192593,I192571);
DFFARX1 I_11149 (I444057,I3035,I192494,I192619,);
nand I_11150 (I192627,I192619,I444048);
not I_11151 (I192644,I192627);
DFFARX1 I_11152 (I192644,I3035,I192494,I192670,);
not I_11153 (I192486,I192670);
nor I_11154 (I192692,I192520,I192627);
nor I_11155 (I192468,I192571,I192692);
DFFARX1 I_11156 (I444060,I3035,I192494,I192732,);
DFFARX1 I_11157 (I192732,I3035,I192494,I192749,);
not I_11158 (I192757,I192749);
not I_11159 (I192774,I192732);
nand I_11160 (I192471,I192774,I192593);
nand I_11161 (I192805,I444042,I444051);
and I_11162 (I192822,I192805,I444045);
DFFARX1 I_11163 (I192822,I3035,I192494,I192848,);
nor I_11164 (I192856,I192848,I192520);
DFFARX1 I_11165 (I192856,I3035,I192494,I192459,);
DFFARX1 I_11166 (I192848,I3035,I192494,I192477,);
nor I_11167 (I192901,I444063,I444051);
not I_11168 (I192918,I192901);
nor I_11169 (I192480,I192757,I192918);
nand I_11170 (I192465,I192774,I192918);
nor I_11171 (I192474,I192520,I192901);
DFFARX1 I_11172 (I192901,I3035,I192494,I192483,);
not I_11173 (I193021,I3042);
DFFARX1 I_11174 (I746034,I3035,I193021,I193047,);
nand I_11175 (I193055,I746013,I746013);
and I_11176 (I193072,I193055,I746040);
DFFARX1 I_11177 (I193072,I3035,I193021,I193098,);
nor I_11178 (I192989,I193098,I193047);
not I_11179 (I193120,I193098);
DFFARX1 I_11180 (I746028,I3035,I193021,I193146,);
nand I_11181 (I193154,I193146,I746031);
not I_11182 (I193171,I193154);
DFFARX1 I_11183 (I193171,I3035,I193021,I193197,);
not I_11184 (I193013,I193197);
nor I_11185 (I193219,I193047,I193154);
nor I_11186 (I192995,I193098,I193219);
DFFARX1 I_11187 (I746022,I3035,I193021,I193259,);
DFFARX1 I_11188 (I193259,I3035,I193021,I193276,);
not I_11189 (I193284,I193276);
not I_11190 (I193301,I193259);
nand I_11191 (I192998,I193301,I193120);
nand I_11192 (I193332,I746019,I746016);
and I_11193 (I193349,I193332,I746037);
DFFARX1 I_11194 (I193349,I3035,I193021,I193375,);
nor I_11195 (I193383,I193375,I193047);
DFFARX1 I_11196 (I193383,I3035,I193021,I192986,);
DFFARX1 I_11197 (I193375,I3035,I193021,I193004,);
nor I_11198 (I193428,I746025,I746016);
not I_11199 (I193445,I193428);
nor I_11200 (I193007,I193284,I193445);
nand I_11201 (I192992,I193301,I193445);
nor I_11202 (I193001,I193047,I193428);
DFFARX1 I_11203 (I193428,I3035,I193021,I193010,);
not I_11204 (I193548,I3042);
DFFARX1 I_11205 (I380508,I3035,I193548,I193574,);
nand I_11206 (I193582,I380499,I380514);
and I_11207 (I193599,I193582,I380520);
DFFARX1 I_11208 (I193599,I3035,I193548,I193625,);
nor I_11209 (I193516,I193625,I193574);
not I_11210 (I193647,I193625);
DFFARX1 I_11211 (I380505,I3035,I193548,I193673,);
nand I_11212 (I193681,I193673,I380499);
not I_11213 (I193698,I193681);
DFFARX1 I_11214 (I193698,I3035,I193548,I193724,);
not I_11215 (I193540,I193724);
nor I_11216 (I193746,I193574,I193681);
nor I_11217 (I193522,I193625,I193746);
DFFARX1 I_11218 (I380502,I3035,I193548,I193786,);
DFFARX1 I_11219 (I193786,I3035,I193548,I193803,);
not I_11220 (I193811,I193803);
not I_11221 (I193828,I193786);
nand I_11222 (I193525,I193828,I193647);
nand I_11223 (I193859,I380496,I380511);
and I_11224 (I193876,I193859,I380496);
DFFARX1 I_11225 (I193876,I3035,I193548,I193902,);
nor I_11226 (I193910,I193902,I193574);
DFFARX1 I_11227 (I193910,I3035,I193548,I193513,);
DFFARX1 I_11228 (I193902,I3035,I193548,I193531,);
nor I_11229 (I193955,I380517,I380511);
not I_11230 (I193972,I193955);
nor I_11231 (I193534,I193811,I193972);
nand I_11232 (I193519,I193828,I193972);
nor I_11233 (I193528,I193574,I193955);
DFFARX1 I_11234 (I193955,I3035,I193548,I193537,);
not I_11235 (I194075,I3042);
DFFARX1 I_11236 (I303637,I3035,I194075,I194101,);
nand I_11237 (I194109,I303622,I303625);
and I_11238 (I194126,I194109,I303640);
DFFARX1 I_11239 (I194126,I3035,I194075,I194152,);
nor I_11240 (I194043,I194152,I194101);
not I_11241 (I194174,I194152);
DFFARX1 I_11242 (I303634,I3035,I194075,I194200,);
nand I_11243 (I194208,I194200,I303625);
not I_11244 (I194225,I194208);
DFFARX1 I_11245 (I194225,I3035,I194075,I194251,);
not I_11246 (I194067,I194251);
nor I_11247 (I194273,I194101,I194208);
nor I_11248 (I194049,I194152,I194273);
DFFARX1 I_11249 (I303631,I3035,I194075,I194313,);
DFFARX1 I_11250 (I194313,I3035,I194075,I194330,);
not I_11251 (I194338,I194330);
not I_11252 (I194355,I194313);
nand I_11253 (I194052,I194355,I194174);
nand I_11254 (I194386,I303646,I303622);
and I_11255 (I194403,I194386,I303643);
DFFARX1 I_11256 (I194403,I3035,I194075,I194429,);
nor I_11257 (I194437,I194429,I194101);
DFFARX1 I_11258 (I194437,I3035,I194075,I194040,);
DFFARX1 I_11259 (I194429,I3035,I194075,I194058,);
nor I_11260 (I194482,I303628,I303622);
not I_11261 (I194499,I194482);
nor I_11262 (I194061,I194338,I194499);
nand I_11263 (I194046,I194355,I194499);
nor I_11264 (I194055,I194101,I194482);
DFFARX1 I_11265 (I194482,I3035,I194075,I194064,);
not I_11266 (I194602,I3042);
DFFARX1 I_11267 (I593098,I3035,I194602,I194628,);
nand I_11268 (I194636,I593113,I593098);
and I_11269 (I194653,I194636,I593116);
DFFARX1 I_11270 (I194653,I3035,I194602,I194679,);
nor I_11271 (I194570,I194679,I194628);
not I_11272 (I194701,I194679);
DFFARX1 I_11273 (I593122,I3035,I194602,I194727,);
nand I_11274 (I194735,I194727,I593104);
not I_11275 (I194752,I194735);
DFFARX1 I_11276 (I194752,I3035,I194602,I194778,);
not I_11277 (I194594,I194778);
nor I_11278 (I194800,I194628,I194735);
nor I_11279 (I194576,I194679,I194800);
DFFARX1 I_11280 (I593101,I3035,I194602,I194840,);
DFFARX1 I_11281 (I194840,I3035,I194602,I194857,);
not I_11282 (I194865,I194857);
not I_11283 (I194882,I194840);
nand I_11284 (I194579,I194882,I194701);
nand I_11285 (I194913,I593101,I593107);
and I_11286 (I194930,I194913,I593119);
DFFARX1 I_11287 (I194930,I3035,I194602,I194956,);
nor I_11288 (I194964,I194956,I194628);
DFFARX1 I_11289 (I194964,I3035,I194602,I194567,);
DFFARX1 I_11290 (I194956,I3035,I194602,I194585,);
nor I_11291 (I195009,I593110,I593107);
not I_11292 (I195026,I195009);
nor I_11293 (I194588,I194865,I195026);
nand I_11294 (I194573,I194882,I195026);
nor I_11295 (I194582,I194628,I195009);
DFFARX1 I_11296 (I195009,I3035,I194602,I194591,);
not I_11297 (I195129,I3042);
DFFARX1 I_11298 (I252753,I3035,I195129,I195155,);
nand I_11299 (I195163,I252765,I252744);
and I_11300 (I195180,I195163,I252768);
DFFARX1 I_11301 (I195180,I3035,I195129,I195206,);
nor I_11302 (I195097,I195206,I195155);
not I_11303 (I195228,I195206);
DFFARX1 I_11304 (I252759,I3035,I195129,I195254,);
nand I_11305 (I195262,I195254,I252741);
not I_11306 (I195279,I195262);
DFFARX1 I_11307 (I195279,I3035,I195129,I195305,);
not I_11308 (I195121,I195305);
nor I_11309 (I195327,I195155,I195262);
nor I_11310 (I195103,I195206,I195327);
DFFARX1 I_11311 (I252756,I3035,I195129,I195367,);
DFFARX1 I_11312 (I195367,I3035,I195129,I195384,);
not I_11313 (I195392,I195384);
not I_11314 (I195409,I195367);
nand I_11315 (I195106,I195409,I195228);
nand I_11316 (I195440,I252741,I252747);
and I_11317 (I195457,I195440,I252750);
DFFARX1 I_11318 (I195457,I3035,I195129,I195483,);
nor I_11319 (I195491,I195483,I195155);
DFFARX1 I_11320 (I195491,I3035,I195129,I195094,);
DFFARX1 I_11321 (I195483,I3035,I195129,I195112,);
nor I_11322 (I195536,I252762,I252747);
not I_11323 (I195553,I195536);
nor I_11324 (I195115,I195392,I195553);
nand I_11325 (I195100,I195409,I195553);
nor I_11326 (I195109,I195155,I195536);
DFFARX1 I_11327 (I195536,I3035,I195129,I195118,);
not I_11328 (I195656,I3042);
DFFARX1 I_11329 (I442464,I3035,I195656,I195682,);
nand I_11330 (I195690,I442467,I442461);
and I_11331 (I195707,I195690,I442473);
DFFARX1 I_11332 (I195707,I3035,I195656,I195733,);
nor I_11333 (I195624,I195733,I195682);
not I_11334 (I195755,I195733);
DFFARX1 I_11335 (I442476,I3035,I195656,I195781,);
nand I_11336 (I195789,I195781,I442467);
not I_11337 (I195806,I195789);
DFFARX1 I_11338 (I195806,I3035,I195656,I195832,);
not I_11339 (I195648,I195832);
nor I_11340 (I195854,I195682,I195789);
nor I_11341 (I195630,I195733,I195854);
DFFARX1 I_11342 (I442479,I3035,I195656,I195894,);
DFFARX1 I_11343 (I195894,I3035,I195656,I195911,);
not I_11344 (I195919,I195911);
not I_11345 (I195936,I195894);
nand I_11346 (I195633,I195936,I195755);
nand I_11347 (I195967,I442461,I442470);
and I_11348 (I195984,I195967,I442464);
DFFARX1 I_11349 (I195984,I3035,I195656,I196010,);
nor I_11350 (I196018,I196010,I195682);
DFFARX1 I_11351 (I196018,I3035,I195656,I195621,);
DFFARX1 I_11352 (I196010,I3035,I195656,I195639,);
nor I_11353 (I196063,I442482,I442470);
not I_11354 (I196080,I196063);
nor I_11355 (I195642,I195919,I196080);
nand I_11356 (I195627,I195936,I196080);
nor I_11357 (I195636,I195682,I196063);
DFFARX1 I_11358 (I196063,I3035,I195656,I195645,);
not I_11359 (I196183,I3042);
DFFARX1 I_11360 (I575758,I3035,I196183,I196209,);
nand I_11361 (I196217,I575773,I575758);
and I_11362 (I196234,I196217,I575776);
DFFARX1 I_11363 (I196234,I3035,I196183,I196260,);
nor I_11364 (I196151,I196260,I196209);
not I_11365 (I196282,I196260);
DFFARX1 I_11366 (I575782,I3035,I196183,I196308,);
nand I_11367 (I196316,I196308,I575764);
not I_11368 (I196333,I196316);
DFFARX1 I_11369 (I196333,I3035,I196183,I196359,);
not I_11370 (I196175,I196359);
nor I_11371 (I196381,I196209,I196316);
nor I_11372 (I196157,I196260,I196381);
DFFARX1 I_11373 (I575761,I3035,I196183,I196421,);
DFFARX1 I_11374 (I196421,I3035,I196183,I196438,);
not I_11375 (I196446,I196438);
not I_11376 (I196463,I196421);
nand I_11377 (I196160,I196463,I196282);
nand I_11378 (I196494,I575761,I575767);
and I_11379 (I196511,I196494,I575779);
DFFARX1 I_11380 (I196511,I3035,I196183,I196537,);
nor I_11381 (I196545,I196537,I196209);
DFFARX1 I_11382 (I196545,I3035,I196183,I196148,);
DFFARX1 I_11383 (I196537,I3035,I196183,I196166,);
nor I_11384 (I196590,I575770,I575767);
not I_11385 (I196607,I196590);
nor I_11386 (I196169,I196446,I196607);
nand I_11387 (I196154,I196463,I196607);
nor I_11388 (I196163,I196209,I196590);
DFFARX1 I_11389 (I196590,I3035,I196183,I196172,);
not I_11390 (I196710,I3042);
DFFARX1 I_11391 (I579226,I3035,I196710,I196736,);
nand I_11392 (I196744,I579241,I579226);
and I_11393 (I196761,I196744,I579244);
DFFARX1 I_11394 (I196761,I3035,I196710,I196787,);
nor I_11395 (I196678,I196787,I196736);
not I_11396 (I196809,I196787);
DFFARX1 I_11397 (I579250,I3035,I196710,I196835,);
nand I_11398 (I196843,I196835,I579232);
not I_11399 (I196860,I196843);
DFFARX1 I_11400 (I196860,I3035,I196710,I196886,);
not I_11401 (I196702,I196886);
nor I_11402 (I196908,I196736,I196843);
nor I_11403 (I196684,I196787,I196908);
DFFARX1 I_11404 (I579229,I3035,I196710,I196948,);
DFFARX1 I_11405 (I196948,I3035,I196710,I196965,);
not I_11406 (I196973,I196965);
not I_11407 (I196990,I196948);
nand I_11408 (I196687,I196990,I196809);
nand I_11409 (I197021,I579229,I579235);
and I_11410 (I197038,I197021,I579247);
DFFARX1 I_11411 (I197038,I3035,I196710,I197064,);
nor I_11412 (I197072,I197064,I196736);
DFFARX1 I_11413 (I197072,I3035,I196710,I196675,);
DFFARX1 I_11414 (I197064,I3035,I196710,I196693,);
nor I_11415 (I197117,I579238,I579235);
not I_11416 (I197134,I197117);
nor I_11417 (I196696,I196973,I197134);
nand I_11418 (I196681,I196990,I197134);
nor I_11419 (I196690,I196736,I197117);
DFFARX1 I_11420 (I197117,I3035,I196710,I196699,);
not I_11421 (I197237,I3042);
DFFARX1 I_11422 (I348140,I3035,I197237,I197263,);
nand I_11423 (I197271,I348131,I348146);
and I_11424 (I197288,I197271,I348152);
DFFARX1 I_11425 (I197288,I3035,I197237,I197314,);
nor I_11426 (I197205,I197314,I197263);
not I_11427 (I197336,I197314);
DFFARX1 I_11428 (I348137,I3035,I197237,I197362,);
nand I_11429 (I197370,I197362,I348131);
not I_11430 (I197387,I197370);
DFFARX1 I_11431 (I197387,I3035,I197237,I197413,);
not I_11432 (I197229,I197413);
nor I_11433 (I197435,I197263,I197370);
nor I_11434 (I197211,I197314,I197435);
DFFARX1 I_11435 (I348134,I3035,I197237,I197475,);
DFFARX1 I_11436 (I197475,I3035,I197237,I197492,);
not I_11437 (I197500,I197492);
not I_11438 (I197517,I197475);
nand I_11439 (I197214,I197517,I197336);
nand I_11440 (I197548,I348128,I348143);
and I_11441 (I197565,I197548,I348128);
DFFARX1 I_11442 (I197565,I3035,I197237,I197591,);
nor I_11443 (I197599,I197591,I197263);
DFFARX1 I_11444 (I197599,I3035,I197237,I197202,);
DFFARX1 I_11445 (I197591,I3035,I197237,I197220,);
nor I_11446 (I197644,I348149,I348143);
not I_11447 (I197661,I197644);
nor I_11448 (I197223,I197500,I197661);
nand I_11449 (I197208,I197517,I197661);
nor I_11450 (I197217,I197263,I197644);
DFFARX1 I_11451 (I197644,I3035,I197237,I197226,);
not I_11452 (I197764,I3042);
DFFARX1 I_11453 (I505789,I3035,I197764,I197790,);
nand I_11454 (I197798,I505786,I505804);
and I_11455 (I197815,I197798,I505795);
DFFARX1 I_11456 (I197815,I3035,I197764,I197841,);
nor I_11457 (I197732,I197841,I197790);
not I_11458 (I197863,I197841);
DFFARX1 I_11459 (I505810,I3035,I197764,I197889,);
nand I_11460 (I197897,I197889,I505792);
not I_11461 (I197914,I197897);
DFFARX1 I_11462 (I197914,I3035,I197764,I197940,);
not I_11463 (I197756,I197940);
nor I_11464 (I197962,I197790,I197897);
nor I_11465 (I197738,I197841,I197962);
DFFARX1 I_11466 (I505798,I3035,I197764,I198002,);
DFFARX1 I_11467 (I198002,I3035,I197764,I198019,);
not I_11468 (I198027,I198019);
not I_11469 (I198044,I198002);
nand I_11470 (I197741,I198044,I197863);
nand I_11471 (I198075,I505786,I505813);
and I_11472 (I198092,I198075,I505801);
DFFARX1 I_11473 (I198092,I3035,I197764,I198118,);
nor I_11474 (I198126,I198118,I197790);
DFFARX1 I_11475 (I198126,I3035,I197764,I197729,);
DFFARX1 I_11476 (I198118,I3035,I197764,I197747,);
nor I_11477 (I198171,I505807,I505813);
not I_11478 (I198188,I198171);
nor I_11479 (I197750,I198027,I198188);
nand I_11480 (I197735,I198044,I198188);
nor I_11481 (I197744,I197790,I198171);
DFFARX1 I_11482 (I198171,I3035,I197764,I197753,);
not I_11483 (I198291,I3042);
DFFARX1 I_11484 (I657240,I3035,I198291,I198317,);
nand I_11485 (I198325,I657222,I657246);
and I_11486 (I198342,I198325,I657237);
DFFARX1 I_11487 (I198342,I3035,I198291,I198368,);
nor I_11488 (I198259,I198368,I198317);
not I_11489 (I198390,I198368);
DFFARX1 I_11490 (I657243,I3035,I198291,I198416,);
nand I_11491 (I198424,I198416,I657231);
not I_11492 (I198441,I198424);
DFFARX1 I_11493 (I198441,I3035,I198291,I198467,);
not I_11494 (I198283,I198467);
nor I_11495 (I198489,I198317,I198424);
nor I_11496 (I198265,I198368,I198489);
DFFARX1 I_11497 (I657222,I3035,I198291,I198529,);
DFFARX1 I_11498 (I198529,I3035,I198291,I198546,);
not I_11499 (I198554,I198546);
not I_11500 (I198571,I198529);
nand I_11501 (I198268,I198571,I198390);
nand I_11502 (I198602,I657228,I657225);
and I_11503 (I198619,I198602,I657234);
DFFARX1 I_11504 (I198619,I3035,I198291,I198645,);
nor I_11505 (I198653,I198645,I198317);
DFFARX1 I_11506 (I198653,I3035,I198291,I198256,);
DFFARX1 I_11507 (I198645,I3035,I198291,I198274,);
nor I_11508 (I198698,I657225,I657225);
not I_11509 (I198715,I198698);
nor I_11510 (I198277,I198554,I198715);
nand I_11511 (I198262,I198571,I198715);
nor I_11512 (I198271,I198317,I198698);
DFFARX1 I_11513 (I198698,I3035,I198291,I198280,);
not I_11514 (I198818,I3042);
DFFARX1 I_11515 (I604080,I3035,I198818,I198844,);
nand I_11516 (I198852,I604095,I604080);
and I_11517 (I198869,I198852,I604098);
DFFARX1 I_11518 (I198869,I3035,I198818,I198895,);
nor I_11519 (I198786,I198895,I198844);
not I_11520 (I198917,I198895);
DFFARX1 I_11521 (I604104,I3035,I198818,I198943,);
nand I_11522 (I198951,I198943,I604086);
not I_11523 (I198968,I198951);
DFFARX1 I_11524 (I198968,I3035,I198818,I198994,);
not I_11525 (I198810,I198994);
nor I_11526 (I199016,I198844,I198951);
nor I_11527 (I198792,I198895,I199016);
DFFARX1 I_11528 (I604083,I3035,I198818,I199056,);
DFFARX1 I_11529 (I199056,I3035,I198818,I199073,);
not I_11530 (I199081,I199073);
not I_11531 (I199098,I199056);
nand I_11532 (I198795,I199098,I198917);
nand I_11533 (I199129,I604083,I604089);
and I_11534 (I199146,I199129,I604101);
DFFARX1 I_11535 (I199146,I3035,I198818,I199172,);
nor I_11536 (I199180,I199172,I198844);
DFFARX1 I_11537 (I199180,I3035,I198818,I198783,);
DFFARX1 I_11538 (I199172,I3035,I198818,I198801,);
nor I_11539 (I199225,I604092,I604089);
not I_11540 (I199242,I199225);
nor I_11541 (I198804,I199081,I199242);
nand I_11542 (I198789,I199098,I199242);
nor I_11543 (I198798,I198844,I199225);
DFFARX1 I_11544 (I199225,I3035,I198818,I198807,);
not I_11545 (I199345,I3042);
DFFARX1 I_11546 (I1500,I3035,I199345,I199371,);
nand I_11547 (I199379,I3004,I1396);
and I_11548 (I199396,I199379,I2516);
DFFARX1 I_11549 (I199396,I3035,I199345,I199422,);
nor I_11550 (I199313,I199422,I199371);
not I_11551 (I199444,I199422);
DFFARX1 I_11552 (I2468,I3035,I199345,I199470,);
nand I_11553 (I199478,I199470,I2556);
not I_11554 (I199495,I199478);
DFFARX1 I_11555 (I199495,I3035,I199345,I199521,);
not I_11556 (I199337,I199521);
nor I_11557 (I199543,I199371,I199478);
nor I_11558 (I199319,I199422,I199543);
DFFARX1 I_11559 (I2892,I3035,I199345,I199583,);
DFFARX1 I_11560 (I199583,I3035,I199345,I199600,);
not I_11561 (I199608,I199600);
not I_11562 (I199625,I199583);
nand I_11563 (I199322,I199625,I199444);
nand I_11564 (I199656,I2100,I2924);
and I_11565 (I199673,I199656,I2844);
DFFARX1 I_11566 (I199673,I3035,I199345,I199699,);
nor I_11567 (I199707,I199699,I199371);
DFFARX1 I_11568 (I199707,I3035,I199345,I199310,);
DFFARX1 I_11569 (I199699,I3035,I199345,I199328,);
nor I_11570 (I199752,I1588,I2924);
not I_11571 (I199769,I199752);
nor I_11572 (I199331,I199608,I199769);
nand I_11573 (I199316,I199625,I199769);
nor I_11574 (I199325,I199371,I199752);
DFFARX1 I_11575 (I199752,I3035,I199345,I199334,);
not I_11576 (I199872,I3042);
DFFARX1 I_11577 (I541965,I3035,I199872,I199898,);
nand I_11578 (I199906,I541962,I541980);
and I_11579 (I199923,I199906,I541971);
DFFARX1 I_11580 (I199923,I3035,I199872,I199949,);
nor I_11581 (I199840,I199949,I199898);
not I_11582 (I199971,I199949);
DFFARX1 I_11583 (I541986,I3035,I199872,I199997,);
nand I_11584 (I200005,I199997,I541968);
not I_11585 (I200022,I200005);
DFFARX1 I_11586 (I200022,I3035,I199872,I200048,);
not I_11587 (I199864,I200048);
nor I_11588 (I200070,I199898,I200005);
nor I_11589 (I199846,I199949,I200070);
DFFARX1 I_11590 (I541974,I3035,I199872,I200110,);
DFFARX1 I_11591 (I200110,I3035,I199872,I200127,);
not I_11592 (I200135,I200127);
not I_11593 (I200152,I200110);
nand I_11594 (I199849,I200152,I199971);
nand I_11595 (I200183,I541962,I541989);
and I_11596 (I200200,I200183,I541977);
DFFARX1 I_11597 (I200200,I3035,I199872,I200226,);
nor I_11598 (I200234,I200226,I199898);
DFFARX1 I_11599 (I200234,I3035,I199872,I199837,);
DFFARX1 I_11600 (I200226,I3035,I199872,I199855,);
nor I_11601 (I200279,I541983,I541989);
not I_11602 (I200296,I200279);
nor I_11603 (I199858,I200135,I200296);
nand I_11604 (I199843,I200152,I200296);
nor I_11605 (I199852,I199898,I200279);
DFFARX1 I_11606 (I200279,I3035,I199872,I199861,);
not I_11607 (I200399,I3042);
DFFARX1 I_11608 (I149109,I3035,I200399,I200425,);
nand I_11609 (I200433,I149109,I149115);
and I_11610 (I200450,I200433,I149133);
DFFARX1 I_11611 (I200450,I3035,I200399,I200476,);
nor I_11612 (I200367,I200476,I200425);
not I_11613 (I200498,I200476);
DFFARX1 I_11614 (I149121,I3035,I200399,I200524,);
nand I_11615 (I200532,I200524,I149118);
not I_11616 (I200549,I200532);
DFFARX1 I_11617 (I200549,I3035,I200399,I200575,);
not I_11618 (I200391,I200575);
nor I_11619 (I200597,I200425,I200532);
nor I_11620 (I200373,I200476,I200597);
DFFARX1 I_11621 (I149127,I3035,I200399,I200637,);
DFFARX1 I_11622 (I200637,I3035,I200399,I200654,);
not I_11623 (I200662,I200654);
not I_11624 (I200679,I200637);
nand I_11625 (I200376,I200679,I200498);
nand I_11626 (I200710,I149112,I149112);
and I_11627 (I200727,I200710,I149124);
DFFARX1 I_11628 (I200727,I3035,I200399,I200753,);
nor I_11629 (I200761,I200753,I200425);
DFFARX1 I_11630 (I200761,I3035,I200399,I200364,);
DFFARX1 I_11631 (I200753,I3035,I200399,I200382,);
nor I_11632 (I200806,I149130,I149112);
not I_11633 (I200823,I200806);
nor I_11634 (I200385,I200662,I200823);
nand I_11635 (I200370,I200679,I200823);
nor I_11636 (I200379,I200425,I200806);
DFFARX1 I_11637 (I200806,I3035,I200399,I200388,);
not I_11638 (I200926,I3042);
DFFARX1 I_11639 (I8859,I3035,I200926,I200952,);
nand I_11640 (I200960,I8883,I8862);
and I_11641 (I200977,I200960,I8859);
DFFARX1 I_11642 (I200977,I3035,I200926,I201003,);
nor I_11643 (I200894,I201003,I200952);
not I_11644 (I201025,I201003);
DFFARX1 I_11645 (I8865,I3035,I200926,I201051,);
nand I_11646 (I201059,I201051,I8874);
not I_11647 (I201076,I201059);
DFFARX1 I_11648 (I201076,I3035,I200926,I201102,);
not I_11649 (I200918,I201102);
nor I_11650 (I201124,I200952,I201059);
nor I_11651 (I200900,I201003,I201124);
DFFARX1 I_11652 (I8868,I3035,I200926,I201164,);
DFFARX1 I_11653 (I201164,I3035,I200926,I201181,);
not I_11654 (I201189,I201181);
not I_11655 (I201206,I201164);
nand I_11656 (I200903,I201206,I201025);
nand I_11657 (I201237,I8880,I8862);
and I_11658 (I201254,I201237,I8871);
DFFARX1 I_11659 (I201254,I3035,I200926,I201280,);
nor I_11660 (I201288,I201280,I200952);
DFFARX1 I_11661 (I201288,I3035,I200926,I200891,);
DFFARX1 I_11662 (I201280,I3035,I200926,I200909,);
nor I_11663 (I201333,I8877,I8862);
not I_11664 (I201350,I201333);
nor I_11665 (I200912,I201189,I201350);
nand I_11666 (I200897,I201206,I201350);
nor I_11667 (I200906,I200952,I201333);
DFFARX1 I_11668 (I201333,I3035,I200926,I200915,);
not I_11669 (I201453,I3042);
DFFARX1 I_11670 (I258737,I3035,I201453,I201479,);
nand I_11671 (I201487,I258749,I258728);
and I_11672 (I201504,I201487,I258752);
DFFARX1 I_11673 (I201504,I3035,I201453,I201530,);
nor I_11674 (I201421,I201530,I201479);
not I_11675 (I201552,I201530);
DFFARX1 I_11676 (I258743,I3035,I201453,I201578,);
nand I_11677 (I201586,I201578,I258725);
not I_11678 (I201603,I201586);
DFFARX1 I_11679 (I201603,I3035,I201453,I201629,);
not I_11680 (I201445,I201629);
nor I_11681 (I201651,I201479,I201586);
nor I_11682 (I201427,I201530,I201651);
DFFARX1 I_11683 (I258740,I3035,I201453,I201691,);
DFFARX1 I_11684 (I201691,I3035,I201453,I201708,);
not I_11685 (I201716,I201708);
not I_11686 (I201733,I201691);
nand I_11687 (I201430,I201733,I201552);
nand I_11688 (I201764,I258725,I258731);
and I_11689 (I201781,I201764,I258734);
DFFARX1 I_11690 (I201781,I3035,I201453,I201807,);
nor I_11691 (I201815,I201807,I201479);
DFFARX1 I_11692 (I201815,I3035,I201453,I201418,);
DFFARX1 I_11693 (I201807,I3035,I201453,I201436,);
nor I_11694 (I201860,I258746,I258731);
not I_11695 (I201877,I201860);
nor I_11696 (I201439,I201716,I201877);
nand I_11697 (I201424,I201733,I201877);
nor I_11698 (I201433,I201479,I201860);
DFFARX1 I_11699 (I201860,I3035,I201453,I201442,);
not I_11700 (I201980,I3042);
DFFARX1 I_11701 (I279944,I3035,I201980,I202006,);
nand I_11702 (I202014,I279944,I279956);
and I_11703 (I202031,I202014,I279941);
DFFARX1 I_11704 (I202031,I3035,I201980,I202057,);
nor I_11705 (I201948,I202057,I202006);
not I_11706 (I202079,I202057);
DFFARX1 I_11707 (I279965,I3035,I201980,I202105,);
nand I_11708 (I202113,I202105,I279962);
not I_11709 (I202130,I202113);
DFFARX1 I_11710 (I202130,I3035,I201980,I202156,);
not I_11711 (I201972,I202156);
nor I_11712 (I202178,I202006,I202113);
nor I_11713 (I201954,I202057,I202178);
DFFARX1 I_11714 (I279953,I3035,I201980,I202218,);
DFFARX1 I_11715 (I202218,I3035,I201980,I202235,);
not I_11716 (I202243,I202235);
not I_11717 (I202260,I202218);
nand I_11718 (I201957,I202260,I202079);
nand I_11719 (I202291,I279941,I279950);
and I_11720 (I202308,I202291,I279959);
DFFARX1 I_11721 (I202308,I3035,I201980,I202334,);
nor I_11722 (I202342,I202334,I202006);
DFFARX1 I_11723 (I202342,I3035,I201980,I201945,);
DFFARX1 I_11724 (I202334,I3035,I201980,I201963,);
nor I_11725 (I202387,I279947,I279950);
not I_11726 (I202404,I202387);
nor I_11727 (I201966,I202243,I202404);
nand I_11728 (I201951,I202260,I202404);
nor I_11729 (I201960,I202006,I202387);
DFFARX1 I_11730 (I202387,I3035,I201980,I201969,);
not I_11731 (I202507,I3042);
DFFARX1 I_11732 (I499329,I3035,I202507,I202533,);
nand I_11733 (I202541,I499326,I499344);
and I_11734 (I202558,I202541,I499335);
DFFARX1 I_11735 (I202558,I3035,I202507,I202584,);
nor I_11736 (I202475,I202584,I202533);
not I_11737 (I202606,I202584);
DFFARX1 I_11738 (I499350,I3035,I202507,I202632,);
nand I_11739 (I202640,I202632,I499332);
not I_11740 (I202657,I202640);
DFFARX1 I_11741 (I202657,I3035,I202507,I202683,);
not I_11742 (I202499,I202683);
nor I_11743 (I202705,I202533,I202640);
nor I_11744 (I202481,I202584,I202705);
DFFARX1 I_11745 (I499338,I3035,I202507,I202745,);
DFFARX1 I_11746 (I202745,I3035,I202507,I202762,);
not I_11747 (I202770,I202762);
not I_11748 (I202787,I202745);
nand I_11749 (I202484,I202787,I202606);
nand I_11750 (I202818,I499326,I499353);
and I_11751 (I202835,I202818,I499341);
DFFARX1 I_11752 (I202835,I3035,I202507,I202861,);
nor I_11753 (I202869,I202861,I202533);
DFFARX1 I_11754 (I202869,I3035,I202507,I202472,);
DFFARX1 I_11755 (I202861,I3035,I202507,I202490,);
nor I_11756 (I202914,I499347,I499353);
not I_11757 (I202931,I202914);
nor I_11758 (I202493,I202770,I202931);
nand I_11759 (I202478,I202787,I202931);
nor I_11760 (I202487,I202533,I202914);
DFFARX1 I_11761 (I202914,I3035,I202507,I202496,);
not I_11762 (I203034,I3042);
DFFARX1 I_11763 (I423492,I3035,I203034,I203060,);
nand I_11764 (I203068,I423495,I423489);
and I_11765 (I203085,I203068,I423501);
DFFARX1 I_11766 (I203085,I3035,I203034,I203111,);
nor I_11767 (I203002,I203111,I203060);
not I_11768 (I203133,I203111);
DFFARX1 I_11769 (I423504,I3035,I203034,I203159,);
nand I_11770 (I203167,I203159,I423495);
not I_11771 (I203184,I203167);
DFFARX1 I_11772 (I203184,I3035,I203034,I203210,);
not I_11773 (I203026,I203210);
nor I_11774 (I203232,I203060,I203167);
nor I_11775 (I203008,I203111,I203232);
DFFARX1 I_11776 (I423507,I3035,I203034,I203272,);
DFFARX1 I_11777 (I203272,I3035,I203034,I203289,);
not I_11778 (I203297,I203289);
not I_11779 (I203314,I203272);
nand I_11780 (I203011,I203314,I203133);
nand I_11781 (I203345,I423489,I423498);
and I_11782 (I203362,I203345,I423492);
DFFARX1 I_11783 (I203362,I3035,I203034,I203388,);
nor I_11784 (I203396,I203388,I203060);
DFFARX1 I_11785 (I203396,I3035,I203034,I202999,);
DFFARX1 I_11786 (I203388,I3035,I203034,I203017,);
nor I_11787 (I203441,I423510,I423498);
not I_11788 (I203458,I203441);
nor I_11789 (I203020,I203297,I203458);
nand I_11790 (I203005,I203314,I203458);
nor I_11791 (I203014,I203060,I203441);
DFFARX1 I_11792 (I203441,I3035,I203034,I203023,);
not I_11793 (I203561,I3042);
DFFARX1 I_11794 (I485763,I3035,I203561,I203587,);
nand I_11795 (I203595,I485760,I485778);
and I_11796 (I203612,I203595,I485769);
DFFARX1 I_11797 (I203612,I3035,I203561,I203638,);
nor I_11798 (I203529,I203638,I203587);
not I_11799 (I203660,I203638);
DFFARX1 I_11800 (I485784,I3035,I203561,I203686,);
nand I_11801 (I203694,I203686,I485766);
not I_11802 (I203711,I203694);
DFFARX1 I_11803 (I203711,I3035,I203561,I203737,);
not I_11804 (I203553,I203737);
nor I_11805 (I203759,I203587,I203694);
nor I_11806 (I203535,I203638,I203759);
DFFARX1 I_11807 (I485772,I3035,I203561,I203799,);
DFFARX1 I_11808 (I203799,I3035,I203561,I203816,);
not I_11809 (I203824,I203816);
not I_11810 (I203841,I203799);
nand I_11811 (I203538,I203841,I203660);
nand I_11812 (I203872,I485760,I485787);
and I_11813 (I203889,I203872,I485775);
DFFARX1 I_11814 (I203889,I3035,I203561,I203915,);
nor I_11815 (I203923,I203915,I203587);
DFFARX1 I_11816 (I203923,I3035,I203561,I203526,);
DFFARX1 I_11817 (I203915,I3035,I203561,I203544,);
nor I_11818 (I203968,I485781,I485787);
not I_11819 (I203985,I203968);
nor I_11820 (I203547,I203824,I203985);
nand I_11821 (I203532,I203841,I203985);
nor I_11822 (I203541,I203587,I203968);
DFFARX1 I_11823 (I203968,I3035,I203561,I203550,);
not I_11824 (I204088,I3042);
DFFARX1 I_11825 (I318087,I3035,I204088,I204114,);
nand I_11826 (I204122,I318072,I318075);
and I_11827 (I204139,I204122,I318090);
DFFARX1 I_11828 (I204139,I3035,I204088,I204165,);
nor I_11829 (I204056,I204165,I204114);
not I_11830 (I204187,I204165);
DFFARX1 I_11831 (I318084,I3035,I204088,I204213,);
nand I_11832 (I204221,I204213,I318075);
not I_11833 (I204238,I204221);
DFFARX1 I_11834 (I204238,I3035,I204088,I204264,);
not I_11835 (I204080,I204264);
nor I_11836 (I204286,I204114,I204221);
nor I_11837 (I204062,I204165,I204286);
DFFARX1 I_11838 (I318081,I3035,I204088,I204326,);
DFFARX1 I_11839 (I204326,I3035,I204088,I204343,);
not I_11840 (I204351,I204343);
not I_11841 (I204368,I204326);
nand I_11842 (I204065,I204368,I204187);
nand I_11843 (I204399,I318096,I318072);
and I_11844 (I204416,I204399,I318093);
DFFARX1 I_11845 (I204416,I3035,I204088,I204442,);
nor I_11846 (I204450,I204442,I204114);
DFFARX1 I_11847 (I204450,I3035,I204088,I204053,);
DFFARX1 I_11848 (I204442,I3035,I204088,I204071,);
nor I_11849 (I204495,I318078,I318072);
not I_11850 (I204512,I204495);
nor I_11851 (I204074,I204351,I204512);
nand I_11852 (I204059,I204368,I204512);
nor I_11853 (I204068,I204114,I204495);
DFFARX1 I_11854 (I204495,I3035,I204088,I204077,);
not I_11855 (I204615,I3042);
DFFARX1 I_11856 (I605814,I3035,I204615,I204641,);
nand I_11857 (I204649,I605829,I605814);
and I_11858 (I204666,I204649,I605832);
DFFARX1 I_11859 (I204666,I3035,I204615,I204692,);
nor I_11860 (I204583,I204692,I204641);
not I_11861 (I204714,I204692);
DFFARX1 I_11862 (I605838,I3035,I204615,I204740,);
nand I_11863 (I204748,I204740,I605820);
not I_11864 (I204765,I204748);
DFFARX1 I_11865 (I204765,I3035,I204615,I204791,);
not I_11866 (I204607,I204791);
nor I_11867 (I204813,I204641,I204748);
nor I_11868 (I204589,I204692,I204813);
DFFARX1 I_11869 (I605817,I3035,I204615,I204853,);
DFFARX1 I_11870 (I204853,I3035,I204615,I204870,);
not I_11871 (I204878,I204870);
not I_11872 (I204895,I204853);
nand I_11873 (I204592,I204895,I204714);
nand I_11874 (I204926,I605817,I605823);
and I_11875 (I204943,I204926,I605835);
DFFARX1 I_11876 (I204943,I3035,I204615,I204969,);
nor I_11877 (I204977,I204969,I204641);
DFFARX1 I_11878 (I204977,I3035,I204615,I204580,);
DFFARX1 I_11879 (I204969,I3035,I204615,I204598,);
nor I_11880 (I205022,I605826,I605823);
not I_11881 (I205039,I205022);
nor I_11882 (I204601,I204878,I205039);
nand I_11883 (I204586,I204895,I205039);
nor I_11884 (I204595,I204641,I205022);
DFFARX1 I_11885 (I205022,I3035,I204615,I204604,);
not I_11886 (I205142,I3042);
DFFARX1 I_11887 (I232625,I3035,I205142,I205168,);
nand I_11888 (I205176,I232637,I232616);
and I_11889 (I205193,I205176,I232640);
DFFARX1 I_11890 (I205193,I3035,I205142,I205219,);
nor I_11891 (I205110,I205219,I205168);
not I_11892 (I205241,I205219);
DFFARX1 I_11893 (I232631,I3035,I205142,I205267,);
nand I_11894 (I205275,I205267,I232613);
not I_11895 (I205292,I205275);
DFFARX1 I_11896 (I205292,I3035,I205142,I205318,);
not I_11897 (I205134,I205318);
nor I_11898 (I205340,I205168,I205275);
nor I_11899 (I205116,I205219,I205340);
DFFARX1 I_11900 (I232628,I3035,I205142,I205380,);
DFFARX1 I_11901 (I205380,I3035,I205142,I205397,);
not I_11902 (I205405,I205397);
not I_11903 (I205422,I205380);
nand I_11904 (I205119,I205422,I205241);
nand I_11905 (I205453,I232613,I232619);
and I_11906 (I205470,I205453,I232622);
DFFARX1 I_11907 (I205470,I3035,I205142,I205496,);
nor I_11908 (I205504,I205496,I205168);
DFFARX1 I_11909 (I205504,I3035,I205142,I205107,);
DFFARX1 I_11910 (I205496,I3035,I205142,I205125,);
nor I_11911 (I205549,I232634,I232619);
not I_11912 (I205566,I205549);
nor I_11913 (I205128,I205405,I205566);
nand I_11914 (I205113,I205422,I205566);
nor I_11915 (I205122,I205168,I205549);
DFFARX1 I_11916 (I205549,I3035,I205142,I205131,);
not I_11917 (I205669,I3042);
DFFARX1 I_11918 (I124714,I3035,I205669,I205695,);
nand I_11919 (I205703,I124714,I124720);
and I_11920 (I205720,I205703,I124738);
DFFARX1 I_11921 (I205720,I3035,I205669,I205746,);
nor I_11922 (I205637,I205746,I205695);
not I_11923 (I205768,I205746);
DFFARX1 I_11924 (I124726,I3035,I205669,I205794,);
nand I_11925 (I205802,I205794,I124723);
not I_11926 (I205819,I205802);
DFFARX1 I_11927 (I205819,I3035,I205669,I205845,);
not I_11928 (I205661,I205845);
nor I_11929 (I205867,I205695,I205802);
nor I_11930 (I205643,I205746,I205867);
DFFARX1 I_11931 (I124732,I3035,I205669,I205907,);
DFFARX1 I_11932 (I205907,I3035,I205669,I205924,);
not I_11933 (I205932,I205924);
not I_11934 (I205949,I205907);
nand I_11935 (I205646,I205949,I205768);
nand I_11936 (I205980,I124717,I124717);
and I_11937 (I205997,I205980,I124729);
DFFARX1 I_11938 (I205997,I3035,I205669,I206023,);
nor I_11939 (I206031,I206023,I205695);
DFFARX1 I_11940 (I206031,I3035,I205669,I205634,);
DFFARX1 I_11941 (I206023,I3035,I205669,I205652,);
nor I_11942 (I206076,I124735,I124717);
not I_11943 (I206093,I206076);
nor I_11944 (I205655,I205932,I206093);
nand I_11945 (I205640,I205949,I206093);
nor I_11946 (I205649,I205695,I206076);
DFFARX1 I_11947 (I206076,I3035,I205669,I205658,);
not I_11948 (I206196,I3042);
DFFARX1 I_11949 (I573446,I3035,I206196,I206222,);
nand I_11950 (I206230,I573461,I573446);
and I_11951 (I206247,I206230,I573464);
DFFARX1 I_11952 (I206247,I3035,I206196,I206273,);
nor I_11953 (I206164,I206273,I206222);
not I_11954 (I206295,I206273);
DFFARX1 I_11955 (I573470,I3035,I206196,I206321,);
nand I_11956 (I206329,I206321,I573452);
not I_11957 (I206346,I206329);
DFFARX1 I_11958 (I206346,I3035,I206196,I206372,);
not I_11959 (I206188,I206372);
nor I_11960 (I206394,I206222,I206329);
nor I_11961 (I206170,I206273,I206394);
DFFARX1 I_11962 (I573449,I3035,I206196,I206434,);
DFFARX1 I_11963 (I206434,I3035,I206196,I206451,);
not I_11964 (I206459,I206451);
not I_11965 (I206476,I206434);
nand I_11966 (I206173,I206476,I206295);
nand I_11967 (I206507,I573449,I573455);
and I_11968 (I206524,I206507,I573467);
DFFARX1 I_11969 (I206524,I3035,I206196,I206550,);
nor I_11970 (I206558,I206550,I206222);
DFFARX1 I_11971 (I206558,I3035,I206196,I206161,);
DFFARX1 I_11972 (I206550,I3035,I206196,I206179,);
nor I_11973 (I206603,I573458,I573455);
not I_11974 (I206620,I206603);
nor I_11975 (I206182,I206459,I206620);
nand I_11976 (I206167,I206476,I206620);
nor I_11977 (I206176,I206222,I206603);
DFFARX1 I_11978 (I206603,I3035,I206196,I206185,);
not I_11979 (I206723,I3042);
DFFARX1 I_11980 (I438775,I3035,I206723,I206749,);
nand I_11981 (I206757,I438778,I438772);
and I_11982 (I206774,I206757,I438784);
DFFARX1 I_11983 (I206774,I3035,I206723,I206800,);
nor I_11984 (I206691,I206800,I206749);
not I_11985 (I206822,I206800);
DFFARX1 I_11986 (I438787,I3035,I206723,I206848,);
nand I_11987 (I206856,I206848,I438778);
not I_11988 (I206873,I206856);
DFFARX1 I_11989 (I206873,I3035,I206723,I206899,);
not I_11990 (I206715,I206899);
nor I_11991 (I206921,I206749,I206856);
nor I_11992 (I206697,I206800,I206921);
DFFARX1 I_11993 (I438790,I3035,I206723,I206961,);
DFFARX1 I_11994 (I206961,I3035,I206723,I206978,);
not I_11995 (I206986,I206978);
not I_11996 (I207003,I206961);
nand I_11997 (I206700,I207003,I206822);
nand I_11998 (I207034,I438772,I438781);
and I_11999 (I207051,I207034,I438775);
DFFARX1 I_12000 (I207051,I3035,I206723,I207077,);
nor I_12001 (I207085,I207077,I206749);
DFFARX1 I_12002 (I207085,I3035,I206723,I206688,);
DFFARX1 I_12003 (I207077,I3035,I206723,I206706,);
nor I_12004 (I207130,I438793,I438781);
not I_12005 (I207147,I207130);
nor I_12006 (I206709,I206986,I207147);
nand I_12007 (I206694,I207003,I207147);
nor I_12008 (I206703,I206749,I207130);
DFFARX1 I_12009 (I207130,I3035,I206723,I206712,);
not I_12010 (I207250,I3042);
DFFARX1 I_12011 (I145539,I3035,I207250,I207276,);
nand I_12012 (I207284,I145539,I145545);
and I_12013 (I207301,I207284,I145563);
DFFARX1 I_12014 (I207301,I3035,I207250,I207327,);
nor I_12015 (I207218,I207327,I207276);
not I_12016 (I207349,I207327);
DFFARX1 I_12017 (I145551,I3035,I207250,I207375,);
nand I_12018 (I207383,I207375,I145548);
not I_12019 (I207400,I207383);
DFFARX1 I_12020 (I207400,I3035,I207250,I207426,);
not I_12021 (I207242,I207426);
nor I_12022 (I207448,I207276,I207383);
nor I_12023 (I207224,I207327,I207448);
DFFARX1 I_12024 (I145557,I3035,I207250,I207488,);
DFFARX1 I_12025 (I207488,I3035,I207250,I207505,);
not I_12026 (I207513,I207505);
not I_12027 (I207530,I207488);
nand I_12028 (I207227,I207530,I207349);
nand I_12029 (I207561,I145542,I145542);
and I_12030 (I207578,I207561,I145554);
DFFARX1 I_12031 (I207578,I3035,I207250,I207604,);
nor I_12032 (I207612,I207604,I207276);
DFFARX1 I_12033 (I207612,I3035,I207250,I207215,);
DFFARX1 I_12034 (I207604,I3035,I207250,I207233,);
nor I_12035 (I207657,I145560,I145542);
not I_12036 (I207674,I207657);
nor I_12037 (I207236,I207513,I207674);
nand I_12038 (I207221,I207530,I207674);
nor I_12039 (I207230,I207276,I207657);
DFFARX1 I_12040 (I207657,I3035,I207250,I207239,);
not I_12041 (I207777,I3042);
DFFARX1 I_12042 (I394380,I3035,I207777,I207803,);
nand I_12043 (I207811,I394371,I394386);
and I_12044 (I207828,I207811,I394392);
DFFARX1 I_12045 (I207828,I3035,I207777,I207854,);
nor I_12046 (I207745,I207854,I207803);
not I_12047 (I207876,I207854);
DFFARX1 I_12048 (I394377,I3035,I207777,I207902,);
nand I_12049 (I207910,I207902,I394371);
not I_12050 (I207927,I207910);
DFFARX1 I_12051 (I207927,I3035,I207777,I207953,);
not I_12052 (I207769,I207953);
nor I_12053 (I207975,I207803,I207910);
nor I_12054 (I207751,I207854,I207975);
DFFARX1 I_12055 (I394374,I3035,I207777,I208015,);
DFFARX1 I_12056 (I208015,I3035,I207777,I208032,);
not I_12057 (I208040,I208032);
not I_12058 (I208057,I208015);
nand I_12059 (I207754,I208057,I207876);
nand I_12060 (I208088,I394368,I394383);
and I_12061 (I208105,I208088,I394368);
DFFARX1 I_12062 (I208105,I3035,I207777,I208131,);
nor I_12063 (I208139,I208131,I207803);
DFFARX1 I_12064 (I208139,I3035,I207777,I207742,);
DFFARX1 I_12065 (I208131,I3035,I207777,I207760,);
nor I_12066 (I208184,I394389,I394383);
not I_12067 (I208201,I208184);
nor I_12068 (I207763,I208040,I208201);
nand I_12069 (I207748,I208057,I208201);
nor I_12070 (I207757,I207803,I208184);
DFFARX1 I_12071 (I208184,I3035,I207777,I207766,);
not I_12072 (I208304,I3042);
DFFARX1 I_12073 (I532921,I3035,I208304,I208330,);
nand I_12074 (I208338,I532918,I532936);
and I_12075 (I208355,I208338,I532927);
DFFARX1 I_12076 (I208355,I3035,I208304,I208381,);
nor I_12077 (I208272,I208381,I208330);
not I_12078 (I208403,I208381);
DFFARX1 I_12079 (I532942,I3035,I208304,I208429,);
nand I_12080 (I208437,I208429,I532924);
not I_12081 (I208454,I208437);
DFFARX1 I_12082 (I208454,I3035,I208304,I208480,);
not I_12083 (I208296,I208480);
nor I_12084 (I208502,I208330,I208437);
nor I_12085 (I208278,I208381,I208502);
DFFARX1 I_12086 (I532930,I3035,I208304,I208542,);
DFFARX1 I_12087 (I208542,I3035,I208304,I208559,);
not I_12088 (I208567,I208559);
not I_12089 (I208584,I208542);
nand I_12090 (I208281,I208584,I208403);
nand I_12091 (I208615,I532918,I532945);
and I_12092 (I208632,I208615,I532933);
DFFARX1 I_12093 (I208632,I3035,I208304,I208658,);
nor I_12094 (I208666,I208658,I208330);
DFFARX1 I_12095 (I208666,I3035,I208304,I208269,);
DFFARX1 I_12096 (I208658,I3035,I208304,I208287,);
nor I_12097 (I208711,I532939,I532945);
not I_12098 (I208728,I208711);
nor I_12099 (I208290,I208567,I208728);
nand I_12100 (I208275,I208584,I208728);
nor I_12101 (I208284,I208330,I208711);
DFFARX1 I_12102 (I208711,I3035,I208304,I208293,);
not I_12103 (I208831,I3042);
DFFARX1 I_12104 (I737704,I3035,I208831,I208857,);
nand I_12105 (I208865,I737683,I737683);
and I_12106 (I208882,I208865,I737710);
DFFARX1 I_12107 (I208882,I3035,I208831,I208908,);
nor I_12108 (I208799,I208908,I208857);
not I_12109 (I208930,I208908);
DFFARX1 I_12110 (I737698,I3035,I208831,I208956,);
nand I_12111 (I208964,I208956,I737701);
not I_12112 (I208981,I208964);
DFFARX1 I_12113 (I208981,I3035,I208831,I209007,);
not I_12114 (I208823,I209007);
nor I_12115 (I209029,I208857,I208964);
nor I_12116 (I208805,I208908,I209029);
DFFARX1 I_12117 (I737692,I3035,I208831,I209069,);
DFFARX1 I_12118 (I209069,I3035,I208831,I209086,);
not I_12119 (I209094,I209086);
not I_12120 (I209111,I209069);
nand I_12121 (I208808,I209111,I208930);
nand I_12122 (I209142,I737689,I737686);
and I_12123 (I209159,I209142,I737707);
DFFARX1 I_12124 (I209159,I3035,I208831,I209185,);
nor I_12125 (I209193,I209185,I208857);
DFFARX1 I_12126 (I209193,I3035,I208831,I208796,);
DFFARX1 I_12127 (I209185,I3035,I208831,I208814,);
nor I_12128 (I209238,I737695,I737686);
not I_12129 (I209255,I209238);
nor I_12130 (I208817,I209094,I209255);
nand I_12131 (I208802,I209111,I209255);
nor I_12132 (I208811,I208857,I209238);
DFFARX1 I_12133 (I209238,I3035,I208831,I208820,);
not I_12134 (I209358,I3042);
DFFARX1 I_12135 (I624310,I3035,I209358,I209384,);
nand I_12136 (I209392,I624325,I624310);
and I_12137 (I209409,I209392,I624328);
DFFARX1 I_12138 (I209409,I3035,I209358,I209435,);
nor I_12139 (I209326,I209435,I209384);
not I_12140 (I209457,I209435);
DFFARX1 I_12141 (I624334,I3035,I209358,I209483,);
nand I_12142 (I209491,I209483,I624316);
not I_12143 (I209508,I209491);
DFFARX1 I_12144 (I209508,I3035,I209358,I209534,);
not I_12145 (I209350,I209534);
nor I_12146 (I209556,I209384,I209491);
nor I_12147 (I209332,I209435,I209556);
DFFARX1 I_12148 (I624313,I3035,I209358,I209596,);
DFFARX1 I_12149 (I209596,I3035,I209358,I209613,);
not I_12150 (I209621,I209613);
not I_12151 (I209638,I209596);
nand I_12152 (I209335,I209638,I209457);
nand I_12153 (I209669,I624313,I624319);
and I_12154 (I209686,I209669,I624331);
DFFARX1 I_12155 (I209686,I3035,I209358,I209712,);
nor I_12156 (I209720,I209712,I209384);
DFFARX1 I_12157 (I209720,I3035,I209358,I209323,);
DFFARX1 I_12158 (I209712,I3035,I209358,I209341,);
nor I_12159 (I209765,I624322,I624319);
not I_12160 (I209782,I209765);
nor I_12161 (I209344,I209621,I209782);
nand I_12162 (I209329,I209638,I209782);
nor I_12163 (I209338,I209384,I209765);
DFFARX1 I_12164 (I209765,I3035,I209358,I209347,);
not I_12165 (I209885,I3042);
DFFARX1 I_12166 (I641072,I3035,I209885,I209911,);
nand I_12167 (I209919,I641087,I641072);
and I_12168 (I209936,I209919,I641090);
DFFARX1 I_12169 (I209936,I3035,I209885,I209962,);
nor I_12170 (I209853,I209962,I209911);
not I_12171 (I209984,I209962);
DFFARX1 I_12172 (I641096,I3035,I209885,I210010,);
nand I_12173 (I210018,I210010,I641078);
not I_12174 (I210035,I210018);
DFFARX1 I_12175 (I210035,I3035,I209885,I210061,);
not I_12176 (I209877,I210061);
nor I_12177 (I210083,I209911,I210018);
nor I_12178 (I209859,I209962,I210083);
DFFARX1 I_12179 (I641075,I3035,I209885,I210123,);
DFFARX1 I_12180 (I210123,I3035,I209885,I210140,);
not I_12181 (I210148,I210140);
not I_12182 (I210165,I210123);
nand I_12183 (I209862,I210165,I209984);
nand I_12184 (I210196,I641075,I641081);
and I_12185 (I210213,I210196,I641093);
DFFARX1 I_12186 (I210213,I3035,I209885,I210239,);
nor I_12187 (I210247,I210239,I209911);
DFFARX1 I_12188 (I210247,I3035,I209885,I209850,);
DFFARX1 I_12189 (I210239,I3035,I209885,I209868,);
nor I_12190 (I210292,I641084,I641081);
not I_12191 (I210309,I210292);
nor I_12192 (I209871,I210148,I210309);
nand I_12193 (I209856,I210165,I210309);
nor I_12194 (I209865,I209911,I210292);
DFFARX1 I_12195 (I210292,I3035,I209885,I209874,);
not I_12196 (I210412,I3042);
DFFARX1 I_12197 (I697839,I3035,I210412,I210438,);
nand I_12198 (I210446,I697818,I697818);
and I_12199 (I210463,I210446,I697845);
DFFARX1 I_12200 (I210463,I3035,I210412,I210489,);
nor I_12201 (I210380,I210489,I210438);
not I_12202 (I210511,I210489);
DFFARX1 I_12203 (I697833,I3035,I210412,I210537,);
nand I_12204 (I210545,I210537,I697836);
not I_12205 (I210562,I210545);
DFFARX1 I_12206 (I210562,I3035,I210412,I210588,);
not I_12207 (I210404,I210588);
nor I_12208 (I210610,I210438,I210545);
nor I_12209 (I210386,I210489,I210610);
DFFARX1 I_12210 (I697827,I3035,I210412,I210650,);
DFFARX1 I_12211 (I210650,I3035,I210412,I210667,);
not I_12212 (I210675,I210667);
not I_12213 (I210692,I210650);
nand I_12214 (I210389,I210692,I210511);
nand I_12215 (I210723,I697824,I697821);
and I_12216 (I210740,I210723,I697842);
DFFARX1 I_12217 (I210740,I3035,I210412,I210766,);
nor I_12218 (I210774,I210766,I210438);
DFFARX1 I_12219 (I210774,I3035,I210412,I210377,);
DFFARX1 I_12220 (I210766,I3035,I210412,I210395,);
nor I_12221 (I210819,I697830,I697821);
not I_12222 (I210836,I210819);
nor I_12223 (I210398,I210675,I210836);
nand I_12224 (I210383,I210692,I210836);
nor I_12225 (I210392,I210438,I210819);
DFFARX1 I_12226 (I210819,I3035,I210412,I210401,);
not I_12227 (I210939,I3042);
DFFARX1 I_12228 (I238065,I3035,I210939,I210965,);
nand I_12229 (I210973,I238077,I238056);
and I_12230 (I210990,I210973,I238080);
DFFARX1 I_12231 (I210990,I3035,I210939,I211016,);
nor I_12232 (I210907,I211016,I210965);
not I_12233 (I211038,I211016);
DFFARX1 I_12234 (I238071,I3035,I210939,I211064,);
nand I_12235 (I211072,I211064,I238053);
not I_12236 (I211089,I211072);
DFFARX1 I_12237 (I211089,I3035,I210939,I211115,);
not I_12238 (I210931,I211115);
nor I_12239 (I211137,I210965,I211072);
nor I_12240 (I210913,I211016,I211137);
DFFARX1 I_12241 (I238068,I3035,I210939,I211177,);
DFFARX1 I_12242 (I211177,I3035,I210939,I211194,);
not I_12243 (I211202,I211194);
not I_12244 (I211219,I211177);
nand I_12245 (I210916,I211219,I211038);
nand I_12246 (I211250,I238053,I238059);
and I_12247 (I211267,I211250,I238062);
DFFARX1 I_12248 (I211267,I3035,I210939,I211293,);
nor I_12249 (I211301,I211293,I210965);
DFFARX1 I_12250 (I211301,I3035,I210939,I210904,);
DFFARX1 I_12251 (I211293,I3035,I210939,I210922,);
nor I_12252 (I211346,I238074,I238059);
not I_12253 (I211363,I211346);
nor I_12254 (I210925,I211202,I211363);
nand I_12255 (I210910,I211219,I211363);
nor I_12256 (I210919,I210965,I211346);
DFFARX1 I_12257 (I211346,I3035,I210939,I210928,);
not I_12258 (I211466,I3042);
DFFARX1 I_12259 (I372416,I3035,I211466,I211492,);
nand I_12260 (I211500,I372407,I372422);
and I_12261 (I211517,I211500,I372428);
DFFARX1 I_12262 (I211517,I3035,I211466,I211543,);
nor I_12263 (I211434,I211543,I211492);
not I_12264 (I211565,I211543);
DFFARX1 I_12265 (I372413,I3035,I211466,I211591,);
nand I_12266 (I211599,I211591,I372407);
not I_12267 (I211616,I211599);
DFFARX1 I_12268 (I211616,I3035,I211466,I211642,);
not I_12269 (I211458,I211642);
nor I_12270 (I211664,I211492,I211599);
nor I_12271 (I211440,I211543,I211664);
DFFARX1 I_12272 (I372410,I3035,I211466,I211704,);
DFFARX1 I_12273 (I211704,I3035,I211466,I211721,);
not I_12274 (I211729,I211721);
not I_12275 (I211746,I211704);
nand I_12276 (I211443,I211746,I211565);
nand I_12277 (I211777,I372404,I372419);
and I_12278 (I211794,I211777,I372404);
DFFARX1 I_12279 (I211794,I3035,I211466,I211820,);
nor I_12280 (I211828,I211820,I211492);
DFFARX1 I_12281 (I211828,I3035,I211466,I211431,);
DFFARX1 I_12282 (I211820,I3035,I211466,I211449,);
nor I_12283 (I211873,I372425,I372419);
not I_12284 (I211890,I211873);
nor I_12285 (I211452,I211729,I211890);
nand I_12286 (I211437,I211746,I211890);
nor I_12287 (I211446,I211492,I211873);
DFFARX1 I_12288 (I211873,I3035,I211466,I211455,);
not I_12289 (I211993,I3042);
DFFARX1 I_12290 (I723424,I3035,I211993,I212019,);
nand I_12291 (I212027,I723403,I723403);
and I_12292 (I212044,I212027,I723430);
DFFARX1 I_12293 (I212044,I3035,I211993,I212070,);
nor I_12294 (I211961,I212070,I212019);
not I_12295 (I212092,I212070);
DFFARX1 I_12296 (I723418,I3035,I211993,I212118,);
nand I_12297 (I212126,I212118,I723421);
not I_12298 (I212143,I212126);
DFFARX1 I_12299 (I212143,I3035,I211993,I212169,);
not I_12300 (I211985,I212169);
nor I_12301 (I212191,I212019,I212126);
nor I_12302 (I211967,I212070,I212191);
DFFARX1 I_12303 (I723412,I3035,I211993,I212231,);
DFFARX1 I_12304 (I212231,I3035,I211993,I212248,);
not I_12305 (I212256,I212248);
not I_12306 (I212273,I212231);
nand I_12307 (I211970,I212273,I212092);
nand I_12308 (I212304,I723409,I723406);
and I_12309 (I212321,I212304,I723427);
DFFARX1 I_12310 (I212321,I3035,I211993,I212347,);
nor I_12311 (I212355,I212347,I212019);
DFFARX1 I_12312 (I212355,I3035,I211993,I211958,);
DFFARX1 I_12313 (I212347,I3035,I211993,I211976,);
nor I_12314 (I212400,I723415,I723406);
not I_12315 (I212417,I212400);
nor I_12316 (I211979,I212256,I212417);
nand I_12317 (I211964,I212273,I212417);
nor I_12318 (I211973,I212019,I212400);
DFFARX1 I_12319 (I212400,I3035,I211993,I211982,);
not I_12320 (I212520,I3042);
DFFARX1 I_12321 (I668120,I3035,I212520,I212546,);
nand I_12322 (I212554,I668102,I668126);
and I_12323 (I212571,I212554,I668117);
DFFARX1 I_12324 (I212571,I3035,I212520,I212597,);
nor I_12325 (I212488,I212597,I212546);
not I_12326 (I212619,I212597);
DFFARX1 I_12327 (I668123,I3035,I212520,I212645,);
nand I_12328 (I212653,I212645,I668111);
not I_12329 (I212670,I212653);
DFFARX1 I_12330 (I212670,I3035,I212520,I212696,);
not I_12331 (I212512,I212696);
nor I_12332 (I212718,I212546,I212653);
nor I_12333 (I212494,I212597,I212718);
DFFARX1 I_12334 (I668102,I3035,I212520,I212758,);
DFFARX1 I_12335 (I212758,I3035,I212520,I212775,);
not I_12336 (I212783,I212775);
not I_12337 (I212800,I212758);
nand I_12338 (I212497,I212800,I212619);
nand I_12339 (I212831,I668108,I668105);
and I_12340 (I212848,I212831,I668114);
DFFARX1 I_12341 (I212848,I3035,I212520,I212874,);
nor I_12342 (I212882,I212874,I212546);
DFFARX1 I_12343 (I212882,I3035,I212520,I212485,);
DFFARX1 I_12344 (I212874,I3035,I212520,I212503,);
nor I_12345 (I212927,I668105,I668105);
not I_12346 (I212944,I212927);
nor I_12347 (I212506,I212783,I212944);
nand I_12348 (I212491,I212800,I212944);
nor I_12349 (I212500,I212546,I212927);
DFFARX1 I_12350 (I212927,I3035,I212520,I212509,);
not I_12351 (I213047,I3042);
DFFARX1 I_12352 (I57346,I3035,I213047,I213073,);
nand I_12353 (I213081,I57358,I57367);
and I_12354 (I213098,I213081,I57346);
DFFARX1 I_12355 (I213098,I3035,I213047,I213124,);
nor I_12356 (I213015,I213124,I213073);
not I_12357 (I213146,I213124);
DFFARX1 I_12358 (I57361,I3035,I213047,I213172,);
nand I_12359 (I213180,I213172,I57349);
not I_12360 (I213197,I213180);
DFFARX1 I_12361 (I213197,I3035,I213047,I213223,);
not I_12362 (I213039,I213223);
nor I_12363 (I213245,I213073,I213180);
nor I_12364 (I213021,I213124,I213245);
DFFARX1 I_12365 (I57352,I3035,I213047,I213285,);
DFFARX1 I_12366 (I213285,I3035,I213047,I213302,);
not I_12367 (I213310,I213302);
not I_12368 (I213327,I213285);
nand I_12369 (I213024,I213327,I213146);
nand I_12370 (I213358,I57343,I57343);
and I_12371 (I213375,I213358,I57355);
DFFARX1 I_12372 (I213375,I3035,I213047,I213401,);
nor I_12373 (I213409,I213401,I213073);
DFFARX1 I_12374 (I213409,I3035,I213047,I213012,);
DFFARX1 I_12375 (I213401,I3035,I213047,I213030,);
nor I_12376 (I213454,I57364,I57343);
not I_12377 (I213471,I213454);
nor I_12378 (I213033,I213310,I213471);
nand I_12379 (I213018,I213327,I213471);
nor I_12380 (I213027,I213073,I213454);
DFFARX1 I_12381 (I213454,I3035,I213047,I213036,);
not I_12382 (I213574,I3042);
DFFARX1 I_12383 (I56292,I3035,I213574,I213600,);
nand I_12384 (I213608,I56304,I56313);
and I_12385 (I213625,I213608,I56292);
DFFARX1 I_12386 (I213625,I3035,I213574,I213651,);
nor I_12387 (I213542,I213651,I213600);
not I_12388 (I213673,I213651);
DFFARX1 I_12389 (I56307,I3035,I213574,I213699,);
nand I_12390 (I213707,I213699,I56295);
not I_12391 (I213724,I213707);
DFFARX1 I_12392 (I213724,I3035,I213574,I213750,);
not I_12393 (I213566,I213750);
nor I_12394 (I213772,I213600,I213707);
nor I_12395 (I213548,I213651,I213772);
DFFARX1 I_12396 (I56298,I3035,I213574,I213812,);
DFFARX1 I_12397 (I213812,I3035,I213574,I213829,);
not I_12398 (I213837,I213829);
not I_12399 (I213854,I213812);
nand I_12400 (I213551,I213854,I213673);
nand I_12401 (I213885,I56289,I56289);
and I_12402 (I213902,I213885,I56301);
DFFARX1 I_12403 (I213902,I3035,I213574,I213928,);
nor I_12404 (I213936,I213928,I213600);
DFFARX1 I_12405 (I213936,I3035,I213574,I213539,);
DFFARX1 I_12406 (I213928,I3035,I213574,I213557,);
nor I_12407 (I213981,I56310,I56289);
not I_12408 (I213998,I213981);
nor I_12409 (I213560,I213837,I213998);
nand I_12410 (I213545,I213854,I213998);
nor I_12411 (I213554,I213600,I213981);
DFFARX1 I_12412 (I213981,I3035,I213574,I213563,);
not I_12413 (I214101,I3042);
DFFARX1 I_12414 (I293629,I3035,I214101,I214127,);
nand I_12415 (I214135,I293629,I293641);
and I_12416 (I214152,I214135,I293626);
DFFARX1 I_12417 (I214152,I3035,I214101,I214178,);
nor I_12418 (I214069,I214178,I214127);
not I_12419 (I214200,I214178);
DFFARX1 I_12420 (I293650,I3035,I214101,I214226,);
nand I_12421 (I214234,I214226,I293647);
not I_12422 (I214251,I214234);
DFFARX1 I_12423 (I214251,I3035,I214101,I214277,);
not I_12424 (I214093,I214277);
nor I_12425 (I214299,I214127,I214234);
nor I_12426 (I214075,I214178,I214299);
DFFARX1 I_12427 (I293638,I3035,I214101,I214339,);
DFFARX1 I_12428 (I214339,I3035,I214101,I214356,);
not I_12429 (I214364,I214356);
not I_12430 (I214381,I214339);
nand I_12431 (I214078,I214381,I214200);
nand I_12432 (I214412,I293626,I293635);
and I_12433 (I214429,I214412,I293644);
DFFARX1 I_12434 (I214429,I3035,I214101,I214455,);
nor I_12435 (I214463,I214455,I214127);
DFFARX1 I_12436 (I214463,I3035,I214101,I214066,);
DFFARX1 I_12437 (I214455,I3035,I214101,I214084,);
nor I_12438 (I214508,I293632,I293635);
not I_12439 (I214525,I214508);
nor I_12440 (I214087,I214364,I214525);
nand I_12441 (I214072,I214381,I214525);
nor I_12442 (I214081,I214127,I214508);
DFFARX1 I_12443 (I214508,I3035,I214101,I214090,);
not I_12444 (I214628,I3042);
DFFARX1 I_12445 (I421911,I3035,I214628,I214654,);
nand I_12446 (I214662,I421914,I421908);
and I_12447 (I214679,I214662,I421920);
DFFARX1 I_12448 (I214679,I3035,I214628,I214705,);
nor I_12449 (I214596,I214705,I214654);
not I_12450 (I214727,I214705);
DFFARX1 I_12451 (I421923,I3035,I214628,I214753,);
nand I_12452 (I214761,I214753,I421914);
not I_12453 (I214778,I214761);
DFFARX1 I_12454 (I214778,I3035,I214628,I214804,);
not I_12455 (I214620,I214804);
nor I_12456 (I214826,I214654,I214761);
nor I_12457 (I214602,I214705,I214826);
DFFARX1 I_12458 (I421926,I3035,I214628,I214866,);
DFFARX1 I_12459 (I214866,I3035,I214628,I214883,);
not I_12460 (I214891,I214883);
not I_12461 (I214908,I214866);
nand I_12462 (I214605,I214908,I214727);
nand I_12463 (I214939,I421908,I421917);
and I_12464 (I214956,I214939,I421911);
DFFARX1 I_12465 (I214956,I3035,I214628,I214982,);
nor I_12466 (I214990,I214982,I214654);
DFFARX1 I_12467 (I214990,I3035,I214628,I214593,);
DFFARX1 I_12468 (I214982,I3035,I214628,I214611,);
nor I_12469 (I215035,I421929,I421917);
not I_12470 (I215052,I215035);
nor I_12471 (I214614,I214891,I215052);
nand I_12472 (I214599,I214908,I215052);
nor I_12473 (I214608,I214654,I215035);
DFFARX1 I_12474 (I215035,I3035,I214628,I214617,);
not I_12475 (I215155,I3042);
DFFARX1 I_12476 (I256561,I3035,I215155,I215181,);
nand I_12477 (I215189,I256573,I256552);
and I_12478 (I215206,I215189,I256576);
DFFARX1 I_12479 (I215206,I3035,I215155,I215232,);
nor I_12480 (I215123,I215232,I215181);
not I_12481 (I215254,I215232);
DFFARX1 I_12482 (I256567,I3035,I215155,I215280,);
nand I_12483 (I215288,I215280,I256549);
not I_12484 (I215305,I215288);
DFFARX1 I_12485 (I215305,I3035,I215155,I215331,);
not I_12486 (I215147,I215331);
nor I_12487 (I215353,I215181,I215288);
nor I_12488 (I215129,I215232,I215353);
DFFARX1 I_12489 (I256564,I3035,I215155,I215393,);
DFFARX1 I_12490 (I215393,I3035,I215155,I215410,);
not I_12491 (I215418,I215410);
not I_12492 (I215435,I215393);
nand I_12493 (I215132,I215435,I215254);
nand I_12494 (I215466,I256549,I256555);
and I_12495 (I215483,I215466,I256558);
DFFARX1 I_12496 (I215483,I3035,I215155,I215509,);
nor I_12497 (I215517,I215509,I215181);
DFFARX1 I_12498 (I215517,I3035,I215155,I215120,);
DFFARX1 I_12499 (I215509,I3035,I215155,I215138,);
nor I_12500 (I215562,I256570,I256555);
not I_12501 (I215579,I215562);
nor I_12502 (I215141,I215418,I215579);
nand I_12503 (I215126,I215435,I215579);
nor I_12504 (I215135,I215181,I215562);
DFFARX1 I_12505 (I215562,I3035,I215155,I215144,);
not I_12506 (I215682,I3042);
DFFARX1 I_12507 (I286489,I3035,I215682,I215708,);
nand I_12508 (I215716,I286489,I286501);
and I_12509 (I215733,I215716,I286486);
DFFARX1 I_12510 (I215733,I3035,I215682,I215759,);
nor I_12511 (I215650,I215759,I215708);
not I_12512 (I215781,I215759);
DFFARX1 I_12513 (I286510,I3035,I215682,I215807,);
nand I_12514 (I215815,I215807,I286507);
not I_12515 (I215832,I215815);
DFFARX1 I_12516 (I215832,I3035,I215682,I215858,);
not I_12517 (I215674,I215858);
nor I_12518 (I215880,I215708,I215815);
nor I_12519 (I215656,I215759,I215880);
DFFARX1 I_12520 (I286498,I3035,I215682,I215920,);
DFFARX1 I_12521 (I215920,I3035,I215682,I215937,);
not I_12522 (I215945,I215937);
not I_12523 (I215962,I215920);
nand I_12524 (I215659,I215962,I215781);
nand I_12525 (I215993,I286486,I286495);
and I_12526 (I216010,I215993,I286504);
DFFARX1 I_12527 (I216010,I3035,I215682,I216036,);
nor I_12528 (I216044,I216036,I215708);
DFFARX1 I_12529 (I216044,I3035,I215682,I215647,);
DFFARX1 I_12530 (I216036,I3035,I215682,I215665,);
nor I_12531 (I216089,I286492,I286495);
not I_12532 (I216106,I216089);
nor I_12533 (I215668,I215945,I216106);
nand I_12534 (I215653,I215962,I216106);
nor I_12535 (I215662,I215708,I216089);
DFFARX1 I_12536 (I216089,I3035,I215682,I215671,);
not I_12537 (I216209,I3042);
DFFARX1 I_12538 (I630090,I3035,I216209,I216235,);
nand I_12539 (I216243,I630105,I630090);
and I_12540 (I216260,I216243,I630108);
DFFARX1 I_12541 (I216260,I3035,I216209,I216286,);
nor I_12542 (I216177,I216286,I216235);
not I_12543 (I216308,I216286);
DFFARX1 I_12544 (I630114,I3035,I216209,I216334,);
nand I_12545 (I216342,I216334,I630096);
not I_12546 (I216359,I216342);
DFFARX1 I_12547 (I216359,I3035,I216209,I216385,);
not I_12548 (I216201,I216385);
nor I_12549 (I216407,I216235,I216342);
nor I_12550 (I216183,I216286,I216407);
DFFARX1 I_12551 (I630093,I3035,I216209,I216447,);
DFFARX1 I_12552 (I216447,I3035,I216209,I216464,);
not I_12553 (I216472,I216464);
not I_12554 (I216489,I216447);
nand I_12555 (I216186,I216489,I216308);
nand I_12556 (I216520,I630093,I630099);
and I_12557 (I216537,I216520,I630111);
DFFARX1 I_12558 (I216537,I3035,I216209,I216563,);
nor I_12559 (I216571,I216563,I216235);
DFFARX1 I_12560 (I216571,I3035,I216209,I216174,);
DFFARX1 I_12561 (I216563,I3035,I216209,I216192,);
nor I_12562 (I216616,I630102,I630099);
not I_12563 (I216633,I216616);
nor I_12564 (I216195,I216472,I216633);
nand I_12565 (I216180,I216489,I216633);
nor I_12566 (I216189,I216235,I216616);
DFFARX1 I_12567 (I216616,I3035,I216209,I216198,);
not I_12568 (I216736,I3042);
DFFARX1 I_12569 (I689843,I3035,I216736,I216762,);
nand I_12570 (I216770,I689840,I689831);
and I_12571 (I216787,I216770,I689828);
DFFARX1 I_12572 (I216787,I3035,I216736,I216813,);
nor I_12573 (I216704,I216813,I216762);
not I_12574 (I216835,I216813);
DFFARX1 I_12575 (I689837,I3035,I216736,I216861,);
nand I_12576 (I216869,I216861,I689846);
not I_12577 (I216886,I216869);
DFFARX1 I_12578 (I216886,I3035,I216736,I216912,);
not I_12579 (I216728,I216912);
nor I_12580 (I216934,I216762,I216869);
nor I_12581 (I216710,I216813,I216934);
DFFARX1 I_12582 (I689849,I3035,I216736,I216974,);
DFFARX1 I_12583 (I216974,I3035,I216736,I216991,);
not I_12584 (I216999,I216991);
not I_12585 (I217016,I216974);
nand I_12586 (I216713,I217016,I216835);
nand I_12587 (I217047,I689828,I689834);
and I_12588 (I217064,I217047,I689852);
DFFARX1 I_12589 (I217064,I3035,I216736,I217090,);
nor I_12590 (I217098,I217090,I216762);
DFFARX1 I_12591 (I217098,I3035,I216736,I216701,);
DFFARX1 I_12592 (I217090,I3035,I216736,I216719,);
nor I_12593 (I217143,I689831,I689834);
not I_12594 (I217160,I217143);
nor I_12595 (I216722,I216999,I217160);
nand I_12596 (I216707,I217016,I217160);
nor I_12597 (I216716,I216762,I217143);
DFFARX1 I_12598 (I217143,I3035,I216736,I216725,);
not I_12599 (I217263,I3042);
DFFARX1 I_12600 (I713309,I3035,I217263,I217289,);
nand I_12601 (I217297,I713288,I713288);
and I_12602 (I217314,I217297,I713315);
DFFARX1 I_12603 (I217314,I3035,I217263,I217340,);
nor I_12604 (I217231,I217340,I217289);
not I_12605 (I217362,I217340);
DFFARX1 I_12606 (I713303,I3035,I217263,I217388,);
nand I_12607 (I217396,I217388,I713306);
not I_12608 (I217413,I217396);
DFFARX1 I_12609 (I217413,I3035,I217263,I217439,);
not I_12610 (I217255,I217439);
nor I_12611 (I217461,I217289,I217396);
nor I_12612 (I217237,I217340,I217461);
DFFARX1 I_12613 (I713297,I3035,I217263,I217501,);
DFFARX1 I_12614 (I217501,I3035,I217263,I217518,);
not I_12615 (I217526,I217518);
not I_12616 (I217543,I217501);
nand I_12617 (I217240,I217543,I217362);
nand I_12618 (I217574,I713294,I713291);
and I_12619 (I217591,I217574,I713312);
DFFARX1 I_12620 (I217591,I3035,I217263,I217617,);
nor I_12621 (I217625,I217617,I217289);
DFFARX1 I_12622 (I217625,I3035,I217263,I217228,);
DFFARX1 I_12623 (I217617,I3035,I217263,I217246,);
nor I_12624 (I217670,I713300,I713291);
not I_12625 (I217687,I217670);
nor I_12626 (I217249,I217526,I217687);
nand I_12627 (I217234,I217543,I217687);
nor I_12628 (I217243,I217289,I217670);
DFFARX1 I_12629 (I217670,I3035,I217263,I217252,);
not I_12630 (I217790,I3042);
DFFARX1 I_12631 (I273969,I3035,I217790,I217816,);
nand I_12632 (I217824,I273981,I273960);
and I_12633 (I217841,I217824,I273984);
DFFARX1 I_12634 (I217841,I3035,I217790,I217867,);
nor I_12635 (I217758,I217867,I217816);
not I_12636 (I217889,I217867);
DFFARX1 I_12637 (I273975,I3035,I217790,I217915,);
nand I_12638 (I217923,I217915,I273957);
not I_12639 (I217940,I217923);
DFFARX1 I_12640 (I217940,I3035,I217790,I217966,);
not I_12641 (I217782,I217966);
nor I_12642 (I217988,I217816,I217923);
nor I_12643 (I217764,I217867,I217988);
DFFARX1 I_12644 (I273972,I3035,I217790,I218028,);
DFFARX1 I_12645 (I218028,I3035,I217790,I218045,);
not I_12646 (I218053,I218045);
not I_12647 (I218070,I218028);
nand I_12648 (I217767,I218070,I217889);
nand I_12649 (I218101,I273957,I273963);
and I_12650 (I218118,I218101,I273966);
DFFARX1 I_12651 (I218118,I3035,I217790,I218144,);
nor I_12652 (I218152,I218144,I217816);
DFFARX1 I_12653 (I218152,I3035,I217790,I217755,);
DFFARX1 I_12654 (I218144,I3035,I217790,I217773,);
nor I_12655 (I218197,I273978,I273963);
not I_12656 (I218214,I218197);
nor I_12657 (I217776,I218053,I218214);
nand I_12658 (I217761,I218070,I218214);
nor I_12659 (I217770,I217816,I218197);
DFFARX1 I_12660 (I218197,I3035,I217790,I217779,);
not I_12661 (I218317,I3042);
DFFARX1 I_12662 (I451423,I3035,I218317,I218343,);
nand I_12663 (I218351,I451426,I451420);
and I_12664 (I218368,I218351,I451432);
DFFARX1 I_12665 (I218368,I3035,I218317,I218394,);
nor I_12666 (I218285,I218394,I218343);
not I_12667 (I218416,I218394);
DFFARX1 I_12668 (I451435,I3035,I218317,I218442,);
nand I_12669 (I218450,I218442,I451426);
not I_12670 (I218467,I218450);
DFFARX1 I_12671 (I218467,I3035,I218317,I218493,);
not I_12672 (I218309,I218493);
nor I_12673 (I218515,I218343,I218450);
nor I_12674 (I218291,I218394,I218515);
DFFARX1 I_12675 (I451438,I3035,I218317,I218555,);
DFFARX1 I_12676 (I218555,I3035,I218317,I218572,);
not I_12677 (I218580,I218572);
not I_12678 (I218597,I218555);
nand I_12679 (I218294,I218597,I218416);
nand I_12680 (I218628,I451420,I451429);
and I_12681 (I218645,I218628,I451423);
DFFARX1 I_12682 (I218645,I3035,I218317,I218671,);
nor I_12683 (I218679,I218671,I218343);
DFFARX1 I_12684 (I218679,I3035,I218317,I218282,);
DFFARX1 I_12685 (I218671,I3035,I218317,I218300,);
nor I_12686 (I218724,I451441,I451429);
not I_12687 (I218741,I218724);
nor I_12688 (I218303,I218580,I218741);
nand I_12689 (I218288,I218597,I218741);
nor I_12690 (I218297,I218343,I218724);
DFFARX1 I_12691 (I218724,I3035,I218317,I218306,);
not I_12692 (I218844,I3042);
DFFARX1 I_12693 (I483825,I3035,I218844,I218870,);
nand I_12694 (I218878,I483822,I483840);
and I_12695 (I218895,I218878,I483831);
DFFARX1 I_12696 (I218895,I3035,I218844,I218921,);
nor I_12697 (I218812,I218921,I218870);
not I_12698 (I218943,I218921);
DFFARX1 I_12699 (I483846,I3035,I218844,I218969,);
nand I_12700 (I218977,I218969,I483828);
not I_12701 (I218994,I218977);
DFFARX1 I_12702 (I218994,I3035,I218844,I219020,);
not I_12703 (I218836,I219020);
nor I_12704 (I219042,I218870,I218977);
nor I_12705 (I218818,I218921,I219042);
DFFARX1 I_12706 (I483834,I3035,I218844,I219082,);
DFFARX1 I_12707 (I219082,I3035,I218844,I219099,);
not I_12708 (I219107,I219099);
not I_12709 (I219124,I219082);
nand I_12710 (I218821,I219124,I218943);
nand I_12711 (I219155,I483822,I483849);
and I_12712 (I219172,I219155,I483837);
DFFARX1 I_12713 (I219172,I3035,I218844,I219198,);
nor I_12714 (I219206,I219198,I218870);
DFFARX1 I_12715 (I219206,I3035,I218844,I218809,);
DFFARX1 I_12716 (I219198,I3035,I218844,I218827,);
nor I_12717 (I219251,I483843,I483849);
not I_12718 (I219268,I219251);
nor I_12719 (I218830,I219107,I219268);
nand I_12720 (I218815,I219124,I219268);
nor I_12721 (I218824,I218870,I219251);
DFFARX1 I_12722 (I219251,I3035,I218844,I218833,);
not I_12723 (I219371,I3042);
DFFARX1 I_12724 (I578648,I3035,I219371,I219397,);
nand I_12725 (I219405,I578663,I578648);
and I_12726 (I219422,I219405,I578666);
DFFARX1 I_12727 (I219422,I3035,I219371,I219448,);
nor I_12728 (I219339,I219448,I219397);
not I_12729 (I219470,I219448);
DFFARX1 I_12730 (I578672,I3035,I219371,I219496,);
nand I_12731 (I219504,I219496,I578654);
not I_12732 (I219521,I219504);
DFFARX1 I_12733 (I219521,I3035,I219371,I219547,);
not I_12734 (I219363,I219547);
nor I_12735 (I219569,I219397,I219504);
nor I_12736 (I219345,I219448,I219569);
DFFARX1 I_12737 (I578651,I3035,I219371,I219609,);
DFFARX1 I_12738 (I219609,I3035,I219371,I219626,);
not I_12739 (I219634,I219626);
not I_12740 (I219651,I219609);
nand I_12741 (I219348,I219651,I219470);
nand I_12742 (I219682,I578651,I578657);
and I_12743 (I219699,I219682,I578669);
DFFARX1 I_12744 (I219699,I3035,I219371,I219725,);
nor I_12745 (I219733,I219725,I219397);
DFFARX1 I_12746 (I219733,I3035,I219371,I219336,);
DFFARX1 I_12747 (I219725,I3035,I219371,I219354,);
nor I_12748 (I219778,I578660,I578657);
not I_12749 (I219795,I219778);
nor I_12750 (I219357,I219634,I219795);
nand I_12751 (I219342,I219651,I219795);
nor I_12752 (I219351,I219397,I219778);
DFFARX1 I_12753 (I219778,I3035,I219371,I219360,);
not I_12754 (I219898,I3042);
DFFARX1 I_12755 (I267985,I3035,I219898,I219924,);
nand I_12756 (I219932,I267997,I267976);
and I_12757 (I219949,I219932,I268000);
DFFARX1 I_12758 (I219949,I3035,I219898,I219975,);
nor I_12759 (I219866,I219975,I219924);
not I_12760 (I219997,I219975);
DFFARX1 I_12761 (I267991,I3035,I219898,I220023,);
nand I_12762 (I220031,I220023,I267973);
not I_12763 (I220048,I220031);
DFFARX1 I_12764 (I220048,I3035,I219898,I220074,);
not I_12765 (I219890,I220074);
nor I_12766 (I220096,I219924,I220031);
nor I_12767 (I219872,I219975,I220096);
DFFARX1 I_12768 (I267988,I3035,I219898,I220136,);
DFFARX1 I_12769 (I220136,I3035,I219898,I220153,);
not I_12770 (I220161,I220153);
not I_12771 (I220178,I220136);
nand I_12772 (I219875,I220178,I219997);
nand I_12773 (I220209,I267973,I267979);
and I_12774 (I220226,I220209,I267982);
DFFARX1 I_12775 (I220226,I3035,I219898,I220252,);
nor I_12776 (I220260,I220252,I219924);
DFFARX1 I_12777 (I220260,I3035,I219898,I219863,);
DFFARX1 I_12778 (I220252,I3035,I219898,I219881,);
nor I_12779 (I220305,I267994,I267979);
not I_12780 (I220322,I220305);
nor I_12781 (I219884,I220161,I220322);
nand I_12782 (I219869,I220178,I220322);
nor I_12783 (I219878,I219924,I220305);
DFFARX1 I_12784 (I220305,I3035,I219898,I219887,);
not I_12785 (I220425,I3042);
DFFARX1 I_12786 (I722829,I3035,I220425,I220451,);
nand I_12787 (I220459,I722808,I722808);
and I_12788 (I220476,I220459,I722835);
DFFARX1 I_12789 (I220476,I3035,I220425,I220502,);
nor I_12790 (I220393,I220502,I220451);
not I_12791 (I220524,I220502);
DFFARX1 I_12792 (I722823,I3035,I220425,I220550,);
nand I_12793 (I220558,I220550,I722826);
not I_12794 (I220575,I220558);
DFFARX1 I_12795 (I220575,I3035,I220425,I220601,);
not I_12796 (I220417,I220601);
nor I_12797 (I220623,I220451,I220558);
nor I_12798 (I220399,I220502,I220623);
DFFARX1 I_12799 (I722817,I3035,I220425,I220663,);
DFFARX1 I_12800 (I220663,I3035,I220425,I220680,);
not I_12801 (I220688,I220680);
not I_12802 (I220705,I220663);
nand I_12803 (I220402,I220705,I220524);
nand I_12804 (I220736,I722814,I722811);
and I_12805 (I220753,I220736,I722832);
DFFARX1 I_12806 (I220753,I3035,I220425,I220779,);
nor I_12807 (I220787,I220779,I220451);
DFFARX1 I_12808 (I220787,I3035,I220425,I220390,);
DFFARX1 I_12809 (I220779,I3035,I220425,I220408,);
nor I_12810 (I220832,I722820,I722811);
not I_12811 (I220849,I220832);
nor I_12812 (I220411,I220688,I220849);
nand I_12813 (I220396,I220705,I220849);
nor I_12814 (I220405,I220451,I220832);
DFFARX1 I_12815 (I220832,I3035,I220425,I220414,);
not I_12816 (I220952,I3042);
DFFARX1 I_12817 (I704384,I3035,I220952,I220978,);
nand I_12818 (I220986,I704363,I704363);
and I_12819 (I221003,I220986,I704390);
DFFARX1 I_12820 (I221003,I3035,I220952,I221029,);
nor I_12821 (I220920,I221029,I220978);
not I_12822 (I221051,I221029);
DFFARX1 I_12823 (I704378,I3035,I220952,I221077,);
nand I_12824 (I221085,I221077,I704381);
not I_12825 (I221102,I221085);
DFFARX1 I_12826 (I221102,I3035,I220952,I221128,);
not I_12827 (I220944,I221128);
nor I_12828 (I221150,I220978,I221085);
nor I_12829 (I220926,I221029,I221150);
DFFARX1 I_12830 (I704372,I3035,I220952,I221190,);
DFFARX1 I_12831 (I221190,I3035,I220952,I221207,);
not I_12832 (I221215,I221207);
not I_12833 (I221232,I221190);
nand I_12834 (I220929,I221232,I221051);
nand I_12835 (I221263,I704369,I704366);
and I_12836 (I221280,I221263,I704387);
DFFARX1 I_12837 (I221280,I3035,I220952,I221306,);
nor I_12838 (I221314,I221306,I220978);
DFFARX1 I_12839 (I221314,I3035,I220952,I220917,);
DFFARX1 I_12840 (I221306,I3035,I220952,I220935,);
nor I_12841 (I221359,I704375,I704366);
not I_12842 (I221376,I221359);
nor I_12843 (I220938,I221215,I221376);
nand I_12844 (I220923,I221232,I221376);
nor I_12845 (I220932,I220978,I221359);
DFFARX1 I_12846 (I221359,I3035,I220952,I220941,);
not I_12847 (I221479,I3042);
DFFARX1 I_12848 (I37320,I3035,I221479,I221505,);
nand I_12849 (I221513,I37332,I37341);
and I_12850 (I221530,I221513,I37320);
DFFARX1 I_12851 (I221530,I3035,I221479,I221556,);
nor I_12852 (I221447,I221556,I221505);
not I_12853 (I221578,I221556);
DFFARX1 I_12854 (I37335,I3035,I221479,I221604,);
nand I_12855 (I221612,I221604,I37323);
not I_12856 (I221629,I221612);
DFFARX1 I_12857 (I221629,I3035,I221479,I221655,);
not I_12858 (I221471,I221655);
nor I_12859 (I221677,I221505,I221612);
nor I_12860 (I221453,I221556,I221677);
DFFARX1 I_12861 (I37326,I3035,I221479,I221717,);
DFFARX1 I_12862 (I221717,I3035,I221479,I221734,);
not I_12863 (I221742,I221734);
not I_12864 (I221759,I221717);
nand I_12865 (I221456,I221759,I221578);
nand I_12866 (I221790,I37317,I37317);
and I_12867 (I221807,I221790,I37329);
DFFARX1 I_12868 (I221807,I3035,I221479,I221833,);
nor I_12869 (I221841,I221833,I221505);
DFFARX1 I_12870 (I221841,I3035,I221479,I221444,);
DFFARX1 I_12871 (I221833,I3035,I221479,I221462,);
nor I_12872 (I221886,I37338,I37317);
not I_12873 (I221903,I221886);
nor I_12874 (I221465,I221742,I221903);
nand I_12875 (I221450,I221759,I221903);
nor I_12876 (I221459,I221505,I221886);
DFFARX1 I_12877 (I221886,I3035,I221479,I221468,);
not I_12878 (I222006,I3042);
DFFARX1 I_12879 (I651800,I3035,I222006,I222032,);
nand I_12880 (I222040,I651782,I651806);
and I_12881 (I222057,I222040,I651797);
DFFARX1 I_12882 (I222057,I3035,I222006,I222083,);
nor I_12883 (I221974,I222083,I222032);
not I_12884 (I222105,I222083);
DFFARX1 I_12885 (I651803,I3035,I222006,I222131,);
nand I_12886 (I222139,I222131,I651791);
not I_12887 (I222156,I222139);
DFFARX1 I_12888 (I222156,I3035,I222006,I222182,);
not I_12889 (I221998,I222182);
nor I_12890 (I222204,I222032,I222139);
nor I_12891 (I221980,I222083,I222204);
DFFARX1 I_12892 (I651782,I3035,I222006,I222244,);
DFFARX1 I_12893 (I222244,I3035,I222006,I222261,);
not I_12894 (I222269,I222261);
not I_12895 (I222286,I222244);
nand I_12896 (I221983,I222286,I222105);
nand I_12897 (I222317,I651788,I651785);
and I_12898 (I222334,I222317,I651794);
DFFARX1 I_12899 (I222334,I3035,I222006,I222360,);
nor I_12900 (I222368,I222360,I222032);
DFFARX1 I_12901 (I222368,I3035,I222006,I221971,);
DFFARX1 I_12902 (I222360,I3035,I222006,I221989,);
nor I_12903 (I222413,I651785,I651785);
not I_12904 (I222430,I222413);
nor I_12905 (I221992,I222269,I222430);
nand I_12906 (I221977,I222286,I222430);
nor I_12907 (I221986,I222032,I222413);
DFFARX1 I_12908 (I222413,I3035,I222006,I221995,);
not I_12909 (I222533,I3042);
DFFARX1 I_12910 (I123524,I3035,I222533,I222559,);
nand I_12911 (I222567,I123524,I123530);
and I_12912 (I222584,I222567,I123548);
DFFARX1 I_12913 (I222584,I3035,I222533,I222610,);
nor I_12914 (I222501,I222610,I222559);
not I_12915 (I222632,I222610);
DFFARX1 I_12916 (I123536,I3035,I222533,I222658,);
nand I_12917 (I222666,I222658,I123533);
not I_12918 (I222683,I222666);
DFFARX1 I_12919 (I222683,I3035,I222533,I222709,);
not I_12920 (I222525,I222709);
nor I_12921 (I222731,I222559,I222666);
nor I_12922 (I222507,I222610,I222731);
DFFARX1 I_12923 (I123542,I3035,I222533,I222771,);
DFFARX1 I_12924 (I222771,I3035,I222533,I222788,);
not I_12925 (I222796,I222788);
not I_12926 (I222813,I222771);
nand I_12927 (I222510,I222813,I222632);
nand I_12928 (I222844,I123527,I123527);
and I_12929 (I222861,I222844,I123539);
DFFARX1 I_12930 (I222861,I3035,I222533,I222887,);
nor I_12931 (I222895,I222887,I222559);
DFFARX1 I_12932 (I222895,I3035,I222533,I222498,);
DFFARX1 I_12933 (I222887,I3035,I222533,I222516,);
nor I_12934 (I222940,I123545,I123527);
not I_12935 (I222957,I222940);
nor I_12936 (I222519,I222796,I222957);
nand I_12937 (I222504,I222813,I222957);
nor I_12938 (I222513,I222559,I222940);
DFFARX1 I_12939 (I222940,I3035,I222533,I222522,);
not I_12940 (I223060,I3042);
DFFARX1 I_12941 (I560512,I3035,I223060,I223086,);
nand I_12942 (I223094,I560509,I560512);
and I_12943 (I223111,I223094,I560521);
DFFARX1 I_12944 (I223111,I3035,I223060,I223137,);
nor I_12945 (I223028,I223137,I223086);
not I_12946 (I223159,I223137);
DFFARX1 I_12947 (I560509,I3035,I223060,I223185,);
nand I_12948 (I223193,I223185,I560527);
not I_12949 (I223210,I223193);
DFFARX1 I_12950 (I223210,I3035,I223060,I223236,);
not I_12951 (I223052,I223236);
nor I_12952 (I223258,I223086,I223193);
nor I_12953 (I223034,I223137,I223258);
DFFARX1 I_12954 (I560515,I3035,I223060,I223298,);
DFFARX1 I_12955 (I223298,I3035,I223060,I223315,);
not I_12956 (I223323,I223315);
not I_12957 (I223340,I223298);
nand I_12958 (I223037,I223340,I223159);
nand I_12959 (I223371,I560524,I560530);
and I_12960 (I223388,I223371,I560515);
DFFARX1 I_12961 (I223388,I3035,I223060,I223414,);
nor I_12962 (I223422,I223414,I223086);
DFFARX1 I_12963 (I223422,I3035,I223060,I223025,);
DFFARX1 I_12964 (I223414,I3035,I223060,I223043,);
nor I_12965 (I223467,I560518,I560530);
not I_12966 (I223484,I223467);
nor I_12967 (I223046,I223323,I223484);
nand I_12968 (I223031,I223340,I223484);
nor I_12969 (I223040,I223086,I223467);
DFFARX1 I_12970 (I223467,I3035,I223060,I223049,);
not I_12971 (I223587,I3042);
DFFARX1 I_12972 (I231537,I3035,I223587,I223613,);
nand I_12973 (I223621,I231549,I231528);
and I_12974 (I223638,I223621,I231552);
DFFARX1 I_12975 (I223638,I3035,I223587,I223664,);
nor I_12976 (I223555,I223664,I223613);
not I_12977 (I223686,I223664);
DFFARX1 I_12978 (I231543,I3035,I223587,I223712,);
nand I_12979 (I223720,I223712,I231525);
not I_12980 (I223737,I223720);
DFFARX1 I_12981 (I223737,I3035,I223587,I223763,);
not I_12982 (I223579,I223763);
nor I_12983 (I223785,I223613,I223720);
nor I_12984 (I223561,I223664,I223785);
DFFARX1 I_12985 (I231540,I3035,I223587,I223825,);
DFFARX1 I_12986 (I223825,I3035,I223587,I223842,);
not I_12987 (I223850,I223842);
not I_12988 (I223867,I223825);
nand I_12989 (I223564,I223867,I223686);
nand I_12990 (I223898,I231525,I231531);
and I_12991 (I223915,I223898,I231534);
DFFARX1 I_12992 (I223915,I3035,I223587,I223941,);
nor I_12993 (I223949,I223941,I223613);
DFFARX1 I_12994 (I223949,I3035,I223587,I223552,);
DFFARX1 I_12995 (I223941,I3035,I223587,I223570,);
nor I_12996 (I223994,I231546,I231531);
not I_12997 (I224011,I223994);
nor I_12998 (I223573,I223850,I224011);
nand I_12999 (I223558,I223867,I224011);
nor I_13000 (I223567,I223613,I223994);
DFFARX1 I_13001 (I223994,I3035,I223587,I223576,);
not I_13002 (I224114,I3042);
DFFARX1 I_13003 (I267441,I3035,I224114,I224140,);
nand I_13004 (I224148,I267453,I267432);
and I_13005 (I224165,I224148,I267456);
DFFARX1 I_13006 (I224165,I3035,I224114,I224191,);
nor I_13007 (I224082,I224191,I224140);
not I_13008 (I224213,I224191);
DFFARX1 I_13009 (I267447,I3035,I224114,I224239,);
nand I_13010 (I224247,I224239,I267429);
not I_13011 (I224264,I224247);
DFFARX1 I_13012 (I224264,I3035,I224114,I224290,);
not I_13013 (I224106,I224290);
nor I_13014 (I224312,I224140,I224247);
nor I_13015 (I224088,I224191,I224312);
DFFARX1 I_13016 (I267444,I3035,I224114,I224352,);
DFFARX1 I_13017 (I224352,I3035,I224114,I224369,);
not I_13018 (I224377,I224369);
not I_13019 (I224394,I224352);
nand I_13020 (I224091,I224394,I224213);
nand I_13021 (I224425,I267429,I267435);
and I_13022 (I224442,I224425,I267438);
DFFARX1 I_13023 (I224442,I3035,I224114,I224468,);
nor I_13024 (I224476,I224468,I224140);
DFFARX1 I_13025 (I224476,I3035,I224114,I224079,);
DFFARX1 I_13026 (I224468,I3035,I224114,I224097,);
nor I_13027 (I224521,I267450,I267435);
not I_13028 (I224538,I224521);
nor I_13029 (I224100,I224377,I224538);
nand I_13030 (I224085,I224394,I224538);
nor I_13031 (I224094,I224140,I224521);
DFFARX1 I_13032 (I224521,I3035,I224114,I224103,);
not I_13033 (I224641,I3042);
DFFARX1 I_13034 (I744844,I3035,I224641,I224667,);
nand I_13035 (I224675,I744823,I744823);
and I_13036 (I224692,I224675,I744850);
DFFARX1 I_13037 (I224692,I3035,I224641,I224718,);
nor I_13038 (I224609,I224718,I224667);
not I_13039 (I224740,I224718);
DFFARX1 I_13040 (I744838,I3035,I224641,I224766,);
nand I_13041 (I224774,I224766,I744841);
not I_13042 (I224791,I224774);
DFFARX1 I_13043 (I224791,I3035,I224641,I224817,);
not I_13044 (I224633,I224817);
nor I_13045 (I224839,I224667,I224774);
nor I_13046 (I224615,I224718,I224839);
DFFARX1 I_13047 (I744832,I3035,I224641,I224879,);
DFFARX1 I_13048 (I224879,I3035,I224641,I224896,);
not I_13049 (I224904,I224896);
not I_13050 (I224921,I224879);
nand I_13051 (I224618,I224921,I224740);
nand I_13052 (I224952,I744829,I744826);
and I_13053 (I224969,I224952,I744847);
DFFARX1 I_13054 (I224969,I3035,I224641,I224995,);
nor I_13055 (I225003,I224995,I224667);
DFFARX1 I_13056 (I225003,I3035,I224641,I224606,);
DFFARX1 I_13057 (I224995,I3035,I224641,I224624,);
nor I_13058 (I225048,I744835,I744826);
not I_13059 (I225065,I225048);
nor I_13060 (I224627,I224904,I225065);
nand I_13061 (I224612,I224921,I225065);
nor I_13062 (I224621,I224667,I225048);
DFFARX1 I_13063 (I225048,I3035,I224641,I224630,);
not I_13064 (I225168,I3042);
DFFARX1 I_13065 (I425600,I3035,I225168,I225194,);
nand I_13066 (I225202,I425603,I425597);
and I_13067 (I225219,I225202,I425609);
DFFARX1 I_13068 (I225219,I3035,I225168,I225245,);
nor I_13069 (I225136,I225245,I225194);
not I_13070 (I225267,I225245);
DFFARX1 I_13071 (I425612,I3035,I225168,I225293,);
nand I_13072 (I225301,I225293,I425603);
not I_13073 (I225318,I225301);
DFFARX1 I_13074 (I225318,I3035,I225168,I225344,);
not I_13075 (I225160,I225344);
nor I_13076 (I225366,I225194,I225301);
nor I_13077 (I225142,I225245,I225366);
DFFARX1 I_13078 (I425615,I3035,I225168,I225406,);
DFFARX1 I_13079 (I225406,I3035,I225168,I225423,);
not I_13080 (I225431,I225423);
not I_13081 (I225448,I225406);
nand I_13082 (I225145,I225448,I225267);
nand I_13083 (I225479,I425597,I425606);
and I_13084 (I225496,I225479,I425600);
DFFARX1 I_13085 (I225496,I3035,I225168,I225522,);
nor I_13086 (I225530,I225522,I225194);
DFFARX1 I_13087 (I225530,I3035,I225168,I225133,);
DFFARX1 I_13088 (I225522,I3035,I225168,I225151,);
nor I_13089 (I225575,I425618,I425606);
not I_13090 (I225592,I225575);
nor I_13091 (I225154,I225431,I225592);
nand I_13092 (I225139,I225448,I225592);
nor I_13093 (I225148,I225194,I225575);
DFFARX1 I_13094 (I225575,I3035,I225168,I225157,);
not I_13095 (I225695,I3042);
DFFARX1 I_13096 (I287084,I3035,I225695,I225721,);
nand I_13097 (I225729,I287084,I287096);
and I_13098 (I225746,I225729,I287081);
DFFARX1 I_13099 (I225746,I3035,I225695,I225772,);
nor I_13100 (I225663,I225772,I225721);
not I_13101 (I225794,I225772);
DFFARX1 I_13102 (I287105,I3035,I225695,I225820,);
nand I_13103 (I225828,I225820,I287102);
not I_13104 (I225845,I225828);
DFFARX1 I_13105 (I225845,I3035,I225695,I225871,);
not I_13106 (I225687,I225871);
nor I_13107 (I225893,I225721,I225828);
nor I_13108 (I225669,I225772,I225893);
DFFARX1 I_13109 (I287093,I3035,I225695,I225933,);
DFFARX1 I_13110 (I225933,I3035,I225695,I225950,);
not I_13111 (I225958,I225950);
not I_13112 (I225975,I225933);
nand I_13113 (I225672,I225975,I225794);
nand I_13114 (I226006,I287081,I287090);
and I_13115 (I226023,I226006,I287099);
DFFARX1 I_13116 (I226023,I3035,I225695,I226049,);
nor I_13117 (I226057,I226049,I225721);
DFFARX1 I_13118 (I226057,I3035,I225695,I225660,);
DFFARX1 I_13119 (I226049,I3035,I225695,I225678,);
nor I_13120 (I226102,I287087,I287090);
not I_13121 (I226119,I226102);
nor I_13122 (I225681,I225958,I226119);
nand I_13123 (I225666,I225975,I226119);
nor I_13124 (I225675,I225721,I226102);
DFFARX1 I_13125 (I226102,I3035,I225695,I225684,);
not I_13126 (I226222,I3042);
DFFARX1 I_13127 (I255473,I3035,I226222,I226248,);
nand I_13128 (I226256,I255485,I255464);
and I_13129 (I226273,I226256,I255488);
DFFARX1 I_13130 (I226273,I3035,I226222,I226299,);
nor I_13131 (I226190,I226299,I226248);
not I_13132 (I226321,I226299);
DFFARX1 I_13133 (I255479,I3035,I226222,I226347,);
nand I_13134 (I226355,I226347,I255461);
not I_13135 (I226372,I226355);
DFFARX1 I_13136 (I226372,I3035,I226222,I226398,);
not I_13137 (I226214,I226398);
nor I_13138 (I226420,I226248,I226355);
nor I_13139 (I226196,I226299,I226420);
DFFARX1 I_13140 (I255476,I3035,I226222,I226460,);
DFFARX1 I_13141 (I226460,I3035,I226222,I226477,);
not I_13142 (I226485,I226477);
not I_13143 (I226502,I226460);
nand I_13144 (I226199,I226502,I226321);
nand I_13145 (I226533,I255461,I255467);
and I_13146 (I226550,I226533,I255470);
DFFARX1 I_13147 (I226550,I3035,I226222,I226576,);
nor I_13148 (I226584,I226576,I226248);
DFFARX1 I_13149 (I226584,I3035,I226222,I226187,);
DFFARX1 I_13150 (I226576,I3035,I226222,I226205,);
nor I_13151 (I226629,I255482,I255467);
not I_13152 (I226646,I226629);
nor I_13153 (I226208,I226485,I226646);
nand I_13154 (I226193,I226502,I226646);
nor I_13155 (I226202,I226248,I226629);
DFFARX1 I_13156 (I226629,I3035,I226222,I226211,);
not I_13157 (I226749,I3042);
DFFARX1 I_13158 (I474084,I3035,I226749,I226775,);
nand I_13159 (I226783,I474087,I474081);
and I_13160 (I226800,I226783,I474093);
DFFARX1 I_13161 (I226800,I3035,I226749,I226826,);
nor I_13162 (I226717,I226826,I226775);
not I_13163 (I226848,I226826);
DFFARX1 I_13164 (I474096,I3035,I226749,I226874,);
nand I_13165 (I226882,I226874,I474087);
not I_13166 (I226899,I226882);
DFFARX1 I_13167 (I226899,I3035,I226749,I226925,);
not I_13168 (I226741,I226925);
nor I_13169 (I226947,I226775,I226882);
nor I_13170 (I226723,I226826,I226947);
DFFARX1 I_13171 (I474099,I3035,I226749,I226987,);
DFFARX1 I_13172 (I226987,I3035,I226749,I227004,);
not I_13173 (I227012,I227004);
not I_13174 (I227029,I226987);
nand I_13175 (I226726,I227029,I226848);
nand I_13176 (I227060,I474081,I474090);
and I_13177 (I227077,I227060,I474084);
DFFARX1 I_13178 (I227077,I3035,I226749,I227103,);
nor I_13179 (I227111,I227103,I226775);
DFFARX1 I_13180 (I227111,I3035,I226749,I226714,);
DFFARX1 I_13181 (I227103,I3035,I226749,I226732,);
nor I_13182 (I227156,I474102,I474090);
not I_13183 (I227173,I227156);
nor I_13184 (I226735,I227012,I227173);
nand I_13185 (I226720,I227029,I227173);
nor I_13186 (I226729,I226775,I227156);
DFFARX1 I_13187 (I227156,I3035,I226749,I226738,);
not I_13188 (I227276,I3042);
DFFARX1 I_13189 (I543257,I3035,I227276,I227302,);
nand I_13190 (I227310,I543254,I543272);
and I_13191 (I227327,I227310,I543263);
DFFARX1 I_13192 (I227327,I3035,I227276,I227353,);
nor I_13193 (I227244,I227353,I227302);
not I_13194 (I227375,I227353);
DFFARX1 I_13195 (I543278,I3035,I227276,I227401,);
nand I_13196 (I227409,I227401,I543260);
not I_13197 (I227426,I227409);
DFFARX1 I_13198 (I227426,I3035,I227276,I227452,);
not I_13199 (I227268,I227452);
nor I_13200 (I227474,I227302,I227409);
nor I_13201 (I227250,I227353,I227474);
DFFARX1 I_13202 (I543266,I3035,I227276,I227514,);
DFFARX1 I_13203 (I227514,I3035,I227276,I227531,);
not I_13204 (I227539,I227531);
not I_13205 (I227556,I227514);
nand I_13206 (I227253,I227556,I227375);
nand I_13207 (I227587,I543254,I543281);
and I_13208 (I227604,I227587,I543269);
DFFARX1 I_13209 (I227604,I3035,I227276,I227630,);
nor I_13210 (I227638,I227630,I227302);
DFFARX1 I_13211 (I227638,I3035,I227276,I227241,);
DFFARX1 I_13212 (I227630,I3035,I227276,I227259,);
nor I_13213 (I227683,I543275,I543281);
not I_13214 (I227700,I227683);
nor I_13215 (I227262,I227539,I227700);
nand I_13216 (I227247,I227556,I227700);
nor I_13217 (I227256,I227302,I227683);
DFFARX1 I_13218 (I227683,I3035,I227276,I227265,);
not I_13219 (I227803,I3042);
DFFARX1 I_13220 (I48914,I3035,I227803,I227829,);
nand I_13221 (I227837,I48926,I48935);
and I_13222 (I227854,I227837,I48914);
DFFARX1 I_13223 (I227854,I3035,I227803,I227880,);
nor I_13224 (I227771,I227880,I227829);
not I_13225 (I227902,I227880);
DFFARX1 I_13226 (I48929,I3035,I227803,I227928,);
nand I_13227 (I227936,I227928,I48917);
not I_13228 (I227953,I227936);
DFFARX1 I_13229 (I227953,I3035,I227803,I227979,);
not I_13230 (I227795,I227979);
nor I_13231 (I228001,I227829,I227936);
nor I_13232 (I227777,I227880,I228001);
DFFARX1 I_13233 (I48920,I3035,I227803,I228041,);
DFFARX1 I_13234 (I228041,I3035,I227803,I228058,);
not I_13235 (I228066,I228058);
not I_13236 (I228083,I228041);
nand I_13237 (I227780,I228083,I227902);
nand I_13238 (I228114,I48911,I48911);
and I_13239 (I228131,I228114,I48923);
DFFARX1 I_13240 (I228131,I3035,I227803,I228157,);
nor I_13241 (I228165,I228157,I227829);
DFFARX1 I_13242 (I228165,I3035,I227803,I227768,);
DFFARX1 I_13243 (I228157,I3035,I227803,I227786,);
nor I_13244 (I228210,I48932,I48911);
not I_13245 (I228227,I228210);
nor I_13246 (I227789,I228066,I228227);
nand I_13247 (I227774,I228083,I228227);
nor I_13248 (I227783,I227829,I228210);
DFFARX1 I_13249 (I228210,I3035,I227803,I227792,);
not I_13250 (I228330,I3042);
DFFARX1 I_13251 (I263089,I3035,I228330,I228356,);
nand I_13252 (I228364,I263101,I263080);
and I_13253 (I228381,I228364,I263104);
DFFARX1 I_13254 (I228381,I3035,I228330,I228407,);
nor I_13255 (I228298,I228407,I228356);
not I_13256 (I228429,I228407);
DFFARX1 I_13257 (I263095,I3035,I228330,I228455,);
nand I_13258 (I228463,I228455,I263077);
not I_13259 (I228480,I228463);
DFFARX1 I_13260 (I228480,I3035,I228330,I228506,);
not I_13261 (I228322,I228506);
nor I_13262 (I228528,I228356,I228463);
nor I_13263 (I228304,I228407,I228528);
DFFARX1 I_13264 (I263092,I3035,I228330,I228568,);
DFFARX1 I_13265 (I228568,I3035,I228330,I228585,);
not I_13266 (I228593,I228585);
not I_13267 (I228610,I228568);
nand I_13268 (I228307,I228610,I228429);
nand I_13269 (I228641,I263077,I263083);
and I_13270 (I228658,I228641,I263086);
DFFARX1 I_13271 (I228658,I3035,I228330,I228684,);
nor I_13272 (I228692,I228684,I228356);
DFFARX1 I_13273 (I228692,I3035,I228330,I228295,);
DFFARX1 I_13274 (I228684,I3035,I228330,I228313,);
nor I_13275 (I228737,I263098,I263083);
not I_13276 (I228754,I228737);
nor I_13277 (I228316,I228593,I228754);
nand I_13278 (I228301,I228610,I228754);
nor I_13279 (I228310,I228356,I228737);
DFFARX1 I_13280 (I228737,I3035,I228330,I228319,);
not I_13281 (I228857,I3042);
DFFARX1 I_13282 (I392646,I3035,I228857,I228883,);
nand I_13283 (I228891,I392637,I392652);
and I_13284 (I228908,I228891,I392658);
DFFARX1 I_13285 (I228908,I3035,I228857,I228934,);
nor I_13286 (I228825,I228934,I228883);
not I_13287 (I228956,I228934);
DFFARX1 I_13288 (I392643,I3035,I228857,I228982,);
nand I_13289 (I228990,I228982,I392637);
not I_13290 (I229007,I228990);
DFFARX1 I_13291 (I229007,I3035,I228857,I229033,);
not I_13292 (I228849,I229033);
nor I_13293 (I229055,I228883,I228990);
nor I_13294 (I228831,I228934,I229055);
DFFARX1 I_13295 (I392640,I3035,I228857,I229095,);
DFFARX1 I_13296 (I229095,I3035,I228857,I229112,);
not I_13297 (I229120,I229112);
not I_13298 (I229137,I229095);
nand I_13299 (I228834,I229137,I228956);
nand I_13300 (I229168,I392634,I392649);
and I_13301 (I229185,I229168,I392634);
DFFARX1 I_13302 (I229185,I3035,I228857,I229211,);
nor I_13303 (I229219,I229211,I228883);
DFFARX1 I_13304 (I229219,I3035,I228857,I228822,);
DFFARX1 I_13305 (I229211,I3035,I228857,I228840,);
nor I_13306 (I229264,I392655,I392649);
not I_13307 (I229281,I229264);
nor I_13308 (I228843,I229120,I229281);
nand I_13309 (I228828,I229137,I229281);
nor I_13310 (I228837,I228883,I229264);
DFFARX1 I_13311 (I229264,I3035,I228857,I228846,);
not I_13312 (I229384,I3042);
DFFARX1 I_13313 (I163495,I3035,I229384,I229410,);
DFFARX1 I_13314 (I229410,I3035,I229384,I229427,);
not I_13315 (I229376,I229427);
not I_13316 (I229449,I229410);
nand I_13317 (I229466,I163474,I163498);
and I_13318 (I229483,I229466,I163501);
DFFARX1 I_13319 (I229483,I3035,I229384,I229509,);
not I_13320 (I229517,I229509);
DFFARX1 I_13321 (I163483,I3035,I229384,I229543,);
and I_13322 (I229551,I229543,I163489);
nand I_13323 (I229568,I229543,I163489);
nand I_13324 (I229355,I229517,I229568);
DFFARX1 I_13325 (I163477,I3035,I229384,I229608,);
nor I_13326 (I229616,I229608,I229551);
DFFARX1 I_13327 (I229616,I3035,I229384,I229349,);
nor I_13328 (I229364,I229608,I229509);
nand I_13329 (I229661,I163486,I163474);
and I_13330 (I229678,I229661,I163480);
DFFARX1 I_13331 (I229678,I3035,I229384,I229704,);
nor I_13332 (I229352,I229704,I229608);
not I_13333 (I229726,I229704);
nor I_13334 (I229743,I229726,I229517);
nor I_13335 (I229760,I229449,I229743);
DFFARX1 I_13336 (I229760,I3035,I229384,I229367,);
nor I_13337 (I229791,I229726,I229608);
nor I_13338 (I229808,I163492,I163474);
nor I_13339 (I229358,I229808,I229791);
not I_13340 (I229839,I229808);
nand I_13341 (I229361,I229568,I229839);
DFFARX1 I_13342 (I229808,I3035,I229384,I229373,);
DFFARX1 I_13343 (I229808,I3035,I229384,I229370,);
not I_13344 (I229928,I3042);
DFFARX1 I_13345 (I647977,I3035,I229928,I229954,);
DFFARX1 I_13346 (I229954,I3035,I229928,I229971,);
not I_13347 (I229920,I229971);
not I_13348 (I229993,I229954);
nand I_13349 (I230010,I647989,I647992);
and I_13350 (I230027,I230010,I647995);
DFFARX1 I_13351 (I230027,I3035,I229928,I230053,);
not I_13352 (I230061,I230053);
DFFARX1 I_13353 (I647980,I3035,I229928,I230087,);
and I_13354 (I230095,I230087,I647986);
nand I_13355 (I230112,I230087,I647986);
nand I_13356 (I229899,I230061,I230112);
DFFARX1 I_13357 (I647974,I3035,I229928,I230152,);
nor I_13358 (I230160,I230152,I230095);
DFFARX1 I_13359 (I230160,I3035,I229928,I229893,);
nor I_13360 (I229908,I230152,I230053);
nand I_13361 (I230205,I647977,I647998);
and I_13362 (I230222,I230205,I647983);
DFFARX1 I_13363 (I230222,I3035,I229928,I230248,);
nor I_13364 (I229896,I230248,I230152);
not I_13365 (I230270,I230248);
nor I_13366 (I230287,I230270,I230061);
nor I_13367 (I230304,I229993,I230287);
DFFARX1 I_13368 (I230304,I3035,I229928,I229911,);
nor I_13369 (I230335,I230270,I230152);
nor I_13370 (I230352,I647974,I647998);
nor I_13371 (I229902,I230352,I230335);
not I_13372 (I230383,I230352);
nand I_13373 (I229905,I230112,I230383);
DFFARX1 I_13374 (I230352,I3035,I229928,I229917,);
DFFARX1 I_13375 (I230352,I3035,I229928,I229914,);
not I_13376 (I230472,I3042);
DFFARX1 I_13377 (I176670,I3035,I230472,I230498,);
DFFARX1 I_13378 (I230498,I3035,I230472,I230515,);
not I_13379 (I230464,I230515);
not I_13380 (I230537,I230498);
nand I_13381 (I230554,I176649,I176673);
and I_13382 (I230571,I230554,I176676);
DFFARX1 I_13383 (I230571,I3035,I230472,I230597,);
not I_13384 (I230605,I230597);
DFFARX1 I_13385 (I176658,I3035,I230472,I230631,);
and I_13386 (I230639,I230631,I176664);
nand I_13387 (I230656,I230631,I176664);
nand I_13388 (I230443,I230605,I230656);
DFFARX1 I_13389 (I176652,I3035,I230472,I230696,);
nor I_13390 (I230704,I230696,I230639);
DFFARX1 I_13391 (I230704,I3035,I230472,I230437,);
nor I_13392 (I230452,I230696,I230597);
nand I_13393 (I230749,I176661,I176649);
and I_13394 (I230766,I230749,I176655);
DFFARX1 I_13395 (I230766,I3035,I230472,I230792,);
nor I_13396 (I230440,I230792,I230696);
not I_13397 (I230814,I230792);
nor I_13398 (I230831,I230814,I230605);
nor I_13399 (I230848,I230537,I230831);
DFFARX1 I_13400 (I230848,I3035,I230472,I230455,);
nor I_13401 (I230879,I230814,I230696);
nor I_13402 (I230896,I176667,I176649);
nor I_13403 (I230446,I230896,I230879);
not I_13404 (I230927,I230896);
nand I_13405 (I230449,I230656,I230927);
DFFARX1 I_13406 (I230896,I3035,I230472,I230461,);
DFFARX1 I_13407 (I230896,I3035,I230472,I230458,);
not I_13408 (I231016,I3042);
DFFARX1 I_13409 (I47336,I3035,I231016,I231042,);
DFFARX1 I_13410 (I231042,I3035,I231016,I231059,);
not I_13411 (I231008,I231059);
not I_13412 (I231081,I231042);
nand I_13413 (I231098,I47351,I47330);
and I_13414 (I231115,I231098,I47333);
DFFARX1 I_13415 (I231115,I3035,I231016,I231141,);
not I_13416 (I231149,I231141);
DFFARX1 I_13417 (I47339,I3035,I231016,I231175,);
and I_13418 (I231183,I231175,I47333);
nand I_13419 (I231200,I231175,I47333);
nand I_13420 (I230987,I231149,I231200);
DFFARX1 I_13421 (I47348,I3035,I231016,I231240,);
nor I_13422 (I231248,I231240,I231183);
DFFARX1 I_13423 (I231248,I3035,I231016,I230981,);
nor I_13424 (I230996,I231240,I231141);
nand I_13425 (I231293,I47330,I47345);
and I_13426 (I231310,I231293,I47342);
DFFARX1 I_13427 (I231310,I3035,I231016,I231336,);
nor I_13428 (I230984,I231336,I231240);
not I_13429 (I231358,I231336);
nor I_13430 (I231375,I231358,I231149);
nor I_13431 (I231392,I231081,I231375);
DFFARX1 I_13432 (I231392,I3035,I231016,I230999,);
nor I_13433 (I231423,I231358,I231240);
nor I_13434 (I231440,I47354,I47345);
nor I_13435 (I230990,I231440,I231423);
not I_13436 (I231471,I231440);
nand I_13437 (I230993,I231200,I231471);
DFFARX1 I_13438 (I231440,I3035,I231016,I231005,);
DFFARX1 I_13439 (I231440,I3035,I231016,I231002,);
not I_13440 (I231560,I3042);
DFFARX1 I_13441 (I54714,I3035,I231560,I231586,);
DFFARX1 I_13442 (I231586,I3035,I231560,I231603,);
not I_13443 (I231552,I231603);
not I_13444 (I231625,I231586);
nand I_13445 (I231642,I54729,I54708);
and I_13446 (I231659,I231642,I54711);
DFFARX1 I_13447 (I231659,I3035,I231560,I231685,);
not I_13448 (I231693,I231685);
DFFARX1 I_13449 (I54717,I3035,I231560,I231719,);
and I_13450 (I231727,I231719,I54711);
nand I_13451 (I231744,I231719,I54711);
nand I_13452 (I231531,I231693,I231744);
DFFARX1 I_13453 (I54726,I3035,I231560,I231784,);
nor I_13454 (I231792,I231784,I231727);
DFFARX1 I_13455 (I231792,I3035,I231560,I231525,);
nor I_13456 (I231540,I231784,I231685);
nand I_13457 (I231837,I54708,I54723);
and I_13458 (I231854,I231837,I54720);
DFFARX1 I_13459 (I231854,I3035,I231560,I231880,);
nor I_13460 (I231528,I231880,I231784);
not I_13461 (I231902,I231880);
nor I_13462 (I231919,I231902,I231693);
nor I_13463 (I231936,I231625,I231919);
DFFARX1 I_13464 (I231936,I3035,I231560,I231543,);
nor I_13465 (I231967,I231902,I231784);
nor I_13466 (I231984,I54732,I54723);
nor I_13467 (I231534,I231984,I231967);
not I_13468 (I232015,I231984);
nand I_13469 (I231537,I231744,I232015);
DFFARX1 I_13470 (I231984,I3035,I231560,I231549,);
DFFARX1 I_13471 (I231984,I3035,I231560,I231546,);
not I_13472 (I232104,I3042);
DFFARX1 I_13473 (I320965,I3035,I232104,I232130,);
DFFARX1 I_13474 (I232130,I3035,I232104,I232147,);
not I_13475 (I232096,I232147);
not I_13476 (I232169,I232130);
nand I_13477 (I232186,I320962,I320983);
and I_13478 (I232203,I232186,I320986);
DFFARX1 I_13479 (I232203,I3035,I232104,I232229,);
not I_13480 (I232237,I232229);
DFFARX1 I_13481 (I320971,I3035,I232104,I232263,);
and I_13482 (I232271,I232263,I320974);
nand I_13483 (I232288,I232263,I320974);
nand I_13484 (I232075,I232237,I232288);
DFFARX1 I_13485 (I320977,I3035,I232104,I232328,);
nor I_13486 (I232336,I232328,I232271);
DFFARX1 I_13487 (I232336,I3035,I232104,I232069,);
nor I_13488 (I232084,I232328,I232229);
nand I_13489 (I232381,I320962,I320968);
and I_13490 (I232398,I232381,I320980);
DFFARX1 I_13491 (I232398,I3035,I232104,I232424,);
nor I_13492 (I232072,I232424,I232328);
not I_13493 (I232446,I232424);
nor I_13494 (I232463,I232446,I232237);
nor I_13495 (I232480,I232169,I232463);
DFFARX1 I_13496 (I232480,I3035,I232104,I232087,);
nor I_13497 (I232511,I232446,I232328);
nor I_13498 (I232528,I320965,I320968);
nor I_13499 (I232078,I232528,I232511);
not I_13500 (I232559,I232528);
nand I_13501 (I232081,I232288,I232559);
DFFARX1 I_13502 (I232528,I3035,I232104,I232093,);
DFFARX1 I_13503 (I232528,I3035,I232104,I232090,);
not I_13504 (I232648,I3042);
DFFARX1 I_13505 (I437730,I3035,I232648,I232674,);
DFFARX1 I_13506 (I232674,I3035,I232648,I232691,);
not I_13507 (I232640,I232691);
not I_13508 (I232713,I232674);
nand I_13509 (I232730,I437724,I437721);
and I_13510 (I232747,I232730,I437736);
DFFARX1 I_13511 (I232747,I3035,I232648,I232773,);
not I_13512 (I232781,I232773);
DFFARX1 I_13513 (I437724,I3035,I232648,I232807,);
and I_13514 (I232815,I232807,I437718);
nand I_13515 (I232832,I232807,I437718);
nand I_13516 (I232619,I232781,I232832);
DFFARX1 I_13517 (I437718,I3035,I232648,I232872,);
nor I_13518 (I232880,I232872,I232815);
DFFARX1 I_13519 (I232880,I3035,I232648,I232613,);
nor I_13520 (I232628,I232872,I232773);
nand I_13521 (I232925,I437733,I437727);
and I_13522 (I232942,I232925,I437721);
DFFARX1 I_13523 (I232942,I3035,I232648,I232968,);
nor I_13524 (I232616,I232968,I232872);
not I_13525 (I232990,I232968);
nor I_13526 (I233007,I232990,I232781);
nor I_13527 (I233024,I232713,I233007);
DFFARX1 I_13528 (I233024,I3035,I232648,I232631,);
nor I_13529 (I233055,I232990,I232872);
nor I_13530 (I233072,I437739,I437727);
nor I_13531 (I232622,I233072,I233055);
not I_13532 (I233103,I233072);
nand I_13533 (I232625,I232832,I233103);
DFFARX1 I_13534 (I233072,I3035,I232648,I232637,);
DFFARX1 I_13535 (I233072,I3035,I232648,I232634,);
not I_13536 (I233192,I3042);
DFFARX1 I_13537 (I459337,I3035,I233192,I233218,);
DFFARX1 I_13538 (I233218,I3035,I233192,I233235,);
not I_13539 (I233184,I233235);
not I_13540 (I233257,I233218);
nand I_13541 (I233274,I459331,I459328);
and I_13542 (I233291,I233274,I459343);
DFFARX1 I_13543 (I233291,I3035,I233192,I233317,);
not I_13544 (I233325,I233317);
DFFARX1 I_13545 (I459331,I3035,I233192,I233351,);
and I_13546 (I233359,I233351,I459325);
nand I_13547 (I233376,I233351,I459325);
nand I_13548 (I233163,I233325,I233376);
DFFARX1 I_13549 (I459325,I3035,I233192,I233416,);
nor I_13550 (I233424,I233416,I233359);
DFFARX1 I_13551 (I233424,I3035,I233192,I233157,);
nor I_13552 (I233172,I233416,I233317);
nand I_13553 (I233469,I459340,I459334);
and I_13554 (I233486,I233469,I459328);
DFFARX1 I_13555 (I233486,I3035,I233192,I233512,);
nor I_13556 (I233160,I233512,I233416);
not I_13557 (I233534,I233512);
nor I_13558 (I233551,I233534,I233325);
nor I_13559 (I233568,I233257,I233551);
DFFARX1 I_13560 (I233568,I3035,I233192,I233175,);
nor I_13561 (I233599,I233534,I233416);
nor I_13562 (I233616,I459346,I459334);
nor I_13563 (I233166,I233616,I233599);
not I_13564 (I233647,I233616);
nand I_13565 (I233169,I233376,I233647);
DFFARX1 I_13566 (I233616,I3035,I233192,I233181,);
DFFARX1 I_13567 (I233616,I3035,I233192,I233178,);
not I_13568 (I233736,I3042);
DFFARX1 I_13569 (I620845,I3035,I233736,I233762,);
DFFARX1 I_13570 (I233762,I3035,I233736,I233779,);
not I_13571 (I233728,I233779);
not I_13572 (I233801,I233762);
nand I_13573 (I233818,I620857,I620845);
and I_13574 (I233835,I233818,I620848);
DFFARX1 I_13575 (I233835,I3035,I233736,I233861,);
not I_13576 (I233869,I233861);
DFFARX1 I_13577 (I620866,I3035,I233736,I233895,);
and I_13578 (I233903,I233895,I620842);
nand I_13579 (I233920,I233895,I620842);
nand I_13580 (I233707,I233869,I233920);
DFFARX1 I_13581 (I620860,I3035,I233736,I233960,);
nor I_13582 (I233968,I233960,I233903);
DFFARX1 I_13583 (I233968,I3035,I233736,I233701,);
nor I_13584 (I233716,I233960,I233861);
nand I_13585 (I234013,I620854,I620851);
and I_13586 (I234030,I234013,I620863);
DFFARX1 I_13587 (I234030,I3035,I233736,I234056,);
nor I_13588 (I233704,I234056,I233960);
not I_13589 (I234078,I234056);
nor I_13590 (I234095,I234078,I233869);
nor I_13591 (I234112,I233801,I234095);
DFFARX1 I_13592 (I234112,I3035,I233736,I233719,);
nor I_13593 (I234143,I234078,I233960);
nor I_13594 (I234160,I620842,I620851);
nor I_13595 (I233710,I234160,I234143);
not I_13596 (I234191,I234160);
nand I_13597 (I233713,I233920,I234191);
DFFARX1 I_13598 (I234160,I3035,I233736,I233725,);
DFFARX1 I_13599 (I234160,I3035,I233736,I233722,);
not I_13600 (I234280,I3042);
DFFARX1 I_13601 (I628937,I3035,I234280,I234306,);
DFFARX1 I_13602 (I234306,I3035,I234280,I234323,);
not I_13603 (I234272,I234323);
not I_13604 (I234345,I234306);
nand I_13605 (I234362,I628949,I628937);
and I_13606 (I234379,I234362,I628940);
DFFARX1 I_13607 (I234379,I3035,I234280,I234405,);
not I_13608 (I234413,I234405);
DFFARX1 I_13609 (I628958,I3035,I234280,I234439,);
and I_13610 (I234447,I234439,I628934);
nand I_13611 (I234464,I234439,I628934);
nand I_13612 (I234251,I234413,I234464);
DFFARX1 I_13613 (I628952,I3035,I234280,I234504,);
nor I_13614 (I234512,I234504,I234447);
DFFARX1 I_13615 (I234512,I3035,I234280,I234245,);
nor I_13616 (I234260,I234504,I234405);
nand I_13617 (I234557,I628946,I628943);
and I_13618 (I234574,I234557,I628955);
DFFARX1 I_13619 (I234574,I3035,I234280,I234600,);
nor I_13620 (I234248,I234600,I234504);
not I_13621 (I234622,I234600);
nor I_13622 (I234639,I234622,I234413);
nor I_13623 (I234656,I234345,I234639);
DFFARX1 I_13624 (I234656,I3035,I234280,I234263,);
nor I_13625 (I234687,I234622,I234504);
nor I_13626 (I234704,I628934,I628943);
nor I_13627 (I234254,I234704,I234687);
not I_13628 (I234735,I234704);
nand I_13629 (I234257,I234464,I234735);
DFFARX1 I_13630 (I234704,I3035,I234280,I234269,);
DFFARX1 I_13631 (I234704,I3035,I234280,I234266,);
not I_13632 (I234824,I3042);
DFFARX1 I_13633 (I488350,I3035,I234824,I234850,);
DFFARX1 I_13634 (I234850,I3035,I234824,I234867,);
not I_13635 (I234816,I234867);
not I_13636 (I234889,I234850);
nand I_13637 (I234906,I488365,I488353);
and I_13638 (I234923,I234906,I488344);
DFFARX1 I_13639 (I234923,I3035,I234824,I234949,);
not I_13640 (I234957,I234949);
DFFARX1 I_13641 (I488356,I3035,I234824,I234983,);
and I_13642 (I234991,I234983,I488347);
nand I_13643 (I235008,I234983,I488347);
nand I_13644 (I234795,I234957,I235008);
DFFARX1 I_13645 (I488362,I3035,I234824,I235048,);
nor I_13646 (I235056,I235048,I234991);
DFFARX1 I_13647 (I235056,I3035,I234824,I234789,);
nor I_13648 (I234804,I235048,I234949);
nand I_13649 (I235101,I488371,I488359);
and I_13650 (I235118,I235101,I488368);
DFFARX1 I_13651 (I235118,I3035,I234824,I235144,);
nor I_13652 (I234792,I235144,I235048);
not I_13653 (I235166,I235144);
nor I_13654 (I235183,I235166,I234957);
nor I_13655 (I235200,I234889,I235183);
DFFARX1 I_13656 (I235200,I3035,I234824,I234807,);
nor I_13657 (I235231,I235166,I235048);
nor I_13658 (I235248,I488344,I488359);
nor I_13659 (I234798,I235248,I235231);
not I_13660 (I235279,I235248);
nand I_13661 (I234801,I235008,I235279);
DFFARX1 I_13662 (I235248,I3035,I234824,I234813,);
DFFARX1 I_13663 (I235248,I3035,I234824,I234810,);
not I_13664 (I235368,I3042);
DFFARX1 I_13665 (I72105,I3035,I235368,I235394,);
DFFARX1 I_13666 (I235394,I3035,I235368,I235411,);
not I_13667 (I235360,I235411);
not I_13668 (I235433,I235394);
nand I_13669 (I235450,I72120,I72099);
and I_13670 (I235467,I235450,I72102);
DFFARX1 I_13671 (I235467,I3035,I235368,I235493,);
not I_13672 (I235501,I235493);
DFFARX1 I_13673 (I72108,I3035,I235368,I235527,);
and I_13674 (I235535,I235527,I72102);
nand I_13675 (I235552,I235527,I72102);
nand I_13676 (I235339,I235501,I235552);
DFFARX1 I_13677 (I72117,I3035,I235368,I235592,);
nor I_13678 (I235600,I235592,I235535);
DFFARX1 I_13679 (I235600,I3035,I235368,I235333,);
nor I_13680 (I235348,I235592,I235493);
nand I_13681 (I235645,I72099,I72114);
and I_13682 (I235662,I235645,I72111);
DFFARX1 I_13683 (I235662,I3035,I235368,I235688,);
nor I_13684 (I235336,I235688,I235592);
not I_13685 (I235710,I235688);
nor I_13686 (I235727,I235710,I235501);
nor I_13687 (I235744,I235433,I235727);
DFFARX1 I_13688 (I235744,I3035,I235368,I235351,);
nor I_13689 (I235775,I235710,I235592);
nor I_13690 (I235792,I72123,I72114);
nor I_13691 (I235342,I235792,I235775);
not I_13692 (I235823,I235792);
nand I_13693 (I235345,I235552,I235823);
DFFARX1 I_13694 (I235792,I3035,I235368,I235357,);
DFFARX1 I_13695 (I235792,I3035,I235368,I235354,);
not I_13696 (I235912,I3042);
DFFARX1 I_13697 (I479306,I3035,I235912,I235938,);
DFFARX1 I_13698 (I235938,I3035,I235912,I235955,);
not I_13699 (I235904,I235955);
not I_13700 (I235977,I235938);
nand I_13701 (I235994,I479321,I479309);
and I_13702 (I236011,I235994,I479300);
DFFARX1 I_13703 (I236011,I3035,I235912,I236037,);
not I_13704 (I236045,I236037);
DFFARX1 I_13705 (I479312,I3035,I235912,I236071,);
and I_13706 (I236079,I236071,I479303);
nand I_13707 (I236096,I236071,I479303);
nand I_13708 (I235883,I236045,I236096);
DFFARX1 I_13709 (I479318,I3035,I235912,I236136,);
nor I_13710 (I236144,I236136,I236079);
DFFARX1 I_13711 (I236144,I3035,I235912,I235877,);
nor I_13712 (I235892,I236136,I236037);
nand I_13713 (I236189,I479327,I479315);
and I_13714 (I236206,I236189,I479324);
DFFARX1 I_13715 (I236206,I3035,I235912,I236232,);
nor I_13716 (I235880,I236232,I236136);
not I_13717 (I236254,I236232);
nor I_13718 (I236271,I236254,I236045);
nor I_13719 (I236288,I235977,I236271);
DFFARX1 I_13720 (I236288,I3035,I235912,I235895,);
nor I_13721 (I236319,I236254,I236136);
nor I_13722 (I236336,I479300,I479315);
nor I_13723 (I235886,I236336,I236319);
not I_13724 (I236367,I236336);
nand I_13725 (I235889,I236096,I236367);
DFFARX1 I_13726 (I236336,I3035,I235912,I235901,);
DFFARX1 I_13727 (I236336,I3035,I235912,I235898,);
not I_13728 (I236456,I3042);
DFFARX1 I_13729 (I209871,I3035,I236456,I236482,);
DFFARX1 I_13730 (I236482,I3035,I236456,I236499,);
not I_13731 (I236448,I236499);
not I_13732 (I236521,I236482);
nand I_13733 (I236538,I209850,I209874);
and I_13734 (I236555,I236538,I209877);
DFFARX1 I_13735 (I236555,I3035,I236456,I236581,);
not I_13736 (I236589,I236581);
DFFARX1 I_13737 (I209859,I3035,I236456,I236615,);
and I_13738 (I236623,I236615,I209865);
nand I_13739 (I236640,I236615,I209865);
nand I_13740 (I236427,I236589,I236640);
DFFARX1 I_13741 (I209853,I3035,I236456,I236680,);
nor I_13742 (I236688,I236680,I236623);
DFFARX1 I_13743 (I236688,I3035,I236456,I236421,);
nor I_13744 (I236436,I236680,I236581);
nand I_13745 (I236733,I209862,I209850);
and I_13746 (I236750,I236733,I209856);
DFFARX1 I_13747 (I236750,I3035,I236456,I236776,);
nor I_13748 (I236424,I236776,I236680);
not I_13749 (I236798,I236776);
nor I_13750 (I236815,I236798,I236589);
nor I_13751 (I236832,I236521,I236815);
DFFARX1 I_13752 (I236832,I3035,I236456,I236439,);
nor I_13753 (I236863,I236798,I236680);
nor I_13754 (I236880,I209868,I209850);
nor I_13755 (I236430,I236880,I236863);
not I_13756 (I236911,I236880);
nand I_13757 (I236433,I236640,I236911);
DFFARX1 I_13758 (I236880,I3035,I236456,I236445,);
DFFARX1 I_13759 (I236880,I3035,I236456,I236442,);
not I_13760 (I237000,I3042);
DFFARX1 I_13761 (I21519,I3035,I237000,I237026,);
DFFARX1 I_13762 (I237026,I3035,I237000,I237043,);
not I_13763 (I236992,I237043);
not I_13764 (I237065,I237026);
nand I_13765 (I237082,I21507,I21522);
and I_13766 (I237099,I237082,I21510);
DFFARX1 I_13767 (I237099,I3035,I237000,I237125,);
not I_13768 (I237133,I237125);
DFFARX1 I_13769 (I21531,I3035,I237000,I237159,);
and I_13770 (I237167,I237159,I21525);
nand I_13771 (I237184,I237159,I21525);
nand I_13772 (I236971,I237133,I237184);
DFFARX1 I_13773 (I21528,I3035,I237000,I237224,);
nor I_13774 (I237232,I237224,I237167);
DFFARX1 I_13775 (I237232,I3035,I237000,I236965,);
nor I_13776 (I236980,I237224,I237125);
nand I_13777 (I237277,I21507,I21510);
and I_13778 (I237294,I237277,I21513);
DFFARX1 I_13779 (I237294,I3035,I237000,I237320,);
nor I_13780 (I236968,I237320,I237224);
not I_13781 (I237342,I237320);
nor I_13782 (I237359,I237342,I237133);
nor I_13783 (I237376,I237065,I237359);
DFFARX1 I_13784 (I237376,I3035,I237000,I236983,);
nor I_13785 (I237407,I237342,I237224);
nor I_13786 (I237424,I21516,I21510);
nor I_13787 (I236974,I237424,I237407);
not I_13788 (I237455,I237424);
nand I_13789 (I236977,I237184,I237455);
DFFARX1 I_13790 (I237424,I3035,I237000,I236989,);
DFFARX1 I_13791 (I237424,I3035,I237000,I236986,);
not I_13792 (I237544,I3042);
DFFARX1 I_13793 (I505146,I3035,I237544,I237570,);
DFFARX1 I_13794 (I237570,I3035,I237544,I237587,);
not I_13795 (I237536,I237587);
not I_13796 (I237609,I237570);
nand I_13797 (I237626,I505161,I505149);
and I_13798 (I237643,I237626,I505140);
DFFARX1 I_13799 (I237643,I3035,I237544,I237669,);
not I_13800 (I237677,I237669);
DFFARX1 I_13801 (I505152,I3035,I237544,I237703,);
and I_13802 (I237711,I237703,I505143);
nand I_13803 (I237728,I237703,I505143);
nand I_13804 (I237515,I237677,I237728);
DFFARX1 I_13805 (I505158,I3035,I237544,I237768,);
nor I_13806 (I237776,I237768,I237711);
DFFARX1 I_13807 (I237776,I3035,I237544,I237509,);
nor I_13808 (I237524,I237768,I237669);
nand I_13809 (I237821,I505167,I505155);
and I_13810 (I237838,I237821,I505164);
DFFARX1 I_13811 (I237838,I3035,I237544,I237864,);
nor I_13812 (I237512,I237864,I237768);
not I_13813 (I237886,I237864);
nor I_13814 (I237903,I237886,I237677);
nor I_13815 (I237920,I237609,I237903);
DFFARX1 I_13816 (I237920,I3035,I237544,I237527,);
nor I_13817 (I237951,I237886,I237768);
nor I_13818 (I237968,I505140,I505155);
nor I_13819 (I237518,I237968,I237951);
not I_13820 (I237999,I237968);
nand I_13821 (I237521,I237728,I237999);
DFFARX1 I_13822 (I237968,I3035,I237544,I237533,);
DFFARX1 I_13823 (I237968,I3035,I237544,I237530,);
not I_13824 (I238088,I3042);
DFFARX1 I_13825 (I365471,I3035,I238088,I238114,);
DFFARX1 I_13826 (I238114,I3035,I238088,I238131,);
not I_13827 (I238080,I238131);
not I_13828 (I238153,I238114);
nand I_13829 (I238170,I365492,I365483);
and I_13830 (I238187,I238170,I365471);
DFFARX1 I_13831 (I238187,I3035,I238088,I238213,);
not I_13832 (I238221,I238213);
DFFARX1 I_13833 (I365477,I3035,I238088,I238247,);
and I_13834 (I238255,I238247,I365474);
nand I_13835 (I238272,I238247,I365474);
nand I_13836 (I238059,I238221,I238272);
DFFARX1 I_13837 (I365468,I3035,I238088,I238312,);
nor I_13838 (I238320,I238312,I238255);
DFFARX1 I_13839 (I238320,I3035,I238088,I238053,);
nor I_13840 (I238068,I238312,I238213);
nand I_13841 (I238365,I365468,I365480);
and I_13842 (I238382,I238365,I365489);
DFFARX1 I_13843 (I238382,I3035,I238088,I238408,);
nor I_13844 (I238056,I238408,I238312);
not I_13845 (I238430,I238408);
nor I_13846 (I238447,I238430,I238221);
nor I_13847 (I238464,I238153,I238447);
DFFARX1 I_13848 (I238464,I3035,I238088,I238071,);
nor I_13849 (I238495,I238430,I238312);
nor I_13850 (I238512,I365486,I365480);
nor I_13851 (I238062,I238512,I238495);
not I_13852 (I238543,I238512);
nand I_13853 (I238065,I238272,I238543);
DFFARX1 I_13854 (I238512,I3035,I238088,I238077,);
DFFARX1 I_13855 (I238512,I3035,I238088,I238074,);
not I_13856 (I238632,I3042);
DFFARX1 I_13857 (I702010,I3035,I238632,I238658,);
DFFARX1 I_13858 (I238658,I3035,I238632,I238675,);
not I_13859 (I238624,I238675);
not I_13860 (I238697,I238658);
nand I_13861 (I238714,I701986,I702007);
and I_13862 (I238731,I238714,I702004);
DFFARX1 I_13863 (I238731,I3035,I238632,I238757,);
not I_13864 (I238765,I238757);
DFFARX1 I_13865 (I701983,I3035,I238632,I238791,);
and I_13866 (I238799,I238791,I701995);
nand I_13867 (I238816,I238791,I701995);
nand I_13868 (I238603,I238765,I238816);
DFFARX1 I_13869 (I701998,I3035,I238632,I238856,);
nor I_13870 (I238864,I238856,I238799);
DFFARX1 I_13871 (I238864,I3035,I238632,I238597,);
nor I_13872 (I238612,I238856,I238757);
nand I_13873 (I238909,I702001,I701989);
and I_13874 (I238926,I238909,I701992);
DFFARX1 I_13875 (I238926,I3035,I238632,I238952,);
nor I_13876 (I238600,I238952,I238856);
not I_13877 (I238974,I238952);
nor I_13878 (I238991,I238974,I238765);
nor I_13879 (I239008,I238697,I238991);
DFFARX1 I_13880 (I239008,I3035,I238632,I238615,);
nor I_13881 (I239039,I238974,I238856);
nor I_13882 (I239056,I701983,I701989);
nor I_13883 (I238606,I239056,I239039);
not I_13884 (I239087,I239056);
nand I_13885 (I238609,I238816,I239087);
DFFARX1 I_13886 (I239056,I3035,I238632,I238621,);
DFFARX1 I_13887 (I239056,I3035,I238632,I238618,);
not I_13888 (I239176,I3042);
DFFARX1 I_13889 (I29945,I3035,I239176,I239202,);
DFFARX1 I_13890 (I239202,I3035,I239176,I239219,);
not I_13891 (I239168,I239219);
not I_13892 (I239241,I239202);
nand I_13893 (I239258,I29960,I29939);
and I_13894 (I239275,I239258,I29942);
DFFARX1 I_13895 (I239275,I3035,I239176,I239301,);
not I_13896 (I239309,I239301);
DFFARX1 I_13897 (I29948,I3035,I239176,I239335,);
and I_13898 (I239343,I239335,I29942);
nand I_13899 (I239360,I239335,I29942);
nand I_13900 (I239147,I239309,I239360);
DFFARX1 I_13901 (I29957,I3035,I239176,I239400,);
nor I_13902 (I239408,I239400,I239343);
DFFARX1 I_13903 (I239408,I3035,I239176,I239141,);
nor I_13904 (I239156,I239400,I239301);
nand I_13905 (I239453,I29939,I29954);
and I_13906 (I239470,I239453,I29951);
DFFARX1 I_13907 (I239470,I3035,I239176,I239496,);
nor I_13908 (I239144,I239496,I239400);
not I_13909 (I239518,I239496);
nor I_13910 (I239535,I239518,I239309);
nor I_13911 (I239552,I239241,I239535);
DFFARX1 I_13912 (I239552,I3035,I239176,I239159,);
nor I_13913 (I239583,I239518,I239400);
nor I_13914 (I239600,I29963,I29954);
nor I_13915 (I239150,I239600,I239583);
not I_13916 (I239631,I239600);
nand I_13917 (I239153,I239360,I239631);
DFFARX1 I_13918 (I239600,I3035,I239176,I239165,);
DFFARX1 I_13919 (I239600,I3035,I239176,I239162,);
not I_13920 (I239720,I3042);
DFFARX1 I_13921 (I341773,I3035,I239720,I239746,);
DFFARX1 I_13922 (I239746,I3035,I239720,I239763,);
not I_13923 (I239712,I239763);
not I_13924 (I239785,I239746);
nand I_13925 (I239802,I341794,I341785);
and I_13926 (I239819,I239802,I341773);
DFFARX1 I_13927 (I239819,I3035,I239720,I239845,);
not I_13928 (I239853,I239845);
DFFARX1 I_13929 (I341779,I3035,I239720,I239879,);
and I_13930 (I239887,I239879,I341776);
nand I_13931 (I239904,I239879,I341776);
nand I_13932 (I239691,I239853,I239904);
DFFARX1 I_13933 (I341770,I3035,I239720,I239944,);
nor I_13934 (I239952,I239944,I239887);
DFFARX1 I_13935 (I239952,I3035,I239720,I239685,);
nor I_13936 (I239700,I239944,I239845);
nand I_13937 (I239997,I341770,I341782);
and I_13938 (I240014,I239997,I341791);
DFFARX1 I_13939 (I240014,I3035,I239720,I240040,);
nor I_13940 (I239688,I240040,I239944);
not I_13941 (I240062,I240040);
nor I_13942 (I240079,I240062,I239853);
nor I_13943 (I240096,I239785,I240079);
DFFARX1 I_13944 (I240096,I3035,I239720,I239703,);
nor I_13945 (I240127,I240062,I239944);
nor I_13946 (I240144,I341788,I341782);
nor I_13947 (I239694,I240144,I240127);
not I_13948 (I240175,I240144);
nand I_13949 (I239697,I239904,I240175);
DFFARX1 I_13950 (I240144,I3035,I239720,I239709,);
DFFARX1 I_13951 (I240144,I3035,I239720,I239706,);
not I_13952 (I240264,I3042);
DFFARX1 I_13953 (I496102,I3035,I240264,I240290,);
DFFARX1 I_13954 (I240290,I3035,I240264,I240307,);
not I_13955 (I240256,I240307);
not I_13956 (I240329,I240290);
nand I_13957 (I240346,I496117,I496105);
and I_13958 (I240363,I240346,I496096);
DFFARX1 I_13959 (I240363,I3035,I240264,I240389,);
not I_13960 (I240397,I240389);
DFFARX1 I_13961 (I496108,I3035,I240264,I240423,);
and I_13962 (I240431,I240423,I496099);
nand I_13963 (I240448,I240423,I496099);
nand I_13964 (I240235,I240397,I240448);
DFFARX1 I_13965 (I496114,I3035,I240264,I240488,);
nor I_13966 (I240496,I240488,I240431);
DFFARX1 I_13967 (I240496,I3035,I240264,I240229,);
nor I_13968 (I240244,I240488,I240389);
nand I_13969 (I240541,I496123,I496111);
and I_13970 (I240558,I240541,I496120);
DFFARX1 I_13971 (I240558,I3035,I240264,I240584,);
nor I_13972 (I240232,I240584,I240488);
not I_13973 (I240606,I240584);
nor I_13974 (I240623,I240606,I240397);
nor I_13975 (I240640,I240329,I240623);
DFFARX1 I_13976 (I240640,I3035,I240264,I240247,);
nor I_13977 (I240671,I240606,I240488);
nor I_13978 (I240688,I496096,I496111);
nor I_13979 (I240238,I240688,I240671);
not I_13980 (I240719,I240688);
nand I_13981 (I240241,I240448,I240719);
DFFARX1 I_13982 (I240688,I3035,I240264,I240253,);
DFFARX1 I_13983 (I240688,I3035,I240264,I240250,);
not I_13984 (I240808,I3042);
DFFARX1 I_13985 (I226735,I3035,I240808,I240834,);
DFFARX1 I_13986 (I240834,I3035,I240808,I240851,);
not I_13987 (I240800,I240851);
not I_13988 (I240873,I240834);
nand I_13989 (I240890,I226714,I226738);
and I_13990 (I240907,I240890,I226741);
DFFARX1 I_13991 (I240907,I3035,I240808,I240933,);
not I_13992 (I240941,I240933);
DFFARX1 I_13993 (I226723,I3035,I240808,I240967,);
and I_13994 (I240975,I240967,I226729);
nand I_13995 (I240992,I240967,I226729);
nand I_13996 (I240779,I240941,I240992);
DFFARX1 I_13997 (I226717,I3035,I240808,I241032,);
nor I_13998 (I241040,I241032,I240975);
DFFARX1 I_13999 (I241040,I3035,I240808,I240773,);
nor I_14000 (I240788,I241032,I240933);
nand I_14001 (I241085,I226726,I226714);
and I_14002 (I241102,I241085,I226720);
DFFARX1 I_14003 (I241102,I3035,I240808,I241128,);
nor I_14004 (I240776,I241128,I241032);
not I_14005 (I241150,I241128);
nor I_14006 (I241167,I241150,I240941);
nor I_14007 (I241184,I240873,I241167);
DFFARX1 I_14008 (I241184,I3035,I240808,I240791,);
nor I_14009 (I241215,I241150,I241032);
nor I_14010 (I241232,I226732,I226714);
nor I_14011 (I240782,I241232,I241215);
not I_14012 (I241263,I241232);
nand I_14013 (I240785,I240992,I241263);
DFFARX1 I_14014 (I241232,I3035,I240808,I240797,);
DFFARX1 I_14015 (I241232,I3035,I240808,I240794,);
not I_14016 (I241352,I3042);
DFFARX1 I_14017 (I516128,I3035,I241352,I241378,);
DFFARX1 I_14018 (I241378,I3035,I241352,I241395,);
not I_14019 (I241344,I241395);
not I_14020 (I241417,I241378);
nand I_14021 (I241434,I516143,I516131);
and I_14022 (I241451,I241434,I516122);
DFFARX1 I_14023 (I241451,I3035,I241352,I241477,);
not I_14024 (I241485,I241477);
DFFARX1 I_14025 (I516134,I3035,I241352,I241511,);
and I_14026 (I241519,I241511,I516125);
nand I_14027 (I241536,I241511,I516125);
nand I_14028 (I241323,I241485,I241536);
DFFARX1 I_14029 (I516140,I3035,I241352,I241576,);
nor I_14030 (I241584,I241576,I241519);
DFFARX1 I_14031 (I241584,I3035,I241352,I241317,);
nor I_14032 (I241332,I241576,I241477);
nand I_14033 (I241629,I516149,I516137);
and I_14034 (I241646,I241629,I516146);
DFFARX1 I_14035 (I241646,I3035,I241352,I241672,);
nor I_14036 (I241320,I241672,I241576);
not I_14037 (I241694,I241672);
nor I_14038 (I241711,I241694,I241485);
nor I_14039 (I241728,I241417,I241711);
DFFARX1 I_14040 (I241728,I3035,I241352,I241335,);
nor I_14041 (I241759,I241694,I241576);
nor I_14042 (I241776,I516122,I516137);
nor I_14043 (I241326,I241776,I241759);
not I_14044 (I241807,I241776);
nand I_14045 (I241329,I241536,I241807);
DFFARX1 I_14046 (I241776,I3035,I241352,I241341,);
DFFARX1 I_14047 (I241776,I3035,I241352,I241338,);
not I_14048 (I241896,I3042);
DFFARX1 I_14049 (I683488,I3035,I241896,I241922,);
DFFARX1 I_14050 (I241922,I3035,I241896,I241939,);
not I_14051 (I241888,I241939);
not I_14052 (I241961,I241922);
nand I_14053 (I241978,I683485,I683482);
and I_14054 (I241995,I241978,I683470);
DFFARX1 I_14055 (I241995,I3035,I241896,I242021,);
not I_14056 (I242029,I242021);
DFFARX1 I_14057 (I683494,I3035,I241896,I242055,);
and I_14058 (I242063,I242055,I683479);
nand I_14059 (I242080,I242055,I683479);
nand I_14060 (I241867,I242029,I242080);
DFFARX1 I_14061 (I683473,I3035,I241896,I242120,);
nor I_14062 (I242128,I242120,I242063);
DFFARX1 I_14063 (I242128,I3035,I241896,I241861,);
nor I_14064 (I241876,I242120,I242021);
nand I_14065 (I242173,I683470,I683476);
and I_14066 (I242190,I242173,I683491);
DFFARX1 I_14067 (I242190,I3035,I241896,I242216,);
nor I_14068 (I241864,I242216,I242120);
not I_14069 (I242238,I242216);
nor I_14070 (I242255,I242238,I242029);
nor I_14071 (I242272,I241961,I242255);
DFFARX1 I_14072 (I242272,I3035,I241896,I241879,);
nor I_14073 (I242303,I242238,I242120);
nor I_14074 (I242320,I683473,I683476);
nor I_14075 (I241870,I242320,I242303);
not I_14076 (I242351,I242320);
nand I_14077 (I241873,I242080,I242351);
DFFARX1 I_14078 (I242320,I3035,I241896,I241885,);
DFFARX1 I_14079 (I242320,I3035,I241896,I241882,);
not I_14080 (I242440,I3042);
DFFARX1 I_14081 (I91998,I3035,I242440,I242466,);
DFFARX1 I_14082 (I242466,I3035,I242440,I242483,);
not I_14083 (I242432,I242483);
not I_14084 (I242505,I242466);
nand I_14085 (I242522,I92010,I91989);
and I_14086 (I242539,I242522,I91992);
DFFARX1 I_14087 (I242539,I3035,I242440,I242565,);
not I_14088 (I242573,I242565);
DFFARX1 I_14089 (I92001,I3035,I242440,I242599,);
and I_14090 (I242607,I242599,I92013);
nand I_14091 (I242624,I242599,I92013);
nand I_14092 (I242411,I242573,I242624);
DFFARX1 I_14093 (I92007,I3035,I242440,I242664,);
nor I_14094 (I242672,I242664,I242607);
DFFARX1 I_14095 (I242672,I3035,I242440,I242405,);
nor I_14096 (I242420,I242664,I242565);
nand I_14097 (I242717,I91995,I91992);
and I_14098 (I242734,I242717,I92004);
DFFARX1 I_14099 (I242734,I3035,I242440,I242760,);
nor I_14100 (I242408,I242760,I242664);
not I_14101 (I242782,I242760);
nor I_14102 (I242799,I242782,I242573);
nor I_14103 (I242816,I242505,I242799);
DFFARX1 I_14104 (I242816,I3035,I242440,I242423,);
nor I_14105 (I242847,I242782,I242664);
nor I_14106 (I242864,I91989,I91992);
nor I_14107 (I242414,I242864,I242847);
not I_14108 (I242895,I242864);
nand I_14109 (I242417,I242624,I242895);
DFFARX1 I_14110 (I242864,I3035,I242440,I242429,);
DFFARX1 I_14111 (I242864,I3035,I242440,I242426,);
not I_14112 (I242984,I3042);
DFFARX1 I_14113 (I2396,I3035,I242984,I243010,);
DFFARX1 I_14114 (I243010,I3035,I242984,I243027,);
not I_14115 (I242976,I243027);
not I_14116 (I243049,I243010);
nand I_14117 (I243066,I1380,I2540);
and I_14118 (I243083,I243066,I1748);
DFFARX1 I_14119 (I243083,I3035,I242984,I243109,);
not I_14120 (I243117,I243109);
DFFARX1 I_14121 (I2812,I3035,I242984,I243143,);
and I_14122 (I243151,I243143,I2388);
nand I_14123 (I243168,I243143,I2388);
nand I_14124 (I242955,I243117,I243168);
DFFARX1 I_14125 (I2644,I3035,I242984,I243208,);
nor I_14126 (I243216,I243208,I243151);
DFFARX1 I_14127 (I243216,I3035,I242984,I242949,);
nor I_14128 (I242964,I243208,I243109);
nand I_14129 (I243261,I2972,I2052);
and I_14130 (I243278,I243261,I3012);
DFFARX1 I_14131 (I243278,I3035,I242984,I243304,);
nor I_14132 (I242952,I243304,I243208);
not I_14133 (I243326,I243304);
nor I_14134 (I243343,I243326,I243117);
nor I_14135 (I243360,I243049,I243343);
DFFARX1 I_14136 (I243360,I3035,I242984,I242967,);
nor I_14137 (I243391,I243326,I243208);
nor I_14138 (I243408,I2036,I2052);
nor I_14139 (I242958,I243408,I243391);
not I_14140 (I243439,I243408);
nand I_14141 (I242961,I243168,I243439);
DFFARX1 I_14142 (I243408,I3035,I242984,I242973,);
DFFARX1 I_14143 (I243408,I3035,I242984,I242970,);
not I_14144 (I243528,I3042);
DFFARX1 I_14145 (I65781,I3035,I243528,I243554,);
DFFARX1 I_14146 (I243554,I3035,I243528,I243571,);
not I_14147 (I243520,I243571);
not I_14148 (I243593,I243554);
nand I_14149 (I243610,I65796,I65775);
and I_14150 (I243627,I243610,I65778);
DFFARX1 I_14151 (I243627,I3035,I243528,I243653,);
not I_14152 (I243661,I243653);
DFFARX1 I_14153 (I65784,I3035,I243528,I243687,);
and I_14154 (I243695,I243687,I65778);
nand I_14155 (I243712,I243687,I65778);
nand I_14156 (I243499,I243661,I243712);
DFFARX1 I_14157 (I65793,I3035,I243528,I243752,);
nor I_14158 (I243760,I243752,I243695);
DFFARX1 I_14159 (I243760,I3035,I243528,I243493,);
nor I_14160 (I243508,I243752,I243653);
nand I_14161 (I243805,I65775,I65790);
and I_14162 (I243822,I243805,I65787);
DFFARX1 I_14163 (I243822,I3035,I243528,I243848,);
nor I_14164 (I243496,I243848,I243752);
not I_14165 (I243870,I243848);
nor I_14166 (I243887,I243870,I243661);
nor I_14167 (I243904,I243593,I243887);
DFFARX1 I_14168 (I243904,I3035,I243528,I243511,);
nor I_14169 (I243935,I243870,I243752);
nor I_14170 (I243952,I65799,I65790);
nor I_14171 (I243502,I243952,I243935);
not I_14172 (I243983,I243952);
nand I_14173 (I243505,I243712,I243983);
DFFARX1 I_14174 (I243952,I3035,I243528,I243517,);
DFFARX1 I_14175 (I243952,I3035,I243528,I243514,);
not I_14176 (I244072,I3042);
DFFARX1 I_14177 (I582697,I3035,I244072,I244098,);
DFFARX1 I_14178 (I244098,I3035,I244072,I244115,);
not I_14179 (I244064,I244115);
not I_14180 (I244137,I244098);
nand I_14181 (I244154,I582709,I582697);
and I_14182 (I244171,I244154,I582700);
DFFARX1 I_14183 (I244171,I3035,I244072,I244197,);
not I_14184 (I244205,I244197);
DFFARX1 I_14185 (I582718,I3035,I244072,I244231,);
and I_14186 (I244239,I244231,I582694);
nand I_14187 (I244256,I244231,I582694);
nand I_14188 (I244043,I244205,I244256);
DFFARX1 I_14189 (I582712,I3035,I244072,I244296,);
nor I_14190 (I244304,I244296,I244239);
DFFARX1 I_14191 (I244304,I3035,I244072,I244037,);
nor I_14192 (I244052,I244296,I244197);
nand I_14193 (I244349,I582706,I582703);
and I_14194 (I244366,I244349,I582715);
DFFARX1 I_14195 (I244366,I3035,I244072,I244392,);
nor I_14196 (I244040,I244392,I244296);
not I_14197 (I244414,I244392);
nor I_14198 (I244431,I244414,I244205);
nor I_14199 (I244448,I244137,I244431);
DFFARX1 I_14200 (I244448,I3035,I244072,I244055,);
nor I_14201 (I244479,I244414,I244296);
nor I_14202 (I244496,I582694,I582703);
nor I_14203 (I244046,I244496,I244479);
not I_14204 (I244527,I244496);
nand I_14205 (I244049,I244256,I244527);
DFFARX1 I_14206 (I244496,I3035,I244072,I244061,);
DFFARX1 I_14207 (I244496,I3035,I244072,I244058,);
not I_14208 (I244616,I3042);
DFFARX1 I_14209 (I607551,I3035,I244616,I244642,);
DFFARX1 I_14210 (I244642,I3035,I244616,I244659,);
not I_14211 (I244608,I244659);
not I_14212 (I244681,I244642);
nand I_14213 (I244698,I607563,I607551);
and I_14214 (I244715,I244698,I607554);
DFFARX1 I_14215 (I244715,I3035,I244616,I244741,);
not I_14216 (I244749,I244741);
DFFARX1 I_14217 (I607572,I3035,I244616,I244775,);
and I_14218 (I244783,I244775,I607548);
nand I_14219 (I244800,I244775,I607548);
nand I_14220 (I244587,I244749,I244800);
DFFARX1 I_14221 (I607566,I3035,I244616,I244840,);
nor I_14222 (I244848,I244840,I244783);
DFFARX1 I_14223 (I244848,I3035,I244616,I244581,);
nor I_14224 (I244596,I244840,I244741);
nand I_14225 (I244893,I607560,I607557);
and I_14226 (I244910,I244893,I607569);
DFFARX1 I_14227 (I244910,I3035,I244616,I244936,);
nor I_14228 (I244584,I244936,I244840);
not I_14229 (I244958,I244936);
nor I_14230 (I244975,I244958,I244749);
nor I_14231 (I244992,I244681,I244975);
DFFARX1 I_14232 (I244992,I3035,I244616,I244599,);
nor I_14233 (I245023,I244958,I244840);
nor I_14234 (I245040,I607548,I607557);
nor I_14235 (I244590,I245040,I245023);
not I_14236 (I245071,I245040);
nand I_14237 (I244593,I244800,I245071);
DFFARX1 I_14238 (I245040,I3035,I244616,I244605,);
DFFARX1 I_14239 (I245040,I3035,I244616,I244602,);
not I_14240 (I245160,I3042);
DFFARX1 I_14241 (I676552,I3035,I245160,I245186,);
DFFARX1 I_14242 (I245186,I3035,I245160,I245203,);
not I_14243 (I245152,I245203);
not I_14244 (I245225,I245186);
nand I_14245 (I245242,I676549,I676546);
and I_14246 (I245259,I245242,I676534);
DFFARX1 I_14247 (I245259,I3035,I245160,I245285,);
not I_14248 (I245293,I245285);
DFFARX1 I_14249 (I676558,I3035,I245160,I245319,);
and I_14250 (I245327,I245319,I676543);
nand I_14251 (I245344,I245319,I676543);
nand I_14252 (I245131,I245293,I245344);
DFFARX1 I_14253 (I676537,I3035,I245160,I245384,);
nor I_14254 (I245392,I245384,I245327);
DFFARX1 I_14255 (I245392,I3035,I245160,I245125,);
nor I_14256 (I245140,I245384,I245285);
nand I_14257 (I245437,I676534,I676540);
and I_14258 (I245454,I245437,I676555);
DFFARX1 I_14259 (I245454,I3035,I245160,I245480,);
nor I_14260 (I245128,I245480,I245384);
not I_14261 (I245502,I245480);
nor I_14262 (I245519,I245502,I245293);
nor I_14263 (I245536,I245225,I245519);
DFFARX1 I_14264 (I245536,I3035,I245160,I245143,);
nor I_14265 (I245567,I245502,I245384);
nor I_14266 (I245584,I676537,I676540);
nor I_14267 (I245134,I245584,I245567);
not I_14268 (I245615,I245584);
nand I_14269 (I245137,I245344,I245615);
DFFARX1 I_14270 (I245584,I3035,I245160,I245149,);
DFFARX1 I_14271 (I245584,I3035,I245160,I245146,);
not I_14272 (I245704,I3042);
DFFARX1 I_14273 (I337727,I3035,I245704,I245730,);
DFFARX1 I_14274 (I245730,I3035,I245704,I245747,);
not I_14275 (I245696,I245747);
not I_14276 (I245769,I245730);
nand I_14277 (I245786,I337724,I337745);
and I_14278 (I245803,I245786,I337748);
DFFARX1 I_14279 (I245803,I3035,I245704,I245829,);
not I_14280 (I245837,I245829);
DFFARX1 I_14281 (I337733,I3035,I245704,I245863,);
and I_14282 (I245871,I245863,I337736);
nand I_14283 (I245888,I245863,I337736);
nand I_14284 (I245675,I245837,I245888);
DFFARX1 I_14285 (I337739,I3035,I245704,I245928,);
nor I_14286 (I245936,I245928,I245871);
DFFARX1 I_14287 (I245936,I3035,I245704,I245669,);
nor I_14288 (I245684,I245928,I245829);
nand I_14289 (I245981,I337724,I337730);
and I_14290 (I245998,I245981,I337742);
DFFARX1 I_14291 (I245998,I3035,I245704,I246024,);
nor I_14292 (I245672,I246024,I245928);
not I_14293 (I246046,I246024);
nor I_14294 (I246063,I246046,I245837);
nor I_14295 (I246080,I245769,I246063);
DFFARX1 I_14296 (I246080,I3035,I245704,I245687,);
nor I_14297 (I246111,I246046,I245928);
nor I_14298 (I246128,I337727,I337730);
nor I_14299 (I245678,I246128,I246111);
not I_14300 (I246159,I246128);
nand I_14301 (I245681,I245888,I246159);
DFFARX1 I_14302 (I246128,I3035,I245704,I245693,);
DFFARX1 I_14303 (I246128,I3035,I245704,I245690,);
not I_14304 (I246248,I3042);
DFFARX1 I_14305 (I147333,I3035,I246248,I246274,);
DFFARX1 I_14306 (I246274,I3035,I246248,I246291,);
not I_14307 (I246240,I246291);
not I_14308 (I246313,I246274);
nand I_14309 (I246330,I147345,I147324);
and I_14310 (I246347,I246330,I147327);
DFFARX1 I_14311 (I246347,I3035,I246248,I246373,);
not I_14312 (I246381,I246373);
DFFARX1 I_14313 (I147336,I3035,I246248,I246407,);
and I_14314 (I246415,I246407,I147348);
nand I_14315 (I246432,I246407,I147348);
nand I_14316 (I246219,I246381,I246432);
DFFARX1 I_14317 (I147342,I3035,I246248,I246472,);
nor I_14318 (I246480,I246472,I246415);
DFFARX1 I_14319 (I246480,I3035,I246248,I246213,);
nor I_14320 (I246228,I246472,I246373);
nand I_14321 (I246525,I147330,I147327);
and I_14322 (I246542,I246525,I147339);
DFFARX1 I_14323 (I246542,I3035,I246248,I246568,);
nor I_14324 (I246216,I246568,I246472);
not I_14325 (I246590,I246568);
nor I_14326 (I246607,I246590,I246381);
nor I_14327 (I246624,I246313,I246607);
DFFARX1 I_14328 (I246624,I3035,I246248,I246231,);
nor I_14329 (I246655,I246590,I246472);
nor I_14330 (I246672,I147324,I147327);
nor I_14331 (I246222,I246672,I246655);
not I_14332 (I246703,I246672);
nand I_14333 (I246225,I246432,I246703);
DFFARX1 I_14334 (I246672,I3035,I246248,I246237,);
DFFARX1 I_14335 (I246672,I3035,I246248,I246234,);
not I_14336 (I246792,I3042);
DFFARX1 I_14337 (I353911,I3035,I246792,I246818,);
DFFARX1 I_14338 (I246818,I3035,I246792,I246835,);
not I_14339 (I246784,I246835);
not I_14340 (I246857,I246818);
nand I_14341 (I246874,I353932,I353923);
and I_14342 (I246891,I246874,I353911);
DFFARX1 I_14343 (I246891,I3035,I246792,I246917,);
not I_14344 (I246925,I246917);
DFFARX1 I_14345 (I353917,I3035,I246792,I246951,);
and I_14346 (I246959,I246951,I353914);
nand I_14347 (I246976,I246951,I353914);
nand I_14348 (I246763,I246925,I246976);
DFFARX1 I_14349 (I353908,I3035,I246792,I247016,);
nor I_14350 (I247024,I247016,I246959);
DFFARX1 I_14351 (I247024,I3035,I246792,I246757,);
nor I_14352 (I246772,I247016,I246917);
nand I_14353 (I247069,I353908,I353920);
and I_14354 (I247086,I247069,I353929);
DFFARX1 I_14355 (I247086,I3035,I246792,I247112,);
nor I_14356 (I246760,I247112,I247016);
not I_14357 (I247134,I247112);
nor I_14358 (I247151,I247134,I246925);
nor I_14359 (I247168,I246857,I247151);
DFFARX1 I_14360 (I247168,I3035,I246792,I246775,);
nor I_14361 (I247199,I247134,I247016);
nor I_14362 (I247216,I353926,I353920);
nor I_14363 (I246766,I247216,I247199);
not I_14364 (I247247,I247216);
nand I_14365 (I246769,I246976,I247247);
DFFARX1 I_14366 (I247216,I3035,I246792,I246781,);
DFFARX1 I_14367 (I247216,I3035,I246792,I246778,);
not I_14368 (I247336,I3042);
DFFARX1 I_14369 (I154009,I3035,I247336,I247362,);
DFFARX1 I_14370 (I247362,I3035,I247336,I247379,);
not I_14371 (I247328,I247379);
not I_14372 (I247401,I247362);
nand I_14373 (I247418,I153988,I154012);
and I_14374 (I247435,I247418,I154015);
DFFARX1 I_14375 (I247435,I3035,I247336,I247461,);
not I_14376 (I247469,I247461);
DFFARX1 I_14377 (I153997,I3035,I247336,I247495,);
and I_14378 (I247503,I247495,I154003);
nand I_14379 (I247520,I247495,I154003);
nand I_14380 (I247307,I247469,I247520);
DFFARX1 I_14381 (I153991,I3035,I247336,I247560,);
nor I_14382 (I247568,I247560,I247503);
DFFARX1 I_14383 (I247568,I3035,I247336,I247301,);
nor I_14384 (I247316,I247560,I247461);
nand I_14385 (I247613,I154000,I153988);
and I_14386 (I247630,I247613,I153994);
DFFARX1 I_14387 (I247630,I3035,I247336,I247656,);
nor I_14388 (I247304,I247656,I247560);
not I_14389 (I247678,I247656);
nor I_14390 (I247695,I247678,I247469);
nor I_14391 (I247712,I247401,I247695);
DFFARX1 I_14392 (I247712,I3035,I247336,I247319,);
nor I_14393 (I247743,I247678,I247560);
nor I_14394 (I247760,I154006,I153988);
nor I_14395 (I247310,I247760,I247743);
not I_14396 (I247791,I247760);
nand I_14397 (I247313,I247520,I247791);
DFFARX1 I_14398 (I247760,I3035,I247336,I247325,);
DFFARX1 I_14399 (I247760,I3035,I247336,I247322,);
not I_14400 (I247880,I3042);
DFFARX1 I_14401 (I320387,I3035,I247880,I247906,);
DFFARX1 I_14402 (I247906,I3035,I247880,I247923,);
not I_14403 (I247872,I247923);
not I_14404 (I247945,I247906);
nand I_14405 (I247962,I320384,I320405);
and I_14406 (I247979,I247962,I320408);
DFFARX1 I_14407 (I247979,I3035,I247880,I248005,);
not I_14408 (I248013,I248005);
DFFARX1 I_14409 (I320393,I3035,I247880,I248039,);
and I_14410 (I248047,I248039,I320396);
nand I_14411 (I248064,I248039,I320396);
nand I_14412 (I247851,I248013,I248064);
DFFARX1 I_14413 (I320399,I3035,I247880,I248104,);
nor I_14414 (I248112,I248104,I248047);
DFFARX1 I_14415 (I248112,I3035,I247880,I247845,);
nor I_14416 (I247860,I248104,I248005);
nand I_14417 (I248157,I320384,I320390);
and I_14418 (I248174,I248157,I320402);
DFFARX1 I_14419 (I248174,I3035,I247880,I248200,);
nor I_14420 (I247848,I248200,I248104);
not I_14421 (I248222,I248200);
nor I_14422 (I248239,I248222,I248013);
nor I_14423 (I248256,I247945,I248239);
DFFARX1 I_14424 (I248256,I3035,I247880,I247863,);
nor I_14425 (I248287,I248222,I248104);
nor I_14426 (I248304,I320387,I320390);
nor I_14427 (I247854,I248304,I248287);
not I_14428 (I248335,I248304);
nand I_14429 (I247857,I248064,I248335);
DFFARX1 I_14430 (I248304,I3035,I247880,I247869,);
DFFARX1 I_14431 (I248304,I3035,I247880,I247866,);
not I_14432 (I248424,I3042);
DFFARX1 I_14433 (I137218,I3035,I248424,I248450,);
DFFARX1 I_14434 (I248450,I3035,I248424,I248467,);
not I_14435 (I248416,I248467);
not I_14436 (I248489,I248450);
nand I_14437 (I248506,I137230,I137209);
and I_14438 (I248523,I248506,I137212);
DFFARX1 I_14439 (I248523,I3035,I248424,I248549,);
not I_14440 (I248557,I248549);
DFFARX1 I_14441 (I137221,I3035,I248424,I248583,);
and I_14442 (I248591,I248583,I137233);
nand I_14443 (I248608,I248583,I137233);
nand I_14444 (I248395,I248557,I248608);
DFFARX1 I_14445 (I137227,I3035,I248424,I248648,);
nor I_14446 (I248656,I248648,I248591);
DFFARX1 I_14447 (I248656,I3035,I248424,I248389,);
nor I_14448 (I248404,I248648,I248549);
nand I_14449 (I248701,I137215,I137212);
and I_14450 (I248718,I248701,I137224);
DFFARX1 I_14451 (I248718,I3035,I248424,I248744,);
nor I_14452 (I248392,I248744,I248648);
not I_14453 (I248766,I248744);
nor I_14454 (I248783,I248766,I248557);
nor I_14455 (I248800,I248489,I248783);
DFFARX1 I_14456 (I248800,I3035,I248424,I248407,);
nor I_14457 (I248831,I248766,I248648);
nor I_14458 (I248848,I137209,I137212);
nor I_14459 (I248398,I248848,I248831);
not I_14460 (I248879,I248848);
nand I_14461 (I248401,I248608,I248879);
DFFARX1 I_14462 (I248848,I3035,I248424,I248413,);
DFFARX1 I_14463 (I248848,I3035,I248424,I248410,);
not I_14464 (I248968,I3042);
DFFARX1 I_14465 (I600615,I3035,I248968,I248994,);
DFFARX1 I_14466 (I248994,I3035,I248968,I249011,);
not I_14467 (I248960,I249011);
not I_14468 (I249033,I248994);
nand I_14469 (I249050,I600627,I600615);
and I_14470 (I249067,I249050,I600618);
DFFARX1 I_14471 (I249067,I3035,I248968,I249093,);
not I_14472 (I249101,I249093);
DFFARX1 I_14473 (I600636,I3035,I248968,I249127,);
and I_14474 (I249135,I249127,I600612);
nand I_14475 (I249152,I249127,I600612);
nand I_14476 (I248939,I249101,I249152);
DFFARX1 I_14477 (I600630,I3035,I248968,I249192,);
nor I_14478 (I249200,I249192,I249135);
DFFARX1 I_14479 (I249200,I3035,I248968,I248933,);
nor I_14480 (I248948,I249192,I249093);
nand I_14481 (I249245,I600624,I600621);
and I_14482 (I249262,I249245,I600633);
DFFARX1 I_14483 (I249262,I3035,I248968,I249288,);
nor I_14484 (I248936,I249288,I249192);
not I_14485 (I249310,I249288);
nor I_14486 (I249327,I249310,I249101);
nor I_14487 (I249344,I249033,I249327);
DFFARX1 I_14488 (I249344,I3035,I248968,I248951,);
nor I_14489 (I249375,I249310,I249192);
nor I_14490 (I249392,I600612,I600621);
nor I_14491 (I248942,I249392,I249375);
not I_14492 (I249423,I249392);
nand I_14493 (I248945,I249152,I249423);
DFFARX1 I_14494 (I249392,I3035,I248968,I248957,);
DFFARX1 I_14495 (I249392,I3035,I248968,I248954,);
not I_14496 (I249512,I3042);
DFFARX1 I_14497 (I561070,I3035,I249512,I249538,);
DFFARX1 I_14498 (I249538,I3035,I249512,I249555,);
not I_14499 (I249504,I249555);
not I_14500 (I249577,I249538);
nand I_14501 (I249594,I561070,I561088);
and I_14502 (I249611,I249594,I561082);
DFFARX1 I_14503 (I249611,I3035,I249512,I249637,);
not I_14504 (I249645,I249637);
DFFARX1 I_14505 (I561076,I3035,I249512,I249671,);
and I_14506 (I249679,I249671,I561085);
nand I_14507 (I249696,I249671,I561085);
nand I_14508 (I249483,I249645,I249696);
DFFARX1 I_14509 (I561073,I3035,I249512,I249736,);
nor I_14510 (I249744,I249736,I249679);
DFFARX1 I_14511 (I249744,I3035,I249512,I249477,);
nor I_14512 (I249492,I249736,I249637);
nand I_14513 (I249789,I561073,I561091);
and I_14514 (I249806,I249789,I561076);
DFFARX1 I_14515 (I249806,I3035,I249512,I249832,);
nor I_14516 (I249480,I249832,I249736);
not I_14517 (I249854,I249832);
nor I_14518 (I249871,I249854,I249645);
nor I_14519 (I249888,I249577,I249871);
DFFARX1 I_14520 (I249888,I3035,I249512,I249495,);
nor I_14521 (I249919,I249854,I249736);
nor I_14522 (I249936,I561079,I561091);
nor I_14523 (I249486,I249936,I249919);
not I_14524 (I249967,I249936);
nand I_14525 (I249489,I249696,I249967);
DFFARX1 I_14526 (I249936,I3035,I249512,I249501,);
DFFARX1 I_14527 (I249936,I3035,I249512,I249498,);
not I_14528 (I250056,I3042);
DFFARX1 I_14529 (I643387,I3035,I250056,I250082,);
DFFARX1 I_14530 (I250082,I3035,I250056,I250099,);
not I_14531 (I250048,I250099);
not I_14532 (I250121,I250082);
nand I_14533 (I250138,I643399,I643387);
and I_14534 (I250155,I250138,I643390);
DFFARX1 I_14535 (I250155,I3035,I250056,I250181,);
not I_14536 (I250189,I250181);
DFFARX1 I_14537 (I643408,I3035,I250056,I250215,);
and I_14538 (I250223,I250215,I643384);
nand I_14539 (I250240,I250215,I643384);
nand I_14540 (I250027,I250189,I250240);
DFFARX1 I_14541 (I643402,I3035,I250056,I250280,);
nor I_14542 (I250288,I250280,I250223);
DFFARX1 I_14543 (I250288,I3035,I250056,I250021,);
nor I_14544 (I250036,I250280,I250181);
nand I_14545 (I250333,I643396,I643393);
and I_14546 (I250350,I250333,I643405);
DFFARX1 I_14547 (I250350,I3035,I250056,I250376,);
nor I_14548 (I250024,I250376,I250280);
not I_14549 (I250398,I250376);
nor I_14550 (I250415,I250398,I250189);
nor I_14551 (I250432,I250121,I250415);
DFFARX1 I_14552 (I250432,I3035,I250056,I250039,);
nor I_14553 (I250463,I250398,I250280);
nor I_14554 (I250480,I643384,I643393);
nor I_14555 (I250030,I250480,I250463);
not I_14556 (I250511,I250480);
nand I_14557 (I250033,I250240,I250511);
DFFARX1 I_14558 (I250480,I3035,I250056,I250045,);
DFFARX1 I_14559 (I250480,I3035,I250056,I250042,);
not I_14560 (I250600,I3042);
DFFARX1 I_14561 (I713910,I3035,I250600,I250626,);
DFFARX1 I_14562 (I250626,I3035,I250600,I250643,);
not I_14563 (I250592,I250643);
not I_14564 (I250665,I250626);
nand I_14565 (I250682,I713886,I713907);
and I_14566 (I250699,I250682,I713904);
DFFARX1 I_14567 (I250699,I3035,I250600,I250725,);
not I_14568 (I250733,I250725);
DFFARX1 I_14569 (I713883,I3035,I250600,I250759,);
and I_14570 (I250767,I250759,I713895);
nand I_14571 (I250784,I250759,I713895);
nand I_14572 (I250571,I250733,I250784);
DFFARX1 I_14573 (I713898,I3035,I250600,I250824,);
nor I_14574 (I250832,I250824,I250767);
DFFARX1 I_14575 (I250832,I3035,I250600,I250565,);
nor I_14576 (I250580,I250824,I250725);
nand I_14577 (I250877,I713901,I713889);
and I_14578 (I250894,I250877,I713892);
DFFARX1 I_14579 (I250894,I3035,I250600,I250920,);
nor I_14580 (I250568,I250920,I250824);
not I_14581 (I250942,I250920);
nor I_14582 (I250959,I250942,I250733);
nor I_14583 (I250976,I250665,I250959);
DFFARX1 I_14584 (I250976,I3035,I250600,I250583,);
nor I_14585 (I251007,I250942,I250824);
nor I_14586 (I251024,I713883,I713889);
nor I_14587 (I250574,I251024,I251007);
not I_14588 (I251055,I251024);
nand I_14589 (I250577,I250784,I251055);
DFFARX1 I_14590 (I251024,I3035,I250600,I250589,);
DFFARX1 I_14591 (I251024,I3035,I250600,I250586,);
not I_14592 (I251144,I3042);
DFFARX1 I_14593 (I7228,I3035,I251144,I251170,);
DFFARX1 I_14594 (I251170,I3035,I251144,I251187,);
not I_14595 (I251136,I251187);
not I_14596 (I251209,I251170);
nand I_14597 (I251226,I7231,I7219);
and I_14598 (I251243,I251226,I7225);
DFFARX1 I_14599 (I251243,I3035,I251144,I251269,);
not I_14600 (I251277,I251269);
DFFARX1 I_14601 (I7213,I3035,I251144,I251303,);
and I_14602 (I251311,I251303,I7210);
nand I_14603 (I251328,I251303,I7210);
nand I_14604 (I251115,I251277,I251328);
DFFARX1 I_14605 (I7216,I3035,I251144,I251368,);
nor I_14606 (I251376,I251368,I251311);
DFFARX1 I_14607 (I251376,I3035,I251144,I251109,);
nor I_14608 (I251124,I251368,I251269);
nand I_14609 (I251421,I7216,I7213);
and I_14610 (I251438,I251421,I7210);
DFFARX1 I_14611 (I251438,I3035,I251144,I251464,);
nor I_14612 (I251112,I251464,I251368);
not I_14613 (I251486,I251464);
nor I_14614 (I251503,I251486,I251277);
nor I_14615 (I251520,I251209,I251503);
DFFARX1 I_14616 (I251520,I3035,I251144,I251127,);
nor I_14617 (I251551,I251486,I251368);
nor I_14618 (I251568,I7222,I7213);
nor I_14619 (I251118,I251568,I251551);
not I_14620 (I251599,I251568);
nand I_14621 (I251121,I251328,I251599);
DFFARX1 I_14622 (I251568,I3035,I251144,I251133,);
DFFARX1 I_14623 (I251568,I3035,I251144,I251130,);
not I_14624 (I251688,I3042);
DFFARX1 I_14625 (I158752,I3035,I251688,I251714,);
DFFARX1 I_14626 (I251714,I3035,I251688,I251731,);
not I_14627 (I251680,I251731);
not I_14628 (I251753,I251714);
nand I_14629 (I251770,I158731,I158755);
and I_14630 (I251787,I251770,I158758);
DFFARX1 I_14631 (I251787,I3035,I251688,I251813,);
not I_14632 (I251821,I251813);
DFFARX1 I_14633 (I158740,I3035,I251688,I251847,);
and I_14634 (I251855,I251847,I158746);
nand I_14635 (I251872,I251847,I158746);
nand I_14636 (I251659,I251821,I251872);
DFFARX1 I_14637 (I158734,I3035,I251688,I251912,);
nor I_14638 (I251920,I251912,I251855);
DFFARX1 I_14639 (I251920,I3035,I251688,I251653,);
nor I_14640 (I251668,I251912,I251813);
nand I_14641 (I251965,I158743,I158731);
and I_14642 (I251982,I251965,I158737);
DFFARX1 I_14643 (I251982,I3035,I251688,I252008,);
nor I_14644 (I251656,I252008,I251912);
not I_14645 (I252030,I252008);
nor I_14646 (I252047,I252030,I251821);
nor I_14647 (I252064,I251753,I252047);
DFFARX1 I_14648 (I252064,I3035,I251688,I251671,);
nor I_14649 (I252095,I252030,I251912);
nor I_14650 (I252112,I158749,I158731);
nor I_14651 (I251662,I252112,I252095);
not I_14652 (I252143,I252112);
nand I_14653 (I251665,I251872,I252143);
DFFARX1 I_14654 (I252112,I3035,I251688,I251677,);
DFFARX1 I_14655 (I252112,I3035,I251688,I251674,);
not I_14656 (I252232,I3042);
DFFARX1 I_14657 (I685222,I3035,I252232,I252258,);
DFFARX1 I_14658 (I252258,I3035,I252232,I252275,);
not I_14659 (I252224,I252275);
not I_14660 (I252297,I252258);
nand I_14661 (I252314,I685219,I685216);
and I_14662 (I252331,I252314,I685204);
DFFARX1 I_14663 (I252331,I3035,I252232,I252357,);
not I_14664 (I252365,I252357);
DFFARX1 I_14665 (I685228,I3035,I252232,I252391,);
and I_14666 (I252399,I252391,I685213);
nand I_14667 (I252416,I252391,I685213);
nand I_14668 (I252203,I252365,I252416);
DFFARX1 I_14669 (I685207,I3035,I252232,I252456,);
nor I_14670 (I252464,I252456,I252399);
DFFARX1 I_14671 (I252464,I3035,I252232,I252197,);
nor I_14672 (I252212,I252456,I252357);
nand I_14673 (I252509,I685204,I685210);
and I_14674 (I252526,I252509,I685225);
DFFARX1 I_14675 (I252526,I3035,I252232,I252552,);
nor I_14676 (I252200,I252552,I252456);
not I_14677 (I252574,I252552);
nor I_14678 (I252591,I252574,I252365);
nor I_14679 (I252608,I252297,I252591);
DFFARX1 I_14680 (I252608,I3035,I252232,I252215,);
nor I_14681 (I252639,I252574,I252456);
nor I_14682 (I252656,I685207,I685210);
nor I_14683 (I252206,I252656,I252639);
not I_14684 (I252687,I252656);
nand I_14685 (I252209,I252416,I252687);
DFFARX1 I_14686 (I252656,I3035,I252232,I252221,);
DFFARX1 I_14687 (I252656,I3035,I252232,I252218,);
not I_14688 (I252776,I3042);
DFFARX1 I_14689 (I132458,I3035,I252776,I252802,);
DFFARX1 I_14690 (I252802,I3035,I252776,I252819,);
not I_14691 (I252768,I252819);
not I_14692 (I252841,I252802);
nand I_14693 (I252858,I132470,I132449);
and I_14694 (I252875,I252858,I132452);
DFFARX1 I_14695 (I252875,I3035,I252776,I252901,);
not I_14696 (I252909,I252901);
DFFARX1 I_14697 (I132461,I3035,I252776,I252935,);
and I_14698 (I252943,I252935,I132473);
nand I_14699 (I252960,I252935,I132473);
nand I_14700 (I252747,I252909,I252960);
DFFARX1 I_14701 (I132467,I3035,I252776,I253000,);
nor I_14702 (I253008,I253000,I252943);
DFFARX1 I_14703 (I253008,I3035,I252776,I252741,);
nor I_14704 (I252756,I253000,I252901);
nand I_14705 (I253053,I132455,I132452);
and I_14706 (I253070,I253053,I132464);
DFFARX1 I_14707 (I253070,I3035,I252776,I253096,);
nor I_14708 (I252744,I253096,I253000);
not I_14709 (I253118,I253096);
nor I_14710 (I253135,I253118,I252909);
nor I_14711 (I253152,I252841,I253135);
DFFARX1 I_14712 (I253152,I3035,I252776,I252759,);
nor I_14713 (I253183,I253118,I253000);
nor I_14714 (I253200,I132449,I132452);
nor I_14715 (I252750,I253200,I253183);
not I_14716 (I253231,I253200);
nand I_14717 (I252753,I252960,I253231);
DFFARX1 I_14718 (I253200,I3035,I252776,I252765,);
DFFARX1 I_14719 (I253200,I3035,I252776,I252762,);
not I_14720 (I253320,I3042);
DFFARX1 I_14721 (I534862,I3035,I253320,I253346,);
DFFARX1 I_14722 (I253346,I3035,I253320,I253363,);
not I_14723 (I253312,I253363);
not I_14724 (I253385,I253346);
nand I_14725 (I253402,I534877,I534865);
and I_14726 (I253419,I253402,I534856);
DFFARX1 I_14727 (I253419,I3035,I253320,I253445,);
not I_14728 (I253453,I253445);
DFFARX1 I_14729 (I534868,I3035,I253320,I253479,);
and I_14730 (I253487,I253479,I534859);
nand I_14731 (I253504,I253479,I534859);
nand I_14732 (I253291,I253453,I253504);
DFFARX1 I_14733 (I534874,I3035,I253320,I253544,);
nor I_14734 (I253552,I253544,I253487);
DFFARX1 I_14735 (I253552,I3035,I253320,I253285,);
nor I_14736 (I253300,I253544,I253445);
nand I_14737 (I253597,I534883,I534871);
and I_14738 (I253614,I253597,I534880);
DFFARX1 I_14739 (I253614,I3035,I253320,I253640,);
nor I_14740 (I253288,I253640,I253544);
not I_14741 (I253662,I253640);
nor I_14742 (I253679,I253662,I253453);
nor I_14743 (I253696,I253385,I253679);
DFFARX1 I_14744 (I253696,I3035,I253320,I253303,);
nor I_14745 (I253727,I253662,I253544);
nor I_14746 (I253744,I534856,I534871);
nor I_14747 (I253294,I253744,I253727);
not I_14748 (I253775,I253744);
nand I_14749 (I253297,I253504,I253775);
DFFARX1 I_14750 (I253744,I3035,I253320,I253309,);
DFFARX1 I_14751 (I253744,I3035,I253320,I253306,);
not I_14752 (I253864,I3042);
DFFARX1 I_14753 (I281729,I3035,I253864,I253890,);
DFFARX1 I_14754 (I253890,I3035,I253864,I253907,);
not I_14755 (I253856,I253907);
not I_14756 (I253929,I253890);
nand I_14757 (I253946,I281732,I281750);
and I_14758 (I253963,I253946,I281738);
DFFARX1 I_14759 (I253963,I3035,I253864,I253989,);
not I_14760 (I253997,I253989);
DFFARX1 I_14761 (I281729,I3035,I253864,I254023,);
and I_14762 (I254031,I254023,I281747);
nand I_14763 (I254048,I254023,I281747);
nand I_14764 (I253835,I253997,I254048);
DFFARX1 I_14765 (I281741,I3035,I253864,I254088,);
nor I_14766 (I254096,I254088,I254031);
DFFARX1 I_14767 (I254096,I3035,I253864,I253829,);
nor I_14768 (I253844,I254088,I253989);
nand I_14769 (I254141,I281744,I281726);
and I_14770 (I254158,I254141,I281735);
DFFARX1 I_14771 (I254158,I3035,I253864,I254184,);
nor I_14772 (I253832,I254184,I254088);
not I_14773 (I254206,I254184);
nor I_14774 (I254223,I254206,I253997);
nor I_14775 (I254240,I253929,I254223);
DFFARX1 I_14776 (I254240,I3035,I253864,I253847,);
nor I_14777 (I254271,I254206,I254088);
nor I_14778 (I254288,I281726,I281726);
nor I_14779 (I253838,I254288,I254271);
not I_14780 (I254319,I254288);
nand I_14781 (I253841,I254048,I254319);
DFFARX1 I_14782 (I254288,I3035,I253864,I253853,);
DFFARX1 I_14783 (I254288,I3035,I253864,I253850,);
not I_14784 (I254408,I3042);
DFFARX1 I_14785 (I623157,I3035,I254408,I254434,);
DFFARX1 I_14786 (I254434,I3035,I254408,I254451,);
not I_14787 (I254400,I254451);
not I_14788 (I254473,I254434);
nand I_14789 (I254490,I623169,I623157);
and I_14790 (I254507,I254490,I623160);
DFFARX1 I_14791 (I254507,I3035,I254408,I254533,);
not I_14792 (I254541,I254533);
DFFARX1 I_14793 (I623178,I3035,I254408,I254567,);
and I_14794 (I254575,I254567,I623154);
nand I_14795 (I254592,I254567,I623154);
nand I_14796 (I254379,I254541,I254592);
DFFARX1 I_14797 (I623172,I3035,I254408,I254632,);
nor I_14798 (I254640,I254632,I254575);
DFFARX1 I_14799 (I254640,I3035,I254408,I254373,);
nor I_14800 (I254388,I254632,I254533);
nand I_14801 (I254685,I623166,I623163);
and I_14802 (I254702,I254685,I623175);
DFFARX1 I_14803 (I254702,I3035,I254408,I254728,);
nor I_14804 (I254376,I254728,I254632);
not I_14805 (I254750,I254728);
nor I_14806 (I254767,I254750,I254541);
nor I_14807 (I254784,I254473,I254767);
DFFARX1 I_14808 (I254784,I3035,I254408,I254391,);
nor I_14809 (I254815,I254750,I254632);
nor I_14810 (I254832,I623154,I623163);
nor I_14811 (I254382,I254832,I254815);
not I_14812 (I254863,I254832);
nand I_14813 (I254385,I254592,I254863);
DFFARX1 I_14814 (I254832,I3035,I254408,I254397,);
DFFARX1 I_14815 (I254832,I3035,I254408,I254394,);
not I_14816 (I254952,I3042);
DFFARX1 I_14817 (I212506,I3035,I254952,I254978,);
DFFARX1 I_14818 (I254978,I3035,I254952,I254995,);
not I_14819 (I254944,I254995);
not I_14820 (I255017,I254978);
nand I_14821 (I255034,I212485,I212509);
and I_14822 (I255051,I255034,I212512);
DFFARX1 I_14823 (I255051,I3035,I254952,I255077,);
not I_14824 (I255085,I255077);
DFFARX1 I_14825 (I212494,I3035,I254952,I255111,);
and I_14826 (I255119,I255111,I212500);
nand I_14827 (I255136,I255111,I212500);
nand I_14828 (I254923,I255085,I255136);
DFFARX1 I_14829 (I212488,I3035,I254952,I255176,);
nor I_14830 (I255184,I255176,I255119);
DFFARX1 I_14831 (I255184,I3035,I254952,I254917,);
nor I_14832 (I254932,I255176,I255077);
nand I_14833 (I255229,I212497,I212485);
and I_14834 (I255246,I255229,I212491);
DFFARX1 I_14835 (I255246,I3035,I254952,I255272,);
nor I_14836 (I254920,I255272,I255176);
not I_14837 (I255294,I255272);
nor I_14838 (I255311,I255294,I255085);
nor I_14839 (I255328,I255017,I255311);
DFFARX1 I_14840 (I255328,I3035,I254952,I254935,);
nor I_14841 (I255359,I255294,I255176);
nor I_14842 (I255376,I212503,I212485);
nor I_14843 (I254926,I255376,I255359);
not I_14844 (I255407,I255376);
nand I_14845 (I254929,I255136,I255407);
DFFARX1 I_14846 (I255376,I3035,I254952,I254941,);
DFFARX1 I_14847 (I255376,I3035,I254952,I254938,);
not I_14848 (I255496,I3042);
DFFARX1 I_14849 (I728785,I3035,I255496,I255522,);
DFFARX1 I_14850 (I255522,I3035,I255496,I255539,);
not I_14851 (I255488,I255539);
not I_14852 (I255561,I255522);
nand I_14853 (I255578,I728761,I728782);
and I_14854 (I255595,I255578,I728779);
DFFARX1 I_14855 (I255595,I3035,I255496,I255621,);
not I_14856 (I255629,I255621);
DFFARX1 I_14857 (I728758,I3035,I255496,I255655,);
and I_14858 (I255663,I255655,I728770);
nand I_14859 (I255680,I255655,I728770);
nand I_14860 (I255467,I255629,I255680);
DFFARX1 I_14861 (I728773,I3035,I255496,I255720,);
nor I_14862 (I255728,I255720,I255663);
DFFARX1 I_14863 (I255728,I3035,I255496,I255461,);
nor I_14864 (I255476,I255720,I255621);
nand I_14865 (I255773,I728776,I728764);
and I_14866 (I255790,I255773,I728767);
DFFARX1 I_14867 (I255790,I3035,I255496,I255816,);
nor I_14868 (I255464,I255816,I255720);
not I_14869 (I255838,I255816);
nor I_14870 (I255855,I255838,I255629);
nor I_14871 (I255872,I255561,I255855);
DFFARX1 I_14872 (I255872,I3035,I255496,I255479,);
nor I_14873 (I255903,I255838,I255720);
nor I_14874 (I255920,I728758,I728764);
nor I_14875 (I255470,I255920,I255903);
not I_14876 (I255951,I255920);
nand I_14877 (I255473,I255680,I255951);
DFFARX1 I_14878 (I255920,I3035,I255496,I255485,);
DFFARX1 I_14879 (I255920,I3035,I255496,I255482,);
not I_14880 (I256040,I3042);
DFFARX1 I_14881 (I224627,I3035,I256040,I256066,);
DFFARX1 I_14882 (I256066,I3035,I256040,I256083,);
not I_14883 (I256032,I256083);
not I_14884 (I256105,I256066);
nand I_14885 (I256122,I224606,I224630);
and I_14886 (I256139,I256122,I224633);
DFFARX1 I_14887 (I256139,I3035,I256040,I256165,);
not I_14888 (I256173,I256165);
DFFARX1 I_14889 (I224615,I3035,I256040,I256199,);
and I_14890 (I256207,I256199,I224621);
nand I_14891 (I256224,I256199,I224621);
nand I_14892 (I256011,I256173,I256224);
DFFARX1 I_14893 (I224609,I3035,I256040,I256264,);
nor I_14894 (I256272,I256264,I256207);
DFFARX1 I_14895 (I256272,I3035,I256040,I256005,);
nor I_14896 (I256020,I256264,I256165);
nand I_14897 (I256317,I224618,I224606);
and I_14898 (I256334,I256317,I224612);
DFFARX1 I_14899 (I256334,I3035,I256040,I256360,);
nor I_14900 (I256008,I256360,I256264);
not I_14901 (I256382,I256360);
nor I_14902 (I256399,I256382,I256173);
nor I_14903 (I256416,I256105,I256399);
DFFARX1 I_14904 (I256416,I3035,I256040,I256023,);
nor I_14905 (I256447,I256382,I256264);
nor I_14906 (I256464,I224624,I224606);
nor I_14907 (I256014,I256464,I256447);
not I_14908 (I256495,I256464);
nand I_14909 (I256017,I256224,I256495);
DFFARX1 I_14910 (I256464,I3035,I256040,I256029,);
DFFARX1 I_14911 (I256464,I3035,I256040,I256026,);
not I_14912 (I256584,I3042);
DFFARX1 I_14913 (I71051,I3035,I256584,I256610,);
DFFARX1 I_14914 (I256610,I3035,I256584,I256627,);
not I_14915 (I256576,I256627);
not I_14916 (I256649,I256610);
nand I_14917 (I256666,I71066,I71045);
and I_14918 (I256683,I256666,I71048);
DFFARX1 I_14919 (I256683,I3035,I256584,I256709,);
not I_14920 (I256717,I256709);
DFFARX1 I_14921 (I71054,I3035,I256584,I256743,);
and I_14922 (I256751,I256743,I71048);
nand I_14923 (I256768,I256743,I71048);
nand I_14924 (I256555,I256717,I256768);
DFFARX1 I_14925 (I71063,I3035,I256584,I256808,);
nor I_14926 (I256816,I256808,I256751);
DFFARX1 I_14927 (I256816,I3035,I256584,I256549,);
nor I_14928 (I256564,I256808,I256709);
nand I_14929 (I256861,I71045,I71060);
and I_14930 (I256878,I256861,I71057);
DFFARX1 I_14931 (I256878,I3035,I256584,I256904,);
nor I_14932 (I256552,I256904,I256808);
not I_14933 (I256926,I256904);
nor I_14934 (I256943,I256926,I256717);
nor I_14935 (I256960,I256649,I256943);
DFFARX1 I_14936 (I256960,I3035,I256584,I256567,);
nor I_14937 (I256991,I256926,I256808);
nor I_14938 (I257008,I71069,I71060);
nor I_14939 (I256558,I257008,I256991);
not I_14940 (I257039,I257008);
nand I_14941 (I256561,I256768,I257039);
DFFARX1 I_14942 (I257008,I3035,I256584,I256573,);
DFFARX1 I_14943 (I257008,I3035,I256584,I256570,);
not I_14944 (I257128,I3042);
DFFARX1 I_14945 (I386279,I3035,I257128,I257154,);
DFFARX1 I_14946 (I257154,I3035,I257128,I257171,);
not I_14947 (I257120,I257171);
not I_14948 (I257193,I257154);
nand I_14949 (I257210,I386300,I386291);
and I_14950 (I257227,I257210,I386279);
DFFARX1 I_14951 (I257227,I3035,I257128,I257253,);
not I_14952 (I257261,I257253);
DFFARX1 I_14953 (I386285,I3035,I257128,I257287,);
and I_14954 (I257295,I257287,I386282);
nand I_14955 (I257312,I257287,I386282);
nand I_14956 (I257099,I257261,I257312);
DFFARX1 I_14957 (I386276,I3035,I257128,I257352,);
nor I_14958 (I257360,I257352,I257295);
DFFARX1 I_14959 (I257360,I3035,I257128,I257093,);
nor I_14960 (I257108,I257352,I257253);
nand I_14961 (I257405,I386276,I386288);
and I_14962 (I257422,I257405,I386297);
DFFARX1 I_14963 (I257422,I3035,I257128,I257448,);
nor I_14964 (I257096,I257448,I257352);
not I_14965 (I257470,I257448);
nor I_14966 (I257487,I257470,I257261);
nor I_14967 (I257504,I257193,I257487);
DFFARX1 I_14968 (I257504,I3035,I257128,I257111,);
nor I_14969 (I257535,I257470,I257352);
nor I_14970 (I257552,I386294,I386288);
nor I_14971 (I257102,I257552,I257535);
not I_14972 (I257583,I257552);
nand I_14973 (I257105,I257312,I257583);
DFFARX1 I_14974 (I257552,I3035,I257128,I257117,);
DFFARX1 I_14975 (I257552,I3035,I257128,I257114,);
not I_14976 (I257672,I3042);
DFFARX1 I_14977 (I523880,I3035,I257672,I257698,);
DFFARX1 I_14978 (I257698,I3035,I257672,I257715,);
not I_14979 (I257664,I257715);
not I_14980 (I257737,I257698);
nand I_14981 (I257754,I523895,I523883);
and I_14982 (I257771,I257754,I523874);
DFFARX1 I_14983 (I257771,I3035,I257672,I257797,);
not I_14984 (I257805,I257797);
DFFARX1 I_14985 (I523886,I3035,I257672,I257831,);
and I_14986 (I257839,I257831,I523877);
nand I_14987 (I257856,I257831,I523877);
nand I_14988 (I257643,I257805,I257856);
DFFARX1 I_14989 (I523892,I3035,I257672,I257896,);
nor I_14990 (I257904,I257896,I257839);
DFFARX1 I_14991 (I257904,I3035,I257672,I257637,);
nor I_14992 (I257652,I257896,I257797);
nand I_14993 (I257949,I523901,I523889);
and I_14994 (I257966,I257949,I523898);
DFFARX1 I_14995 (I257966,I3035,I257672,I257992,);
nor I_14996 (I257640,I257992,I257896);
not I_14997 (I258014,I257992);
nor I_14998 (I258031,I258014,I257805);
nor I_14999 (I258048,I257737,I258031);
DFFARX1 I_15000 (I258048,I3035,I257672,I257655,);
nor I_15001 (I258079,I258014,I257896);
nor I_15002 (I258096,I523874,I523889);
nor I_15003 (I257646,I258096,I258079);
not I_15004 (I258127,I258096);
nand I_15005 (I257649,I257856,I258127);
DFFARX1 I_15006 (I258096,I3035,I257672,I257661,);
DFFARX1 I_15007 (I258096,I3035,I257672,I257658,);
not I_15008 (I258216,I3042);
DFFARX1 I_15009 (I167184,I3035,I258216,I258242,);
DFFARX1 I_15010 (I258242,I3035,I258216,I258259,);
not I_15011 (I258208,I258259);
not I_15012 (I258281,I258242);
nand I_15013 (I258298,I167163,I167187);
and I_15014 (I258315,I258298,I167190);
DFFARX1 I_15015 (I258315,I3035,I258216,I258341,);
not I_15016 (I258349,I258341);
DFFARX1 I_15017 (I167172,I3035,I258216,I258375,);
and I_15018 (I258383,I258375,I167178);
nand I_15019 (I258400,I258375,I167178);
nand I_15020 (I258187,I258349,I258400);
DFFARX1 I_15021 (I167166,I3035,I258216,I258440,);
nor I_15022 (I258448,I258440,I258383);
DFFARX1 I_15023 (I258448,I3035,I258216,I258181,);
nor I_15024 (I258196,I258440,I258341);
nand I_15025 (I258493,I167175,I167163);
and I_15026 (I258510,I258493,I167169);
DFFARX1 I_15027 (I258510,I3035,I258216,I258536,);
nor I_15028 (I258184,I258536,I258440);
not I_15029 (I258558,I258536);
nor I_15030 (I258575,I258558,I258349);
nor I_15031 (I258592,I258281,I258575);
DFFARX1 I_15032 (I258592,I3035,I258216,I258199,);
nor I_15033 (I258623,I258558,I258440);
nor I_15034 (I258640,I167181,I167163);
nor I_15035 (I258190,I258640,I258623);
not I_15036 (I258671,I258640);
nand I_15037 (I258193,I258400,I258671);
DFFARX1 I_15038 (I258640,I3035,I258216,I258205,);
DFFARX1 I_15039 (I258640,I3035,I258216,I258202,);
not I_15040 (I258760,I3042);
DFFARX1 I_15041 (I465134,I3035,I258760,I258786,);
DFFARX1 I_15042 (I258786,I3035,I258760,I258803,);
not I_15043 (I258752,I258803);
not I_15044 (I258825,I258786);
nand I_15045 (I258842,I465128,I465125);
and I_15046 (I258859,I258842,I465140);
DFFARX1 I_15047 (I258859,I3035,I258760,I258885,);
not I_15048 (I258893,I258885);
DFFARX1 I_15049 (I465128,I3035,I258760,I258919,);
and I_15050 (I258927,I258919,I465122);
nand I_15051 (I258944,I258919,I465122);
nand I_15052 (I258731,I258893,I258944);
DFFARX1 I_15053 (I465122,I3035,I258760,I258984,);
nor I_15054 (I258992,I258984,I258927);
DFFARX1 I_15055 (I258992,I3035,I258760,I258725,);
nor I_15056 (I258740,I258984,I258885);
nand I_15057 (I259037,I465137,I465131);
and I_15058 (I259054,I259037,I465125);
DFFARX1 I_15059 (I259054,I3035,I258760,I259080,);
nor I_15060 (I258728,I259080,I258984);
not I_15061 (I259102,I259080);
nor I_15062 (I259119,I259102,I258893);
nor I_15063 (I259136,I258825,I259119);
DFFARX1 I_15064 (I259136,I3035,I258760,I258743,);
nor I_15065 (I259167,I259102,I258984);
nor I_15066 (I259184,I465143,I465131);
nor I_15067 (I258734,I259184,I259167);
not I_15068 (I259215,I259184);
nand I_15069 (I258737,I258944,I259215);
DFFARX1 I_15070 (I259184,I3035,I258760,I258749,);
DFFARX1 I_15071 (I259184,I3035,I258760,I258746,);
not I_15072 (I259304,I3042);
DFFARX1 I_15073 (I657769,I3035,I259304,I259330,);
DFFARX1 I_15074 (I259330,I3035,I259304,I259347,);
not I_15075 (I259296,I259347);
not I_15076 (I259369,I259330);
nand I_15077 (I259386,I657781,I657784);
and I_15078 (I259403,I259386,I657787);
DFFARX1 I_15079 (I259403,I3035,I259304,I259429,);
not I_15080 (I259437,I259429);
DFFARX1 I_15081 (I657772,I3035,I259304,I259463,);
and I_15082 (I259471,I259463,I657778);
nand I_15083 (I259488,I259463,I657778);
nand I_15084 (I259275,I259437,I259488);
DFFARX1 I_15085 (I657766,I3035,I259304,I259528,);
nor I_15086 (I259536,I259528,I259471);
DFFARX1 I_15087 (I259536,I3035,I259304,I259269,);
nor I_15088 (I259284,I259528,I259429);
nand I_15089 (I259581,I657769,I657790);
and I_15090 (I259598,I259581,I657775);
DFFARX1 I_15091 (I259598,I3035,I259304,I259624,);
nor I_15092 (I259272,I259624,I259528);
not I_15093 (I259646,I259624);
nor I_15094 (I259663,I259646,I259437);
nor I_15095 (I259680,I259369,I259663);
DFFARX1 I_15096 (I259680,I3035,I259304,I259287,);
nor I_15097 (I259711,I259646,I259528);
nor I_15098 (I259728,I657766,I657790);
nor I_15099 (I259278,I259728,I259711);
not I_15100 (I259759,I259728);
nand I_15101 (I259281,I259488,I259759);
DFFARX1 I_15102 (I259728,I3035,I259304,I259293,);
DFFARX1 I_15103 (I259728,I3035,I259304,I259290,);
not I_15104 (I259848,I3042);
DFFARX1 I_15105 (I179305,I3035,I259848,I259874,);
DFFARX1 I_15106 (I259874,I3035,I259848,I259891,);
not I_15107 (I259840,I259891);
not I_15108 (I259913,I259874);
nand I_15109 (I259930,I179284,I179308);
and I_15110 (I259947,I259930,I179311);
DFFARX1 I_15111 (I259947,I3035,I259848,I259973,);
not I_15112 (I259981,I259973);
DFFARX1 I_15113 (I179293,I3035,I259848,I260007,);
and I_15114 (I260015,I260007,I179299);
nand I_15115 (I260032,I260007,I179299);
nand I_15116 (I259819,I259981,I260032);
DFFARX1 I_15117 (I179287,I3035,I259848,I260072,);
nor I_15118 (I260080,I260072,I260015);
DFFARX1 I_15119 (I260080,I3035,I259848,I259813,);
nor I_15120 (I259828,I260072,I259973);
nand I_15121 (I260125,I179296,I179284);
and I_15122 (I260142,I260125,I179290);
DFFARX1 I_15123 (I260142,I3035,I259848,I260168,);
nor I_15124 (I259816,I260168,I260072);
not I_15125 (I260190,I260168);
nor I_15126 (I260207,I260190,I259981);
nor I_15127 (I260224,I259913,I260207);
DFFARX1 I_15128 (I260224,I3035,I259848,I259831,);
nor I_15129 (I260255,I260190,I260072);
nor I_15130 (I260272,I179302,I179284);
nor I_15131 (I259822,I260272,I260255);
not I_15132 (I260303,I260272);
nand I_15133 (I259825,I260032,I260303);
DFFARX1 I_15134 (I260272,I3035,I259848,I259837,);
DFFARX1 I_15135 (I260272,I3035,I259848,I259834,);
not I_15136 (I260392,I3042);
DFFARX1 I_15137 (I567241,I3035,I260392,I260418,);
DFFARX1 I_15138 (I260418,I3035,I260392,I260435,);
not I_15139 (I260384,I260435);
not I_15140 (I260457,I260418);
nand I_15141 (I260474,I567241,I567259);
and I_15142 (I260491,I260474,I567253);
DFFARX1 I_15143 (I260491,I3035,I260392,I260517,);
not I_15144 (I260525,I260517);
DFFARX1 I_15145 (I567247,I3035,I260392,I260551,);
and I_15146 (I260559,I260551,I567256);
nand I_15147 (I260576,I260551,I567256);
nand I_15148 (I260363,I260525,I260576);
DFFARX1 I_15149 (I567244,I3035,I260392,I260616,);
nor I_15150 (I260624,I260616,I260559);
DFFARX1 I_15151 (I260624,I3035,I260392,I260357,);
nor I_15152 (I260372,I260616,I260517);
nand I_15153 (I260669,I567244,I567262);
and I_15154 (I260686,I260669,I567247);
DFFARX1 I_15155 (I260686,I3035,I260392,I260712,);
nor I_15156 (I260360,I260712,I260616);
not I_15157 (I260734,I260712);
nor I_15158 (I260751,I260734,I260525);
nor I_15159 (I260768,I260457,I260751);
DFFARX1 I_15160 (I260768,I3035,I260392,I260375,);
nor I_15161 (I260799,I260734,I260616);
nor I_15162 (I260816,I567250,I567262);
nor I_15163 (I260366,I260816,I260799);
not I_15164 (I260847,I260816);
nand I_15165 (I260369,I260576,I260847);
DFFARX1 I_15166 (I260816,I3035,I260392,I260381,);
DFFARX1 I_15167 (I260816,I3035,I260392,I260378,);
not I_15168 (I260936,I3042);
DFFARX1 I_15169 (I315185,I3035,I260936,I260962,);
DFFARX1 I_15170 (I260962,I3035,I260936,I260979,);
not I_15171 (I260928,I260979);
not I_15172 (I261001,I260962);
nand I_15173 (I261018,I315182,I315203);
and I_15174 (I261035,I261018,I315206);
DFFARX1 I_15175 (I261035,I3035,I260936,I261061,);
not I_15176 (I261069,I261061);
DFFARX1 I_15177 (I315191,I3035,I260936,I261095,);
and I_15178 (I261103,I261095,I315194);
nand I_15179 (I261120,I261095,I315194);
nand I_15180 (I260907,I261069,I261120);
DFFARX1 I_15181 (I315197,I3035,I260936,I261160,);
nor I_15182 (I261168,I261160,I261103);
DFFARX1 I_15183 (I261168,I3035,I260936,I260901,);
nor I_15184 (I260916,I261160,I261061);
nand I_15185 (I261213,I315182,I315188);
and I_15186 (I261230,I261213,I315200);
DFFARX1 I_15187 (I261230,I3035,I260936,I261256,);
nor I_15188 (I260904,I261256,I261160);
not I_15189 (I261278,I261256);
nor I_15190 (I261295,I261278,I261069);
nor I_15191 (I261312,I261001,I261295);
DFFARX1 I_15192 (I261312,I3035,I260936,I260919,);
nor I_15193 (I261343,I261278,I261160);
nor I_15194 (I261360,I315185,I315188);
nor I_15195 (I260910,I261360,I261343);
not I_15196 (I261391,I261360);
nand I_15197 (I260913,I261120,I261391);
DFFARX1 I_15198 (I261360,I3035,I260936,I260925,);
DFFARX1 I_15199 (I261360,I3035,I260936,I260922,);
not I_15200 (I261480,I3042);
DFFARX1 I_15201 (I347553,I3035,I261480,I261506,);
DFFARX1 I_15202 (I261506,I3035,I261480,I261523,);
not I_15203 (I261472,I261523);
not I_15204 (I261545,I261506);
nand I_15205 (I261562,I347574,I347565);
and I_15206 (I261579,I261562,I347553);
DFFARX1 I_15207 (I261579,I3035,I261480,I261605,);
not I_15208 (I261613,I261605);
DFFARX1 I_15209 (I347559,I3035,I261480,I261639,);
and I_15210 (I261647,I261639,I347556);
nand I_15211 (I261664,I261639,I347556);
nand I_15212 (I261451,I261613,I261664);
DFFARX1 I_15213 (I347550,I3035,I261480,I261704,);
nor I_15214 (I261712,I261704,I261647);
DFFARX1 I_15215 (I261712,I3035,I261480,I261445,);
nor I_15216 (I261460,I261704,I261605);
nand I_15217 (I261757,I347550,I347562);
and I_15218 (I261774,I261757,I347571);
DFFARX1 I_15219 (I261774,I3035,I261480,I261800,);
nor I_15220 (I261448,I261800,I261704);
not I_15221 (I261822,I261800);
nor I_15222 (I261839,I261822,I261613);
nor I_15223 (I261856,I261545,I261839);
DFFARX1 I_15224 (I261856,I3035,I261480,I261463,);
nor I_15225 (I261887,I261822,I261704);
nor I_15226 (I261904,I347568,I347562);
nor I_15227 (I261454,I261904,I261887);
not I_15228 (I261935,I261904);
nand I_15229 (I261457,I261664,I261935);
DFFARX1 I_15230 (I261904,I3035,I261480,I261469,);
DFFARX1 I_15231 (I261904,I3035,I261480,I261466,);
not I_15232 (I262024,I3042);
DFFARX1 I_15233 (I378187,I3035,I262024,I262050,);
DFFARX1 I_15234 (I262050,I3035,I262024,I262067,);
not I_15235 (I262016,I262067);
not I_15236 (I262089,I262050);
nand I_15237 (I262106,I378208,I378199);
and I_15238 (I262123,I262106,I378187);
DFFARX1 I_15239 (I262123,I3035,I262024,I262149,);
not I_15240 (I262157,I262149);
DFFARX1 I_15241 (I378193,I3035,I262024,I262183,);
and I_15242 (I262191,I262183,I378190);
nand I_15243 (I262208,I262183,I378190);
nand I_15244 (I261995,I262157,I262208);
DFFARX1 I_15245 (I378184,I3035,I262024,I262248,);
nor I_15246 (I262256,I262248,I262191);
DFFARX1 I_15247 (I262256,I3035,I262024,I261989,);
nor I_15248 (I262004,I262248,I262149);
nand I_15249 (I262301,I378184,I378196);
and I_15250 (I262318,I262301,I378205);
DFFARX1 I_15251 (I262318,I3035,I262024,I262344,);
nor I_15252 (I261992,I262344,I262248);
not I_15253 (I262366,I262344);
nor I_15254 (I262383,I262366,I262157);
nor I_15255 (I262400,I262089,I262383);
DFFARX1 I_15256 (I262400,I3035,I262024,I262007,);
nor I_15257 (I262431,I262366,I262248);
nor I_15258 (I262448,I378202,I378196);
nor I_15259 (I261998,I262448,I262431);
not I_15260 (I262479,I262448);
nand I_15261 (I262001,I262208,I262479);
DFFARX1 I_15262 (I262448,I3035,I262024,I262013,);
DFFARX1 I_15263 (I262448,I3035,I262024,I262010,);
not I_15264 (I262568,I3042);
DFFARX1 I_15265 (I650153,I3035,I262568,I262594,);
DFFARX1 I_15266 (I262594,I3035,I262568,I262611,);
not I_15267 (I262560,I262611);
not I_15268 (I262633,I262594);
nand I_15269 (I262650,I650165,I650168);
and I_15270 (I262667,I262650,I650171);
DFFARX1 I_15271 (I262667,I3035,I262568,I262693,);
not I_15272 (I262701,I262693);
DFFARX1 I_15273 (I650156,I3035,I262568,I262727,);
and I_15274 (I262735,I262727,I650162);
nand I_15275 (I262752,I262727,I650162);
nand I_15276 (I262539,I262701,I262752);
DFFARX1 I_15277 (I650150,I3035,I262568,I262792,);
nor I_15278 (I262800,I262792,I262735);
DFFARX1 I_15279 (I262800,I3035,I262568,I262533,);
nor I_15280 (I262548,I262792,I262693);
nand I_15281 (I262845,I650153,I650174);
and I_15282 (I262862,I262845,I650159);
DFFARX1 I_15283 (I262862,I3035,I262568,I262888,);
nor I_15284 (I262536,I262888,I262792);
not I_15285 (I262910,I262888);
nor I_15286 (I262927,I262910,I262701);
nor I_15287 (I262944,I262633,I262927);
DFFARX1 I_15288 (I262944,I3035,I262568,I262551,);
nor I_15289 (I262975,I262910,I262792);
nor I_15290 (I262992,I650150,I650174);
nor I_15291 (I262542,I262992,I262975);
not I_15292 (I263023,I262992);
nand I_15293 (I262545,I262752,I263023);
DFFARX1 I_15294 (I262992,I3035,I262568,I262557,);
DFFARX1 I_15295 (I262992,I3035,I262568,I262554,);
not I_15296 (I263112,I3042);
DFFARX1 I_15297 (I569485,I3035,I263112,I263138,);
DFFARX1 I_15298 (I263138,I3035,I263112,I263155,);
not I_15299 (I263104,I263155);
not I_15300 (I263177,I263138);
nand I_15301 (I263194,I569485,I569503);
and I_15302 (I263211,I263194,I569497);
DFFARX1 I_15303 (I263211,I3035,I263112,I263237,);
not I_15304 (I263245,I263237);
DFFARX1 I_15305 (I569491,I3035,I263112,I263271,);
and I_15306 (I263279,I263271,I569500);
nand I_15307 (I263296,I263271,I569500);
nand I_15308 (I263083,I263245,I263296);
DFFARX1 I_15309 (I569488,I3035,I263112,I263336,);
nor I_15310 (I263344,I263336,I263279);
DFFARX1 I_15311 (I263344,I3035,I263112,I263077,);
nor I_15312 (I263092,I263336,I263237);
nand I_15313 (I263389,I569488,I569506);
and I_15314 (I263406,I263389,I569491);
DFFARX1 I_15315 (I263406,I3035,I263112,I263432,);
nor I_15316 (I263080,I263432,I263336);
not I_15317 (I263454,I263432);
nor I_15318 (I263471,I263454,I263245);
nor I_15319 (I263488,I263177,I263471);
DFFARX1 I_15320 (I263488,I3035,I263112,I263095,);
nor I_15321 (I263519,I263454,I263336);
nor I_15322 (I263536,I569494,I569506);
nor I_15323 (I263086,I263536,I263519);
not I_15324 (I263567,I263536);
nand I_15325 (I263089,I263296,I263567);
DFFARX1 I_15326 (I263536,I3035,I263112,I263101,);
DFFARX1 I_15327 (I263536,I3035,I263112,I263098,);
not I_15328 (I263656,I3042);
DFFARX1 I_15329 (I20465,I3035,I263656,I263682,);
DFFARX1 I_15330 (I263682,I3035,I263656,I263699,);
not I_15331 (I263648,I263699);
not I_15332 (I263721,I263682);
nand I_15333 (I263738,I20453,I20468);
and I_15334 (I263755,I263738,I20456);
DFFARX1 I_15335 (I263755,I3035,I263656,I263781,);
not I_15336 (I263789,I263781);
DFFARX1 I_15337 (I20477,I3035,I263656,I263815,);
and I_15338 (I263823,I263815,I20471);
nand I_15339 (I263840,I263815,I20471);
nand I_15340 (I263627,I263789,I263840);
DFFARX1 I_15341 (I20474,I3035,I263656,I263880,);
nor I_15342 (I263888,I263880,I263823);
DFFARX1 I_15343 (I263888,I3035,I263656,I263621,);
nor I_15344 (I263636,I263880,I263781);
nand I_15345 (I263933,I20453,I20456);
and I_15346 (I263950,I263933,I20459);
DFFARX1 I_15347 (I263950,I3035,I263656,I263976,);
nor I_15348 (I263624,I263976,I263880);
not I_15349 (I263998,I263976);
nor I_15350 (I264015,I263998,I263789);
nor I_15351 (I264032,I263721,I264015);
DFFARX1 I_15352 (I264032,I3035,I263656,I263639,);
nor I_15353 (I264063,I263998,I263880);
nor I_15354 (I264080,I20462,I20456);
nor I_15355 (I263630,I264080,I264063);
not I_15356 (I264111,I264080);
nand I_15357 (I263633,I263840,I264111);
DFFARX1 I_15358 (I264080,I3035,I263656,I263645,);
DFFARX1 I_15359 (I264080,I3035,I263656,I263642,);
not I_15360 (I264200,I3042);
DFFARX1 I_15361 (I332525,I3035,I264200,I264226,);
DFFARX1 I_15362 (I264226,I3035,I264200,I264243,);
not I_15363 (I264192,I264243);
not I_15364 (I264265,I264226);
nand I_15365 (I264282,I332522,I332543);
and I_15366 (I264299,I264282,I332546);
DFFARX1 I_15367 (I264299,I3035,I264200,I264325,);
not I_15368 (I264333,I264325);
DFFARX1 I_15369 (I332531,I3035,I264200,I264359,);
and I_15370 (I264367,I264359,I332534);
nand I_15371 (I264384,I264359,I332534);
nand I_15372 (I264171,I264333,I264384);
DFFARX1 I_15373 (I332537,I3035,I264200,I264424,);
nor I_15374 (I264432,I264424,I264367);
DFFARX1 I_15375 (I264432,I3035,I264200,I264165,);
nor I_15376 (I264180,I264424,I264325);
nand I_15377 (I264477,I332522,I332528);
and I_15378 (I264494,I264477,I332540);
DFFARX1 I_15379 (I264494,I3035,I264200,I264520,);
nor I_15380 (I264168,I264520,I264424);
not I_15381 (I264542,I264520);
nor I_15382 (I264559,I264542,I264333);
nor I_15383 (I264576,I264265,I264559);
DFFARX1 I_15384 (I264576,I3035,I264200,I264183,);
nor I_15385 (I264607,I264542,I264424);
nor I_15386 (I264624,I332525,I332528);
nor I_15387 (I264174,I264624,I264607);
not I_15388 (I264655,I264624);
nand I_15389 (I264177,I264384,I264655);
DFFARX1 I_15390 (I264624,I3035,I264200,I264189,);
DFFARX1 I_15391 (I264624,I3035,I264200,I264186,);
not I_15392 (I264744,I3042);
DFFARX1 I_15393 (I398417,I3035,I264744,I264770,);
DFFARX1 I_15394 (I264770,I3035,I264744,I264787,);
not I_15395 (I264736,I264787);
not I_15396 (I264809,I264770);
nand I_15397 (I264826,I398438,I398429);
and I_15398 (I264843,I264826,I398417);
DFFARX1 I_15399 (I264843,I3035,I264744,I264869,);
not I_15400 (I264877,I264869);
DFFARX1 I_15401 (I398423,I3035,I264744,I264903,);
and I_15402 (I264911,I264903,I398420);
nand I_15403 (I264928,I264903,I398420);
nand I_15404 (I264715,I264877,I264928);
DFFARX1 I_15405 (I398414,I3035,I264744,I264968,);
nor I_15406 (I264976,I264968,I264911);
DFFARX1 I_15407 (I264976,I3035,I264744,I264709,);
nor I_15408 (I264724,I264968,I264869);
nand I_15409 (I265021,I398414,I398426);
and I_15410 (I265038,I265021,I398435);
DFFARX1 I_15411 (I265038,I3035,I264744,I265064,);
nor I_15412 (I264712,I265064,I264968);
not I_15413 (I265086,I265064);
nor I_15414 (I265103,I265086,I264877);
nor I_15415 (I265120,I264809,I265103);
DFFARX1 I_15416 (I265120,I3035,I264744,I264727,);
nor I_15417 (I265151,I265086,I264968);
nor I_15418 (I265168,I398432,I398426);
nor I_15419 (I264718,I265168,I265151);
not I_15420 (I265199,I265168);
nand I_15421 (I264721,I264928,I265199);
DFFARX1 I_15422 (I265168,I3035,I264744,I264733,);
DFFARX1 I_15423 (I265168,I3035,I264744,I264730,);
not I_15424 (I265288,I3042);
DFFARX1 I_15425 (I696116,I3035,I265288,I265314,);
DFFARX1 I_15426 (I265314,I3035,I265288,I265331,);
not I_15427 (I265280,I265331);
not I_15428 (I265353,I265314);
nand I_15429 (I265370,I696122,I696125);
and I_15430 (I265387,I265370,I696101);
DFFARX1 I_15431 (I265387,I3035,I265288,I265413,);
not I_15432 (I265421,I265413);
DFFARX1 I_15433 (I696128,I3035,I265288,I265447,);
and I_15434 (I265455,I265447,I696110);
nand I_15435 (I265472,I265447,I696110);
nand I_15436 (I265259,I265421,I265472);
DFFARX1 I_15437 (I696107,I3035,I265288,I265512,);
nor I_15438 (I265520,I265512,I265455);
DFFARX1 I_15439 (I265520,I3035,I265288,I265253,);
nor I_15440 (I265268,I265512,I265413);
nand I_15441 (I265565,I696104,I696113);
and I_15442 (I265582,I265565,I696119);
DFFARX1 I_15443 (I265582,I3035,I265288,I265608,);
nor I_15444 (I265256,I265608,I265512);
not I_15445 (I265630,I265608);
nor I_15446 (I265647,I265630,I265421);
nor I_15447 (I265664,I265353,I265647);
DFFARX1 I_15448 (I265664,I3035,I265288,I265271,);
nor I_15449 (I265695,I265630,I265512);
nor I_15450 (I265712,I696101,I696113);
nor I_15451 (I265262,I265712,I265695);
not I_15452 (I265743,I265712);
nand I_15453 (I265265,I265472,I265743);
DFFARX1 I_15454 (I265712,I3035,I265288,I265277,);
DFFARX1 I_15455 (I265712,I3035,I265288,I265274,);
not I_15456 (I265832,I3042);
DFFARX1 I_15457 (I718670,I3035,I265832,I265858,);
DFFARX1 I_15458 (I265858,I3035,I265832,I265875,);
not I_15459 (I265824,I265875);
not I_15460 (I265897,I265858);
nand I_15461 (I265914,I718646,I718667);
and I_15462 (I265931,I265914,I718664);
DFFARX1 I_15463 (I265931,I3035,I265832,I265957,);
not I_15464 (I265965,I265957);
DFFARX1 I_15465 (I718643,I3035,I265832,I265991,);
and I_15466 (I265999,I265991,I718655);
nand I_15467 (I266016,I265991,I718655);
nand I_15468 (I265803,I265965,I266016);
DFFARX1 I_15469 (I718658,I3035,I265832,I266056,);
nor I_15470 (I266064,I266056,I265999);
DFFARX1 I_15471 (I266064,I3035,I265832,I265797,);
nor I_15472 (I265812,I266056,I265957);
nand I_15473 (I266109,I718661,I718649);
and I_15474 (I266126,I266109,I718652);
DFFARX1 I_15475 (I266126,I3035,I265832,I266152,);
nor I_15476 (I265800,I266152,I266056);
not I_15477 (I266174,I266152);
nor I_15478 (I266191,I266174,I265965);
nor I_15479 (I266208,I265897,I266191);
DFFARX1 I_15480 (I266208,I3035,I265832,I265815,);
nor I_15481 (I266239,I266174,I266056);
nor I_15482 (I266256,I718643,I718649);
nor I_15483 (I265806,I266256,I266239);
not I_15484 (I266287,I266256);
nand I_15485 (I265809,I266016,I266287);
DFFARX1 I_15486 (I266256,I3035,I265832,I265821,);
DFFARX1 I_15487 (I266256,I3035,I265832,I265818,);
not I_15488 (I266376,I3042);
DFFARX1 I_15489 (I719265,I3035,I266376,I266402,);
DFFARX1 I_15490 (I266402,I3035,I266376,I266419,);
not I_15491 (I266368,I266419);
not I_15492 (I266441,I266402);
nand I_15493 (I266458,I719241,I719262);
and I_15494 (I266475,I266458,I719259);
DFFARX1 I_15495 (I266475,I3035,I266376,I266501,);
not I_15496 (I266509,I266501);
DFFARX1 I_15497 (I719238,I3035,I266376,I266535,);
and I_15498 (I266543,I266535,I719250);
nand I_15499 (I266560,I266535,I719250);
nand I_15500 (I266347,I266509,I266560);
DFFARX1 I_15501 (I719253,I3035,I266376,I266600,);
nor I_15502 (I266608,I266600,I266543);
DFFARX1 I_15503 (I266608,I3035,I266376,I266341,);
nor I_15504 (I266356,I266600,I266501);
nand I_15505 (I266653,I719256,I719244);
and I_15506 (I266670,I266653,I719247);
DFFARX1 I_15507 (I266670,I3035,I266376,I266696,);
nor I_15508 (I266344,I266696,I266600);
not I_15509 (I266718,I266696);
nor I_15510 (I266735,I266718,I266509);
nor I_15511 (I266752,I266441,I266735);
DFFARX1 I_15512 (I266752,I3035,I266376,I266359,);
nor I_15513 (I266783,I266718,I266600);
nor I_15514 (I266800,I719238,I719244);
nor I_15515 (I266350,I266800,I266783);
not I_15516 (I266831,I266800);
nand I_15517 (I266353,I266560,I266831);
DFFARX1 I_15518 (I266800,I3035,I266376,I266365,);
DFFARX1 I_15519 (I266800,I3035,I266376,I266362,);
not I_15520 (I266920,I3042);
DFFARX1 I_15521 (I30999,I3035,I266920,I266946,);
DFFARX1 I_15522 (I266946,I3035,I266920,I266963,);
not I_15523 (I266912,I266963);
not I_15524 (I266985,I266946);
nand I_15525 (I267002,I31014,I30993);
and I_15526 (I267019,I267002,I30996);
DFFARX1 I_15527 (I267019,I3035,I266920,I267045,);
not I_15528 (I267053,I267045);
DFFARX1 I_15529 (I31002,I3035,I266920,I267079,);
and I_15530 (I267087,I267079,I30996);
nand I_15531 (I267104,I267079,I30996);
nand I_15532 (I266891,I267053,I267104);
DFFARX1 I_15533 (I31011,I3035,I266920,I267144,);
nor I_15534 (I267152,I267144,I267087);
DFFARX1 I_15535 (I267152,I3035,I266920,I266885,);
nor I_15536 (I266900,I267144,I267045);
nand I_15537 (I267197,I30993,I31008);
and I_15538 (I267214,I267197,I31005);
DFFARX1 I_15539 (I267214,I3035,I266920,I267240,);
nor I_15540 (I266888,I267240,I267144);
not I_15541 (I267262,I267240);
nor I_15542 (I267279,I267262,I267053);
nor I_15543 (I267296,I266985,I267279);
DFFARX1 I_15544 (I267296,I3035,I266920,I266903,);
nor I_15545 (I267327,I267262,I267144);
nor I_15546 (I267344,I31017,I31008);
nor I_15547 (I266894,I267344,I267327);
not I_15548 (I267375,I267344);
nand I_15549 (I266897,I267104,I267375);
DFFARX1 I_15550 (I267344,I3035,I266920,I266909,);
DFFARX1 I_15551 (I267344,I3035,I266920,I266906,);
not I_15552 (I267464,I3042);
DFFARX1 I_15553 (I703200,I3035,I267464,I267490,);
DFFARX1 I_15554 (I267490,I3035,I267464,I267507,);
not I_15555 (I267456,I267507);
not I_15556 (I267529,I267490);
nand I_15557 (I267546,I703176,I703197);
and I_15558 (I267563,I267546,I703194);
DFFARX1 I_15559 (I267563,I3035,I267464,I267589,);
not I_15560 (I267597,I267589);
DFFARX1 I_15561 (I703173,I3035,I267464,I267623,);
and I_15562 (I267631,I267623,I703185);
nand I_15563 (I267648,I267623,I703185);
nand I_15564 (I267435,I267597,I267648);
DFFARX1 I_15565 (I703188,I3035,I267464,I267688,);
nor I_15566 (I267696,I267688,I267631);
DFFARX1 I_15567 (I267696,I3035,I267464,I267429,);
nor I_15568 (I267444,I267688,I267589);
nand I_15569 (I267741,I703191,I703179);
and I_15570 (I267758,I267741,I703182);
DFFARX1 I_15571 (I267758,I3035,I267464,I267784,);
nor I_15572 (I267432,I267784,I267688);
not I_15573 (I267806,I267784);
nor I_15574 (I267823,I267806,I267597);
nor I_15575 (I267840,I267529,I267823);
DFFARX1 I_15576 (I267840,I3035,I267464,I267447,);
nor I_15577 (I267871,I267806,I267688);
nor I_15578 (I267888,I703173,I703179);
nor I_15579 (I267438,I267888,I267871);
not I_15580 (I267919,I267888);
nand I_15581 (I267441,I267648,I267919);
DFFARX1 I_15582 (I267888,I3035,I267464,I267453,);
DFFARX1 I_15583 (I267888,I3035,I267464,I267450,);
not I_15584 (I268008,I3042);
DFFARX1 I_15585 (I166130,I3035,I268008,I268034,);
DFFARX1 I_15586 (I268034,I3035,I268008,I268051,);
not I_15587 (I268000,I268051);
not I_15588 (I268073,I268034);
nand I_15589 (I268090,I166109,I166133);
and I_15590 (I268107,I268090,I166136);
DFFARX1 I_15591 (I268107,I3035,I268008,I268133,);
not I_15592 (I268141,I268133);
DFFARX1 I_15593 (I166118,I3035,I268008,I268167,);
and I_15594 (I268175,I268167,I166124);
nand I_15595 (I268192,I268167,I166124);
nand I_15596 (I267979,I268141,I268192);
DFFARX1 I_15597 (I166112,I3035,I268008,I268232,);
nor I_15598 (I268240,I268232,I268175);
DFFARX1 I_15599 (I268240,I3035,I268008,I267973,);
nor I_15600 (I267988,I268232,I268133);
nand I_15601 (I268285,I166121,I166109);
and I_15602 (I268302,I268285,I166115);
DFFARX1 I_15603 (I268302,I3035,I268008,I268328,);
nor I_15604 (I267976,I268328,I268232);
not I_15605 (I268350,I268328);
nor I_15606 (I268367,I268350,I268141);
nor I_15607 (I268384,I268073,I268367);
DFFARX1 I_15608 (I268384,I3035,I268008,I267991,);
nor I_15609 (I268415,I268350,I268232);
nor I_15610 (I268432,I166127,I166109);
nor I_15611 (I267982,I268432,I268415);
not I_15612 (I268463,I268432);
nand I_15613 (I267985,I268192,I268463);
DFFARX1 I_15614 (I268432,I3035,I268008,I267997,);
DFFARX1 I_15615 (I268432,I3035,I268008,I267994,);
not I_15616 (I268552,I3042);
DFFARX1 I_15617 (I688112,I3035,I268552,I268578,);
DFFARX1 I_15618 (I268578,I3035,I268552,I268595,);
not I_15619 (I268544,I268595);
not I_15620 (I268617,I268578);
nand I_15621 (I268634,I688109,I688106);
and I_15622 (I268651,I268634,I688094);
DFFARX1 I_15623 (I268651,I3035,I268552,I268677,);
not I_15624 (I268685,I268677);
DFFARX1 I_15625 (I688118,I3035,I268552,I268711,);
and I_15626 (I268719,I268711,I688103);
nand I_15627 (I268736,I268711,I688103);
nand I_15628 (I268523,I268685,I268736);
DFFARX1 I_15629 (I688097,I3035,I268552,I268776,);
nor I_15630 (I268784,I268776,I268719);
DFFARX1 I_15631 (I268784,I3035,I268552,I268517,);
nor I_15632 (I268532,I268776,I268677);
nand I_15633 (I268829,I688094,I688100);
and I_15634 (I268846,I268829,I688115);
DFFARX1 I_15635 (I268846,I3035,I268552,I268872,);
nor I_15636 (I268520,I268872,I268776);
not I_15637 (I268894,I268872);
nor I_15638 (I268911,I268894,I268685);
nor I_15639 (I268928,I268617,I268911);
DFFARX1 I_15640 (I268928,I3035,I268552,I268535,);
nor I_15641 (I268959,I268894,I268776);
nor I_15642 (I268976,I688097,I688100);
nor I_15643 (I268526,I268976,I268959);
not I_15644 (I269007,I268976);
nand I_15645 (I268529,I268736,I269007);
DFFARX1 I_15646 (I268976,I3035,I268552,I268541,);
DFFARX1 I_15647 (I268976,I3035,I268552,I268538,);
not I_15648 (I269096,I3042);
DFFARX1 I_15649 (I493518,I3035,I269096,I269122,);
DFFARX1 I_15650 (I269122,I3035,I269096,I269139,);
not I_15651 (I269088,I269139);
not I_15652 (I269161,I269122);
nand I_15653 (I269178,I493533,I493521);
and I_15654 (I269195,I269178,I493512);
DFFARX1 I_15655 (I269195,I3035,I269096,I269221,);
not I_15656 (I269229,I269221);
DFFARX1 I_15657 (I493524,I3035,I269096,I269255,);
and I_15658 (I269263,I269255,I493515);
nand I_15659 (I269280,I269255,I493515);
nand I_15660 (I269067,I269229,I269280);
DFFARX1 I_15661 (I493530,I3035,I269096,I269320,);
nor I_15662 (I269328,I269320,I269263);
DFFARX1 I_15663 (I269328,I3035,I269096,I269061,);
nor I_15664 (I269076,I269320,I269221);
nand I_15665 (I269373,I493539,I493527);
and I_15666 (I269390,I269373,I493536);
DFFARX1 I_15667 (I269390,I3035,I269096,I269416,);
nor I_15668 (I269064,I269416,I269320);
not I_15669 (I269438,I269416);
nor I_15670 (I269455,I269438,I269229);
nor I_15671 (I269472,I269161,I269455);
DFFARX1 I_15672 (I269472,I3035,I269096,I269079,);
nor I_15673 (I269503,I269438,I269320);
nor I_15674 (I269520,I493512,I493527);
nor I_15675 (I269070,I269520,I269503);
not I_15676 (I269551,I269520);
nand I_15677 (I269073,I269280,I269551);
DFFARX1 I_15678 (I269520,I3035,I269096,I269085,);
DFFARX1 I_15679 (I269520,I3035,I269096,I269082,);
not I_15680 (I269640,I3042);
DFFARX1 I_15681 (I557143,I3035,I269640,I269666,);
DFFARX1 I_15682 (I269666,I3035,I269640,I269683,);
not I_15683 (I269632,I269683);
not I_15684 (I269705,I269666);
nand I_15685 (I269722,I557143,I557161);
and I_15686 (I269739,I269722,I557155);
DFFARX1 I_15687 (I269739,I3035,I269640,I269765,);
not I_15688 (I269773,I269765);
DFFARX1 I_15689 (I557149,I3035,I269640,I269799,);
and I_15690 (I269807,I269799,I557158);
nand I_15691 (I269824,I269799,I557158);
nand I_15692 (I269611,I269773,I269824);
DFFARX1 I_15693 (I557146,I3035,I269640,I269864,);
nor I_15694 (I269872,I269864,I269807);
DFFARX1 I_15695 (I269872,I3035,I269640,I269605,);
nor I_15696 (I269620,I269864,I269765);
nand I_15697 (I269917,I557146,I557164);
and I_15698 (I269934,I269917,I557149);
DFFARX1 I_15699 (I269934,I3035,I269640,I269960,);
nor I_15700 (I269608,I269960,I269864);
not I_15701 (I269982,I269960);
nor I_15702 (I269999,I269982,I269773);
nor I_15703 (I270016,I269705,I269999);
DFFARX1 I_15704 (I270016,I3035,I269640,I269623,);
nor I_15705 (I270047,I269982,I269864);
nor I_15706 (I270064,I557152,I557164);
nor I_15707 (I269614,I270064,I270047);
not I_15708 (I270095,I270064);
nand I_15709 (I269617,I269824,I270095);
DFFARX1 I_15710 (I270064,I3035,I269640,I269629,);
DFFARX1 I_15711 (I270064,I3035,I269640,I269626,);
not I_15712 (I270184,I3042);
DFFARX1 I_15713 (I640497,I3035,I270184,I270210,);
DFFARX1 I_15714 (I270210,I3035,I270184,I270227,);
not I_15715 (I270176,I270227);
not I_15716 (I270249,I270210);
nand I_15717 (I270266,I640509,I640497);
and I_15718 (I270283,I270266,I640500);
DFFARX1 I_15719 (I270283,I3035,I270184,I270309,);
not I_15720 (I270317,I270309);
DFFARX1 I_15721 (I640518,I3035,I270184,I270343,);
and I_15722 (I270351,I270343,I640494);
nand I_15723 (I270368,I270343,I640494);
nand I_15724 (I270155,I270317,I270368);
DFFARX1 I_15725 (I640512,I3035,I270184,I270408,);
nor I_15726 (I270416,I270408,I270351);
DFFARX1 I_15727 (I270416,I3035,I270184,I270149,);
nor I_15728 (I270164,I270408,I270309);
nand I_15729 (I270461,I640506,I640503);
and I_15730 (I270478,I270461,I640515);
DFFARX1 I_15731 (I270478,I3035,I270184,I270504,);
nor I_15732 (I270152,I270504,I270408);
not I_15733 (I270526,I270504);
nor I_15734 (I270543,I270526,I270317);
nor I_15735 (I270560,I270249,I270543);
DFFARX1 I_15736 (I270560,I3035,I270184,I270167,);
nor I_15737 (I270591,I270526,I270408);
nor I_15738 (I270608,I640494,I640503);
nor I_15739 (I270158,I270608,I270591);
not I_15740 (I270639,I270608);
nand I_15741 (I270161,I270368,I270639);
DFFARX1 I_15742 (I270608,I3035,I270184,I270173,);
DFFARX1 I_15743 (I270608,I3035,I270184,I270170,);
not I_15744 (I270728,I3042);
DFFARX1 I_15745 (I354489,I3035,I270728,I270754,);
DFFARX1 I_15746 (I270754,I3035,I270728,I270771,);
not I_15747 (I270720,I270771);
not I_15748 (I270793,I270754);
nand I_15749 (I270810,I354510,I354501);
and I_15750 (I270827,I270810,I354489);
DFFARX1 I_15751 (I270827,I3035,I270728,I270853,);
not I_15752 (I270861,I270853);
DFFARX1 I_15753 (I354495,I3035,I270728,I270887,);
and I_15754 (I270895,I270887,I354492);
nand I_15755 (I270912,I270887,I354492);
nand I_15756 (I270699,I270861,I270912);
DFFARX1 I_15757 (I354486,I3035,I270728,I270952,);
nor I_15758 (I270960,I270952,I270895);
DFFARX1 I_15759 (I270960,I3035,I270728,I270693,);
nor I_15760 (I270708,I270952,I270853);
nand I_15761 (I271005,I354486,I354498);
and I_15762 (I271022,I271005,I354507);
DFFARX1 I_15763 (I271022,I3035,I270728,I271048,);
nor I_15764 (I270696,I271048,I270952);
not I_15765 (I271070,I271048);
nor I_15766 (I271087,I271070,I270861);
nor I_15767 (I271104,I270793,I271087);
DFFARX1 I_15768 (I271104,I3035,I270728,I270711,);
nor I_15769 (I271135,I271070,I270952);
nor I_15770 (I271152,I354504,I354498);
nor I_15771 (I270702,I271152,I271135);
not I_15772 (I271183,I271152);
nand I_15773 (I270705,I270912,I271183);
DFFARX1 I_15774 (I271152,I3035,I270728,I270717,);
DFFARX1 I_15775 (I271152,I3035,I270728,I270714,);
not I_15776 (I271272,I3042);
DFFARX1 I_15777 (I310561,I3035,I271272,I271298,);
DFFARX1 I_15778 (I271298,I3035,I271272,I271315,);
not I_15779 (I271264,I271315);
not I_15780 (I271337,I271298);
nand I_15781 (I271354,I310558,I310579);
and I_15782 (I271371,I271354,I310582);
DFFARX1 I_15783 (I271371,I3035,I271272,I271397,);
not I_15784 (I271405,I271397);
DFFARX1 I_15785 (I310567,I3035,I271272,I271431,);
and I_15786 (I271439,I271431,I310570);
nand I_15787 (I271456,I271431,I310570);
nand I_15788 (I271243,I271405,I271456);
DFFARX1 I_15789 (I310573,I3035,I271272,I271496,);
nor I_15790 (I271504,I271496,I271439);
DFFARX1 I_15791 (I271504,I3035,I271272,I271237,);
nor I_15792 (I271252,I271496,I271397);
nand I_15793 (I271549,I310558,I310564);
and I_15794 (I271566,I271549,I310576);
DFFARX1 I_15795 (I271566,I3035,I271272,I271592,);
nor I_15796 (I271240,I271592,I271496);
not I_15797 (I271614,I271592);
nor I_15798 (I271631,I271614,I271405);
nor I_15799 (I271648,I271337,I271631);
DFFARX1 I_15800 (I271648,I3035,I271272,I271255,);
nor I_15801 (I271679,I271614,I271496);
nor I_15802 (I271696,I310561,I310564);
nor I_15803 (I271246,I271696,I271679);
not I_15804 (I271727,I271696);
nand I_15805 (I271249,I271456,I271727);
DFFARX1 I_15806 (I271696,I3035,I271272,I271261,);
DFFARX1 I_15807 (I271696,I3035,I271272,I271258,);
not I_15808 (I271816,I3042);
DFFARX1 I_15809 (I144953,I3035,I271816,I271842,);
DFFARX1 I_15810 (I271842,I3035,I271816,I271859,);
not I_15811 (I271808,I271859);
not I_15812 (I271881,I271842);
nand I_15813 (I271898,I144965,I144944);
and I_15814 (I271915,I271898,I144947);
DFFARX1 I_15815 (I271915,I3035,I271816,I271941,);
not I_15816 (I271949,I271941);
DFFARX1 I_15817 (I144956,I3035,I271816,I271975,);
and I_15818 (I271983,I271975,I144968);
nand I_15819 (I272000,I271975,I144968);
nand I_15820 (I271787,I271949,I272000);
DFFARX1 I_15821 (I144962,I3035,I271816,I272040,);
nor I_15822 (I272048,I272040,I271983);
DFFARX1 I_15823 (I272048,I3035,I271816,I271781,);
nor I_15824 (I271796,I272040,I271941);
nand I_15825 (I272093,I144950,I144947);
and I_15826 (I272110,I272093,I144959);
DFFARX1 I_15827 (I272110,I3035,I271816,I272136,);
nor I_15828 (I271784,I272136,I272040);
not I_15829 (I272158,I272136);
nor I_15830 (I272175,I272158,I271949);
nor I_15831 (I272192,I271881,I272175);
DFFARX1 I_15832 (I272192,I3035,I271816,I271799,);
nor I_15833 (I272223,I272158,I272040);
nor I_15834 (I272240,I144944,I144947);
nor I_15835 (I271790,I272240,I272223);
not I_15836 (I272271,I272240);
nand I_15837 (I271793,I272000,I272271);
DFFARX1 I_15838 (I272240,I3035,I271816,I271805,);
DFFARX1 I_15839 (I272240,I3035,I271816,I271802,);
not I_15840 (I272360,I3042);
DFFARX1 I_15841 (I456702,I3035,I272360,I272386,);
DFFARX1 I_15842 (I272386,I3035,I272360,I272403,);
not I_15843 (I272352,I272403);
not I_15844 (I272425,I272386);
nand I_15845 (I272442,I456696,I456693);
and I_15846 (I272459,I272442,I456708);
DFFARX1 I_15847 (I272459,I3035,I272360,I272485,);
not I_15848 (I272493,I272485);
DFFARX1 I_15849 (I456696,I3035,I272360,I272519,);
and I_15850 (I272527,I272519,I456690);
nand I_15851 (I272544,I272519,I456690);
nand I_15852 (I272331,I272493,I272544);
DFFARX1 I_15853 (I456690,I3035,I272360,I272584,);
nor I_15854 (I272592,I272584,I272527);
DFFARX1 I_15855 (I272592,I3035,I272360,I272325,);
nor I_15856 (I272340,I272584,I272485);
nand I_15857 (I272637,I456705,I456699);
and I_15858 (I272654,I272637,I456693);
DFFARX1 I_15859 (I272654,I3035,I272360,I272680,);
nor I_15860 (I272328,I272680,I272584);
not I_15861 (I272702,I272680);
nor I_15862 (I272719,I272702,I272493);
nor I_15863 (I272736,I272425,I272719);
DFFARX1 I_15864 (I272736,I3035,I272360,I272343,);
nor I_15865 (I272767,I272702,I272584);
nor I_15866 (I272784,I456711,I456699);
nor I_15867 (I272334,I272784,I272767);
not I_15868 (I272815,I272784);
nand I_15869 (I272337,I272544,I272815);
DFFARX1 I_15870 (I272784,I3035,I272360,I272349,);
DFFARX1 I_15871 (I272784,I3035,I272360,I272346,);
not I_15872 (I272904,I3042);
DFFARX1 I_15873 (I98543,I3035,I272904,I272930,);
DFFARX1 I_15874 (I272930,I3035,I272904,I272947,);
not I_15875 (I272896,I272947);
not I_15876 (I272969,I272930);
nand I_15877 (I272986,I98555,I98534);
and I_15878 (I273003,I272986,I98537);
DFFARX1 I_15879 (I273003,I3035,I272904,I273029,);
not I_15880 (I273037,I273029);
DFFARX1 I_15881 (I98546,I3035,I272904,I273063,);
and I_15882 (I273071,I273063,I98558);
nand I_15883 (I273088,I273063,I98558);
nand I_15884 (I272875,I273037,I273088);
DFFARX1 I_15885 (I98552,I3035,I272904,I273128,);
nor I_15886 (I273136,I273128,I273071);
DFFARX1 I_15887 (I273136,I3035,I272904,I272869,);
nor I_15888 (I272884,I273128,I273029);
nand I_15889 (I273181,I98540,I98537);
and I_15890 (I273198,I273181,I98549);
DFFARX1 I_15891 (I273198,I3035,I272904,I273224,);
nor I_15892 (I272872,I273224,I273128);
not I_15893 (I273246,I273224);
nor I_15894 (I273263,I273246,I273037);
nor I_15895 (I273280,I272969,I273263);
DFFARX1 I_15896 (I273280,I3035,I272904,I272887,);
nor I_15897 (I273311,I273246,I273128);
nor I_15898 (I273328,I98534,I98537);
nor I_15899 (I272878,I273328,I273311);
not I_15900 (I273359,I273328);
nand I_15901 (I272881,I273088,I273359);
DFFARX1 I_15902 (I273328,I3035,I272904,I272893,);
DFFARX1 I_15903 (I273328,I3035,I272904,I272890,);
not I_15904 (I273448,I3042);
DFFARX1 I_15905 (I401307,I3035,I273448,I273474,);
DFFARX1 I_15906 (I273474,I3035,I273448,I273491,);
not I_15907 (I273440,I273491);
not I_15908 (I273513,I273474);
nand I_15909 (I273530,I401328,I401319);
and I_15910 (I273547,I273530,I401307);
DFFARX1 I_15911 (I273547,I3035,I273448,I273573,);
not I_15912 (I273581,I273573);
DFFARX1 I_15913 (I401313,I3035,I273448,I273607,);
and I_15914 (I273615,I273607,I401310);
nand I_15915 (I273632,I273607,I401310);
nand I_15916 (I273419,I273581,I273632);
DFFARX1 I_15917 (I401304,I3035,I273448,I273672,);
nor I_15918 (I273680,I273672,I273615);
DFFARX1 I_15919 (I273680,I3035,I273448,I273413,);
nor I_15920 (I273428,I273672,I273573);
nand I_15921 (I273725,I401304,I401316);
and I_15922 (I273742,I273725,I401325);
DFFARX1 I_15923 (I273742,I3035,I273448,I273768,);
nor I_15924 (I273416,I273768,I273672);
not I_15925 (I273790,I273768);
nor I_15926 (I273807,I273790,I273581);
nor I_15927 (I273824,I273513,I273807);
DFFARX1 I_15928 (I273824,I3035,I273448,I273431,);
nor I_15929 (I273855,I273790,I273672);
nor I_15930 (I273872,I401322,I401316);
nor I_15931 (I273422,I273872,I273855);
not I_15932 (I273903,I273872);
nand I_15933 (I273425,I273632,I273903);
DFFARX1 I_15934 (I273872,I3035,I273448,I273437,);
DFFARX1 I_15935 (I273872,I3035,I273448,I273434,);
not I_15936 (I273992,I3042);
DFFARX1 I_15937 (I478660,I3035,I273992,I274018,);
DFFARX1 I_15938 (I274018,I3035,I273992,I274035,);
not I_15939 (I273984,I274035);
not I_15940 (I274057,I274018);
nand I_15941 (I274074,I478675,I478663);
and I_15942 (I274091,I274074,I478654);
DFFARX1 I_15943 (I274091,I3035,I273992,I274117,);
not I_15944 (I274125,I274117);
DFFARX1 I_15945 (I478666,I3035,I273992,I274151,);
and I_15946 (I274159,I274151,I478657);
nand I_15947 (I274176,I274151,I478657);
nand I_15948 (I273963,I274125,I274176);
DFFARX1 I_15949 (I478672,I3035,I273992,I274216,);
nor I_15950 (I274224,I274216,I274159);
DFFARX1 I_15951 (I274224,I3035,I273992,I273957,);
nor I_15952 (I273972,I274216,I274117);
nand I_15953 (I274269,I478681,I478669);
and I_15954 (I274286,I274269,I478678);
DFFARX1 I_15955 (I274286,I3035,I273992,I274312,);
nor I_15956 (I273960,I274312,I274216);
not I_15957 (I274334,I274312);
nor I_15958 (I274351,I274334,I274125);
nor I_15959 (I274368,I274057,I274351);
DFFARX1 I_15960 (I274368,I3035,I273992,I273975,);
nor I_15961 (I274399,I274334,I274216);
nor I_15962 (I274416,I478654,I478669);
nor I_15963 (I273966,I274416,I274399);
not I_15964 (I274447,I274416);
nand I_15965 (I273969,I274176,I274447);
DFFARX1 I_15966 (I274416,I3035,I273992,I273981,);
DFFARX1 I_15967 (I274416,I3035,I273992,I273978,);
not I_15968 (I274536,I3042);
DFFARX1 I_15969 (I602349,I3035,I274536,I274562,);
DFFARX1 I_15970 (I274562,I3035,I274536,I274579,);
not I_15971 (I274528,I274579);
not I_15972 (I274601,I274562);
nand I_15973 (I274618,I602361,I602349);
and I_15974 (I274635,I274618,I602352);
DFFARX1 I_15975 (I274635,I3035,I274536,I274661,);
not I_15976 (I274669,I274661);
DFFARX1 I_15977 (I602370,I3035,I274536,I274695,);
and I_15978 (I274703,I274695,I602346);
nand I_15979 (I274720,I274695,I602346);
nand I_15980 (I274507,I274669,I274720);
DFFARX1 I_15981 (I602364,I3035,I274536,I274760,);
nor I_15982 (I274768,I274760,I274703);
DFFARX1 I_15983 (I274768,I3035,I274536,I274501,);
nor I_15984 (I274516,I274760,I274661);
nand I_15985 (I274813,I602358,I602355);
and I_15986 (I274830,I274813,I602367);
DFFARX1 I_15987 (I274830,I3035,I274536,I274856,);
nor I_15988 (I274504,I274856,I274760);
not I_15989 (I274878,I274856);
nor I_15990 (I274895,I274878,I274669);
nor I_15991 (I274912,I274601,I274895);
DFFARX1 I_15992 (I274912,I3035,I274536,I274519,);
nor I_15993 (I274943,I274878,I274760);
nor I_15994 (I274960,I602346,I602355);
nor I_15995 (I274510,I274960,I274943);
not I_15996 (I274991,I274960);
nand I_15997 (I274513,I274720,I274991);
DFFARX1 I_15998 (I274960,I3035,I274536,I274525,);
DFFARX1 I_15999 (I274960,I3035,I274536,I274522,);
not I_16000 (I275080,I3042);
DFFARX1 I_16001 (I610441,I3035,I275080,I275106,);
DFFARX1 I_16002 (I275106,I3035,I275080,I275123,);
not I_16003 (I275072,I275123);
not I_16004 (I275145,I275106);
nand I_16005 (I275162,I610453,I610441);
and I_16006 (I275179,I275162,I610444);
DFFARX1 I_16007 (I275179,I3035,I275080,I275205,);
not I_16008 (I275213,I275205);
DFFARX1 I_16009 (I610462,I3035,I275080,I275239,);
and I_16010 (I275247,I275239,I610438);
nand I_16011 (I275264,I275239,I610438);
nand I_16012 (I275051,I275213,I275264);
DFFARX1 I_16013 (I610456,I3035,I275080,I275304,);
nor I_16014 (I275312,I275304,I275247);
DFFARX1 I_16015 (I275312,I3035,I275080,I275045,);
nor I_16016 (I275060,I275304,I275205);
nand I_16017 (I275357,I610450,I610447);
and I_16018 (I275374,I275357,I610459);
DFFARX1 I_16019 (I275374,I3035,I275080,I275400,);
nor I_16020 (I275048,I275400,I275304);
not I_16021 (I275422,I275400);
nor I_16022 (I275439,I275422,I275213);
nor I_16023 (I275456,I275145,I275439);
DFFARX1 I_16024 (I275456,I3035,I275080,I275063,);
nor I_16025 (I275487,I275422,I275304);
nor I_16026 (I275504,I610438,I610447);
nor I_16027 (I275054,I275504,I275487);
not I_16028 (I275535,I275504);
nand I_16029 (I275057,I275264,I275535);
DFFARX1 I_16030 (I275504,I3035,I275080,I275069,);
DFFARX1 I_16031 (I275504,I3035,I275080,I275066,);
not I_16032 (I275624,I3042);
DFFARX1 I_16033 (I656681,I3035,I275624,I275650,);
DFFARX1 I_16034 (I275650,I3035,I275624,I275667,);
not I_16035 (I275616,I275667);
not I_16036 (I275689,I275650);
nand I_16037 (I275706,I656693,I656696);
and I_16038 (I275723,I275706,I656699);
DFFARX1 I_16039 (I275723,I3035,I275624,I275749,);
not I_16040 (I275757,I275749);
DFFARX1 I_16041 (I656684,I3035,I275624,I275783,);
and I_16042 (I275791,I275783,I656690);
nand I_16043 (I275808,I275783,I656690);
nand I_16044 (I275595,I275757,I275808);
DFFARX1 I_16045 (I656678,I3035,I275624,I275848,);
nor I_16046 (I275856,I275848,I275791);
DFFARX1 I_16047 (I275856,I3035,I275624,I275589,);
nor I_16048 (I275604,I275848,I275749);
nand I_16049 (I275901,I656681,I656702);
and I_16050 (I275918,I275901,I656687);
DFFARX1 I_16051 (I275918,I3035,I275624,I275944,);
nor I_16052 (I275592,I275944,I275848);
not I_16053 (I275966,I275944);
nor I_16054 (I275983,I275966,I275757);
nor I_16055 (I276000,I275689,I275983);
DFFARX1 I_16056 (I276000,I3035,I275624,I275607,);
nor I_16057 (I276031,I275966,I275848);
nor I_16058 (I276048,I656678,I656702);
nor I_16059 (I275598,I276048,I276031);
not I_16060 (I276079,I276048);
nand I_16061 (I275601,I275808,I276079);
DFFARX1 I_16062 (I276048,I3035,I275624,I275613,);
DFFARX1 I_16063 (I276048,I3035,I275624,I275610,);
not I_16064 (I276168,I3042);
DFFARX1 I_16065 (I20992,I3035,I276168,I276194,);
DFFARX1 I_16066 (I276194,I3035,I276168,I276211,);
not I_16067 (I276160,I276211);
not I_16068 (I276233,I276194);
nand I_16069 (I276250,I20980,I20995);
and I_16070 (I276267,I276250,I20983);
DFFARX1 I_16071 (I276267,I3035,I276168,I276293,);
not I_16072 (I276301,I276293);
DFFARX1 I_16073 (I21004,I3035,I276168,I276327,);
and I_16074 (I276335,I276327,I20998);
nand I_16075 (I276352,I276327,I20998);
nand I_16076 (I276139,I276301,I276352);
DFFARX1 I_16077 (I21001,I3035,I276168,I276392,);
nor I_16078 (I276400,I276392,I276335);
DFFARX1 I_16079 (I276400,I3035,I276168,I276133,);
nor I_16080 (I276148,I276392,I276293);
nand I_16081 (I276445,I20980,I20983);
and I_16082 (I276462,I276445,I20986);
DFFARX1 I_16083 (I276462,I3035,I276168,I276488,);
nor I_16084 (I276136,I276488,I276392);
not I_16085 (I276510,I276488);
nor I_16086 (I276527,I276510,I276301);
nor I_16087 (I276544,I276233,I276527);
DFFARX1 I_16088 (I276544,I3035,I276168,I276151,);
nor I_16089 (I276575,I276510,I276392);
nor I_16090 (I276592,I20989,I20983);
nor I_16091 (I276142,I276592,I276575);
not I_16092 (I276623,I276592);
nand I_16093 (I276145,I276352,I276623);
DFFARX1 I_16094 (I276592,I3035,I276168,I276157,);
DFFARX1 I_16095 (I276592,I3035,I276168,I276154,);
not I_16096 (I276712,I3042);
DFFARX1 I_16097 (I122343,I3035,I276712,I276738,);
DFFARX1 I_16098 (I276738,I3035,I276712,I276755,);
not I_16099 (I276704,I276755);
not I_16100 (I276777,I276738);
nand I_16101 (I276794,I122355,I122334);
and I_16102 (I276811,I276794,I122337);
DFFARX1 I_16103 (I276811,I3035,I276712,I276837,);
not I_16104 (I276845,I276837);
DFFARX1 I_16105 (I122346,I3035,I276712,I276871,);
and I_16106 (I276879,I276871,I122358);
nand I_16107 (I276896,I276871,I122358);
nand I_16108 (I276683,I276845,I276896);
DFFARX1 I_16109 (I122352,I3035,I276712,I276936,);
nor I_16110 (I276944,I276936,I276879);
DFFARX1 I_16111 (I276944,I3035,I276712,I276677,);
nor I_16112 (I276692,I276936,I276837);
nand I_16113 (I276989,I122340,I122337);
and I_16114 (I277006,I276989,I122349);
DFFARX1 I_16115 (I277006,I3035,I276712,I277032,);
nor I_16116 (I276680,I277032,I276936);
not I_16117 (I277054,I277032);
nor I_16118 (I277071,I277054,I276845);
nor I_16119 (I277088,I276777,I277071);
DFFARX1 I_16120 (I277088,I3035,I276712,I276695,);
nor I_16121 (I277119,I277054,I276936);
nor I_16122 (I277136,I122334,I122337);
nor I_16123 (I276686,I277136,I277119);
not I_16124 (I277167,I277136);
nand I_16125 (I276689,I276896,I277167);
DFFARX1 I_16126 (I277136,I3035,I276712,I276701,);
DFFARX1 I_16127 (I277136,I3035,I276712,I276698,);
not I_16128 (I277256,I3042);
DFFARX1 I_16129 (I158225,I3035,I277256,I277282,);
DFFARX1 I_16130 (I277282,I3035,I277256,I277299,);
not I_16131 (I277248,I277299);
not I_16132 (I277321,I277282);
nand I_16133 (I277338,I158204,I158228);
and I_16134 (I277355,I277338,I158231);
DFFARX1 I_16135 (I277355,I3035,I277256,I277381,);
not I_16136 (I277389,I277381);
DFFARX1 I_16137 (I158213,I3035,I277256,I277415,);
and I_16138 (I277423,I277415,I158219);
nand I_16139 (I277440,I277415,I158219);
nand I_16140 (I277227,I277389,I277440);
DFFARX1 I_16141 (I158207,I3035,I277256,I277480,);
nor I_16142 (I277488,I277480,I277423);
DFFARX1 I_16143 (I277488,I3035,I277256,I277221,);
nor I_16144 (I277236,I277480,I277381);
nand I_16145 (I277533,I158216,I158204);
and I_16146 (I277550,I277533,I158210);
DFFARX1 I_16147 (I277550,I3035,I277256,I277576,);
nor I_16148 (I277224,I277576,I277480);
not I_16149 (I277598,I277576);
nor I_16150 (I277615,I277598,I277389);
nor I_16151 (I277632,I277321,I277615);
DFFARX1 I_16152 (I277632,I3035,I277256,I277239,);
nor I_16153 (I277663,I277598,I277480);
nor I_16154 (I277680,I158222,I158204);
nor I_16155 (I277230,I277680,I277663);
not I_16156 (I277711,I277680);
nand I_16157 (I277233,I277440,I277711);
DFFARX1 I_16158 (I277680,I3035,I277256,I277245,);
DFFARX1 I_16159 (I277680,I3035,I277256,I277242,);
not I_16160 (I277800,I3042);
DFFARX1 I_16161 (I51552,I3035,I277800,I277826,);
DFFARX1 I_16162 (I277826,I3035,I277800,I277843,);
not I_16163 (I277792,I277843);
not I_16164 (I277865,I277826);
nand I_16165 (I277882,I51567,I51546);
and I_16166 (I277899,I277882,I51549);
DFFARX1 I_16167 (I277899,I3035,I277800,I277925,);
not I_16168 (I277933,I277925);
DFFARX1 I_16169 (I51555,I3035,I277800,I277959,);
and I_16170 (I277967,I277959,I51549);
nand I_16171 (I277984,I277959,I51549);
nand I_16172 (I277771,I277933,I277984);
DFFARX1 I_16173 (I51564,I3035,I277800,I278024,);
nor I_16174 (I278032,I278024,I277967);
DFFARX1 I_16175 (I278032,I3035,I277800,I277765,);
nor I_16176 (I277780,I278024,I277925);
nand I_16177 (I278077,I51546,I51561);
and I_16178 (I278094,I278077,I51558);
DFFARX1 I_16179 (I278094,I3035,I277800,I278120,);
nor I_16180 (I277768,I278120,I278024);
not I_16181 (I278142,I278120);
nor I_16182 (I278159,I278142,I277933);
nor I_16183 (I278176,I277865,I278159);
DFFARX1 I_16184 (I278176,I3035,I277800,I277783,);
nor I_16185 (I278207,I278142,I278024);
nor I_16186 (I278224,I51570,I51561);
nor I_16187 (I277774,I278224,I278207);
not I_16188 (I278255,I278224);
nand I_16189 (I277777,I277984,I278255);
DFFARX1 I_16190 (I278224,I3035,I277800,I277789,);
DFFARX1 I_16191 (I278224,I3035,I277800,I277786,);
not I_16192 (I278344,I3042);
DFFARX1 I_16193 (I219884,I3035,I278344,I278370,);
DFFARX1 I_16194 (I278370,I3035,I278344,I278387,);
not I_16195 (I278336,I278387);
not I_16196 (I278409,I278370);
nand I_16197 (I278426,I219863,I219887);
and I_16198 (I278443,I278426,I219890);
DFFARX1 I_16199 (I278443,I3035,I278344,I278469,);
not I_16200 (I278477,I278469);
DFFARX1 I_16201 (I219872,I3035,I278344,I278503,);
and I_16202 (I278511,I278503,I219878);
nand I_16203 (I278528,I278503,I219878);
nand I_16204 (I278315,I278477,I278528);
DFFARX1 I_16205 (I219866,I3035,I278344,I278568,);
nor I_16206 (I278576,I278568,I278511);
DFFARX1 I_16207 (I278576,I3035,I278344,I278309,);
nor I_16208 (I278324,I278568,I278469);
nand I_16209 (I278621,I219875,I219863);
and I_16210 (I278638,I278621,I219869);
DFFARX1 I_16211 (I278638,I3035,I278344,I278664,);
nor I_16212 (I278312,I278664,I278568);
not I_16213 (I278686,I278664);
nor I_16214 (I278703,I278686,I278477);
nor I_16215 (I278720,I278409,I278703);
DFFARX1 I_16216 (I278720,I3035,I278344,I278327,);
nor I_16217 (I278751,I278686,I278568);
nor I_16218 (I278768,I219881,I219863);
nor I_16219 (I278318,I278768,I278751);
not I_16220 (I278799,I278768);
nand I_16221 (I278321,I278528,I278799);
DFFARX1 I_16222 (I278768,I3035,I278344,I278333,);
DFFARX1 I_16223 (I278768,I3035,I278344,I278330,);
not I_16224 (I278888,I3042);
DFFARX1 I_16225 (I712720,I3035,I278888,I278914,);
DFFARX1 I_16226 (I278914,I3035,I278888,I278931,);
not I_16227 (I278880,I278931);
not I_16228 (I278953,I278914);
nand I_16229 (I278970,I712696,I712717);
and I_16230 (I278987,I278970,I712714);
DFFARX1 I_16231 (I278987,I3035,I278888,I279013,);
not I_16232 (I279021,I279013);
DFFARX1 I_16233 (I712693,I3035,I278888,I279047,);
and I_16234 (I279055,I279047,I712705);
nand I_16235 (I279072,I279047,I712705);
nand I_16236 (I278859,I279021,I279072);
DFFARX1 I_16237 (I712708,I3035,I278888,I279112,);
nor I_16238 (I279120,I279112,I279055);
DFFARX1 I_16239 (I279120,I3035,I278888,I278853,);
nor I_16240 (I278868,I279112,I279013);
nand I_16241 (I279165,I712711,I712699);
and I_16242 (I279182,I279165,I712702);
DFFARX1 I_16243 (I279182,I3035,I278888,I279208,);
nor I_16244 (I278856,I279208,I279112);
not I_16245 (I279230,I279208);
nor I_16246 (I279247,I279230,I279021);
nor I_16247 (I279264,I278953,I279247);
DFFARX1 I_16248 (I279264,I3035,I278888,I278871,);
nor I_16249 (I279295,I279230,I279112);
nor I_16250 (I279312,I712693,I712699);
nor I_16251 (I278862,I279312,I279295);
not I_16252 (I279343,I279312);
nand I_16253 (I278865,I279072,I279343);
DFFARX1 I_16254 (I279312,I3035,I278888,I278877,);
DFFARX1 I_16255 (I279312,I3035,I278888,I278874,);
not I_16256 (I279432,I3042);
DFFARX1 I_16257 (I490288,I3035,I279432,I279458,);
DFFARX1 I_16258 (I279458,I3035,I279432,I279475,);
not I_16259 (I279424,I279475);
not I_16260 (I279497,I279458);
nand I_16261 (I279514,I490303,I490291);
and I_16262 (I279531,I279514,I490282);
DFFARX1 I_16263 (I279531,I3035,I279432,I279557,);
not I_16264 (I279565,I279557);
DFFARX1 I_16265 (I490294,I3035,I279432,I279591,);
and I_16266 (I279599,I279591,I490285);
nand I_16267 (I279616,I279591,I490285);
nand I_16268 (I279403,I279565,I279616);
DFFARX1 I_16269 (I490300,I3035,I279432,I279656,);
nor I_16270 (I279664,I279656,I279599);
DFFARX1 I_16271 (I279664,I3035,I279432,I279397,);
nor I_16272 (I279412,I279656,I279557);
nand I_16273 (I279709,I490309,I490297);
and I_16274 (I279726,I279709,I490306);
DFFARX1 I_16275 (I279726,I3035,I279432,I279752,);
nor I_16276 (I279400,I279752,I279656);
not I_16277 (I279774,I279752);
nor I_16278 (I279791,I279774,I279565);
nor I_16279 (I279808,I279497,I279791);
DFFARX1 I_16280 (I279808,I3035,I279432,I279415,);
nor I_16281 (I279839,I279774,I279656);
nor I_16282 (I279856,I490282,I490297);
nor I_16283 (I279406,I279856,I279839);
not I_16284 (I279887,I279856);
nand I_16285 (I279409,I279616,I279887);
DFFARX1 I_16286 (I279856,I3035,I279432,I279421,);
DFFARX1 I_16287 (I279856,I3035,I279432,I279418,);
not I_16288 (I279973,I3042);
DFFARX1 I_16289 (I443524,I3035,I279973,I279999,);
DFFARX1 I_16290 (I279999,I3035,I279973,I280016,);
not I_16291 (I279965,I280016);
DFFARX1 I_16292 (I443521,I3035,I279973,I280047,);
not I_16293 (I280055,I443521);
nor I_16294 (I280072,I279999,I280055);
not I_16295 (I280089,I443518);
not I_16296 (I280106,I443533);
nand I_16297 (I280123,I280106,I443518);
nor I_16298 (I280140,I280055,I280123);
nor I_16299 (I280157,I280047,I280140);
DFFARX1 I_16300 (I280106,I3035,I279973,I279962,);
nor I_16301 (I280188,I443533,I443527);
nand I_16302 (I280205,I280188,I443515);
nor I_16303 (I280222,I280205,I280089);
nand I_16304 (I279947,I280222,I443521);
DFFARX1 I_16305 (I280205,I3035,I279973,I279959,);
nand I_16306 (I280267,I280089,I443533);
nor I_16307 (I280284,I280089,I443533);
nand I_16308 (I279953,I280072,I280284);
not I_16309 (I280315,I443536);
nor I_16310 (I280332,I280315,I280267);
DFFARX1 I_16311 (I280332,I3035,I279973,I279941,);
nor I_16312 (I280363,I280315,I443515);
and I_16313 (I280380,I280363,I443530);
or I_16314 (I280397,I280380,I443518);
DFFARX1 I_16315 (I280397,I3035,I279973,I280423,);
nor I_16316 (I280431,I280423,I280047);
nor I_16317 (I279950,I279999,I280431);
not I_16318 (I280462,I280423);
nor I_16319 (I280479,I280462,I280157);
DFFARX1 I_16320 (I280479,I3035,I279973,I279956,);
nand I_16321 (I280510,I280462,I280089);
nor I_16322 (I279944,I280315,I280510);
not I_16323 (I280568,I3042);
DFFARX1 I_16324 (I645136,I3035,I280568,I280594,);
DFFARX1 I_16325 (I280594,I3035,I280568,I280611,);
not I_16326 (I280560,I280611);
DFFARX1 I_16327 (I645118,I3035,I280568,I280642,);
not I_16328 (I280650,I645124);
nor I_16329 (I280667,I280594,I280650);
not I_16330 (I280684,I645139);
not I_16331 (I280701,I645130);
nand I_16332 (I280718,I280701,I645139);
nor I_16333 (I280735,I280650,I280718);
nor I_16334 (I280752,I280642,I280735);
DFFARX1 I_16335 (I280701,I3035,I280568,I280557,);
nor I_16336 (I280783,I645130,I645142);
nand I_16337 (I280800,I280783,I645121);
nor I_16338 (I280817,I280800,I280684);
nand I_16339 (I280542,I280817,I645124);
DFFARX1 I_16340 (I280800,I3035,I280568,I280554,);
nand I_16341 (I280862,I280684,I645130);
nor I_16342 (I280879,I280684,I645130);
nand I_16343 (I280548,I280667,I280879);
not I_16344 (I280910,I645127);
nor I_16345 (I280927,I280910,I280862);
DFFARX1 I_16346 (I280927,I3035,I280568,I280536,);
nor I_16347 (I280958,I280910,I645133);
and I_16348 (I280975,I280958,I645118);
or I_16349 (I280992,I280975,I645121);
DFFARX1 I_16350 (I280992,I3035,I280568,I281018,);
nor I_16351 (I281026,I281018,I280642);
nor I_16352 (I280545,I280594,I281026);
not I_16353 (I281057,I281018);
nor I_16354 (I281074,I281057,I280752);
DFFARX1 I_16355 (I281074,I3035,I280568,I280551,);
nand I_16356 (I281105,I281057,I280684);
nor I_16357 (I280539,I280910,I281105);
not I_16358 (I281163,I3042);
DFFARX1 I_16359 (I206176,I3035,I281163,I281189,);
DFFARX1 I_16360 (I281189,I3035,I281163,I281206,);
not I_16361 (I281155,I281206);
DFFARX1 I_16362 (I206164,I3035,I281163,I281237,);
not I_16363 (I281245,I206167);
nor I_16364 (I281262,I281189,I281245);
not I_16365 (I281279,I206170);
not I_16366 (I281296,I206182);
nand I_16367 (I281313,I281296,I206170);
nor I_16368 (I281330,I281245,I281313);
nor I_16369 (I281347,I281237,I281330);
DFFARX1 I_16370 (I281296,I3035,I281163,I281152,);
nor I_16371 (I281378,I206182,I206173);
nand I_16372 (I281395,I281378,I206161);
nor I_16373 (I281412,I281395,I281279);
nand I_16374 (I281137,I281412,I206167);
DFFARX1 I_16375 (I281395,I3035,I281163,I281149,);
nand I_16376 (I281457,I281279,I206182);
nor I_16377 (I281474,I281279,I206182);
nand I_16378 (I281143,I281262,I281474);
not I_16379 (I281505,I206179);
nor I_16380 (I281522,I281505,I281457);
DFFARX1 I_16381 (I281522,I3035,I281163,I281131,);
nor I_16382 (I281553,I281505,I206185);
and I_16383 (I281570,I281553,I206188);
or I_16384 (I281587,I281570,I206161);
DFFARX1 I_16385 (I281587,I3035,I281163,I281613,);
nor I_16386 (I281621,I281613,I281237);
nor I_16387 (I281140,I281189,I281621);
not I_16388 (I281652,I281613);
nor I_16389 (I281669,I281652,I281347);
DFFARX1 I_16390 (I281669,I3035,I281163,I281146,);
nand I_16391 (I281700,I281652,I281279);
nor I_16392 (I281134,I281505,I281700);
not I_16393 (I281758,I3042);
DFFARX1 I_16394 (I572886,I3035,I281758,I281784,);
DFFARX1 I_16395 (I281784,I3035,I281758,I281801,);
not I_16396 (I281750,I281801);
DFFARX1 I_16397 (I572868,I3035,I281758,I281832,);
not I_16398 (I281840,I572874);
nor I_16399 (I281857,I281784,I281840);
not I_16400 (I281874,I572889);
not I_16401 (I281891,I572880);
nand I_16402 (I281908,I281891,I572889);
nor I_16403 (I281925,I281840,I281908);
nor I_16404 (I281942,I281832,I281925);
DFFARX1 I_16405 (I281891,I3035,I281758,I281747,);
nor I_16406 (I281973,I572880,I572892);
nand I_16407 (I281990,I281973,I572871);
nor I_16408 (I282007,I281990,I281874);
nand I_16409 (I281732,I282007,I572874);
DFFARX1 I_16410 (I281990,I3035,I281758,I281744,);
nand I_16411 (I282052,I281874,I572880);
nor I_16412 (I282069,I281874,I572880);
nand I_16413 (I281738,I281857,I282069);
not I_16414 (I282100,I572877);
nor I_16415 (I282117,I282100,I282052);
DFFARX1 I_16416 (I282117,I3035,I281758,I281726,);
nor I_16417 (I282148,I282100,I572883);
and I_16418 (I282165,I282148,I572868);
or I_16419 (I282182,I282165,I572871);
DFFARX1 I_16420 (I282182,I3035,I281758,I282208,);
nor I_16421 (I282216,I282208,I281832);
nor I_16422 (I281735,I281784,I282216);
not I_16423 (I282247,I282208);
nor I_16424 (I282264,I282247,I281942);
DFFARX1 I_16425 (I282264,I3035,I281758,I281741,);
nand I_16426 (I282295,I282247,I281874);
nor I_16427 (I281729,I282100,I282295);
not I_16428 (I282353,I3042);
DFFARX1 I_16429 (I319809,I3035,I282353,I282379,);
DFFARX1 I_16430 (I282379,I3035,I282353,I282396,);
not I_16431 (I282345,I282396);
DFFARX1 I_16432 (I319821,I3035,I282353,I282427,);
not I_16433 (I282435,I319806);
nor I_16434 (I282452,I282379,I282435);
not I_16435 (I282469,I319824);
not I_16436 (I282486,I319815);
nand I_16437 (I282503,I282486,I319824);
nor I_16438 (I282520,I282435,I282503);
nor I_16439 (I282537,I282427,I282520);
DFFARX1 I_16440 (I282486,I3035,I282353,I282342,);
nor I_16441 (I282568,I319815,I319827);
nand I_16442 (I282585,I282568,I319830);
nor I_16443 (I282602,I282585,I282469);
nand I_16444 (I282327,I282602,I319806);
DFFARX1 I_16445 (I282585,I3035,I282353,I282339,);
nand I_16446 (I282647,I282469,I319815);
nor I_16447 (I282664,I282469,I319815);
nand I_16448 (I282333,I282452,I282664);
not I_16449 (I282695,I319806);
nor I_16450 (I282712,I282695,I282647);
DFFARX1 I_16451 (I282712,I3035,I282353,I282321,);
nor I_16452 (I282743,I282695,I319818);
and I_16453 (I282760,I282743,I319812);
or I_16454 (I282777,I282760,I319809);
DFFARX1 I_16455 (I282777,I3035,I282353,I282803,);
nor I_16456 (I282811,I282803,I282427);
nor I_16457 (I282330,I282379,I282811);
not I_16458 (I282842,I282803);
nor I_16459 (I282859,I282842,I282537);
DFFARX1 I_16460 (I282859,I3035,I282353,I282336,);
nand I_16461 (I282890,I282842,I282469);
nor I_16462 (I282324,I282695,I282890);
not I_16463 (I282948,I3042);
DFFARX1 I_16464 (I358541,I3035,I282948,I282974,);
DFFARX1 I_16465 (I282974,I3035,I282948,I282991,);
not I_16466 (I282940,I282991);
DFFARX1 I_16467 (I358535,I3035,I282948,I283022,);
not I_16468 (I283030,I358532);
nor I_16469 (I283047,I282974,I283030);
not I_16470 (I283064,I358544);
not I_16471 (I283081,I358547);
nand I_16472 (I283098,I283081,I358544);
nor I_16473 (I283115,I283030,I283098);
nor I_16474 (I283132,I283022,I283115);
DFFARX1 I_16475 (I283081,I3035,I282948,I282937,);
nor I_16476 (I283163,I358547,I358556);
nand I_16477 (I283180,I283163,I358550);
nor I_16478 (I283197,I283180,I283064);
nand I_16479 (I282922,I283197,I358532);
DFFARX1 I_16480 (I283180,I3035,I282948,I282934,);
nand I_16481 (I283242,I283064,I358547);
nor I_16482 (I283259,I283064,I358547);
nand I_16483 (I282928,I283047,I283259);
not I_16484 (I283290,I358538);
nor I_16485 (I283307,I283290,I283242);
DFFARX1 I_16486 (I283307,I3035,I282948,I282916,);
nor I_16487 (I283338,I283290,I358553);
and I_16488 (I283355,I283338,I358532);
or I_16489 (I283372,I283355,I358535);
DFFARX1 I_16490 (I283372,I3035,I282948,I283398,);
nor I_16491 (I283406,I283398,I283022);
nor I_16492 (I282925,I282974,I283406);
not I_16493 (I283437,I283398);
nor I_16494 (I283454,I283437,I283132);
DFFARX1 I_16495 (I283454,I3035,I282948,I282931,);
nand I_16496 (I283485,I283437,I283064);
nor I_16497 (I282919,I283290,I283485);
not I_16498 (I283543,I3042);
DFFARX1 I_16499 (I238597,I3035,I283543,I283569,);
DFFARX1 I_16500 (I283569,I3035,I283543,I283586,);
not I_16501 (I283535,I283586);
DFFARX1 I_16502 (I238621,I3035,I283543,I283617,);
not I_16503 (I283625,I238600);
nor I_16504 (I283642,I283569,I283625);
not I_16505 (I283659,I238606);
not I_16506 (I283676,I238612);
nand I_16507 (I283693,I283676,I238606);
nor I_16508 (I283710,I283625,I283693);
nor I_16509 (I283727,I283617,I283710);
DFFARX1 I_16510 (I283676,I3035,I283543,I283532,);
nor I_16511 (I283758,I238612,I238624);
nand I_16512 (I283775,I283758,I238618);
nor I_16513 (I283792,I283775,I283659);
nand I_16514 (I283517,I283792,I238600);
DFFARX1 I_16515 (I283775,I3035,I283543,I283529,);
nand I_16516 (I283837,I283659,I238612);
nor I_16517 (I283854,I283659,I238612);
nand I_16518 (I283523,I283642,I283854);
not I_16519 (I283885,I238603);
nor I_16520 (I283902,I283885,I283837);
DFFARX1 I_16521 (I283902,I3035,I283543,I283511,);
nor I_16522 (I283933,I283885,I238597);
and I_16523 (I283950,I283933,I238615);
or I_16524 (I283967,I283950,I238609);
DFFARX1 I_16525 (I283967,I3035,I283543,I283993,);
nor I_16526 (I284001,I283993,I283617);
nor I_16527 (I283520,I283569,I284001);
not I_16528 (I284032,I283993);
nor I_16529 (I284049,I284032,I283727);
DFFARX1 I_16530 (I284049,I3035,I283543,I283526,);
nand I_16531 (I284080,I284032,I283659);
nor I_16532 (I283514,I283885,I284080);
not I_16533 (I284138,I3042);
DFFARX1 I_16534 (I263621,I3035,I284138,I284164,);
DFFARX1 I_16535 (I284164,I3035,I284138,I284181,);
not I_16536 (I284130,I284181);
DFFARX1 I_16537 (I263645,I3035,I284138,I284212,);
not I_16538 (I284220,I263624);
nor I_16539 (I284237,I284164,I284220);
not I_16540 (I284254,I263630);
not I_16541 (I284271,I263636);
nand I_16542 (I284288,I284271,I263630);
nor I_16543 (I284305,I284220,I284288);
nor I_16544 (I284322,I284212,I284305);
DFFARX1 I_16545 (I284271,I3035,I284138,I284127,);
nor I_16546 (I284353,I263636,I263648);
nand I_16547 (I284370,I284353,I263642);
nor I_16548 (I284387,I284370,I284254);
nand I_16549 (I284112,I284387,I263624);
DFFARX1 I_16550 (I284370,I3035,I284138,I284124,);
nand I_16551 (I284432,I284254,I263636);
nor I_16552 (I284449,I284254,I263636);
nand I_16553 (I284118,I284237,I284449);
not I_16554 (I284480,I263627);
nor I_16555 (I284497,I284480,I284432);
DFFARX1 I_16556 (I284497,I3035,I284138,I284106,);
nor I_16557 (I284528,I284480,I263621);
and I_16558 (I284545,I284528,I263639);
or I_16559 (I284562,I284545,I263633);
DFFARX1 I_16560 (I284562,I3035,I284138,I284588,);
nor I_16561 (I284596,I284588,I284212);
nor I_16562 (I284115,I284164,I284596);
not I_16563 (I284627,I284588);
nor I_16564 (I284644,I284627,I284322);
DFFARX1 I_16565 (I284644,I3035,I284138,I284121,);
nand I_16566 (I284675,I284627,I284254);
nor I_16567 (I284109,I284480,I284675);
not I_16568 (I284733,I3042);
DFFARX1 I_16569 (I260357,I3035,I284733,I284759,);
DFFARX1 I_16570 (I284759,I3035,I284733,I284776,);
not I_16571 (I284725,I284776);
DFFARX1 I_16572 (I260381,I3035,I284733,I284807,);
not I_16573 (I284815,I260360);
nor I_16574 (I284832,I284759,I284815);
not I_16575 (I284849,I260366);
not I_16576 (I284866,I260372);
nand I_16577 (I284883,I284866,I260366);
nor I_16578 (I284900,I284815,I284883);
nor I_16579 (I284917,I284807,I284900);
DFFARX1 I_16580 (I284866,I3035,I284733,I284722,);
nor I_16581 (I284948,I260372,I260384);
nand I_16582 (I284965,I284948,I260378);
nor I_16583 (I284982,I284965,I284849);
nand I_16584 (I284707,I284982,I260360);
DFFARX1 I_16585 (I284965,I3035,I284733,I284719,);
nand I_16586 (I285027,I284849,I260372);
nor I_16587 (I285044,I284849,I260372);
nand I_16588 (I284713,I284832,I285044);
not I_16589 (I285075,I260363);
nor I_16590 (I285092,I285075,I285027);
DFFARX1 I_16591 (I285092,I3035,I284733,I284701,);
nor I_16592 (I285123,I285075,I260357);
and I_16593 (I285140,I285123,I260375);
or I_16594 (I285157,I285140,I260369);
DFFARX1 I_16595 (I285157,I3035,I284733,I285183,);
nor I_16596 (I285191,I285183,I284807);
nor I_16597 (I284710,I284759,I285191);
not I_16598 (I285222,I285183);
nor I_16599 (I285239,I285222,I284917);
DFFARX1 I_16600 (I285239,I3035,I284733,I284716,);
nand I_16601 (I285270,I285222,I284849);
nor I_16602 (I284704,I285075,I285270);
not I_16603 (I285328,I3042);
DFFARX1 I_16604 (I106269,I3035,I285328,I285354,);
DFFARX1 I_16605 (I285354,I3035,I285328,I285371,);
not I_16606 (I285320,I285371);
DFFARX1 I_16607 (I106293,I3035,I285328,I285402,);
not I_16608 (I285410,I106287);
nor I_16609 (I285427,I285354,I285410);
not I_16610 (I285444,I106281);
not I_16611 (I285461,I106278);
nand I_16612 (I285478,I285461,I106281);
nor I_16613 (I285495,I285410,I285478);
nor I_16614 (I285512,I285402,I285495);
DFFARX1 I_16615 (I285461,I3035,I285328,I285317,);
nor I_16616 (I285543,I106278,I106272);
nand I_16617 (I285560,I285543,I106290);
nor I_16618 (I285577,I285560,I285444);
nand I_16619 (I285302,I285577,I106287);
DFFARX1 I_16620 (I285560,I3035,I285328,I285314,);
nand I_16621 (I285622,I285444,I106278);
nor I_16622 (I285639,I285444,I106278);
nand I_16623 (I285308,I285427,I285639);
not I_16624 (I285670,I106284);
nor I_16625 (I285687,I285670,I285622);
DFFARX1 I_16626 (I285687,I3035,I285328,I285296,);
nor I_16627 (I285718,I285670,I106269);
and I_16628 (I285735,I285718,I106275);
or I_16629 (I285752,I285735,I106272);
DFFARX1 I_16630 (I285752,I3035,I285328,I285778,);
nor I_16631 (I285786,I285778,I285402);
nor I_16632 (I285305,I285354,I285786);
not I_16633 (I285817,I285778);
nor I_16634 (I285834,I285817,I285512);
DFFARX1 I_16635 (I285834,I3035,I285328,I285311,);
nand I_16636 (I285865,I285817,I285444);
nor I_16637 (I285299,I285670,I285865);
not I_16638 (I285923,I3042);
DFFARX1 I_16639 (I205649,I3035,I285923,I285949,);
DFFARX1 I_16640 (I285949,I3035,I285923,I285966,);
not I_16641 (I285915,I285966);
DFFARX1 I_16642 (I205637,I3035,I285923,I285997,);
not I_16643 (I286005,I205640);
nor I_16644 (I286022,I285949,I286005);
not I_16645 (I286039,I205643);
not I_16646 (I286056,I205655);
nand I_16647 (I286073,I286056,I205643);
nor I_16648 (I286090,I286005,I286073);
nor I_16649 (I286107,I285997,I286090);
DFFARX1 I_16650 (I286056,I3035,I285923,I285912,);
nor I_16651 (I286138,I205655,I205646);
nand I_16652 (I286155,I286138,I205634);
nor I_16653 (I286172,I286155,I286039);
nand I_16654 (I285897,I286172,I205640);
DFFARX1 I_16655 (I286155,I3035,I285923,I285909,);
nand I_16656 (I286217,I286039,I205655);
nor I_16657 (I286234,I286039,I205655);
nand I_16658 (I285903,I286022,I286234);
not I_16659 (I286265,I205652);
nor I_16660 (I286282,I286265,I286217);
DFFARX1 I_16661 (I286282,I3035,I285923,I285891,);
nor I_16662 (I286313,I286265,I205658);
and I_16663 (I286330,I286313,I205661);
or I_16664 (I286347,I286330,I205634);
DFFARX1 I_16665 (I286347,I3035,I285923,I286373,);
nor I_16666 (I286381,I286373,I285997);
nor I_16667 (I285900,I285949,I286381);
not I_16668 (I286412,I286373);
nor I_16669 (I286429,I286412,I286107);
DFFARX1 I_16670 (I286429,I3035,I285923,I285906,);
nand I_16671 (I286460,I286412,I286039);
nor I_16672 (I285894,I286265,I286460);
not I_16673 (I286518,I3042);
DFFARX1 I_16674 (I303047,I3035,I286518,I286544,);
DFFARX1 I_16675 (I286544,I3035,I286518,I286561,);
not I_16676 (I286510,I286561);
DFFARX1 I_16677 (I303059,I3035,I286518,I286592,);
not I_16678 (I286600,I303044);
nor I_16679 (I286617,I286544,I286600);
not I_16680 (I286634,I303062);
not I_16681 (I286651,I303053);
nand I_16682 (I286668,I286651,I303062);
nor I_16683 (I286685,I286600,I286668);
nor I_16684 (I286702,I286592,I286685);
DFFARX1 I_16685 (I286651,I3035,I286518,I286507,);
nor I_16686 (I286733,I303053,I303065);
nand I_16687 (I286750,I286733,I303068);
nor I_16688 (I286767,I286750,I286634);
nand I_16689 (I286492,I286767,I303044);
DFFARX1 I_16690 (I286750,I3035,I286518,I286504,);
nand I_16691 (I286812,I286634,I303053);
nor I_16692 (I286829,I286634,I303053);
nand I_16693 (I286498,I286617,I286829);
not I_16694 (I286860,I303044);
nor I_16695 (I286877,I286860,I286812);
DFFARX1 I_16696 (I286877,I3035,I286518,I286486,);
nor I_16697 (I286908,I286860,I303056);
and I_16698 (I286925,I286908,I303050);
or I_16699 (I286942,I286925,I303047);
DFFARX1 I_16700 (I286942,I3035,I286518,I286968,);
nor I_16701 (I286976,I286968,I286592);
nor I_16702 (I286495,I286544,I286976);
not I_16703 (I287007,I286968);
nor I_16704 (I287024,I287007,I286702);
DFFARX1 I_16705 (I287024,I3035,I286518,I286501,);
nand I_16706 (I287055,I287007,I286634);
nor I_16707 (I286489,I286860,I287055);
not I_16708 (I287113,I3042);
DFFARX1 I_16709 (I43123,I3035,I287113,I287139,);
DFFARX1 I_16710 (I287139,I3035,I287113,I287156,);
not I_16711 (I287105,I287156);
DFFARX1 I_16712 (I43135,I3035,I287113,I287187,);
not I_16713 (I287195,I43126);
nor I_16714 (I287212,I287139,I287195);
not I_16715 (I287229,I43117);
not I_16716 (I287246,I43114);
nand I_16717 (I287263,I287246,I43117);
nor I_16718 (I287280,I287195,I287263);
nor I_16719 (I287297,I287187,I287280);
DFFARX1 I_16720 (I287246,I3035,I287113,I287102,);
nor I_16721 (I287328,I43114,I43114);
nand I_16722 (I287345,I287328,I43132);
nor I_16723 (I287362,I287345,I287229);
nand I_16724 (I287087,I287362,I43126);
DFFARX1 I_16725 (I287345,I3035,I287113,I287099,);
nand I_16726 (I287407,I287229,I43114);
nor I_16727 (I287424,I287229,I43114);
nand I_16728 (I287093,I287212,I287424);
not I_16729 (I287455,I43138);
nor I_16730 (I287472,I287455,I287407);
DFFARX1 I_16731 (I287472,I3035,I287113,I287081,);
nor I_16732 (I287503,I287455,I43117);
and I_16733 (I287520,I287503,I43120);
or I_16734 (I287537,I287520,I43129);
DFFARX1 I_16735 (I287537,I3035,I287113,I287563,);
nor I_16736 (I287571,I287563,I287187);
nor I_16737 (I287090,I287139,I287571);
not I_16738 (I287602,I287563);
nor I_16739 (I287619,I287602,I287297);
DFFARX1 I_16740 (I287619,I3035,I287113,I287096,);
nand I_16741 (I287650,I287602,I287229);
nor I_16742 (I287084,I287455,I287650);
not I_16743 (I287708,I3042);
DFFARX1 I_16744 (I717453,I3035,I287708,I287734,);
DFFARX1 I_16745 (I287734,I3035,I287708,I287751,);
not I_16746 (I287700,I287751);
DFFARX1 I_16747 (I717459,I3035,I287708,I287782,);
not I_16748 (I287790,I717474);
nor I_16749 (I287807,I287734,I287790);
not I_16750 (I287824,I717465);
not I_16751 (I287841,I717462);
nand I_16752 (I287858,I287841,I717465);
nor I_16753 (I287875,I287790,I287858);
nor I_16754 (I287892,I287782,I287875);
DFFARX1 I_16755 (I287841,I3035,I287708,I287697,);
nor I_16756 (I287923,I717462,I717453);
nand I_16757 (I287940,I287923,I717477);
nor I_16758 (I287957,I287940,I287824);
nand I_16759 (I287682,I287957,I717474);
DFFARX1 I_16760 (I287940,I3035,I287708,I287694,);
nand I_16761 (I288002,I287824,I717462);
nor I_16762 (I288019,I287824,I717462);
nand I_16763 (I287688,I287807,I288019);
not I_16764 (I288050,I717471);
nor I_16765 (I288067,I288050,I288002);
DFFARX1 I_16766 (I288067,I3035,I287708,I287676,);
nor I_16767 (I288098,I288050,I717456);
and I_16768 (I288115,I288098,I717468);
or I_16769 (I288132,I288115,I717480);
DFFARX1 I_16770 (I288132,I3035,I287708,I288158,);
nor I_16771 (I288166,I288158,I287782);
nor I_16772 (I287685,I287734,I288166);
not I_16773 (I288197,I288158);
nor I_16774 (I288214,I288197,I287892);
DFFARX1 I_16775 (I288214,I3035,I287708,I287691,);
nand I_16776 (I288245,I288197,I287824);
nor I_16777 (I287679,I288050,I288245);
not I_16778 (I288303,I3042);
DFFARX1 I_16779 (I1956,I3035,I288303,I288329,);
DFFARX1 I_16780 (I288329,I3035,I288303,I288346,);
not I_16781 (I288295,I288346);
DFFARX1 I_16782 (I2324,I3035,I288303,I288377,);
not I_16783 (I288385,I1604);
nor I_16784 (I288402,I288329,I288385);
not I_16785 (I288419,I1852);
not I_16786 (I288436,I2108);
nand I_16787 (I288453,I288436,I1852);
nor I_16788 (I288470,I288385,I288453);
nor I_16789 (I288487,I288377,I288470);
DFFARX1 I_16790 (I288436,I3035,I288303,I288292,);
nor I_16791 (I288518,I2108,I2228);
nand I_16792 (I288535,I288518,I2500);
nor I_16793 (I288552,I288535,I288419);
nand I_16794 (I288277,I288552,I1604);
DFFARX1 I_16795 (I288535,I3035,I288303,I288289,);
nand I_16796 (I288597,I288419,I2108);
nor I_16797 (I288614,I288419,I2108);
nand I_16798 (I288283,I288402,I288614);
not I_16799 (I288645,I2828);
nor I_16800 (I288662,I288645,I288597);
DFFARX1 I_16801 (I288662,I3035,I288303,I288271,);
nor I_16802 (I288693,I288645,I1988);
and I_16803 (I288710,I288693,I1364);
or I_16804 (I288727,I288710,I1860);
DFFARX1 I_16805 (I288727,I3035,I288303,I288753,);
nor I_16806 (I288761,I288753,I288377);
nor I_16807 (I288280,I288329,I288761);
not I_16808 (I288792,I288753);
nor I_16809 (I288809,I288792,I288487);
DFFARX1 I_16810 (I288809,I3035,I288303,I288286,);
nand I_16811 (I288840,I288792,I288419);
nor I_16812 (I288274,I288645,I288840);
not I_16813 (I288898,I3042);
DFFARX1 I_16814 (I522597,I3035,I288898,I288924,);
DFFARX1 I_16815 (I288924,I3035,I288898,I288941,);
not I_16816 (I288890,I288941);
DFFARX1 I_16817 (I522585,I3035,I288898,I288972,);
not I_16818 (I288980,I522582);
nor I_16819 (I288997,I288924,I288980);
not I_16820 (I289014,I522594);
not I_16821 (I289031,I522591);
nand I_16822 (I289048,I289031,I522594);
nor I_16823 (I289065,I288980,I289048);
nor I_16824 (I289082,I288972,I289065);
DFFARX1 I_16825 (I289031,I3035,I288898,I288887,);
nor I_16826 (I289113,I522591,I522600);
nand I_16827 (I289130,I289113,I522603);
nor I_16828 (I289147,I289130,I289014);
nand I_16829 (I288872,I289147,I522582);
DFFARX1 I_16830 (I289130,I3035,I288898,I288884,);
nand I_16831 (I289192,I289014,I522591);
nor I_16832 (I289209,I289014,I522591);
nand I_16833 (I288878,I288997,I289209);
not I_16834 (I289240,I522606);
nor I_16835 (I289257,I289240,I289192);
DFFARX1 I_16836 (I289257,I3035,I288898,I288866,);
nor I_16837 (I289288,I289240,I522609);
and I_16838 (I289305,I289288,I522588);
or I_16839 (I289322,I289305,I522582);
DFFARX1 I_16840 (I289322,I3035,I288898,I289348,);
nor I_16841 (I289356,I289348,I288972);
nor I_16842 (I288875,I288924,I289356);
not I_16843 (I289387,I289348);
nor I_16844 (I289404,I289387,I289082);
DFFARX1 I_16845 (I289404,I3035,I288898,I288881,);
nand I_16846 (I289435,I289387,I289014);
nor I_16847 (I288869,I289240,I289435);
not I_16848 (I289493,I3042);
DFFARX1 I_16849 (I264709,I3035,I289493,I289519,);
DFFARX1 I_16850 (I289519,I3035,I289493,I289536,);
not I_16851 (I289485,I289536);
DFFARX1 I_16852 (I264733,I3035,I289493,I289567,);
not I_16853 (I289575,I264712);
nor I_16854 (I289592,I289519,I289575);
not I_16855 (I289609,I264718);
not I_16856 (I289626,I264724);
nand I_16857 (I289643,I289626,I264718);
nor I_16858 (I289660,I289575,I289643);
nor I_16859 (I289677,I289567,I289660);
DFFARX1 I_16860 (I289626,I3035,I289493,I289482,);
nor I_16861 (I289708,I264724,I264736);
nand I_16862 (I289725,I289708,I264730);
nor I_16863 (I289742,I289725,I289609);
nand I_16864 (I289467,I289742,I264712);
DFFARX1 I_16865 (I289725,I3035,I289493,I289479,);
nand I_16866 (I289787,I289609,I264724);
nor I_16867 (I289804,I289609,I264724);
nand I_16868 (I289473,I289592,I289804);
not I_16869 (I289835,I264715);
nor I_16870 (I289852,I289835,I289787);
DFFARX1 I_16871 (I289852,I3035,I289493,I289461,);
nor I_16872 (I289883,I289835,I264709);
and I_16873 (I289900,I289883,I264727);
or I_16874 (I289917,I289900,I264721);
DFFARX1 I_16875 (I289917,I3035,I289493,I289943,);
nor I_16876 (I289951,I289943,I289567);
nor I_16877 (I289470,I289519,I289951);
not I_16878 (I289982,I289943);
nor I_16879 (I289999,I289982,I289677);
DFFARX1 I_16880 (I289999,I3035,I289493,I289476,);
nand I_16881 (I290030,I289982,I289609);
nor I_16882 (I289464,I289835,I290030);
not I_16883 (I290088,I3042);
DFFARX1 I_16884 (I382239,I3035,I290088,I290114,);
DFFARX1 I_16885 (I290114,I3035,I290088,I290131,);
not I_16886 (I290080,I290131);
DFFARX1 I_16887 (I382233,I3035,I290088,I290162,);
not I_16888 (I290170,I382230);
nor I_16889 (I290187,I290114,I290170);
not I_16890 (I290204,I382242);
not I_16891 (I290221,I382245);
nand I_16892 (I290238,I290221,I382242);
nor I_16893 (I290255,I290170,I290238);
nor I_16894 (I290272,I290162,I290255);
DFFARX1 I_16895 (I290221,I3035,I290088,I290077,);
nor I_16896 (I290303,I382245,I382254);
nand I_16897 (I290320,I290303,I382248);
nor I_16898 (I290337,I290320,I290204);
nand I_16899 (I290062,I290337,I382230);
DFFARX1 I_16900 (I290320,I3035,I290088,I290074,);
nand I_16901 (I290382,I290204,I382245);
nor I_16902 (I290399,I290204,I382245);
nand I_16903 (I290068,I290187,I290399);
not I_16904 (I290430,I382236);
nor I_16905 (I290447,I290430,I290382);
DFFARX1 I_16906 (I290447,I3035,I290088,I290056,);
nor I_16907 (I290478,I290430,I382251);
and I_16908 (I290495,I290478,I382230);
or I_16909 (I290512,I290495,I382233);
DFFARX1 I_16910 (I290512,I3035,I290088,I290538,);
nor I_16911 (I290546,I290538,I290162);
nor I_16912 (I290065,I290114,I290546);
not I_16913 (I290577,I290538);
nor I_16914 (I290594,I290577,I290272);
DFFARX1 I_16915 (I290594,I3035,I290088,I290071,);
nand I_16916 (I290625,I290577,I290204);
nor I_16917 (I290059,I290430,I290625);
not I_16918 (I290683,I3042);
DFFARX1 I_16919 (I2756,I3035,I290683,I290709,);
DFFARX1 I_16920 (I290709,I3035,I290683,I290726,);
not I_16921 (I290675,I290726);
DFFARX1 I_16922 (I2156,I3035,I290683,I290757,);
not I_16923 (I290765,I1828);
nor I_16924 (I290782,I290709,I290765);
not I_16925 (I290799,I2276);
not I_16926 (I290816,I1772);
nand I_16927 (I290833,I290816,I2276);
nor I_16928 (I290850,I290765,I290833);
nor I_16929 (I290867,I290757,I290850);
DFFARX1 I_16930 (I290816,I3035,I290683,I290672,);
nor I_16931 (I290898,I1772,I2316);
nand I_16932 (I290915,I290898,I1628);
nor I_16933 (I290932,I290915,I290799);
nand I_16934 (I290657,I290932,I1828);
DFFARX1 I_16935 (I290915,I3035,I290683,I290669,);
nand I_16936 (I290977,I290799,I1772);
nor I_16937 (I290994,I290799,I1772);
nand I_16938 (I290663,I290782,I290994);
not I_16939 (I291025,I2572);
nor I_16940 (I291042,I291025,I290977);
DFFARX1 I_16941 (I291042,I3035,I290683,I290651,);
nor I_16942 (I291073,I291025,I2436);
and I_16943 (I291090,I291073,I2788);
or I_16944 (I291107,I291090,I2748);
DFFARX1 I_16945 (I291107,I3035,I290683,I291133,);
nor I_16946 (I291141,I291133,I290757);
nor I_16947 (I290660,I290709,I291141);
not I_16948 (I291172,I291133);
nor I_16949 (I291189,I291172,I290867);
DFFARX1 I_16950 (I291189,I3035,I290683,I290666,);
nand I_16951 (I291220,I291172,I290799);
nor I_16952 (I290654,I291025,I291220);
not I_16953 (I291278,I3042);
DFFARX1 I_16954 (I612190,I3035,I291278,I291304,);
DFFARX1 I_16955 (I291304,I3035,I291278,I291321,);
not I_16956 (I291270,I291321);
DFFARX1 I_16957 (I612172,I3035,I291278,I291352,);
not I_16958 (I291360,I612178);
nor I_16959 (I291377,I291304,I291360);
not I_16960 (I291394,I612193);
not I_16961 (I291411,I612184);
nand I_16962 (I291428,I291411,I612193);
nor I_16963 (I291445,I291360,I291428);
nor I_16964 (I291462,I291352,I291445);
DFFARX1 I_16965 (I291411,I3035,I291278,I291267,);
nor I_16966 (I291493,I612184,I612196);
nand I_16967 (I291510,I291493,I612175);
nor I_16968 (I291527,I291510,I291394);
nand I_16969 (I291252,I291527,I612178);
DFFARX1 I_16970 (I291510,I3035,I291278,I291264,);
nand I_16971 (I291572,I291394,I612184);
nor I_16972 (I291589,I291394,I612184);
nand I_16973 (I291258,I291377,I291589);
not I_16974 (I291620,I612181);
nor I_16975 (I291637,I291620,I291572);
DFFARX1 I_16976 (I291637,I3035,I291278,I291246,);
nor I_16977 (I291668,I291620,I612187);
and I_16978 (I291685,I291668,I612172);
or I_16979 (I291702,I291685,I612175);
DFFARX1 I_16980 (I291702,I3035,I291278,I291728,);
nor I_16981 (I291736,I291728,I291352);
nor I_16982 (I291255,I291304,I291736);
not I_16983 (I291767,I291728);
nor I_16984 (I291784,I291767,I291462);
DFFARX1 I_16985 (I291784,I3035,I291278,I291261,);
nand I_16986 (I291815,I291767,I291394);
nor I_16987 (I291249,I291620,I291815);
not I_16988 (I291873,I3042);
DFFARX1 I_16989 (I746608,I3035,I291873,I291899,);
DFFARX1 I_16990 (I291899,I3035,I291873,I291916,);
not I_16991 (I291865,I291916);
DFFARX1 I_16992 (I746614,I3035,I291873,I291947,);
not I_16993 (I291955,I746629);
nor I_16994 (I291972,I291899,I291955);
not I_16995 (I291989,I746620);
not I_16996 (I292006,I746617);
nand I_16997 (I292023,I292006,I746620);
nor I_16998 (I292040,I291955,I292023);
nor I_16999 (I292057,I291947,I292040);
DFFARX1 I_17000 (I292006,I3035,I291873,I291862,);
nor I_17001 (I292088,I746617,I746608);
nand I_17002 (I292105,I292088,I746632);
nor I_17003 (I292122,I292105,I291989);
nand I_17004 (I291847,I292122,I746629);
DFFARX1 I_17005 (I292105,I3035,I291873,I291859,);
nand I_17006 (I292167,I291989,I746617);
nor I_17007 (I292184,I291989,I746617);
nand I_17008 (I291853,I291972,I292184);
not I_17009 (I292215,I746626);
nor I_17010 (I292232,I292215,I292167);
DFFARX1 I_17011 (I292232,I3035,I291873,I291841,);
nor I_17012 (I292263,I292215,I746611);
and I_17013 (I292280,I292263,I746623);
or I_17014 (I292297,I292280,I746635);
DFFARX1 I_17015 (I292297,I3035,I291873,I292323,);
nor I_17016 (I292331,I292323,I291947);
nor I_17017 (I291850,I291899,I292331);
not I_17018 (I292362,I292323);
nor I_17019 (I292379,I292362,I292057);
DFFARX1 I_17020 (I292379,I3035,I291873,I291856,);
nand I_17021 (I292410,I292362,I291989);
nor I_17022 (I291844,I292215,I292410);
not I_17023 (I292468,I3042);
DFFARX1 I_17024 (I432984,I3035,I292468,I292494,);
DFFARX1 I_17025 (I292494,I3035,I292468,I292511,);
not I_17026 (I292460,I292511);
DFFARX1 I_17027 (I432981,I3035,I292468,I292542,);
not I_17028 (I292550,I432981);
nor I_17029 (I292567,I292494,I292550);
not I_17030 (I292584,I432978);
not I_17031 (I292601,I432993);
nand I_17032 (I292618,I292601,I432978);
nor I_17033 (I292635,I292550,I292618);
nor I_17034 (I292652,I292542,I292635);
DFFARX1 I_17035 (I292601,I3035,I292468,I292457,);
nor I_17036 (I292683,I432993,I432987);
nand I_17037 (I292700,I292683,I432975);
nor I_17038 (I292717,I292700,I292584);
nand I_17039 (I292442,I292717,I432981);
DFFARX1 I_17040 (I292700,I3035,I292468,I292454,);
nand I_17041 (I292762,I292584,I432993);
nor I_17042 (I292779,I292584,I432993);
nand I_17043 (I292448,I292567,I292779);
not I_17044 (I292810,I432996);
nor I_17045 (I292827,I292810,I292762);
DFFARX1 I_17046 (I292827,I3035,I292468,I292436,);
nor I_17047 (I292858,I292810,I432975);
and I_17048 (I292875,I292858,I432990);
or I_17049 (I292892,I292875,I432978);
DFFARX1 I_17050 (I292892,I3035,I292468,I292918,);
nor I_17051 (I292926,I292918,I292542);
nor I_17052 (I292445,I292494,I292926);
not I_17053 (I292957,I292918);
nor I_17054 (I292974,I292957,I292652);
DFFARX1 I_17055 (I292974,I3035,I292468,I292451,);
nand I_17056 (I293005,I292957,I292584);
nor I_17057 (I292439,I292810,I293005);
not I_17058 (I293063,I3042);
DFFARX1 I_17059 (I735303,I3035,I293063,I293089,);
DFFARX1 I_17060 (I293089,I3035,I293063,I293106,);
not I_17061 (I293055,I293106);
DFFARX1 I_17062 (I735309,I3035,I293063,I293137,);
not I_17063 (I293145,I735324);
nor I_17064 (I293162,I293089,I293145);
not I_17065 (I293179,I735315);
not I_17066 (I293196,I735312);
nand I_17067 (I293213,I293196,I735315);
nor I_17068 (I293230,I293145,I293213);
nor I_17069 (I293247,I293137,I293230);
DFFARX1 I_17070 (I293196,I3035,I293063,I293052,);
nor I_17071 (I293278,I735312,I735303);
nand I_17072 (I293295,I293278,I735327);
nor I_17073 (I293312,I293295,I293179);
nand I_17074 (I293037,I293312,I735324);
DFFARX1 I_17075 (I293295,I3035,I293063,I293049,);
nand I_17076 (I293357,I293179,I735312);
nor I_17077 (I293374,I293179,I735312);
nand I_17078 (I293043,I293162,I293374);
not I_17079 (I293405,I735321);
nor I_17080 (I293422,I293405,I293357);
DFFARX1 I_17081 (I293422,I3035,I293063,I293031,);
nor I_17082 (I293453,I293405,I735306);
and I_17083 (I293470,I293453,I735318);
or I_17084 (I293487,I293470,I735330);
DFFARX1 I_17085 (I293487,I3035,I293063,I293513,);
nor I_17086 (I293521,I293513,I293137);
nor I_17087 (I293040,I293089,I293521);
not I_17088 (I293552,I293513);
nor I_17089 (I293569,I293552,I293247);
DFFARX1 I_17090 (I293569,I3035,I293063,I293046,);
nand I_17091 (I293600,I293552,I293179);
nor I_17092 (I293034,I293405,I293600);
not I_17093 (I293658,I3042);
DFFARX1 I_17094 (I507093,I3035,I293658,I293684,);
DFFARX1 I_17095 (I293684,I3035,I293658,I293701,);
not I_17096 (I293650,I293701);
DFFARX1 I_17097 (I507081,I3035,I293658,I293732,);
not I_17098 (I293740,I507078);
nor I_17099 (I293757,I293684,I293740);
not I_17100 (I293774,I507090);
not I_17101 (I293791,I507087);
nand I_17102 (I293808,I293791,I507090);
nor I_17103 (I293825,I293740,I293808);
nor I_17104 (I293842,I293732,I293825);
DFFARX1 I_17105 (I293791,I3035,I293658,I293647,);
nor I_17106 (I293873,I507087,I507096);
nand I_17107 (I293890,I293873,I507099);
nor I_17108 (I293907,I293890,I293774);
nand I_17109 (I293632,I293907,I507078);
DFFARX1 I_17110 (I293890,I3035,I293658,I293644,);
nand I_17111 (I293952,I293774,I507087);
nor I_17112 (I293969,I293774,I507087);
nand I_17113 (I293638,I293757,I293969);
not I_17114 (I294000,I507102);
nor I_17115 (I294017,I294000,I293952);
DFFARX1 I_17116 (I294017,I3035,I293658,I293626,);
nor I_17117 (I294048,I294000,I507105);
and I_17118 (I294065,I294048,I507084);
or I_17119 (I294082,I294065,I507078);
DFFARX1 I_17120 (I294082,I3035,I293658,I294108,);
nor I_17121 (I294116,I294108,I293732);
nor I_17122 (I293635,I293684,I294116);
not I_17123 (I294147,I294108);
nor I_17124 (I294164,I294147,I293842);
DFFARX1 I_17125 (I294164,I3035,I293658,I293641,);
nand I_17126 (I294195,I294147,I293774);
nor I_17127 (I293629,I294000,I294195);
not I_17128 (I294253,I3042);
DFFARX1 I_17129 (I697223,I3035,I294253,I294279,);
DFFARX1 I_17130 (I294279,I3035,I294253,I294296,);
not I_17131 (I294245,I294296);
DFFARX1 I_17132 (I697229,I3035,I294253,I294327,);
not I_17133 (I294335,I697244);
nor I_17134 (I294352,I294279,I294335);
not I_17135 (I294369,I697235);
not I_17136 (I294386,I697232);
nand I_17137 (I294403,I294386,I697235);
nor I_17138 (I294420,I294335,I294403);
nor I_17139 (I294437,I294327,I294420);
DFFARX1 I_17140 (I294386,I3035,I294253,I294242,);
nor I_17141 (I294468,I697232,I697223);
nand I_17142 (I294485,I294468,I697247);
nor I_17143 (I294502,I294485,I294369);
nand I_17144 (I294227,I294502,I697244);
DFFARX1 I_17145 (I294485,I3035,I294253,I294239,);
nand I_17146 (I294547,I294369,I697232);
nor I_17147 (I294564,I294369,I697232);
nand I_17148 (I294233,I294352,I294564);
not I_17149 (I294595,I697241);
nor I_17150 (I294612,I294595,I294547);
DFFARX1 I_17151 (I294612,I3035,I294253,I294221,);
nor I_17152 (I294643,I294595,I697226);
and I_17153 (I294660,I294643,I697238);
or I_17154 (I294677,I294660,I697250);
DFFARX1 I_17155 (I294677,I3035,I294253,I294703,);
nor I_17156 (I294711,I294703,I294327);
nor I_17157 (I294230,I294279,I294711);
not I_17158 (I294742,I294703);
nor I_17159 (I294759,I294742,I294437);
DFFARX1 I_17160 (I294759,I3035,I294253,I294236,);
nand I_17161 (I294790,I294742,I294369);
nor I_17162 (I294224,I294595,I294790);
not I_17163 (I294848,I3042);
DFFARX1 I_17164 (I539393,I3035,I294848,I294874,);
DFFARX1 I_17165 (I294874,I3035,I294848,I294891,);
not I_17166 (I294840,I294891);
DFFARX1 I_17167 (I539381,I3035,I294848,I294922,);
not I_17168 (I294930,I539378);
nor I_17169 (I294947,I294874,I294930);
not I_17170 (I294964,I539390);
not I_17171 (I294981,I539387);
nand I_17172 (I294998,I294981,I539390);
nor I_17173 (I295015,I294930,I294998);
nor I_17174 (I295032,I294922,I295015);
DFFARX1 I_17175 (I294981,I3035,I294848,I294837,);
nor I_17176 (I295063,I539387,I539396);
nand I_17177 (I295080,I295063,I539399);
nor I_17178 (I295097,I295080,I294964);
nand I_17179 (I294822,I295097,I539378);
DFFARX1 I_17180 (I295080,I3035,I294848,I294834,);
nand I_17181 (I295142,I294964,I539387);
nor I_17182 (I295159,I294964,I539387);
nand I_17183 (I294828,I294947,I295159);
not I_17184 (I295190,I539402);
nor I_17185 (I295207,I295190,I295142);
DFFARX1 I_17186 (I295207,I3035,I294848,I294816,);
nor I_17187 (I295238,I295190,I539405);
and I_17188 (I295255,I295238,I539384);
or I_17189 (I295272,I295255,I539378);
DFFARX1 I_17190 (I295272,I3035,I294848,I295298,);
nor I_17191 (I295306,I295298,I294922);
nor I_17192 (I294825,I294874,I295306);
not I_17193 (I295337,I295298);
nor I_17194 (I295354,I295337,I295032);
DFFARX1 I_17195 (I295354,I3035,I294848,I294831,);
nand I_17196 (I295385,I295337,I294964);
nor I_17197 (I294819,I295190,I295385);
not I_17198 (I295443,I3042);
DFFARX1 I_17199 (I587336,I3035,I295443,I295469,);
DFFARX1 I_17200 (I295469,I3035,I295443,I295486,);
not I_17201 (I295435,I295486);
DFFARX1 I_17202 (I587318,I3035,I295443,I295517,);
not I_17203 (I295525,I587324);
nor I_17204 (I295542,I295469,I295525);
not I_17205 (I295559,I587339);
not I_17206 (I295576,I587330);
nand I_17207 (I295593,I295576,I587339);
nor I_17208 (I295610,I295525,I295593);
nor I_17209 (I295627,I295517,I295610);
DFFARX1 I_17210 (I295576,I3035,I295443,I295432,);
nor I_17211 (I295658,I587330,I587342);
nand I_17212 (I295675,I295658,I587321);
nor I_17213 (I295692,I295675,I295559);
nand I_17214 (I295417,I295692,I587324);
DFFARX1 I_17215 (I295675,I3035,I295443,I295429,);
nand I_17216 (I295737,I295559,I587330);
nor I_17217 (I295754,I295559,I587330);
nand I_17218 (I295423,I295542,I295754);
not I_17219 (I295785,I587327);
nor I_17220 (I295802,I295785,I295737);
DFFARX1 I_17221 (I295802,I3035,I295443,I295411,);
nor I_17222 (I295833,I295785,I587333);
and I_17223 (I295850,I295833,I587318);
or I_17224 (I295867,I295850,I587321);
DFFARX1 I_17225 (I295867,I3035,I295443,I295893,);
nor I_17226 (I295901,I295893,I295517);
nor I_17227 (I295420,I295469,I295901);
not I_17228 (I295932,I295893);
nor I_17229 (I295949,I295932,I295627);
DFFARX1 I_17230 (I295949,I3035,I295443,I295426,);
nand I_17231 (I295980,I295932,I295559);
nor I_17232 (I295414,I295785,I295980);
not I_17233 (I296038,I3042);
DFFARX1 I_17234 (I513553,I3035,I296038,I296064,);
DFFARX1 I_17235 (I296064,I3035,I296038,I296081,);
not I_17236 (I296030,I296081);
DFFARX1 I_17237 (I513541,I3035,I296038,I296112,);
not I_17238 (I296120,I513538);
nor I_17239 (I296137,I296064,I296120);
not I_17240 (I296154,I513550);
not I_17241 (I296171,I513547);
nand I_17242 (I296188,I296171,I513550);
nor I_17243 (I296205,I296120,I296188);
nor I_17244 (I296222,I296112,I296205);
DFFARX1 I_17245 (I296171,I3035,I296038,I296027,);
nor I_17246 (I296253,I513547,I513556);
nand I_17247 (I296270,I296253,I513559);
nor I_17248 (I296287,I296270,I296154);
nand I_17249 (I296012,I296287,I513538);
DFFARX1 I_17250 (I296270,I3035,I296038,I296024,);
nand I_17251 (I296332,I296154,I513547);
nor I_17252 (I296349,I296154,I513547);
nand I_17253 (I296018,I296137,I296349);
not I_17254 (I296380,I513562);
nor I_17255 (I296397,I296380,I296332);
DFFARX1 I_17256 (I296397,I3035,I296038,I296006,);
nor I_17257 (I296428,I296380,I513565);
and I_17258 (I296445,I296428,I513544);
or I_17259 (I296462,I296445,I513538);
DFFARX1 I_17260 (I296462,I3035,I296038,I296488,);
nor I_17261 (I296496,I296488,I296112);
nor I_17262 (I296015,I296064,I296496);
not I_17263 (I296527,I296488);
nor I_17264 (I296544,I296527,I296222);
DFFARX1 I_17265 (I296544,I3035,I296038,I296021,);
nand I_17266 (I296575,I296527,I296154);
nor I_17267 (I296009,I296380,I296575);
not I_17268 (I296633,I3042);
DFFARX1 I_17269 (I404781,I3035,I296633,I296659,);
DFFARX1 I_17270 (I296659,I3035,I296633,I296676,);
not I_17271 (I296625,I296676);
DFFARX1 I_17272 (I404775,I3035,I296633,I296707,);
not I_17273 (I296715,I404772);
nor I_17274 (I296732,I296659,I296715);
not I_17275 (I296749,I404784);
not I_17276 (I296766,I404787);
nand I_17277 (I296783,I296766,I404784);
nor I_17278 (I296800,I296715,I296783);
nor I_17279 (I296817,I296707,I296800);
DFFARX1 I_17280 (I296766,I3035,I296633,I296622,);
nor I_17281 (I296848,I404787,I404796);
nand I_17282 (I296865,I296848,I404790);
nor I_17283 (I296882,I296865,I296749);
nand I_17284 (I296607,I296882,I404772);
DFFARX1 I_17285 (I296865,I3035,I296633,I296619,);
nand I_17286 (I296927,I296749,I404787);
nor I_17287 (I296944,I296749,I404787);
nand I_17288 (I296613,I296732,I296944);
not I_17289 (I296975,I404778);
nor I_17290 (I296992,I296975,I296927);
DFFARX1 I_17291 (I296992,I3035,I296633,I296601,);
nor I_17292 (I297023,I296975,I404793);
and I_17293 (I297040,I297023,I404772);
or I_17294 (I297057,I297040,I404775);
DFFARX1 I_17295 (I297057,I3035,I296633,I297083,);
nor I_17296 (I297091,I297083,I296707);
nor I_17297 (I296610,I296659,I297091);
not I_17298 (I297122,I297083);
nor I_17299 (I297139,I297122,I296817);
DFFARX1 I_17300 (I297139,I3035,I296633,I296616,);
nand I_17301 (I297170,I297122,I296749);
nor I_17302 (I296604,I296975,I297170);
not I_17303 (I297228,I3042);
DFFARX1 I_17304 (I422971,I3035,I297228,I297254,);
DFFARX1 I_17305 (I297254,I3035,I297228,I297271,);
not I_17306 (I297220,I297271);
DFFARX1 I_17307 (I422968,I3035,I297228,I297302,);
not I_17308 (I297310,I422968);
nor I_17309 (I297327,I297254,I297310);
not I_17310 (I297344,I422965);
not I_17311 (I297361,I422980);
nand I_17312 (I297378,I297361,I422965);
nor I_17313 (I297395,I297310,I297378);
nor I_17314 (I297412,I297302,I297395);
DFFARX1 I_17315 (I297361,I3035,I297228,I297217,);
nor I_17316 (I297443,I422980,I422974);
nand I_17317 (I297460,I297443,I422962);
nor I_17318 (I297477,I297460,I297344);
nand I_17319 (I297202,I297477,I422968);
DFFARX1 I_17320 (I297460,I3035,I297228,I297214,);
nand I_17321 (I297522,I297344,I422980);
nor I_17322 (I297539,I297344,I422980);
nand I_17323 (I297208,I297327,I297539);
not I_17324 (I297570,I422983);
nor I_17325 (I297587,I297570,I297522);
DFFARX1 I_17326 (I297587,I3035,I297228,I297196,);
nor I_17327 (I297618,I297570,I422962);
and I_17328 (I297635,I297618,I422977);
or I_17329 (I297652,I297635,I422965);
DFFARX1 I_17330 (I297652,I3035,I297228,I297678,);
nor I_17331 (I297686,I297678,I297302);
nor I_17332 (I297205,I297254,I297686);
not I_17333 (I297717,I297678);
nor I_17334 (I297734,I297717,I297412);
DFFARX1 I_17335 (I297734,I3035,I297228,I297211,);
nand I_17336 (I297765,I297717,I297344);
nor I_17337 (I297199,I297570,I297765);
not I_17338 (I297823,I3042);
DFFARX1 I_17339 (I626062,I3035,I297823,I297849,);
DFFARX1 I_17340 (I297849,I3035,I297823,I297866,);
not I_17341 (I297815,I297866);
DFFARX1 I_17342 (I626044,I3035,I297823,I297897,);
not I_17343 (I297905,I626050);
nor I_17344 (I297922,I297849,I297905);
not I_17345 (I297939,I626065);
not I_17346 (I297956,I626056);
nand I_17347 (I297973,I297956,I626065);
nor I_17348 (I297990,I297905,I297973);
nor I_17349 (I298007,I297897,I297990);
DFFARX1 I_17350 (I297956,I3035,I297823,I297812,);
nor I_17351 (I298038,I626056,I626068);
nand I_17352 (I298055,I298038,I626047);
nor I_17353 (I298072,I298055,I297939);
nand I_17354 (I297797,I298072,I626050);
DFFARX1 I_17355 (I298055,I3035,I297823,I297809,);
nand I_17356 (I298117,I297939,I626056);
nor I_17357 (I298134,I297939,I626056);
nand I_17358 (I297803,I297922,I298134);
not I_17359 (I298165,I626053);
nor I_17360 (I298182,I298165,I298117);
DFFARX1 I_17361 (I298182,I3035,I297823,I297791,);
nor I_17362 (I298213,I298165,I626059);
and I_17363 (I298230,I298213,I626044);
or I_17364 (I298247,I298230,I626047);
DFFARX1 I_17365 (I298247,I3035,I297823,I298273,);
nor I_17366 (I298281,I298273,I297897);
nor I_17367 (I297800,I297849,I298281);
not I_17368 (I298312,I298273);
nor I_17369 (I298329,I298312,I298007);
DFFARX1 I_17370 (I298329,I3035,I297823,I297806,);
nand I_17371 (I298360,I298312,I297939);
nor I_17372 (I297794,I298165,I298360);
not I_17373 (I298418,I3042);
DFFARX1 I_17374 (I299579,I3035,I298418,I298444,);
DFFARX1 I_17375 (I298444,I3035,I298418,I298461,);
not I_17376 (I298410,I298461);
DFFARX1 I_17377 (I299591,I3035,I298418,I298492,);
not I_17378 (I298500,I299576);
nor I_17379 (I298517,I298444,I298500);
not I_17380 (I298534,I299594);
not I_17381 (I298551,I299585);
nand I_17382 (I298568,I298551,I299594);
nor I_17383 (I298585,I298500,I298568);
nor I_17384 (I298602,I298492,I298585);
DFFARX1 I_17385 (I298551,I3035,I298418,I298407,);
nor I_17386 (I298633,I299585,I299597);
nand I_17387 (I298650,I298633,I299600);
nor I_17388 (I298667,I298650,I298534);
nand I_17389 (I298392,I298667,I299576);
DFFARX1 I_17390 (I298650,I3035,I298418,I298404,);
nand I_17391 (I298712,I298534,I299585);
nor I_17392 (I298729,I298534,I299585);
nand I_17393 (I298398,I298517,I298729);
not I_17394 (I298760,I299576);
nor I_17395 (I298777,I298760,I298712);
DFFARX1 I_17396 (I298777,I3035,I298418,I298386,);
nor I_17397 (I298808,I298760,I299588);
and I_17398 (I298825,I298808,I299582);
or I_17399 (I298842,I298825,I299579);
DFFARX1 I_17400 (I298842,I3035,I298418,I298868,);
nor I_17401 (I298876,I298868,I298492);
nor I_17402 (I298395,I298444,I298876);
not I_17403 (I298907,I298868);
nor I_17404 (I298924,I298907,I298602);
DFFARX1 I_17405 (I298924,I3035,I298418,I298401,);
nand I_17406 (I298955,I298907,I298534);
nor I_17407 (I298389,I298760,I298955);
not I_17408 (I299013,I3042);
DFFARX1 I_17409 (I185096,I3035,I299013,I299039,);
DFFARX1 I_17410 (I299039,I3035,I299013,I299056,);
not I_17411 (I299005,I299056);
DFFARX1 I_17412 (I185084,I3035,I299013,I299087,);
not I_17413 (I299095,I185087);
nor I_17414 (I299112,I299039,I299095);
not I_17415 (I299129,I185090);
not I_17416 (I299146,I185102);
nand I_17417 (I299163,I299146,I185090);
nor I_17418 (I299180,I299095,I299163);
nor I_17419 (I299197,I299087,I299180);
DFFARX1 I_17420 (I299146,I3035,I299013,I299002,);
nor I_17421 (I299228,I185102,I185093);
nand I_17422 (I299245,I299228,I185081);
nor I_17423 (I299262,I299245,I299129);
nand I_17424 (I298987,I299262,I185087);
DFFARX1 I_17425 (I299245,I3035,I299013,I298999,);
nand I_17426 (I299307,I299129,I185102);
nor I_17427 (I299324,I299129,I185102);
nand I_17428 (I298993,I299112,I299324);
not I_17429 (I299355,I185099);
nor I_17430 (I299372,I299355,I299307);
DFFARX1 I_17431 (I299372,I3035,I299013,I298981,);
nor I_17432 (I299403,I299355,I185105);
and I_17433 (I299420,I299403,I185108);
or I_17434 (I299437,I299420,I185081);
DFFARX1 I_17435 (I299437,I3035,I299013,I299463,);
nor I_17436 (I299471,I299463,I299087);
nor I_17437 (I298990,I299039,I299471);
not I_17438 (I299502,I299463);
nor I_17439 (I299519,I299502,I299197);
DFFARX1 I_17440 (I299519,I3035,I299013,I298996,);
nand I_17441 (I299550,I299502,I299129);
nor I_17442 (I298984,I299355,I299550);
not I_17443 (I299608,I3042);
DFFARX1 I_17444 (I385698,I3035,I299608,I299634,);
not I_17445 (I299642,I299634);
DFFARX1 I_17446 (I385710,I3035,I299608,I299668,);
not I_17447 (I299676,I385701);
nand I_17448 (I299693,I299676,I385704);
not I_17449 (I299710,I299693);
nor I_17450 (I299727,I299710,I385707);
nor I_17451 (I299744,I299642,I299727);
DFFARX1 I_17452 (I299744,I3035,I299608,I299594,);
not I_17453 (I299775,I385707);
nand I_17454 (I299792,I299775,I299710);
and I_17455 (I299809,I299775,I385701);
nand I_17456 (I299826,I299809,I385713);
nor I_17457 (I299591,I299826,I299775);
and I_17458 (I299582,I299668,I299826);
not I_17459 (I299871,I299826);
nand I_17460 (I299585,I299668,I299871);
nor I_17461 (I299579,I299634,I299826);
not I_17462 (I299916,I385719);
nor I_17463 (I299933,I299916,I385701);
nand I_17464 (I299950,I299933,I299775);
nor I_17465 (I299588,I299693,I299950);
nor I_17466 (I299981,I299916,I385698);
and I_17467 (I299998,I299981,I385716);
or I_17468 (I300015,I299998,I385722);
DFFARX1 I_17469 (I300015,I3035,I299608,I300041,);
nor I_17470 (I300049,I300041,I299792);
DFFARX1 I_17471 (I300049,I3035,I299608,I299576,);
DFFARX1 I_17472 (I300041,I3035,I299608,I299600,);
not I_17473 (I300094,I300041);
nor I_17474 (I300111,I300094,I299668);
nor I_17475 (I300128,I299933,I300111);
DFFARX1 I_17476 (I300128,I3035,I299608,I299597,);
not I_17477 (I300186,I3042);
DFFARX1 I_17478 (I634714,I3035,I300186,I300212,);
not I_17479 (I300220,I300212);
DFFARX1 I_17480 (I634720,I3035,I300186,I300246,);
not I_17481 (I300254,I634714);
nand I_17482 (I300271,I300254,I634717);
not I_17483 (I300288,I300271);
nor I_17484 (I300305,I300288,I634735);
nor I_17485 (I300322,I300220,I300305);
DFFARX1 I_17486 (I300322,I3035,I300186,I300172,);
not I_17487 (I300353,I634735);
nand I_17488 (I300370,I300353,I300288);
and I_17489 (I300387,I300353,I634738);
nand I_17490 (I300404,I300387,I634717);
nor I_17491 (I300169,I300404,I300353);
and I_17492 (I300160,I300246,I300404);
not I_17493 (I300449,I300404);
nand I_17494 (I300163,I300246,I300449);
nor I_17495 (I300157,I300212,I300404);
not I_17496 (I300494,I634723);
nor I_17497 (I300511,I300494,I634738);
nand I_17498 (I300528,I300511,I300353);
nor I_17499 (I300166,I300271,I300528);
nor I_17500 (I300559,I300494,I634729);
and I_17501 (I300576,I300559,I634726);
or I_17502 (I300593,I300576,I634732);
DFFARX1 I_17503 (I300593,I3035,I300186,I300619,);
nor I_17504 (I300627,I300619,I300370);
DFFARX1 I_17505 (I300627,I3035,I300186,I300154,);
DFFARX1 I_17506 (I300619,I3035,I300186,I300178,);
not I_17507 (I300672,I300619);
nor I_17508 (I300689,I300672,I300246);
nor I_17509 (I300706,I300511,I300689);
DFFARX1 I_17510 (I300706,I3035,I300186,I300175,);
not I_17511 (I300764,I3042);
DFFARX1 I_17512 (I244049,I3035,I300764,I300790,);
not I_17513 (I300798,I300790);
DFFARX1 I_17514 (I244061,I3035,I300764,I300824,);
not I_17515 (I300832,I244037);
nand I_17516 (I300849,I300832,I244064);
not I_17517 (I300866,I300849);
nor I_17518 (I300883,I300866,I244052);
nor I_17519 (I300900,I300798,I300883);
DFFARX1 I_17520 (I300900,I3035,I300764,I300750,);
not I_17521 (I300931,I244052);
nand I_17522 (I300948,I300931,I300866);
and I_17523 (I300965,I300931,I244037);
nand I_17524 (I300982,I300965,I244040);
nor I_17525 (I300747,I300982,I300931);
and I_17526 (I300738,I300824,I300982);
not I_17527 (I301027,I300982);
nand I_17528 (I300741,I300824,I301027);
nor I_17529 (I300735,I300790,I300982);
not I_17530 (I301072,I244046);
nor I_17531 (I301089,I301072,I244037);
nand I_17532 (I301106,I301089,I300931);
nor I_17533 (I300744,I300849,I301106);
nor I_17534 (I301137,I301072,I244055);
and I_17535 (I301154,I301137,I244043);
or I_17536 (I301171,I301154,I244058);
DFFARX1 I_17537 (I301171,I3035,I300764,I301197,);
nor I_17538 (I301205,I301197,I300948);
DFFARX1 I_17539 (I301205,I3035,I300764,I300732,);
DFFARX1 I_17540 (I301197,I3035,I300764,I300756,);
not I_17541 (I301250,I301197);
nor I_17542 (I301267,I301250,I300824);
nor I_17543 (I301284,I301089,I301267);
DFFARX1 I_17544 (I301284,I3035,I300764,I300753,);
not I_17545 (I301342,I3042);
DFFARX1 I_17546 (I468817,I3035,I301342,I301368,);
not I_17547 (I301376,I301368);
DFFARX1 I_17548 (I468817,I3035,I301342,I301402,);
not I_17549 (I301410,I468814);
nand I_17550 (I301427,I301410,I468829);
not I_17551 (I301444,I301427);
nor I_17552 (I301461,I301444,I468823);
nor I_17553 (I301478,I301376,I301461);
DFFARX1 I_17554 (I301478,I3035,I301342,I301328,);
not I_17555 (I301509,I468823);
nand I_17556 (I301526,I301509,I301444);
and I_17557 (I301543,I301509,I468820);
nand I_17558 (I301560,I301543,I468811);
nor I_17559 (I301325,I301560,I301509);
and I_17560 (I301316,I301402,I301560);
not I_17561 (I301605,I301560);
nand I_17562 (I301319,I301402,I301605);
nor I_17563 (I301313,I301368,I301560);
not I_17564 (I301650,I468832);
nor I_17565 (I301667,I301650,I468820);
nand I_17566 (I301684,I301667,I301509);
nor I_17567 (I301322,I301427,I301684);
nor I_17568 (I301715,I301650,I468811);
and I_17569 (I301732,I301715,I468814);
or I_17570 (I301749,I301732,I468826);
DFFARX1 I_17571 (I301749,I3035,I301342,I301775,);
nor I_17572 (I301783,I301775,I301526);
DFFARX1 I_17573 (I301783,I3035,I301342,I301310,);
DFFARX1 I_17574 (I301775,I3035,I301342,I301334,);
not I_17575 (I301828,I301775);
nor I_17576 (I301845,I301828,I301402);
nor I_17577 (I301862,I301667,I301845);
DFFARX1 I_17578 (I301862,I3035,I301342,I301331,);
not I_17579 (I301920,I3042);
DFFARX1 I_17580 (I637026,I3035,I301920,I301946,);
not I_17581 (I301954,I301946);
DFFARX1 I_17582 (I637032,I3035,I301920,I301980,);
not I_17583 (I301988,I637026);
nand I_17584 (I302005,I301988,I637029);
not I_17585 (I302022,I302005);
nor I_17586 (I302039,I302022,I637047);
nor I_17587 (I302056,I301954,I302039);
DFFARX1 I_17588 (I302056,I3035,I301920,I301906,);
not I_17589 (I302087,I637047);
nand I_17590 (I302104,I302087,I302022);
and I_17591 (I302121,I302087,I637050);
nand I_17592 (I302138,I302121,I637029);
nor I_17593 (I301903,I302138,I302087);
and I_17594 (I301894,I301980,I302138);
not I_17595 (I302183,I302138);
nand I_17596 (I301897,I301980,I302183);
nor I_17597 (I301891,I301946,I302138);
not I_17598 (I302228,I637035);
nor I_17599 (I302245,I302228,I637050);
nand I_17600 (I302262,I302245,I302087);
nor I_17601 (I301900,I302005,I302262);
nor I_17602 (I302293,I302228,I637041);
and I_17603 (I302310,I302293,I637038);
or I_17604 (I302327,I302310,I637044);
DFFARX1 I_17605 (I302327,I3035,I301920,I302353,);
nor I_17606 (I302361,I302353,I302104);
DFFARX1 I_17607 (I302361,I3035,I301920,I301888,);
DFFARX1 I_17608 (I302353,I3035,I301920,I301912,);
not I_17609 (I302406,I302353);
nor I_17610 (I302423,I302406,I301980);
nor I_17611 (I302440,I302245,I302423);
DFFARX1 I_17612 (I302440,I3035,I301920,I301909,);
not I_17613 (I302498,I3042);
DFFARX1 I_17614 (I108664,I3035,I302498,I302524,);
not I_17615 (I302532,I302524);
DFFARX1 I_17616 (I108649,I3035,I302498,I302558,);
not I_17617 (I302566,I108667);
nand I_17618 (I302583,I302566,I108652);
not I_17619 (I302600,I302583);
nor I_17620 (I302617,I302600,I108649);
nor I_17621 (I302634,I302532,I302617);
DFFARX1 I_17622 (I302634,I3035,I302498,I302484,);
not I_17623 (I302665,I108649);
nand I_17624 (I302682,I302665,I302600);
and I_17625 (I302699,I302665,I108652);
nand I_17626 (I302716,I302699,I108673);
nor I_17627 (I302481,I302716,I302665);
and I_17628 (I302472,I302558,I302716);
not I_17629 (I302761,I302716);
nand I_17630 (I302475,I302558,I302761);
nor I_17631 (I302469,I302524,I302716);
not I_17632 (I302806,I108661);
nor I_17633 (I302823,I302806,I108652);
nand I_17634 (I302840,I302823,I302665);
nor I_17635 (I302478,I302583,I302840);
nor I_17636 (I302871,I302806,I108655);
and I_17637 (I302888,I302871,I108670);
or I_17638 (I302905,I302888,I108658);
DFFARX1 I_17639 (I302905,I3035,I302498,I302931,);
nor I_17640 (I302939,I302931,I302682);
DFFARX1 I_17641 (I302939,I3035,I302498,I302466,);
DFFARX1 I_17642 (I302931,I3035,I302498,I302490,);
not I_17643 (I302984,I302931);
nor I_17644 (I303001,I302984,I302558);
nor I_17645 (I303018,I302823,I303001);
DFFARX1 I_17646 (I303018,I3035,I302498,I302487,);
not I_17647 (I303076,I3042);
DFFARX1 I_17648 (I653976,I3035,I303076,I303102,);
not I_17649 (I303110,I303102);
DFFARX1 I_17650 (I653970,I3035,I303076,I303136,);
not I_17651 (I303144,I653979);
nand I_17652 (I303161,I303144,I653958);
not I_17653 (I303178,I303161);
nor I_17654 (I303195,I303178,I653967);
nor I_17655 (I303212,I303110,I303195);
DFFARX1 I_17656 (I303212,I3035,I303076,I303062,);
not I_17657 (I303243,I653967);
nand I_17658 (I303260,I303243,I303178);
and I_17659 (I303277,I303243,I653982);
nand I_17660 (I303294,I303277,I653961);
nor I_17661 (I303059,I303294,I303243);
and I_17662 (I303050,I303136,I303294);
not I_17663 (I303339,I303294);
nand I_17664 (I303053,I303136,I303339);
nor I_17665 (I303047,I303102,I303294);
not I_17666 (I303384,I653964);
nor I_17667 (I303401,I303384,I653982);
nand I_17668 (I303418,I303401,I303243);
nor I_17669 (I303056,I303161,I303418);
nor I_17670 (I303449,I303384,I653973);
and I_17671 (I303466,I303449,I653961);
or I_17672 (I303483,I303466,I653958);
DFFARX1 I_17673 (I303483,I3035,I303076,I303509,);
nor I_17674 (I303517,I303509,I303260);
DFFARX1 I_17675 (I303517,I3035,I303076,I303044,);
DFFARX1 I_17676 (I303509,I3035,I303076,I303068,);
not I_17677 (I303562,I303509);
nor I_17678 (I303579,I303562,I303136);
nor I_17679 (I303596,I303401,I303579);
DFFARX1 I_17680 (I303596,I3035,I303076,I303065,);
not I_17681 (I303654,I3042);
DFFARX1 I_17682 (I60529,I3035,I303654,I303680,);
not I_17683 (I303688,I303680);
DFFARX1 I_17684 (I60508,I3035,I303654,I303714,);
not I_17685 (I303722,I60505);
nand I_17686 (I303739,I303722,I60520);
not I_17687 (I303756,I303739);
nor I_17688 (I303773,I303756,I60508);
nor I_17689 (I303790,I303688,I303773);
DFFARX1 I_17690 (I303790,I3035,I303654,I303640,);
not I_17691 (I303821,I60508);
nand I_17692 (I303838,I303821,I303756);
and I_17693 (I303855,I303821,I60511);
nand I_17694 (I303872,I303855,I60526);
nor I_17695 (I303637,I303872,I303821);
and I_17696 (I303628,I303714,I303872);
not I_17697 (I303917,I303872);
nand I_17698 (I303631,I303714,I303917);
nor I_17699 (I303625,I303680,I303872);
not I_17700 (I303962,I60517);
nor I_17701 (I303979,I303962,I60511);
nand I_17702 (I303996,I303979,I303821);
nor I_17703 (I303634,I303739,I303996);
nor I_17704 (I304027,I303962,I60505);
and I_17705 (I304044,I304027,I60514);
or I_17706 (I304061,I304044,I60523);
DFFARX1 I_17707 (I304061,I3035,I303654,I304087,);
nor I_17708 (I304095,I304087,I303838);
DFFARX1 I_17709 (I304095,I3035,I303654,I303622,);
DFFARX1 I_17710 (I304087,I3035,I303654,I303646,);
not I_17711 (I304140,I304087);
nor I_17712 (I304157,I304140,I303714);
nor I_17713 (I304174,I303979,I304157);
DFFARX1 I_17714 (I304174,I3035,I303654,I303643,);
not I_17715 (I304232,I3042);
DFFARX1 I_17716 (I344660,I3035,I304232,I304258,);
not I_17717 (I304266,I304258);
DFFARX1 I_17718 (I344672,I3035,I304232,I304292,);
not I_17719 (I304300,I344663);
nand I_17720 (I304317,I304300,I344666);
not I_17721 (I304334,I304317);
nor I_17722 (I304351,I304334,I344669);
nor I_17723 (I304368,I304266,I304351);
DFFARX1 I_17724 (I304368,I3035,I304232,I304218,);
not I_17725 (I304399,I344669);
nand I_17726 (I304416,I304399,I304334);
and I_17727 (I304433,I304399,I344663);
nand I_17728 (I304450,I304433,I344675);
nor I_17729 (I304215,I304450,I304399);
and I_17730 (I304206,I304292,I304450);
not I_17731 (I304495,I304450);
nand I_17732 (I304209,I304292,I304495);
nor I_17733 (I304203,I304258,I304450);
not I_17734 (I304540,I344681);
nor I_17735 (I304557,I304540,I344663);
nand I_17736 (I304574,I304557,I304399);
nor I_17737 (I304212,I304317,I304574);
nor I_17738 (I304605,I304540,I344660);
and I_17739 (I304622,I304605,I344678);
or I_17740 (I304639,I304622,I344684);
DFFARX1 I_17741 (I304639,I3035,I304232,I304665,);
nor I_17742 (I304673,I304665,I304416);
DFFARX1 I_17743 (I304673,I3035,I304232,I304200,);
DFFARX1 I_17744 (I304665,I3035,I304232,I304224,);
not I_17745 (I304718,I304665);
nor I_17746 (I304735,I304718,I304292);
nor I_17747 (I304752,I304557,I304735);
DFFARX1 I_17748 (I304752,I3035,I304232,I304221,);
not I_17749 (I304810,I3042);
DFFARX1 I_17750 (I654520,I3035,I304810,I304836,);
not I_17751 (I304844,I304836);
DFFARX1 I_17752 (I654514,I3035,I304810,I304870,);
not I_17753 (I304878,I654523);
nand I_17754 (I304895,I304878,I654502);
not I_17755 (I304912,I304895);
nor I_17756 (I304929,I304912,I654511);
nor I_17757 (I304946,I304844,I304929);
DFFARX1 I_17758 (I304946,I3035,I304810,I304796,);
not I_17759 (I304977,I654511);
nand I_17760 (I304994,I304977,I304912);
and I_17761 (I305011,I304977,I654526);
nand I_17762 (I305028,I305011,I654505);
nor I_17763 (I304793,I305028,I304977);
and I_17764 (I304784,I304870,I305028);
not I_17765 (I305073,I305028);
nand I_17766 (I304787,I304870,I305073);
nor I_17767 (I304781,I304836,I305028);
not I_17768 (I305118,I654508);
nor I_17769 (I305135,I305118,I654526);
nand I_17770 (I305152,I305135,I304977);
nor I_17771 (I304790,I304895,I305152);
nor I_17772 (I305183,I305118,I654517);
and I_17773 (I305200,I305183,I654505);
or I_17774 (I305217,I305200,I654502);
DFFARX1 I_17775 (I305217,I3035,I304810,I305243,);
nor I_17776 (I305251,I305243,I304994);
DFFARX1 I_17777 (I305251,I3035,I304810,I304778,);
DFFARX1 I_17778 (I305243,I3035,I304810,I304802,);
not I_17779 (I305296,I305243);
nor I_17780 (I305313,I305296,I304870);
nor I_17781 (I305330,I305135,I305313);
DFFARX1 I_17782 (I305330,I3035,I304810,I304799,);
not I_17783 (I305388,I3042);
DFFARX1 I_17784 (I196154,I3035,I305388,I305414,);
not I_17785 (I305422,I305414);
DFFARX1 I_17786 (I196169,I3035,I305388,I305448,);
not I_17787 (I305456,I196172);
nand I_17788 (I305473,I305456,I196151);
not I_17789 (I305490,I305473);
nor I_17790 (I305507,I305490,I196175);
nor I_17791 (I305524,I305422,I305507);
DFFARX1 I_17792 (I305524,I3035,I305388,I305374,);
not I_17793 (I305555,I196175);
nand I_17794 (I305572,I305555,I305490);
and I_17795 (I305589,I305555,I196157);
nand I_17796 (I305606,I305589,I196148);
nor I_17797 (I305371,I305606,I305555);
and I_17798 (I305362,I305448,I305606);
not I_17799 (I305651,I305606);
nand I_17800 (I305365,I305448,I305651);
nor I_17801 (I305359,I305414,I305606);
not I_17802 (I305696,I196148);
nor I_17803 (I305713,I305696,I196157);
nand I_17804 (I305730,I305713,I305555);
nor I_17805 (I305368,I305473,I305730);
nor I_17806 (I305761,I305696,I196163);
and I_17807 (I305778,I305761,I196166);
or I_17808 (I305795,I305778,I196160);
DFFARX1 I_17809 (I305795,I3035,I305388,I305821,);
nor I_17810 (I305829,I305821,I305572);
DFFARX1 I_17811 (I305829,I3035,I305388,I305356,);
DFFARX1 I_17812 (I305821,I3035,I305388,I305380,);
not I_17813 (I305874,I305821);
nor I_17814 (I305891,I305874,I305448);
nor I_17815 (I305908,I305713,I305891);
DFFARX1 I_17816 (I305908,I3035,I305388,I305377,);
not I_17817 (I305966,I3042);
DFFARX1 I_17818 (I416910,I3035,I305966,I305992,);
not I_17819 (I306000,I305992);
DFFARX1 I_17820 (I416922,I3035,I305966,I306026,);
not I_17821 (I306034,I416913);
nand I_17822 (I306051,I306034,I416916);
not I_17823 (I306068,I306051);
nor I_17824 (I306085,I306068,I416919);
nor I_17825 (I306102,I306000,I306085);
DFFARX1 I_17826 (I306102,I3035,I305966,I305952,);
not I_17827 (I306133,I416919);
nand I_17828 (I306150,I306133,I306068);
and I_17829 (I306167,I306133,I416913);
nand I_17830 (I306184,I306167,I416925);
nor I_17831 (I305949,I306184,I306133);
and I_17832 (I305940,I306026,I306184);
not I_17833 (I306229,I306184);
nand I_17834 (I305943,I306026,I306229);
nor I_17835 (I305937,I305992,I306184);
not I_17836 (I306274,I416931);
nor I_17837 (I306291,I306274,I416913);
nand I_17838 (I306308,I306291,I306133);
nor I_17839 (I305946,I306051,I306308);
nor I_17840 (I306339,I306274,I416910);
and I_17841 (I306356,I306339,I416928);
or I_17842 (I306373,I306356,I416934);
DFFARX1 I_17843 (I306373,I3035,I305966,I306399,);
nor I_17844 (I306407,I306399,I306150);
DFFARX1 I_17845 (I306407,I3035,I305966,I305934,);
DFFARX1 I_17846 (I306399,I3035,I305966,I305958,);
not I_17847 (I306452,I306399);
nor I_17848 (I306469,I306452,I306026);
nor I_17849 (I306486,I306291,I306469);
DFFARX1 I_17850 (I306486,I3035,I305966,I305955,);
not I_17851 (I306544,I3042);
DFFARX1 I_17852 (I201951,I3035,I306544,I306570,);
not I_17853 (I306578,I306570);
DFFARX1 I_17854 (I201966,I3035,I306544,I306604,);
not I_17855 (I306612,I201969);
nand I_17856 (I306629,I306612,I201948);
not I_17857 (I306646,I306629);
nor I_17858 (I306663,I306646,I201972);
nor I_17859 (I306680,I306578,I306663);
DFFARX1 I_17860 (I306680,I3035,I306544,I306530,);
not I_17861 (I306711,I201972);
nand I_17862 (I306728,I306711,I306646);
and I_17863 (I306745,I306711,I201954);
nand I_17864 (I306762,I306745,I201945);
nor I_17865 (I306527,I306762,I306711);
and I_17866 (I306518,I306604,I306762);
not I_17867 (I306807,I306762);
nand I_17868 (I306521,I306604,I306807);
nor I_17869 (I306515,I306570,I306762);
not I_17870 (I306852,I201945);
nor I_17871 (I306869,I306852,I201954);
nand I_17872 (I306886,I306869,I306711);
nor I_17873 (I306524,I306629,I306886);
nor I_17874 (I306917,I306852,I201960);
and I_17875 (I306934,I306917,I201963);
or I_17876 (I306951,I306934,I201957);
DFFARX1 I_17877 (I306951,I3035,I306544,I306977,);
nor I_17878 (I306985,I306977,I306728);
DFFARX1 I_17879 (I306985,I3035,I306544,I306512,);
DFFARX1 I_17880 (I306977,I3035,I306544,I306536,);
not I_17881 (I307030,I306977);
nor I_17882 (I307047,I307030,I306604);
nor I_17883 (I307064,I306869,I307047);
DFFARX1 I_17884 (I307064,I3035,I306544,I306533,);
not I_17885 (I307122,I3042);
DFFARX1 I_17886 (I502562,I3035,I307122,I307148,);
not I_17887 (I307156,I307148);
DFFARX1 I_17888 (I502559,I3035,I307122,I307182,);
not I_17889 (I307190,I502556);
nand I_17890 (I307207,I307190,I502583);
not I_17891 (I307224,I307207);
nor I_17892 (I307241,I307224,I502571);
nor I_17893 (I307258,I307156,I307241);
DFFARX1 I_17894 (I307258,I3035,I307122,I307108,);
not I_17895 (I307289,I502571);
nand I_17896 (I307306,I307289,I307224);
and I_17897 (I307323,I307289,I502577);
nand I_17898 (I307340,I307323,I502568);
nor I_17899 (I307105,I307340,I307289);
and I_17900 (I307096,I307182,I307340);
not I_17901 (I307385,I307340);
nand I_17902 (I307099,I307182,I307385);
nor I_17903 (I307093,I307148,I307340);
not I_17904 (I307430,I502565);
nor I_17905 (I307447,I307430,I502577);
nand I_17906 (I307464,I307447,I307289);
nor I_17907 (I307102,I307207,I307464);
nor I_17908 (I307495,I307430,I502580);
and I_17909 (I307512,I307495,I502574);
or I_17910 (I307529,I307512,I502556);
DFFARX1 I_17911 (I307529,I3035,I307122,I307555,);
nor I_17912 (I307563,I307555,I307306);
DFFARX1 I_17913 (I307563,I3035,I307122,I307090,);
DFFARX1 I_17914 (I307555,I3035,I307122,I307114,);
not I_17915 (I307608,I307555);
nor I_17916 (I307625,I307608,I307182);
nor I_17917 (I307642,I307447,I307625);
DFFARX1 I_17918 (I307642,I3035,I307122,I307111,);
not I_17919 (I307700,I3042);
DFFARX1 I_17920 (I716858,I3035,I307700,I307726,);
not I_17921 (I307734,I307726);
DFFARX1 I_17922 (I716858,I3035,I307700,I307760,);
not I_17923 (I307768,I716882);
nand I_17924 (I307785,I307768,I716864);
not I_17925 (I307802,I307785);
nor I_17926 (I307819,I307802,I716879);
nor I_17927 (I307836,I307734,I307819);
DFFARX1 I_17928 (I307836,I3035,I307700,I307686,);
not I_17929 (I307867,I716879);
nand I_17930 (I307884,I307867,I307802);
and I_17931 (I307901,I307867,I716861);
nand I_17932 (I307918,I307901,I716870);
nor I_17933 (I307683,I307918,I307867);
and I_17934 (I307674,I307760,I307918);
not I_17935 (I307963,I307918);
nand I_17936 (I307677,I307760,I307963);
nor I_17937 (I307671,I307726,I307918);
not I_17938 (I308008,I716867);
nor I_17939 (I308025,I308008,I716861);
nand I_17940 (I308042,I308025,I307867);
nor I_17941 (I307680,I307785,I308042);
nor I_17942 (I308073,I308008,I716876);
and I_17943 (I308090,I308073,I716885);
or I_17944 (I308107,I308090,I716873);
DFFARX1 I_17945 (I308107,I3035,I307700,I308133,);
nor I_17946 (I308141,I308133,I307884);
DFFARX1 I_17947 (I308141,I3035,I307700,I307668,);
DFFARX1 I_17948 (I308133,I3035,I307700,I307692,);
not I_17949 (I308186,I308133);
nor I_17950 (I308203,I308186,I307760);
nor I_17951 (I308220,I308025,I308203);
DFFARX1 I_17952 (I308220,I3035,I307700,I307689,);
not I_17953 (I308278,I3042);
DFFARX1 I_17954 (I379918,I3035,I308278,I308304,);
not I_17955 (I308312,I308304);
DFFARX1 I_17956 (I379930,I3035,I308278,I308338,);
not I_17957 (I308346,I379921);
nand I_17958 (I308363,I308346,I379924);
not I_17959 (I308380,I308363);
nor I_17960 (I308397,I308380,I379927);
nor I_17961 (I308414,I308312,I308397);
DFFARX1 I_17962 (I308414,I3035,I308278,I308264,);
not I_17963 (I308445,I379927);
nand I_17964 (I308462,I308445,I308380);
and I_17965 (I308479,I308445,I379921);
nand I_17966 (I308496,I308479,I379933);
nor I_17967 (I308261,I308496,I308445);
and I_17968 (I308252,I308338,I308496);
not I_17969 (I308541,I308496);
nand I_17970 (I308255,I308338,I308541);
nor I_17971 (I308249,I308304,I308496);
not I_17972 (I308586,I379939);
nor I_17973 (I308603,I308586,I379921);
nand I_17974 (I308620,I308603,I308445);
nor I_17975 (I308258,I308363,I308620);
nor I_17976 (I308651,I308586,I379918);
and I_17977 (I308668,I308651,I379936);
or I_17978 (I308685,I308668,I379942);
DFFARX1 I_17979 (I308685,I3035,I308278,I308711,);
nor I_17980 (I308719,I308711,I308462);
DFFARX1 I_17981 (I308719,I3035,I308278,I308246,);
DFFARX1 I_17982 (I308711,I3035,I308278,I308270,);
not I_17983 (I308764,I308711);
nor I_17984 (I308781,I308764,I308338);
nor I_17985 (I308798,I308603,I308781);
DFFARX1 I_17986 (I308798,I3035,I308278,I308267,);
not I_17987 (I308856,I3042);
DFFARX1 I_17988 (I678280,I3035,I308856,I308882,);
not I_17989 (I308890,I308882);
DFFARX1 I_17990 (I678292,I3035,I308856,I308916,);
not I_17991 (I308924,I678283);
nand I_17992 (I308941,I308924,I678271);
not I_17993 (I308958,I308941);
nor I_17994 (I308975,I308958,I678268);
nor I_17995 (I308992,I308890,I308975);
DFFARX1 I_17996 (I308992,I3035,I308856,I308842,);
not I_17997 (I309023,I678268);
nand I_17998 (I309040,I309023,I308958);
and I_17999 (I309057,I309023,I678274);
nand I_18000 (I309074,I309057,I678271);
nor I_18001 (I308839,I309074,I309023);
and I_18002 (I308830,I308916,I309074);
not I_18003 (I309119,I309074);
nand I_18004 (I308833,I308916,I309119);
nor I_18005 (I308827,I308882,I309074);
not I_18006 (I309164,I678289);
nor I_18007 (I309181,I309164,I678274);
nand I_18008 (I309198,I309181,I309023);
nor I_18009 (I308836,I308941,I309198);
nor I_18010 (I309229,I309164,I678277);
and I_18011 (I309246,I309229,I678268);
or I_18012 (I309263,I309246,I678286);
DFFARX1 I_18013 (I309263,I3035,I308856,I309289,);
nor I_18014 (I309297,I309289,I309040);
DFFARX1 I_18015 (I309297,I3035,I308856,I308824,);
DFFARX1 I_18016 (I309289,I3035,I308856,I308848,);
not I_18017 (I309342,I309289);
nor I_18018 (I309359,I309342,I308916);
nor I_18019 (I309376,I309181,I309359);
DFFARX1 I_18020 (I309376,I3035,I308856,I308845,);
not I_18021 (I309434,I3042);
DFFARX1 I_18022 (I227247,I3035,I309434,I309460,);
not I_18023 (I309468,I309460);
DFFARX1 I_18024 (I227262,I3035,I309434,I309494,);
not I_18025 (I309502,I227265);
nand I_18026 (I309519,I309502,I227244);
not I_18027 (I309536,I309519);
nor I_18028 (I309553,I309536,I227268);
nor I_18029 (I309570,I309468,I309553);
DFFARX1 I_18030 (I309570,I3035,I309434,I309420,);
not I_18031 (I309601,I227268);
nand I_18032 (I309618,I309601,I309536);
and I_18033 (I309635,I309601,I227250);
nand I_18034 (I309652,I309635,I227241);
nor I_18035 (I309417,I309652,I309601);
and I_18036 (I309408,I309494,I309652);
not I_18037 (I309697,I309652);
nand I_18038 (I309411,I309494,I309697);
nor I_18039 (I309405,I309460,I309652);
not I_18040 (I309742,I227241);
nor I_18041 (I309759,I309742,I227250);
nand I_18042 (I309776,I309759,I309601);
nor I_18043 (I309414,I309519,I309776);
nor I_18044 (I309807,I309742,I227256);
and I_18045 (I309824,I309807,I227259);
or I_18046 (I309841,I309824,I227253);
DFFARX1 I_18047 (I309841,I3035,I309434,I309867,);
nor I_18048 (I309875,I309867,I309618);
DFFARX1 I_18049 (I309875,I3035,I309434,I309402,);
DFFARX1 I_18050 (I309867,I3035,I309434,I309426,);
not I_18051 (I309920,I309867);
nor I_18052 (I309937,I309920,I309494);
nor I_18053 (I309954,I309759,I309937);
DFFARX1 I_18054 (I309954,I3035,I309434,I309423,);
not I_18055 (I310012,I3042);
DFFARX1 I_18056 (I478014,I3035,I310012,I310038,);
not I_18057 (I310046,I310038);
DFFARX1 I_18058 (I478011,I3035,I310012,I310072,);
not I_18059 (I310080,I478008);
nand I_18060 (I310097,I310080,I478035);
not I_18061 (I310114,I310097);
nor I_18062 (I310131,I310114,I478023);
nor I_18063 (I310148,I310046,I310131);
DFFARX1 I_18064 (I310148,I3035,I310012,I309998,);
not I_18065 (I310179,I478023);
nand I_18066 (I310196,I310179,I310114);
and I_18067 (I310213,I310179,I478029);
nand I_18068 (I310230,I310213,I478020);
nor I_18069 (I309995,I310230,I310179);
and I_18070 (I309986,I310072,I310230);
not I_18071 (I310275,I310230);
nand I_18072 (I309989,I310072,I310275);
nor I_18073 (I309983,I310038,I310230);
not I_18074 (I310320,I478017);
nor I_18075 (I310337,I310320,I478029);
nand I_18076 (I310354,I310337,I310179);
nor I_18077 (I309992,I310097,I310354);
nor I_18078 (I310385,I310320,I478032);
and I_18079 (I310402,I310385,I478026);
or I_18080 (I310419,I310402,I478008);
DFFARX1 I_18081 (I310419,I3035,I310012,I310445,);
nor I_18082 (I310453,I310445,I310196);
DFFARX1 I_18083 (I310453,I3035,I310012,I309980,);
DFFARX1 I_18084 (I310445,I3035,I310012,I310004,);
not I_18085 (I310498,I310445);
nor I_18086 (I310515,I310498,I310072);
nor I_18087 (I310532,I310337,I310515);
DFFARX1 I_18088 (I310532,I3035,I310012,I310001,);
not I_18089 (I310590,I3042);
DFFARX1 I_18090 (I721618,I3035,I310590,I310616,);
not I_18091 (I310624,I310616);
DFFARX1 I_18092 (I721618,I3035,I310590,I310650,);
not I_18093 (I310658,I721642);
nand I_18094 (I310675,I310658,I721624);
not I_18095 (I310692,I310675);
nor I_18096 (I310709,I310692,I721639);
nor I_18097 (I310726,I310624,I310709);
DFFARX1 I_18098 (I310726,I3035,I310590,I310576,);
not I_18099 (I310757,I721639);
nand I_18100 (I310774,I310757,I310692);
and I_18101 (I310791,I310757,I721621);
nand I_18102 (I310808,I310791,I721630);
nor I_18103 (I310573,I310808,I310757);
and I_18104 (I310564,I310650,I310808);
not I_18105 (I310853,I310808);
nand I_18106 (I310567,I310650,I310853);
nor I_18107 (I310561,I310616,I310808);
not I_18108 (I310898,I721627);
nor I_18109 (I310915,I310898,I721621);
nand I_18110 (I310932,I310915,I310757);
nor I_18111 (I310570,I310675,I310932);
nor I_18112 (I310963,I310898,I721636);
and I_18113 (I310980,I310963,I721645);
or I_18114 (I310997,I310980,I721633);
DFFARX1 I_18115 (I310997,I3035,I310590,I311023,);
nor I_18116 (I311031,I311023,I310774);
DFFARX1 I_18117 (I311031,I3035,I310590,I310558,);
DFFARX1 I_18118 (I311023,I3035,I310590,I310582,);
not I_18119 (I311076,I311023);
nor I_18120 (I311093,I311076,I310650);
nor I_18121 (I311110,I310915,I311093);
DFFARX1 I_18122 (I311110,I3035,I310590,I310579,);
not I_18123 (I311168,I3042);
DFFARX1 I_18124 (I506438,I3035,I311168,I311194,);
not I_18125 (I311202,I311194);
DFFARX1 I_18126 (I506435,I3035,I311168,I311228,);
not I_18127 (I311236,I506432);
nand I_18128 (I311253,I311236,I506459);
not I_18129 (I311270,I311253);
nor I_18130 (I311287,I311270,I506447);
nor I_18131 (I311304,I311202,I311287);
DFFARX1 I_18132 (I311304,I3035,I311168,I311154,);
not I_18133 (I311335,I506447);
nand I_18134 (I311352,I311335,I311270);
and I_18135 (I311369,I311335,I506453);
nand I_18136 (I311386,I311369,I506444);
nor I_18137 (I311151,I311386,I311335);
and I_18138 (I311142,I311228,I311386);
not I_18139 (I311431,I311386);
nand I_18140 (I311145,I311228,I311431);
nor I_18141 (I311139,I311194,I311386);
not I_18142 (I311476,I506441);
nor I_18143 (I311493,I311476,I506453);
nand I_18144 (I311510,I311493,I311335);
nor I_18145 (I311148,I311253,I311510);
nor I_18146 (I311541,I311476,I506456);
and I_18147 (I311558,I311541,I506450);
or I_18148 (I311575,I311558,I506432);
DFFARX1 I_18149 (I311575,I3035,I311168,I311601,);
nor I_18150 (I311609,I311601,I311352);
DFFARX1 I_18151 (I311609,I3035,I311168,I311136,);
DFFARX1 I_18152 (I311601,I3035,I311168,I311160,);
not I_18153 (I311654,I311601);
nor I_18154 (I311671,I311654,I311228);
nor I_18155 (I311688,I311493,I311671);
DFFARX1 I_18156 (I311688,I3035,I311168,I311157,);
not I_18157 (I311746,I3042);
DFFARX1 I_18158 (I490934,I3035,I311746,I311772,);
not I_18159 (I311780,I311772);
DFFARX1 I_18160 (I490931,I3035,I311746,I311806,);
not I_18161 (I311814,I490928);
nand I_18162 (I311831,I311814,I490955);
not I_18163 (I311848,I311831);
nor I_18164 (I311865,I311848,I490943);
nor I_18165 (I311882,I311780,I311865);
DFFARX1 I_18166 (I311882,I3035,I311746,I311732,);
not I_18167 (I311913,I490943);
nand I_18168 (I311930,I311913,I311848);
and I_18169 (I311947,I311913,I490949);
nand I_18170 (I311964,I311947,I490940);
nor I_18171 (I311729,I311964,I311913);
and I_18172 (I311720,I311806,I311964);
not I_18173 (I312009,I311964);
nand I_18174 (I311723,I311806,I312009);
nor I_18175 (I311717,I311772,I311964);
not I_18176 (I312054,I490937);
nor I_18177 (I312071,I312054,I490949);
nand I_18178 (I312088,I312071,I311913);
nor I_18179 (I311726,I311831,I312088);
nor I_18180 (I312119,I312054,I490952);
and I_18181 (I312136,I312119,I490946);
or I_18182 (I312153,I312136,I490928);
DFFARX1 I_18183 (I312153,I3035,I311746,I312179,);
nor I_18184 (I312187,I312179,I311930);
DFFARX1 I_18185 (I312187,I3035,I311746,I311714,);
DFFARX1 I_18186 (I312179,I3035,I311746,I311738,);
not I_18187 (I312232,I312179);
nor I_18188 (I312249,I312232,I311806);
nor I_18189 (I312266,I312071,I312249);
DFFARX1 I_18190 (I312266,I3035,I311746,I311735,);
not I_18191 (I312324,I3042);
DFFARX1 I_18192 (I105689,I3035,I312324,I312350,);
not I_18193 (I312358,I312350);
DFFARX1 I_18194 (I105674,I3035,I312324,I312384,);
not I_18195 (I312392,I105692);
nand I_18196 (I312409,I312392,I105677);
not I_18197 (I312426,I312409);
nor I_18198 (I312443,I312426,I105674);
nor I_18199 (I312460,I312358,I312443);
DFFARX1 I_18200 (I312460,I3035,I312324,I312310,);
not I_18201 (I312491,I105674);
nand I_18202 (I312508,I312491,I312426);
and I_18203 (I312525,I312491,I105677);
nand I_18204 (I312542,I312525,I105698);
nor I_18205 (I312307,I312542,I312491);
and I_18206 (I312298,I312384,I312542);
not I_18207 (I312587,I312542);
nand I_18208 (I312301,I312384,I312587);
nor I_18209 (I312295,I312350,I312542);
not I_18210 (I312632,I105686);
nor I_18211 (I312649,I312632,I105677);
nand I_18212 (I312666,I312649,I312491);
nor I_18213 (I312304,I312409,I312666);
nor I_18214 (I312697,I312632,I105680);
and I_18215 (I312714,I312697,I105695);
or I_18216 (I312731,I312714,I105683);
DFFARX1 I_18217 (I312731,I3035,I312324,I312757,);
nor I_18218 (I312765,I312757,I312508);
DFFARX1 I_18219 (I312765,I3035,I312324,I312292,);
DFFARX1 I_18220 (I312757,I3035,I312324,I312316,);
not I_18221 (I312810,I312757);
nor I_18222 (I312827,I312810,I312384);
nor I_18223 (I312844,I312649,I312827);
DFFARX1 I_18224 (I312844,I3035,I312324,I312313,);
not I_18225 (I312902,I3042);
DFFARX1 I_18226 (I246769,I3035,I312902,I312928,);
not I_18227 (I312936,I312928);
DFFARX1 I_18228 (I246781,I3035,I312902,I312962,);
not I_18229 (I312970,I246757);
nand I_18230 (I312987,I312970,I246784);
not I_18231 (I313004,I312987);
nor I_18232 (I313021,I313004,I246772);
nor I_18233 (I313038,I312936,I313021);
DFFARX1 I_18234 (I313038,I3035,I312902,I312888,);
not I_18235 (I313069,I246772);
nand I_18236 (I313086,I313069,I313004);
and I_18237 (I313103,I313069,I246757);
nand I_18238 (I313120,I313103,I246760);
nor I_18239 (I312885,I313120,I313069);
and I_18240 (I312876,I312962,I313120);
not I_18241 (I313165,I313120);
nand I_18242 (I312879,I312962,I313165);
nor I_18243 (I312873,I312928,I313120);
not I_18244 (I313210,I246766);
nor I_18245 (I313227,I313210,I246757);
nand I_18246 (I313244,I313227,I313069);
nor I_18247 (I312882,I312987,I313244);
nor I_18248 (I313275,I313210,I246775);
and I_18249 (I313292,I313275,I246763);
or I_18250 (I313309,I313292,I246778);
DFFARX1 I_18251 (I313309,I3035,I312902,I313335,);
nor I_18252 (I313343,I313335,I313086);
DFFARX1 I_18253 (I313343,I3035,I312902,I312870,);
DFFARX1 I_18254 (I313335,I3035,I312902,I312894,);
not I_18255 (I313388,I313335);
nor I_18256 (I313405,I313388,I312962);
nor I_18257 (I313422,I313227,I313405);
DFFARX1 I_18258 (I313422,I3035,I312902,I312891,);
not I_18259 (I313480,I3042);
DFFARX1 I_18260 (I115804,I3035,I313480,I313506,);
not I_18261 (I313514,I313506);
DFFARX1 I_18262 (I115789,I3035,I313480,I313540,);
not I_18263 (I313548,I115807);
nand I_18264 (I313565,I313548,I115792);
not I_18265 (I313582,I313565);
nor I_18266 (I313599,I313582,I115789);
nor I_18267 (I313616,I313514,I313599);
DFFARX1 I_18268 (I313616,I3035,I313480,I313466,);
not I_18269 (I313647,I115789);
nand I_18270 (I313664,I313647,I313582);
and I_18271 (I313681,I313647,I115792);
nand I_18272 (I313698,I313681,I115813);
nor I_18273 (I313463,I313698,I313647);
and I_18274 (I313454,I313540,I313698);
not I_18275 (I313743,I313698);
nand I_18276 (I313457,I313540,I313743);
nor I_18277 (I313451,I313506,I313698);
not I_18278 (I313788,I115801);
nor I_18279 (I313805,I313788,I115792);
nand I_18280 (I313822,I313805,I313647);
nor I_18281 (I313460,I313565,I313822);
nor I_18282 (I313853,I313788,I115795);
and I_18283 (I313870,I313853,I115810);
or I_18284 (I313887,I313870,I115798);
DFFARX1 I_18285 (I313887,I3035,I313480,I313913,);
nor I_18286 (I313921,I313913,I313664);
DFFARX1 I_18287 (I313921,I3035,I313480,I313448,);
DFFARX1 I_18288 (I313913,I3035,I313480,I313472,);
not I_18289 (I313966,I313913);
nor I_18290 (I313983,I313966,I313540);
nor I_18291 (I314000,I313805,I313983);
DFFARX1 I_18292 (I314000,I3035,I313480,I313469,);
not I_18293 (I314058,I3042);
DFFARX1 I_18294 (I415754,I3035,I314058,I314084,);
not I_18295 (I314092,I314084);
DFFARX1 I_18296 (I415766,I3035,I314058,I314118,);
not I_18297 (I314126,I415757);
nand I_18298 (I314143,I314126,I415760);
not I_18299 (I314160,I314143);
nor I_18300 (I314177,I314160,I415763);
nor I_18301 (I314194,I314092,I314177);
DFFARX1 I_18302 (I314194,I3035,I314058,I314044,);
not I_18303 (I314225,I415763);
nand I_18304 (I314242,I314225,I314160);
and I_18305 (I314259,I314225,I415757);
nand I_18306 (I314276,I314259,I415769);
nor I_18307 (I314041,I314276,I314225);
and I_18308 (I314032,I314118,I314276);
not I_18309 (I314321,I314276);
nand I_18310 (I314035,I314118,I314321);
nor I_18311 (I314029,I314084,I314276);
not I_18312 (I314366,I415775);
nor I_18313 (I314383,I314366,I415757);
nand I_18314 (I314400,I314383,I314225);
nor I_18315 (I314038,I314143,I314400);
nor I_18316 (I314431,I314366,I415754);
and I_18317 (I314448,I314431,I415772);
or I_18318 (I314465,I314448,I415778);
DFFARX1 I_18319 (I314465,I3035,I314058,I314491,);
nor I_18320 (I314499,I314491,I314242);
DFFARX1 I_18321 (I314499,I3035,I314058,I314026,);
DFFARX1 I_18322 (I314491,I3035,I314058,I314050,);
not I_18323 (I314544,I314491);
nor I_18324 (I314561,I314544,I314118);
nor I_18325 (I314578,I314383,I314561);
DFFARX1 I_18326 (I314578,I3035,I314058,I314047,);
not I_18327 (I314636,I3042);
DFFARX1 I_18328 (I298984,I3035,I314636,I314662,);
not I_18329 (I314670,I314662);
DFFARX1 I_18330 (I298996,I3035,I314636,I314696,);
not I_18331 (I314704,I299002);
nand I_18332 (I314721,I314704,I298993);
not I_18333 (I314738,I314721);
nor I_18334 (I314755,I314738,I298999);
nor I_18335 (I314772,I314670,I314755);
DFFARX1 I_18336 (I314772,I3035,I314636,I314622,);
not I_18337 (I314803,I298999);
nand I_18338 (I314820,I314803,I314738);
and I_18339 (I314837,I314803,I298990);
nand I_18340 (I314854,I314837,I298981);
nor I_18341 (I314619,I314854,I314803);
and I_18342 (I314610,I314696,I314854);
not I_18343 (I314899,I314854);
nand I_18344 (I314613,I314696,I314899);
nor I_18345 (I314607,I314662,I314854);
not I_18346 (I314944,I298987);
nor I_18347 (I314961,I314944,I298990);
nand I_18348 (I314978,I314961,I314803);
nor I_18349 (I314616,I314721,I314978);
nor I_18350 (I315009,I314944,I298984);
and I_18351 (I315026,I315009,I298981);
or I_18352 (I315043,I315026,I299005);
DFFARX1 I_18353 (I315043,I3035,I314636,I315069,);
nor I_18354 (I315077,I315069,I314820);
DFFARX1 I_18355 (I315077,I3035,I314636,I314604,);
DFFARX1 I_18356 (I315069,I3035,I314636,I314628,);
not I_18357 (I315122,I315069);
nor I_18358 (I315139,I315122,I314696);
nor I_18359 (I315156,I314961,I315139);
DFFARX1 I_18360 (I315156,I3035,I314636,I314625,);
not I_18361 (I315214,I3042);
DFFARX1 I_18362 (I665400,I3035,I315214,I315240,);
not I_18363 (I315248,I315240);
DFFARX1 I_18364 (I665394,I3035,I315214,I315274,);
not I_18365 (I315282,I665403);
nand I_18366 (I315299,I315282,I665382);
not I_18367 (I315316,I315299);
nor I_18368 (I315333,I315316,I665391);
nor I_18369 (I315350,I315248,I315333);
DFFARX1 I_18370 (I315350,I3035,I315214,I315200,);
not I_18371 (I315381,I665391);
nand I_18372 (I315398,I315381,I315316);
and I_18373 (I315415,I315381,I665406);
nand I_18374 (I315432,I315415,I665385);
nor I_18375 (I315197,I315432,I315381);
and I_18376 (I315188,I315274,I315432);
not I_18377 (I315477,I315432);
nand I_18378 (I315191,I315274,I315477);
nor I_18379 (I315185,I315240,I315432);
not I_18380 (I315522,I665388);
nor I_18381 (I315539,I315522,I665406);
nand I_18382 (I315556,I315539,I315381);
nor I_18383 (I315194,I315299,I315556);
nor I_18384 (I315587,I315522,I665397);
and I_18385 (I315604,I315587,I665385);
or I_18386 (I315621,I315604,I665382);
DFFARX1 I_18387 (I315621,I3035,I315214,I315647,);
nor I_18388 (I315655,I315647,I315398);
DFFARX1 I_18389 (I315655,I3035,I315214,I315182,);
DFFARX1 I_18390 (I315647,I3035,I315214,I315206,);
not I_18391 (I315700,I315647);
nor I_18392 (I315717,I315700,I315274);
nor I_18393 (I315734,I315539,I315717);
DFFARX1 I_18394 (I315734,I3035,I315214,I315203,);
not I_18395 (I315792,I3042);
DFFARX1 I_18396 (I359688,I3035,I315792,I315818,);
not I_18397 (I315826,I315818);
DFFARX1 I_18398 (I359700,I3035,I315792,I315852,);
not I_18399 (I315860,I359691);
nand I_18400 (I315877,I315860,I359694);
not I_18401 (I315894,I315877);
nor I_18402 (I315911,I315894,I359697);
nor I_18403 (I315928,I315826,I315911);
DFFARX1 I_18404 (I315928,I3035,I315792,I315778,);
not I_18405 (I315959,I359697);
nand I_18406 (I315976,I315959,I315894);
and I_18407 (I315993,I315959,I359691);
nand I_18408 (I316010,I315993,I359703);
nor I_18409 (I315775,I316010,I315959);
and I_18410 (I315766,I315852,I316010);
not I_18411 (I316055,I316010);
nand I_18412 (I315769,I315852,I316055);
nor I_18413 (I315763,I315818,I316010);
not I_18414 (I316100,I359709);
nor I_18415 (I316117,I316100,I359691);
nand I_18416 (I316134,I316117,I315959);
nor I_18417 (I315772,I315877,I316134);
nor I_18418 (I316165,I316100,I359688);
and I_18419 (I316182,I316165,I359706);
or I_18420 (I316199,I316182,I359712);
DFFARX1 I_18421 (I316199,I3035,I315792,I316225,);
nor I_18422 (I316233,I316225,I315976);
DFFARX1 I_18423 (I316233,I3035,I315792,I315760,);
DFFARX1 I_18424 (I316225,I3035,I315792,I315784,);
not I_18425 (I316278,I316225);
nor I_18426 (I316295,I316278,I315852);
nor I_18427 (I316312,I316117,I316295);
DFFARX1 I_18428 (I316312,I3035,I315792,I315781,);
not I_18429 (I316370,I3042);
DFFARX1 I_18430 (I343504,I3035,I316370,I316396,);
not I_18431 (I316404,I316396);
DFFARX1 I_18432 (I343516,I3035,I316370,I316430,);
not I_18433 (I316438,I343507);
nand I_18434 (I316455,I316438,I343510);
not I_18435 (I316472,I316455);
nor I_18436 (I316489,I316472,I343513);
nor I_18437 (I316506,I316404,I316489);
DFFARX1 I_18438 (I316506,I3035,I316370,I316356,);
not I_18439 (I316537,I343513);
nand I_18440 (I316554,I316537,I316472);
and I_18441 (I316571,I316537,I343507);
nand I_18442 (I316588,I316571,I343519);
nor I_18443 (I316353,I316588,I316537);
and I_18444 (I316344,I316430,I316588);
not I_18445 (I316633,I316588);
nand I_18446 (I316347,I316430,I316633);
nor I_18447 (I316341,I316396,I316588);
not I_18448 (I316678,I343525);
nor I_18449 (I316695,I316678,I343507);
nand I_18450 (I316712,I316695,I316537);
nor I_18451 (I316350,I316455,I316712);
nor I_18452 (I316743,I316678,I343504);
and I_18453 (I316760,I316743,I343522);
or I_18454 (I316777,I316760,I343528);
DFFARX1 I_18455 (I316777,I3035,I316370,I316803,);
nor I_18456 (I316811,I316803,I316554);
DFFARX1 I_18457 (I316811,I3035,I316370,I316338,);
DFFARX1 I_18458 (I316803,I3035,I316370,I316362,);
not I_18459 (I316856,I316803);
nor I_18460 (I316873,I316856,I316430);
nor I_18461 (I316890,I316695,I316873);
DFFARX1 I_18462 (I316890,I3035,I316370,I316359,);
not I_18463 (I316948,I3042);
DFFARX1 I_18464 (I627778,I3035,I316948,I316974,);
not I_18465 (I316982,I316974);
DFFARX1 I_18466 (I627784,I3035,I316948,I317008,);
not I_18467 (I317016,I627778);
nand I_18468 (I317033,I317016,I627781);
not I_18469 (I317050,I317033);
nor I_18470 (I317067,I317050,I627799);
nor I_18471 (I317084,I316982,I317067);
DFFARX1 I_18472 (I317084,I3035,I316948,I316934,);
not I_18473 (I317115,I627799);
nand I_18474 (I317132,I317115,I317050);
and I_18475 (I317149,I317115,I627802);
nand I_18476 (I317166,I317149,I627781);
nor I_18477 (I316931,I317166,I317115);
and I_18478 (I316922,I317008,I317166);
not I_18479 (I317211,I317166);
nand I_18480 (I316925,I317008,I317211);
nor I_18481 (I316919,I316974,I317166);
not I_18482 (I317256,I627787);
nor I_18483 (I317273,I317256,I627802);
nand I_18484 (I317290,I317273,I317115);
nor I_18485 (I316928,I317033,I317290);
nor I_18486 (I317321,I317256,I627793);
and I_18487 (I317338,I317321,I627790);
or I_18488 (I317355,I317338,I627796);
DFFARX1 I_18489 (I317355,I3035,I316948,I317381,);
nor I_18490 (I317389,I317381,I317132);
DFFARX1 I_18491 (I317389,I3035,I316948,I316916,);
DFFARX1 I_18492 (I317381,I3035,I316948,I316940,);
not I_18493 (I317434,I317381);
nor I_18494 (I317451,I317434,I317008);
nor I_18495 (I317468,I317273,I317451);
DFFARX1 I_18496 (I317468,I3035,I316948,I316937,);
not I_18497 (I317526,I3042);
DFFARX1 I_18498 (I419222,I3035,I317526,I317552,);
not I_18499 (I317560,I317552);
DFFARX1 I_18500 (I419234,I3035,I317526,I317586,);
not I_18501 (I317594,I419225);
nand I_18502 (I317611,I317594,I419228);
not I_18503 (I317628,I317611);
nor I_18504 (I317645,I317628,I419231);
nor I_18505 (I317662,I317560,I317645);
DFFARX1 I_18506 (I317662,I3035,I317526,I317512,);
not I_18507 (I317693,I419231);
nand I_18508 (I317710,I317693,I317628);
and I_18509 (I317727,I317693,I419225);
nand I_18510 (I317744,I317727,I419237);
nor I_18511 (I317509,I317744,I317693);
and I_18512 (I317500,I317586,I317744);
not I_18513 (I317789,I317744);
nand I_18514 (I317503,I317586,I317789);
nor I_18515 (I317497,I317552,I317744);
not I_18516 (I317834,I419243);
nor I_18517 (I317851,I317834,I419225);
nand I_18518 (I317868,I317851,I317693);
nor I_18519 (I317506,I317611,I317868);
nor I_18520 (I317899,I317834,I419222);
and I_18521 (I317916,I317899,I419240);
or I_18522 (I317933,I317916,I419246);
DFFARX1 I_18523 (I317933,I3035,I317526,I317959,);
nor I_18524 (I317967,I317959,I317710);
DFFARX1 I_18525 (I317967,I3035,I317526,I317494,);
DFFARX1 I_18526 (I317959,I3035,I317526,I317518,);
not I_18527 (I318012,I317959);
nor I_18528 (I318029,I318012,I317586);
nor I_18529 (I318046,I317851,I318029);
DFFARX1 I_18530 (I318046,I3035,I317526,I317515,);
not I_18531 (I318104,I3042);
DFFARX1 I_18532 (I65272,I3035,I318104,I318130,);
not I_18533 (I318138,I318130);
DFFARX1 I_18534 (I65251,I3035,I318104,I318164,);
not I_18535 (I318172,I65248);
nand I_18536 (I318189,I318172,I65263);
not I_18537 (I318206,I318189);
nor I_18538 (I318223,I318206,I65251);
nor I_18539 (I318240,I318138,I318223);
DFFARX1 I_18540 (I318240,I3035,I318104,I318090,);
not I_18541 (I318271,I65251);
nand I_18542 (I318288,I318271,I318206);
and I_18543 (I318305,I318271,I65254);
nand I_18544 (I318322,I318305,I65269);
nor I_18545 (I318087,I318322,I318271);
and I_18546 (I318078,I318164,I318322);
not I_18547 (I318367,I318322);
nand I_18548 (I318081,I318164,I318367);
nor I_18549 (I318075,I318130,I318322);
not I_18550 (I318412,I65260);
nor I_18551 (I318429,I318412,I65254);
nand I_18552 (I318446,I318429,I318271);
nor I_18553 (I318084,I318189,I318446);
nor I_18554 (I318477,I318412,I65248);
and I_18555 (I318494,I318477,I65257);
or I_18556 (I318511,I318494,I65266);
DFFARX1 I_18557 (I318511,I3035,I318104,I318537,);
nor I_18558 (I318545,I318537,I318288);
DFFARX1 I_18559 (I318545,I3035,I318104,I318072,);
DFFARX1 I_18560 (I318537,I3035,I318104,I318096,);
not I_18561 (I318590,I318537);
nor I_18562 (I318607,I318590,I318164);
nor I_18563 (I318624,I318429,I318607);
DFFARX1 I_18564 (I318624,I3035,I318104,I318093,);
not I_18565 (I318682,I3042);
DFFARX1 I_18566 (I96764,I3035,I318682,I318708,);
not I_18567 (I318716,I318708);
DFFARX1 I_18568 (I96749,I3035,I318682,I318742,);
not I_18569 (I318750,I96767);
nand I_18570 (I318767,I318750,I96752);
not I_18571 (I318784,I318767);
nor I_18572 (I318801,I318784,I96749);
nor I_18573 (I318818,I318716,I318801);
DFFARX1 I_18574 (I318818,I3035,I318682,I318668,);
not I_18575 (I318849,I96749);
nand I_18576 (I318866,I318849,I318784);
and I_18577 (I318883,I318849,I96752);
nand I_18578 (I318900,I318883,I96773);
nor I_18579 (I318665,I318900,I318849);
and I_18580 (I318656,I318742,I318900);
not I_18581 (I318945,I318900);
nand I_18582 (I318659,I318742,I318945);
nor I_18583 (I318653,I318708,I318900);
not I_18584 (I318990,I96761);
nor I_18585 (I319007,I318990,I96752);
nand I_18586 (I319024,I319007,I318849);
nor I_18587 (I318662,I318767,I319024);
nor I_18588 (I319055,I318990,I96755);
and I_18589 (I319072,I319055,I96770);
or I_18590 (I319089,I319072,I96758);
DFFARX1 I_18591 (I319089,I3035,I318682,I319115,);
nor I_18592 (I319123,I319115,I318866);
DFFARX1 I_18593 (I319123,I3035,I318682,I318650,);
DFFARX1 I_18594 (I319115,I3035,I318682,I318674,);
not I_18595 (I319168,I319115);
nor I_18596 (I319185,I319168,I318742);
nor I_18597 (I319202,I319007,I319185);
DFFARX1 I_18598 (I319202,I3035,I318682,I318671,);
not I_18599 (I319260,I3042);
DFFARX1 I_18600 (I362578,I3035,I319260,I319286,);
not I_18601 (I319294,I319286);
DFFARX1 I_18602 (I362590,I3035,I319260,I319320,);
not I_18603 (I319328,I362581);
nand I_18604 (I319345,I319328,I362584);
not I_18605 (I319362,I319345);
nor I_18606 (I319379,I319362,I362587);
nor I_18607 (I319396,I319294,I319379);
DFFARX1 I_18608 (I319396,I3035,I319260,I319246,);
not I_18609 (I319427,I362587);
nand I_18610 (I319444,I319427,I319362);
and I_18611 (I319461,I319427,I362581);
nand I_18612 (I319478,I319461,I362593);
nor I_18613 (I319243,I319478,I319427);
and I_18614 (I319234,I319320,I319478);
not I_18615 (I319523,I319478);
nand I_18616 (I319237,I319320,I319523);
nor I_18617 (I319231,I319286,I319478);
not I_18618 (I319568,I362599);
nor I_18619 (I319585,I319568,I362581);
nand I_18620 (I319602,I319585,I319427);
nor I_18621 (I319240,I319345,I319602);
nor I_18622 (I319633,I319568,I362578);
and I_18623 (I319650,I319633,I362596);
or I_18624 (I319667,I319650,I362602);
DFFARX1 I_18625 (I319667,I3035,I319260,I319693,);
nor I_18626 (I319701,I319693,I319444);
DFFARX1 I_18627 (I319701,I3035,I319260,I319228,);
DFFARX1 I_18628 (I319693,I3035,I319260,I319252,);
not I_18629 (I319746,I319693);
nor I_18630 (I319763,I319746,I319320);
nor I_18631 (I319780,I319585,I319763);
DFFARX1 I_18632 (I319780,I3035,I319260,I319249,);
not I_18633 (I319838,I3042);
DFFARX1 I_18634 (I353330,I3035,I319838,I319864,);
not I_18635 (I319872,I319864);
DFFARX1 I_18636 (I353342,I3035,I319838,I319898,);
not I_18637 (I319906,I353333);
nand I_18638 (I319923,I319906,I353336);
not I_18639 (I319940,I319923);
nor I_18640 (I319957,I319940,I353339);
nor I_18641 (I319974,I319872,I319957);
DFFARX1 I_18642 (I319974,I3035,I319838,I319824,);
not I_18643 (I320005,I353339);
nand I_18644 (I320022,I320005,I319940);
and I_18645 (I320039,I320005,I353333);
nand I_18646 (I320056,I320039,I353345);
nor I_18647 (I319821,I320056,I320005);
and I_18648 (I319812,I319898,I320056);
not I_18649 (I320101,I320056);
nand I_18650 (I319815,I319898,I320101);
nor I_18651 (I319809,I319864,I320056);
not I_18652 (I320146,I353351);
nor I_18653 (I320163,I320146,I353333);
nand I_18654 (I320180,I320163,I320005);
nor I_18655 (I319818,I319923,I320180);
nor I_18656 (I320211,I320146,I353330);
and I_18657 (I320228,I320211,I353348);
or I_18658 (I320245,I320228,I353354);
DFFARX1 I_18659 (I320245,I3035,I319838,I320271,);
nor I_18660 (I320279,I320271,I320022);
DFFARX1 I_18661 (I320279,I3035,I319838,I319806,);
DFFARX1 I_18662 (I320271,I3035,I319838,I319830,);
not I_18663 (I320324,I320271);
nor I_18664 (I320341,I320324,I319898);
nor I_18665 (I320358,I320163,I320341);
DFFARX1 I_18666 (I320358,I3035,I319838,I319827,);
not I_18667 (I320416,I3042);
DFFARX1 I_18668 (I244593,I3035,I320416,I320442,);
not I_18669 (I320450,I320442);
DFFARX1 I_18670 (I244605,I3035,I320416,I320476,);
not I_18671 (I320484,I244581);
nand I_18672 (I320501,I320484,I244608);
not I_18673 (I320518,I320501);
nor I_18674 (I320535,I320518,I244596);
nor I_18675 (I320552,I320450,I320535);
DFFARX1 I_18676 (I320552,I3035,I320416,I320402,);
not I_18677 (I320583,I244596);
nand I_18678 (I320600,I320583,I320518);
and I_18679 (I320617,I320583,I244581);
nand I_18680 (I320634,I320617,I244584);
nor I_18681 (I320399,I320634,I320583);
and I_18682 (I320390,I320476,I320634);
not I_18683 (I320679,I320634);
nand I_18684 (I320393,I320476,I320679);
nor I_18685 (I320387,I320442,I320634);
not I_18686 (I320724,I244590);
nor I_18687 (I320741,I320724,I244581);
nand I_18688 (I320758,I320741,I320583);
nor I_18689 (I320396,I320501,I320758);
nor I_18690 (I320789,I320724,I244599);
and I_18691 (I320806,I320789,I244587);
or I_18692 (I320823,I320806,I244602);
DFFARX1 I_18693 (I320823,I3035,I320416,I320849,);
nor I_18694 (I320857,I320849,I320600);
DFFARX1 I_18695 (I320857,I3035,I320416,I320384,);
DFFARX1 I_18696 (I320849,I3035,I320416,I320408,);
not I_18697 (I320902,I320849);
nor I_18698 (I320919,I320902,I320476);
nor I_18699 (I320936,I320741,I320919);
DFFARX1 I_18700 (I320936,I3035,I320416,I320405,);
not I_18701 (I320994,I3042);
DFFARX1 I_18702 (I339458,I3035,I320994,I321020,);
not I_18703 (I321028,I321020);
DFFARX1 I_18704 (I339470,I3035,I320994,I321054,);
not I_18705 (I321062,I339461);
nand I_18706 (I321079,I321062,I339464);
not I_18707 (I321096,I321079);
nor I_18708 (I321113,I321096,I339467);
nor I_18709 (I321130,I321028,I321113);
DFFARX1 I_18710 (I321130,I3035,I320994,I320980,);
not I_18711 (I321161,I339467);
nand I_18712 (I321178,I321161,I321096);
and I_18713 (I321195,I321161,I339461);
nand I_18714 (I321212,I321195,I339473);
nor I_18715 (I320977,I321212,I321161);
and I_18716 (I320968,I321054,I321212);
not I_18717 (I321257,I321212);
nand I_18718 (I320971,I321054,I321257);
nor I_18719 (I320965,I321020,I321212);
not I_18720 (I321302,I339479);
nor I_18721 (I321319,I321302,I339461);
nand I_18722 (I321336,I321319,I321161);
nor I_18723 (I320974,I321079,I321336);
nor I_18724 (I321367,I321302,I339458);
and I_18725 (I321384,I321367,I339476);
or I_18726 (I321401,I321384,I339482);
DFFARX1 I_18727 (I321401,I3035,I320994,I321427,);
nor I_18728 (I321435,I321427,I321178);
DFFARX1 I_18729 (I321435,I3035,I320994,I320962,);
DFFARX1 I_18730 (I321427,I3035,I320994,I320986,);
not I_18731 (I321480,I321427);
nor I_18732 (I321497,I321480,I321054);
nor I_18733 (I321514,I321319,I321497);
DFFARX1 I_18734 (I321514,I3035,I320994,I320983,);
not I_18735 (I321572,I3042);
DFFARX1 I_18736 (I257649,I3035,I321572,I321598,);
not I_18737 (I321606,I321598);
DFFARX1 I_18738 (I257661,I3035,I321572,I321632,);
not I_18739 (I321640,I257637);
nand I_18740 (I321657,I321640,I257664);
not I_18741 (I321674,I321657);
nor I_18742 (I321691,I321674,I257652);
nor I_18743 (I321708,I321606,I321691);
DFFARX1 I_18744 (I321708,I3035,I321572,I321558,);
not I_18745 (I321739,I257652);
nand I_18746 (I321756,I321739,I321674);
and I_18747 (I321773,I321739,I257637);
nand I_18748 (I321790,I321773,I257640);
nor I_18749 (I321555,I321790,I321739);
and I_18750 (I321546,I321632,I321790);
not I_18751 (I321835,I321790);
nand I_18752 (I321549,I321632,I321835);
nor I_18753 (I321543,I321598,I321790);
not I_18754 (I321880,I257646);
nor I_18755 (I321897,I321880,I257637);
nand I_18756 (I321914,I321897,I321739);
nor I_18757 (I321552,I321657,I321914);
nor I_18758 (I321945,I321880,I257655);
and I_18759 (I321962,I321945,I257643);
or I_18760 (I321979,I321962,I257658);
DFFARX1 I_18761 (I321979,I3035,I321572,I322005,);
nor I_18762 (I322013,I322005,I321756);
DFFARX1 I_18763 (I322013,I3035,I321572,I321540,);
DFFARX1 I_18764 (I322005,I3035,I321572,I321564,);
not I_18765 (I322058,I322005);
nor I_18766 (I322075,I322058,I321632);
nor I_18767 (I322092,I321897,I322075);
DFFARX1 I_18768 (I322092,I3035,I321572,I321561,);
not I_18769 (I322150,I3042);
DFFARX1 I_18770 (I582116,I3035,I322150,I322176,);
not I_18771 (I322184,I322176);
DFFARX1 I_18772 (I582122,I3035,I322150,I322210,);
not I_18773 (I322218,I582116);
nand I_18774 (I322235,I322218,I582119);
not I_18775 (I322252,I322235);
nor I_18776 (I322269,I322252,I582137);
nor I_18777 (I322286,I322184,I322269);
DFFARX1 I_18778 (I322286,I3035,I322150,I322136,);
not I_18779 (I322317,I582137);
nand I_18780 (I322334,I322317,I322252);
and I_18781 (I322351,I322317,I582140);
nand I_18782 (I322368,I322351,I582119);
nor I_18783 (I322133,I322368,I322317);
and I_18784 (I322124,I322210,I322368);
not I_18785 (I322413,I322368);
nand I_18786 (I322127,I322210,I322413);
nor I_18787 (I322121,I322176,I322368);
not I_18788 (I322458,I582125);
nor I_18789 (I322475,I322458,I582140);
nand I_18790 (I322492,I322475,I322317);
nor I_18791 (I322130,I322235,I322492);
nor I_18792 (I322523,I322458,I582131);
and I_18793 (I322540,I322523,I582128);
or I_18794 (I322557,I322540,I582134);
DFFARX1 I_18795 (I322557,I3035,I322150,I322583,);
nor I_18796 (I322591,I322583,I322334);
DFFARX1 I_18797 (I322591,I3035,I322150,I322118,);
DFFARX1 I_18798 (I322583,I3035,I322150,I322142,);
not I_18799 (I322636,I322583);
nor I_18800 (I322653,I322636,I322210);
nor I_18801 (I322670,I322475,I322653);
DFFARX1 I_18802 (I322670,I3035,I322150,I322139,);
not I_18803 (I322728,I3042);
DFFARX1 I_18804 (I422441,I3035,I322728,I322754,);
not I_18805 (I322762,I322754);
DFFARX1 I_18806 (I422441,I3035,I322728,I322788,);
not I_18807 (I322796,I422438);
nand I_18808 (I322813,I322796,I422453);
not I_18809 (I322830,I322813);
nor I_18810 (I322847,I322830,I422447);
nor I_18811 (I322864,I322762,I322847);
DFFARX1 I_18812 (I322864,I3035,I322728,I322714,);
not I_18813 (I322895,I422447);
nand I_18814 (I322912,I322895,I322830);
and I_18815 (I322929,I322895,I422444);
nand I_18816 (I322946,I322929,I422435);
nor I_18817 (I322711,I322946,I322895);
and I_18818 (I322702,I322788,I322946);
not I_18819 (I322991,I322946);
nand I_18820 (I322705,I322788,I322991);
nor I_18821 (I322699,I322754,I322946);
not I_18822 (I323036,I422456);
nor I_18823 (I323053,I323036,I422444);
nand I_18824 (I323070,I323053,I322895);
nor I_18825 (I322708,I322813,I323070);
nor I_18826 (I323101,I323036,I422435);
and I_18827 (I323118,I323101,I422438);
or I_18828 (I323135,I323118,I422450);
DFFARX1 I_18829 (I323135,I3035,I322728,I323161,);
nor I_18830 (I323169,I323161,I322912);
DFFARX1 I_18831 (I323169,I3035,I322728,I322696,);
DFFARX1 I_18832 (I323161,I3035,I322728,I322720,);
not I_18833 (I323214,I323161);
nor I_18834 (I323231,I323214,I322788);
nor I_18835 (I323248,I323053,I323231);
DFFARX1 I_18836 (I323248,I3035,I322728,I322717,);
not I_18837 (I323306,I3042);
DFFARX1 I_18838 (I435089,I3035,I323306,I323332,);
not I_18839 (I323340,I323332);
DFFARX1 I_18840 (I435089,I3035,I323306,I323366,);
not I_18841 (I323374,I435086);
nand I_18842 (I323391,I323374,I435101);
not I_18843 (I323408,I323391);
nor I_18844 (I323425,I323408,I435095);
nor I_18845 (I323442,I323340,I323425);
DFFARX1 I_18846 (I323442,I3035,I323306,I323292,);
not I_18847 (I323473,I435095);
nand I_18848 (I323490,I323473,I323408);
and I_18849 (I323507,I323473,I435092);
nand I_18850 (I323524,I323507,I435083);
nor I_18851 (I323289,I323524,I323473);
and I_18852 (I323280,I323366,I323524);
not I_18853 (I323569,I323524);
nand I_18854 (I323283,I323366,I323569);
nor I_18855 (I323277,I323332,I323524);
not I_18856 (I323614,I435104);
nor I_18857 (I323631,I323614,I435092);
nand I_18858 (I323648,I323631,I323473);
nor I_18859 (I323286,I323391,I323648);
nor I_18860 (I323679,I323614,I435083);
and I_18861 (I323696,I323679,I435086);
or I_18862 (I323713,I323696,I435098);
DFFARX1 I_18863 (I323713,I3035,I323306,I323739,);
nor I_18864 (I323747,I323739,I323490);
DFFARX1 I_18865 (I323747,I3035,I323306,I323274,);
DFFARX1 I_18866 (I323739,I3035,I323306,I323298,);
not I_18867 (I323792,I323739);
nor I_18868 (I323809,I323792,I323366);
nor I_18869 (I323826,I323631,I323809);
DFFARX1 I_18870 (I323826,I3035,I323306,I323295,);
not I_18871 (I323884,I3042);
DFFARX1 I_18872 (I515482,I3035,I323884,I323910,);
not I_18873 (I323918,I323910);
DFFARX1 I_18874 (I515479,I3035,I323884,I323944,);
not I_18875 (I323952,I515476);
nand I_18876 (I323969,I323952,I515503);
not I_18877 (I323986,I323969);
nor I_18878 (I324003,I323986,I515491);
nor I_18879 (I324020,I323918,I324003);
DFFARX1 I_18880 (I324020,I3035,I323884,I323870,);
not I_18881 (I324051,I515491);
nand I_18882 (I324068,I324051,I323986);
and I_18883 (I324085,I324051,I515497);
nand I_18884 (I324102,I324085,I515488);
nor I_18885 (I323867,I324102,I324051);
and I_18886 (I323858,I323944,I324102);
not I_18887 (I324147,I324102);
nand I_18888 (I323861,I323944,I324147);
nor I_18889 (I323855,I323910,I324102);
not I_18890 (I324192,I515485);
nor I_18891 (I324209,I324192,I515497);
nand I_18892 (I324226,I324209,I324051);
nor I_18893 (I323864,I323969,I324226);
nor I_18894 (I324257,I324192,I515500);
and I_18895 (I324274,I324257,I515494);
or I_18896 (I324291,I324274,I515476);
DFFARX1 I_18897 (I324291,I3035,I323884,I324317,);
nor I_18898 (I324325,I324317,I324068);
DFFARX1 I_18899 (I324325,I3035,I323884,I323852,);
DFFARX1 I_18900 (I324317,I3035,I323884,I323876,);
not I_18901 (I324370,I324317);
nor I_18902 (I324387,I324370,I323944);
nor I_18903 (I324404,I324209,I324387);
DFFARX1 I_18904 (I324404,I3035,I323884,I323873,);
not I_18905 (I324462,I3042);
DFFARX1 I_18906 (I434562,I3035,I324462,I324488,);
not I_18907 (I324496,I324488);
DFFARX1 I_18908 (I434562,I3035,I324462,I324522,);
not I_18909 (I324530,I434559);
nand I_18910 (I324547,I324530,I434574);
not I_18911 (I324564,I324547);
nor I_18912 (I324581,I324564,I434568);
nor I_18913 (I324598,I324496,I324581);
DFFARX1 I_18914 (I324598,I3035,I324462,I324448,);
not I_18915 (I324629,I434568);
nand I_18916 (I324646,I324629,I324564);
and I_18917 (I324663,I324629,I434565);
nand I_18918 (I324680,I324663,I434556);
nor I_18919 (I324445,I324680,I324629);
and I_18920 (I324436,I324522,I324680);
not I_18921 (I324725,I324680);
nand I_18922 (I324439,I324522,I324725);
nor I_18923 (I324433,I324488,I324680);
not I_18924 (I324770,I434577);
nor I_18925 (I324787,I324770,I434565);
nand I_18926 (I324804,I324787,I324629);
nor I_18927 (I324442,I324547,I324804);
nor I_18928 (I324835,I324770,I434556);
and I_18929 (I324852,I324835,I434559);
or I_18930 (I324869,I324852,I434571);
DFFARX1 I_18931 (I324869,I3035,I324462,I324895,);
nor I_18932 (I324903,I324895,I324646);
DFFARX1 I_18933 (I324903,I3035,I324462,I324430,);
DFFARX1 I_18934 (I324895,I3035,I324462,I324454,);
not I_18935 (I324948,I324895);
nor I_18936 (I324965,I324948,I324522);
nor I_18937 (I324982,I324787,I324965);
DFFARX1 I_18938 (I324982,I3035,I324462,I324451,);
not I_18939 (I325040,I3042);
DFFARX1 I_18940 (I349284,I3035,I325040,I325066,);
not I_18941 (I325074,I325066);
DFFARX1 I_18942 (I349296,I3035,I325040,I325100,);
not I_18943 (I325108,I349287);
nand I_18944 (I325125,I325108,I349290);
not I_18945 (I325142,I325125);
nor I_18946 (I325159,I325142,I349293);
nor I_18947 (I325176,I325074,I325159);
DFFARX1 I_18948 (I325176,I3035,I325040,I325026,);
not I_18949 (I325207,I349293);
nand I_18950 (I325224,I325207,I325142);
and I_18951 (I325241,I325207,I349287);
nand I_18952 (I325258,I325241,I349299);
nor I_18953 (I325023,I325258,I325207);
and I_18954 (I325014,I325100,I325258);
not I_18955 (I325303,I325258);
nand I_18956 (I325017,I325100,I325303);
nor I_18957 (I325011,I325066,I325258);
not I_18958 (I325348,I349305);
nor I_18959 (I325365,I325348,I349287);
nand I_18960 (I325382,I325365,I325207);
nor I_18961 (I325020,I325125,I325382);
nor I_18962 (I325413,I325348,I349284);
and I_18963 (I325430,I325413,I349302);
or I_18964 (I325447,I325430,I349308);
DFFARX1 I_18965 (I325447,I3035,I325040,I325473,);
nor I_18966 (I325481,I325473,I325224);
DFFARX1 I_18967 (I325481,I3035,I325040,I325008,);
DFFARX1 I_18968 (I325473,I3035,I325040,I325032,);
not I_18969 (I325526,I325473);
nor I_18970 (I325543,I325526,I325100);
nor I_18971 (I325560,I325365,I325543);
DFFARX1 I_18972 (I325560,I3035,I325040,I325029,);
not I_18973 (I325618,I3042);
DFFARX1 I_18974 (I456169,I3035,I325618,I325644,);
not I_18975 (I325652,I325644);
DFFARX1 I_18976 (I456169,I3035,I325618,I325678,);
not I_18977 (I325686,I456166);
nand I_18978 (I325703,I325686,I456181);
not I_18979 (I325720,I325703);
nor I_18980 (I325737,I325720,I456175);
nor I_18981 (I325754,I325652,I325737);
DFFARX1 I_18982 (I325754,I3035,I325618,I325604,);
not I_18983 (I325785,I456175);
nand I_18984 (I325802,I325785,I325720);
and I_18985 (I325819,I325785,I456172);
nand I_18986 (I325836,I325819,I456163);
nor I_18987 (I325601,I325836,I325785);
and I_18988 (I325592,I325678,I325836);
not I_18989 (I325881,I325836);
nand I_18990 (I325595,I325678,I325881);
nor I_18991 (I325589,I325644,I325836);
not I_18992 (I325926,I456184);
nor I_18993 (I325943,I325926,I456172);
nand I_18994 (I325960,I325943,I325785);
nor I_18995 (I325598,I325703,I325960);
nor I_18996 (I325991,I325926,I456163);
and I_18997 (I326008,I325991,I456166);
or I_18998 (I326025,I326008,I456178);
DFFARX1 I_18999 (I326025,I3035,I325618,I326051,);
nor I_19000 (I326059,I326051,I325802);
DFFARX1 I_19001 (I326059,I3035,I325618,I325586,);
DFFARX1 I_19002 (I326051,I3035,I325618,I325610,);
not I_19003 (I326104,I326051);
nor I_19004 (I326121,I326104,I325678);
nor I_19005 (I326138,I325943,I326121);
DFFARX1 I_19006 (I326138,I3035,I325618,I325607,);
not I_19007 (I326196,I3042);
DFFARX1 I_19008 (I341192,I3035,I326196,I326222,);
not I_19009 (I326230,I326222);
DFFARX1 I_19010 (I341204,I3035,I326196,I326256,);
not I_19011 (I326264,I341195);
nand I_19012 (I326281,I326264,I341198);
not I_19013 (I326298,I326281);
nor I_19014 (I326315,I326298,I341201);
nor I_19015 (I326332,I326230,I326315);
DFFARX1 I_19016 (I326332,I3035,I326196,I326182,);
not I_19017 (I326363,I341201);
nand I_19018 (I326380,I326363,I326298);
and I_19019 (I326397,I326363,I341195);
nand I_19020 (I326414,I326397,I341207);
nor I_19021 (I326179,I326414,I326363);
and I_19022 (I326170,I326256,I326414);
not I_19023 (I326459,I326414);
nand I_19024 (I326173,I326256,I326459);
nor I_19025 (I326167,I326222,I326414);
not I_19026 (I326504,I341213);
nor I_19027 (I326521,I326504,I341195);
nand I_19028 (I326538,I326521,I326363);
nor I_19029 (I326176,I326281,I326538);
nor I_19030 (I326569,I326504,I341192);
and I_19031 (I326586,I326569,I341210);
or I_19032 (I326603,I326586,I341216);
DFFARX1 I_19033 (I326603,I3035,I326196,I326629,);
nor I_19034 (I326637,I326629,I326380);
DFFARX1 I_19035 (I326637,I3035,I326196,I326164,);
DFFARX1 I_19036 (I326629,I3035,I326196,I326188,);
not I_19037 (I326682,I326629);
nor I_19038 (I326699,I326682,I326256);
nor I_19039 (I326716,I326521,I326699);
DFFARX1 I_19040 (I326716,I3035,I326196,I326185,);
not I_19041 (I326774,I3042);
DFFARX1 I_19042 (I1908,I3035,I326774,I326800,);
not I_19043 (I326808,I326800);
DFFARX1 I_19044 (I2612,I3035,I326774,I326834,);
not I_19045 (I326842,I2132);
nand I_19046 (I326859,I326842,I1548);
not I_19047 (I326876,I326859);
nor I_19048 (I326893,I326876,I2716);
nor I_19049 (I326910,I326808,I326893);
DFFARX1 I_19050 (I326910,I3035,I326774,I326760,);
not I_19051 (I326941,I2716);
nand I_19052 (I326958,I326941,I326876);
and I_19053 (I326975,I326941,I2060);
nand I_19054 (I326992,I326975,I2284);
nor I_19055 (I326757,I326992,I326941);
and I_19056 (I326748,I326834,I326992);
not I_19057 (I327037,I326992);
nand I_19058 (I326751,I326834,I327037);
nor I_19059 (I326745,I326800,I326992);
not I_19060 (I327082,I2796);
nor I_19061 (I327099,I327082,I2060);
nand I_19062 (I327116,I327099,I326941);
nor I_19063 (I326754,I326859,I327116);
nor I_19064 (I327147,I327082,I1468);
and I_19065 (I327164,I327147,I1716);
or I_19066 (I327181,I327164,I2124);
DFFARX1 I_19067 (I327181,I3035,I326774,I327207,);
nor I_19068 (I327215,I327207,I326958);
DFFARX1 I_19069 (I327215,I3035,I326774,I326742,);
DFFARX1 I_19070 (I327207,I3035,I326774,I326766,);
not I_19071 (I327260,I327207);
nor I_19072 (I327277,I327260,I326834);
nor I_19073 (I327294,I327099,I327277);
DFFARX1 I_19074 (I327294,I3035,I326774,I326763,);
not I_19075 (I327352,I3042);
DFFARX1 I_19076 (I470925,I3035,I327352,I327378,);
not I_19077 (I327386,I327378);
DFFARX1 I_19078 (I470925,I3035,I327352,I327412,);
not I_19079 (I327420,I470922);
nand I_19080 (I327437,I327420,I470937);
not I_19081 (I327454,I327437);
nor I_19082 (I327471,I327454,I470931);
nor I_19083 (I327488,I327386,I327471);
DFFARX1 I_19084 (I327488,I3035,I327352,I327338,);
not I_19085 (I327519,I470931);
nand I_19086 (I327536,I327519,I327454);
and I_19087 (I327553,I327519,I470928);
nand I_19088 (I327570,I327553,I470919);
nor I_19089 (I327335,I327570,I327519);
and I_19090 (I327326,I327412,I327570);
not I_19091 (I327615,I327570);
nand I_19092 (I327329,I327412,I327615);
nor I_19093 (I327323,I327378,I327570);
not I_19094 (I327660,I470940);
nor I_19095 (I327677,I327660,I470928);
nand I_19096 (I327694,I327677,I327519);
nor I_19097 (I327332,I327437,I327694);
nor I_19098 (I327725,I327660,I470919);
and I_19099 (I327742,I327725,I470922);
or I_19100 (I327759,I327742,I470934);
DFFARX1 I_19101 (I327759,I3035,I327352,I327785,);
nor I_19102 (I327793,I327785,I327536);
DFFARX1 I_19103 (I327793,I3035,I327352,I327320,);
DFFARX1 I_19104 (I327785,I3035,I327352,I327344,);
not I_19105 (I327838,I327785);
nor I_19106 (I327855,I327838,I327412);
nor I_19107 (I327872,I327677,I327855);
DFFARX1 I_19108 (I327872,I3035,I327352,I327341,);
not I_19109 (I327930,I3042);
DFFARX1 I_19110 (I587896,I3035,I327930,I327956,);
not I_19111 (I327964,I327956);
DFFARX1 I_19112 (I587902,I3035,I327930,I327990,);
not I_19113 (I327998,I587896);
nand I_19114 (I328015,I327998,I587899);
not I_19115 (I328032,I328015);
nor I_19116 (I328049,I328032,I587917);
nor I_19117 (I328066,I327964,I328049);
DFFARX1 I_19118 (I328066,I3035,I327930,I327916,);
not I_19119 (I328097,I587917);
nand I_19120 (I328114,I328097,I328032);
and I_19121 (I328131,I328097,I587920);
nand I_19122 (I328148,I328131,I587899);
nor I_19123 (I327913,I328148,I328097);
and I_19124 (I327904,I327990,I328148);
not I_19125 (I328193,I328148);
nand I_19126 (I327907,I327990,I328193);
nor I_19127 (I327901,I327956,I328148);
not I_19128 (I328238,I587905);
nor I_19129 (I328255,I328238,I587920);
nand I_19130 (I328272,I328255,I328097);
nor I_19131 (I327910,I328015,I328272);
nor I_19132 (I328303,I328238,I587911);
and I_19133 (I328320,I328303,I587908);
or I_19134 (I328337,I328320,I587914);
DFFARX1 I_19135 (I328337,I3035,I327930,I328363,);
nor I_19136 (I328371,I328363,I328114);
DFFARX1 I_19137 (I328371,I3035,I327930,I327898,);
DFFARX1 I_19138 (I328363,I3035,I327930,I327922,);
not I_19139 (I328416,I328363);
nor I_19140 (I328433,I328416,I327990);
nor I_19141 (I328450,I328255,I328433);
DFFARX1 I_19142 (I328450,I3035,I327930,I327919,);
not I_19143 (I328508,I3042);
DFFARX1 I_19144 (I359110,I3035,I328508,I328534,);
not I_19145 (I328542,I328534);
DFFARX1 I_19146 (I359122,I3035,I328508,I328568,);
not I_19147 (I328576,I359113);
nand I_19148 (I328593,I328576,I359116);
not I_19149 (I328610,I328593);
nor I_19150 (I328627,I328610,I359119);
nor I_19151 (I328644,I328542,I328627);
DFFARX1 I_19152 (I328644,I3035,I328508,I328494,);
not I_19153 (I328675,I359119);
nand I_19154 (I328692,I328675,I328610);
and I_19155 (I328709,I328675,I359113);
nand I_19156 (I328726,I328709,I359125);
nor I_19157 (I328491,I328726,I328675);
and I_19158 (I328482,I328568,I328726);
not I_19159 (I328771,I328726);
nand I_19160 (I328485,I328568,I328771);
nor I_19161 (I328479,I328534,I328726);
not I_19162 (I328816,I359131);
nor I_19163 (I328833,I328816,I359113);
nand I_19164 (I328850,I328833,I328675);
nor I_19165 (I328488,I328593,I328850);
nor I_19166 (I328881,I328816,I359110);
and I_19167 (I328898,I328881,I359128);
or I_19168 (I328915,I328898,I359134);
DFFARX1 I_19169 (I328915,I3035,I328508,I328941,);
nor I_19170 (I328949,I328941,I328692);
DFFARX1 I_19171 (I328949,I3035,I328508,I328476,);
DFFARX1 I_19172 (I328941,I3035,I328508,I328500,);
not I_19173 (I328994,I328941);
nor I_19174 (I329011,I328994,I328568);
nor I_19175 (I329028,I328833,I329011);
DFFARX1 I_19176 (I329028,I3035,I328508,I328497,);
not I_19177 (I329086,I3042);
DFFARX1 I_19178 (I147934,I3035,I329086,I329112,);
not I_19179 (I329120,I329112);
DFFARX1 I_19180 (I147919,I3035,I329086,I329146,);
not I_19181 (I329154,I147937);
nand I_19182 (I329171,I329154,I147922);
not I_19183 (I329188,I329171);
nor I_19184 (I329205,I329188,I147919);
nor I_19185 (I329222,I329120,I329205);
DFFARX1 I_19186 (I329222,I3035,I329086,I329072,);
not I_19187 (I329253,I147919);
nand I_19188 (I329270,I329253,I329188);
and I_19189 (I329287,I329253,I147922);
nand I_19190 (I329304,I329287,I147943);
nor I_19191 (I329069,I329304,I329253);
and I_19192 (I329060,I329146,I329304);
not I_19193 (I329349,I329304);
nand I_19194 (I329063,I329146,I329349);
nor I_19195 (I329057,I329112,I329304);
not I_19196 (I329394,I147931);
nor I_19197 (I329411,I329394,I147922);
nand I_19198 (I329428,I329411,I329253);
nor I_19199 (I329066,I329171,I329428);
nor I_19200 (I329459,I329394,I147925);
and I_19201 (I329476,I329459,I147940);
or I_19202 (I329493,I329476,I147928);
DFFARX1 I_19203 (I329493,I3035,I329086,I329519,);
nor I_19204 (I329527,I329519,I329270);
DFFARX1 I_19205 (I329527,I3035,I329086,I329054,);
DFFARX1 I_19206 (I329519,I3035,I329086,I329078,);
not I_19207 (I329572,I329519);
nor I_19208 (I329589,I329572,I329146);
nor I_19209 (I329606,I329411,I329589);
DFFARX1 I_19210 (I329606,I3035,I329086,I329075,);
not I_19211 (I329664,I3042);
DFFARX1 I_19212 (I24672,I3035,I329664,I329690,);
not I_19213 (I329698,I329690);
DFFARX1 I_19214 (I24675,I3035,I329664,I329724,);
not I_19215 (I329732,I24669);
nand I_19216 (I329749,I329732,I24693);
not I_19217 (I329766,I329749);
nor I_19218 (I329783,I329766,I24672);
nor I_19219 (I329800,I329698,I329783);
DFFARX1 I_19220 (I329800,I3035,I329664,I329650,);
not I_19221 (I329831,I24672);
nand I_19222 (I329848,I329831,I329766);
and I_19223 (I329865,I329831,I24687);
nand I_19224 (I329882,I329865,I24681);
nor I_19225 (I329647,I329882,I329831);
and I_19226 (I329638,I329724,I329882);
not I_19227 (I329927,I329882);
nand I_19228 (I329641,I329724,I329927);
nor I_19229 (I329635,I329690,I329882);
not I_19230 (I329972,I24690);
nor I_19231 (I329989,I329972,I24687);
nand I_19232 (I330006,I329989,I329831);
nor I_19233 (I329644,I329749,I330006);
nor I_19234 (I330037,I329972,I24669);
and I_19235 (I330054,I330037,I24678);
or I_19236 (I330071,I330054,I24684);
DFFARX1 I_19237 (I330071,I3035,I329664,I330097,);
nor I_19238 (I330105,I330097,I329848);
DFFARX1 I_19239 (I330105,I3035,I329664,I329632,);
DFFARX1 I_19240 (I330097,I3035,I329664,I329656,);
not I_19241 (I330150,I330097);
nor I_19242 (I330167,I330150,I329724);
nor I_19243 (I330184,I329989,I330167);
DFFARX1 I_19244 (I330184,I3035,I329664,I329653,);
not I_19245 (I330242,I3042);
DFFARX1 I_19246 (I680592,I3035,I330242,I330268,);
not I_19247 (I330276,I330268);
DFFARX1 I_19248 (I680604,I3035,I330242,I330302,);
not I_19249 (I330310,I680595);
nand I_19250 (I330327,I330310,I680583);
not I_19251 (I330344,I330327);
nor I_19252 (I330361,I330344,I680580);
nor I_19253 (I330378,I330276,I330361);
DFFARX1 I_19254 (I330378,I3035,I330242,I330228,);
not I_19255 (I330409,I680580);
nand I_19256 (I330426,I330409,I330344);
and I_19257 (I330443,I330409,I680586);
nand I_19258 (I330460,I330443,I680583);
nor I_19259 (I330225,I330460,I330409);
and I_19260 (I330216,I330302,I330460);
not I_19261 (I330505,I330460);
nand I_19262 (I330219,I330302,I330505);
nor I_19263 (I330213,I330268,I330460);
not I_19264 (I330550,I680601);
nor I_19265 (I330567,I330550,I680586);
nand I_19266 (I330584,I330567,I330409);
nor I_19267 (I330222,I330327,I330584);
nor I_19268 (I330615,I330550,I680589);
and I_19269 (I330632,I330615,I680580);
or I_19270 (I330649,I330632,I680598);
DFFARX1 I_19271 (I330649,I3035,I330242,I330675,);
nor I_19272 (I330683,I330675,I330426);
DFFARX1 I_19273 (I330683,I3035,I330242,I330210,);
DFFARX1 I_19274 (I330675,I3035,I330242,I330234,);
not I_19275 (I330728,I330675);
nor I_19276 (I330745,I330728,I330302);
nor I_19277 (I330762,I330567,I330745);
DFFARX1 I_19278 (I330762,I3035,I330242,I330231,);
not I_19279 (I330820,I3042);
DFFARX1 I_19280 (I561652,I3035,I330820,I330846,);
not I_19281 (I330854,I330846);
DFFARX1 I_19282 (I561643,I3035,I330820,I330880,);
not I_19283 (I330888,I561637);
nand I_19284 (I330905,I330888,I561649);
not I_19285 (I330922,I330905);
nor I_19286 (I330939,I330922,I561640);
nor I_19287 (I330956,I330854,I330939);
DFFARX1 I_19288 (I330956,I3035,I330820,I330806,);
not I_19289 (I330987,I561640);
nand I_19290 (I331004,I330987,I330922);
and I_19291 (I331021,I330987,I561646);
nand I_19292 (I331038,I331021,I561631);
nor I_19293 (I330803,I331038,I330987);
and I_19294 (I330794,I330880,I331038);
not I_19295 (I331083,I331038);
nand I_19296 (I330797,I330880,I331083);
nor I_19297 (I330791,I330846,I331038);
not I_19298 (I331128,I561631);
nor I_19299 (I331145,I331128,I561646);
nand I_19300 (I331162,I331145,I330987);
nor I_19301 (I330800,I330905,I331162);
nor I_19302 (I331193,I331128,I561634);
and I_19303 (I331210,I331193,I561637);
or I_19304 (I331227,I331210,I561634);
DFFARX1 I_19305 (I331227,I3035,I330820,I331253,);
nor I_19306 (I331261,I331253,I331004);
DFFARX1 I_19307 (I331261,I3035,I330820,I330788,);
DFFARX1 I_19308 (I331253,I3035,I330820,I330812,);
not I_19309 (I331306,I331253);
nor I_19310 (I331323,I331306,I330880);
nor I_19311 (I331340,I331145,I331323);
DFFARX1 I_19312 (I331340,I3035,I330820,I330809,);
not I_19313 (I331398,I3042);
DFFARX1 I_19314 (I634136,I3035,I331398,I331424,);
not I_19315 (I331432,I331424);
DFFARX1 I_19316 (I634142,I3035,I331398,I331458,);
not I_19317 (I331466,I634136);
nand I_19318 (I331483,I331466,I634139);
not I_19319 (I331500,I331483);
nor I_19320 (I331517,I331500,I634157);
nor I_19321 (I331534,I331432,I331517);
DFFARX1 I_19322 (I331534,I3035,I331398,I331384,);
not I_19323 (I331565,I634157);
nand I_19324 (I331582,I331565,I331500);
and I_19325 (I331599,I331565,I634160);
nand I_19326 (I331616,I331599,I634139);
nor I_19327 (I331381,I331616,I331565);
and I_19328 (I331372,I331458,I331616);
not I_19329 (I331661,I331616);
nand I_19330 (I331375,I331458,I331661);
nor I_19331 (I331369,I331424,I331616);
not I_19332 (I331706,I634145);
nor I_19333 (I331723,I331706,I634160);
nand I_19334 (I331740,I331723,I331565);
nor I_19335 (I331378,I331483,I331740);
nor I_19336 (I331771,I331706,I634151);
and I_19337 (I331788,I331771,I634148);
or I_19338 (I331805,I331788,I634154);
DFFARX1 I_19339 (I331805,I3035,I331398,I331831,);
nor I_19340 (I331839,I331831,I331582);
DFFARX1 I_19341 (I331839,I3035,I331398,I331366,);
DFFARX1 I_19342 (I331831,I3035,I331398,I331390,);
not I_19343 (I331884,I331831);
nor I_19344 (I331901,I331884,I331458);
nor I_19345 (I331918,I331723,I331901);
DFFARX1 I_19346 (I331918,I3035,I331398,I331387,);
not I_19347 (I331976,I3042);
DFFARX1 I_19348 (I254929,I3035,I331976,I332002,);
not I_19349 (I332010,I332002);
DFFARX1 I_19350 (I254941,I3035,I331976,I332036,);
not I_19351 (I332044,I254917);
nand I_19352 (I332061,I332044,I254944);
not I_19353 (I332078,I332061);
nor I_19354 (I332095,I332078,I254932);
nor I_19355 (I332112,I332010,I332095);
DFFARX1 I_19356 (I332112,I3035,I331976,I331962,);
not I_19357 (I332143,I254932);
nand I_19358 (I332160,I332143,I332078);
and I_19359 (I332177,I332143,I254917);
nand I_19360 (I332194,I332177,I254920);
nor I_19361 (I331959,I332194,I332143);
and I_19362 (I331950,I332036,I332194);
not I_19363 (I332239,I332194);
nand I_19364 (I331953,I332036,I332239);
nor I_19365 (I331947,I332002,I332194);
not I_19366 (I332284,I254926);
nor I_19367 (I332301,I332284,I254917);
nand I_19368 (I332318,I332301,I332143);
nor I_19369 (I331956,I332061,I332318);
nor I_19370 (I332349,I332284,I254935);
and I_19371 (I332366,I332349,I254923);
or I_19372 (I332383,I332366,I254938);
DFFARX1 I_19373 (I332383,I3035,I331976,I332409,);
nor I_19374 (I332417,I332409,I332160);
DFFARX1 I_19375 (I332417,I3035,I331976,I331944,);
DFFARX1 I_19376 (I332409,I3035,I331976,I331968,);
not I_19377 (I332462,I332409);
nor I_19378 (I332479,I332462,I332036);
nor I_19379 (I332496,I332301,I332479);
DFFARX1 I_19380 (I332496,I3035,I331976,I331965,);
not I_19381 (I332554,I3042);
DFFARX1 I_19382 (I508376,I3035,I332554,I332580,);
not I_19383 (I332588,I332580);
DFFARX1 I_19384 (I508373,I3035,I332554,I332614,);
not I_19385 (I332622,I508370);
nand I_19386 (I332639,I332622,I508397);
not I_19387 (I332656,I332639);
nor I_19388 (I332673,I332656,I508385);
nor I_19389 (I332690,I332588,I332673);
DFFARX1 I_19390 (I332690,I3035,I332554,I332540,);
not I_19391 (I332721,I508385);
nand I_19392 (I332738,I332721,I332656);
and I_19393 (I332755,I332721,I508391);
nand I_19394 (I332772,I332755,I508382);
nor I_19395 (I332537,I332772,I332721);
and I_19396 (I332528,I332614,I332772);
not I_19397 (I332817,I332772);
nand I_19398 (I332531,I332614,I332817);
nor I_19399 (I332525,I332580,I332772);
not I_19400 (I332862,I508379);
nor I_19401 (I332879,I332862,I508391);
nand I_19402 (I332896,I332879,I332721);
nor I_19403 (I332534,I332639,I332896);
nor I_19404 (I332927,I332862,I508394);
and I_19405 (I332944,I332927,I508388);
or I_19406 (I332961,I332944,I508370);
DFFARX1 I_19407 (I332961,I3035,I332554,I332987,);
nor I_19408 (I332995,I332987,I332738);
DFFARX1 I_19409 (I332995,I3035,I332554,I332522,);
DFFARX1 I_19410 (I332987,I3035,I332554,I332546,);
not I_19411 (I333040,I332987);
nor I_19412 (I333057,I333040,I332614);
nor I_19413 (I333074,I332879,I333057);
DFFARX1 I_19414 (I333074,I3035,I332554,I332543,);
not I_19415 (I333132,I3042);
DFFARX1 I_19416 (I437197,I3035,I333132,I333158,);
not I_19417 (I333166,I333158);
DFFARX1 I_19418 (I437197,I3035,I333132,I333192,);
not I_19419 (I333200,I437194);
nand I_19420 (I333217,I333200,I437209);
not I_19421 (I333234,I333217);
nor I_19422 (I333251,I333234,I437203);
nor I_19423 (I333268,I333166,I333251);
DFFARX1 I_19424 (I333268,I3035,I333132,I333118,);
not I_19425 (I333299,I437203);
nand I_19426 (I333316,I333299,I333234);
and I_19427 (I333333,I333299,I437200);
nand I_19428 (I333350,I333333,I437191);
nor I_19429 (I333115,I333350,I333299);
and I_19430 (I333106,I333192,I333350);
not I_19431 (I333395,I333350);
nand I_19432 (I333109,I333192,I333395);
nor I_19433 (I333103,I333158,I333350);
not I_19434 (I333440,I437212);
nor I_19435 (I333457,I333440,I437200);
nand I_19436 (I333474,I333457,I333299);
nor I_19437 (I333112,I333217,I333474);
nor I_19438 (I333505,I333440,I437191);
and I_19439 (I333522,I333505,I437194);
or I_19440 (I333539,I333522,I437206);
DFFARX1 I_19441 (I333539,I3035,I333132,I333565,);
nor I_19442 (I333573,I333565,I333316);
DFFARX1 I_19443 (I333573,I3035,I333132,I333100,);
DFFARX1 I_19444 (I333565,I3035,I333132,I333124,);
not I_19445 (I333618,I333565);
nor I_19446 (I333635,I333618,I333192);
nor I_19447 (I333652,I333457,I333635);
DFFARX1 I_19448 (I333652,I3035,I333132,I333121,);
not I_19449 (I333710,I3042);
DFFARX1 I_19450 (I466709,I3035,I333710,I333736,);
not I_19451 (I333744,I333736);
DFFARX1 I_19452 (I466709,I3035,I333710,I333770,);
not I_19453 (I333778,I466706);
nand I_19454 (I333795,I333778,I466721);
not I_19455 (I333812,I333795);
nor I_19456 (I333829,I333812,I466715);
nor I_19457 (I333846,I333744,I333829);
DFFARX1 I_19458 (I333846,I3035,I333710,I333696,);
not I_19459 (I333877,I466715);
nand I_19460 (I333894,I333877,I333812);
and I_19461 (I333911,I333877,I466712);
nand I_19462 (I333928,I333911,I466703);
nor I_19463 (I333693,I333928,I333877);
and I_19464 (I333684,I333770,I333928);
not I_19465 (I333973,I333928);
nand I_19466 (I333687,I333770,I333973);
nor I_19467 (I333681,I333736,I333928);
not I_19468 (I334018,I466724);
nor I_19469 (I334035,I334018,I466712);
nand I_19470 (I334052,I334035,I333877);
nor I_19471 (I333690,I333795,I334052);
nor I_19472 (I334083,I334018,I466703);
and I_19473 (I334100,I334083,I466706);
or I_19474 (I334117,I334100,I466718);
DFFARX1 I_19475 (I334117,I3035,I333710,I334143,);
nor I_19476 (I334151,I334143,I333894);
DFFARX1 I_19477 (I334151,I3035,I333710,I333678,);
DFFARX1 I_19478 (I334143,I3035,I333710,I333702,);
not I_19479 (I334196,I334143);
nor I_19480 (I334213,I334196,I333770);
nor I_19481 (I334230,I334035,I334213);
DFFARX1 I_19482 (I334230,I3035,I333710,I333699,);
not I_19483 (I334288,I3042);
DFFARX1 I_19484 (I424549,I3035,I334288,I334314,);
not I_19485 (I334322,I334314);
DFFARX1 I_19486 (I424549,I3035,I334288,I334348,);
not I_19487 (I334356,I424546);
nand I_19488 (I334373,I334356,I424561);
not I_19489 (I334390,I334373);
nor I_19490 (I334407,I334390,I424555);
nor I_19491 (I334424,I334322,I334407);
DFFARX1 I_19492 (I334424,I3035,I334288,I334274,);
not I_19493 (I334455,I424555);
nand I_19494 (I334472,I334455,I334390);
and I_19495 (I334489,I334455,I424552);
nand I_19496 (I334506,I334489,I424543);
nor I_19497 (I334271,I334506,I334455);
and I_19498 (I334262,I334348,I334506);
not I_19499 (I334551,I334506);
nand I_19500 (I334265,I334348,I334551);
nor I_19501 (I334259,I334314,I334506);
not I_19502 (I334596,I424564);
nor I_19503 (I334613,I334596,I424552);
nand I_19504 (I334630,I334613,I334455);
nor I_19505 (I334268,I334373,I334630);
nor I_19506 (I334661,I334596,I424543);
and I_19507 (I334678,I334661,I424546);
or I_19508 (I334695,I334678,I424558);
DFFARX1 I_19509 (I334695,I3035,I334288,I334721,);
nor I_19510 (I334729,I334721,I334472);
DFFARX1 I_19511 (I334729,I3035,I334288,I334256,);
DFFARX1 I_19512 (I334721,I3035,I334288,I334280,);
not I_19513 (I334774,I334721);
nor I_19514 (I334791,I334774,I334348);
nor I_19515 (I334808,I334613,I334791);
DFFARX1 I_19516 (I334808,I3035,I334288,I334277,);
not I_19517 (I334866,I3042);
DFFARX1 I_19518 (I376450,I3035,I334866,I334892,);
not I_19519 (I334900,I334892);
DFFARX1 I_19520 (I376462,I3035,I334866,I334926,);
not I_19521 (I334934,I376453);
nand I_19522 (I334951,I334934,I376456);
not I_19523 (I334968,I334951);
nor I_19524 (I334985,I334968,I376459);
nor I_19525 (I335002,I334900,I334985);
DFFARX1 I_19526 (I335002,I3035,I334866,I334852,);
not I_19527 (I335033,I376459);
nand I_19528 (I335050,I335033,I334968);
and I_19529 (I335067,I335033,I376453);
nand I_19530 (I335084,I335067,I376465);
nor I_19531 (I334849,I335084,I335033);
and I_19532 (I334840,I334926,I335084);
not I_19533 (I335129,I335084);
nand I_19534 (I334843,I334926,I335129);
nor I_19535 (I334837,I334892,I335084);
not I_19536 (I335174,I376471);
nor I_19537 (I335191,I335174,I376453);
nand I_19538 (I335208,I335191,I335033);
nor I_19539 (I334846,I334951,I335208);
nor I_19540 (I335239,I335174,I376450);
and I_19541 (I335256,I335239,I376468);
or I_19542 (I335273,I335256,I376474);
DFFARX1 I_19543 (I335273,I3035,I334866,I335299,);
nor I_19544 (I335307,I335299,I335050);
DFFARX1 I_19545 (I335307,I3035,I334866,I334834,);
DFFARX1 I_19546 (I335299,I3035,I334866,I334858,);
not I_19547 (I335352,I335299);
nor I_19548 (I335369,I335352,I334926);
nor I_19549 (I335386,I335191,I335369);
DFFARX1 I_19550 (I335386,I3035,I334866,I334855,);
not I_19551 (I335444,I3042);
DFFARX1 I_19552 (I42611,I3035,I335444,I335470,);
not I_19553 (I335478,I335470);
DFFARX1 I_19554 (I42590,I3035,I335444,I335504,);
not I_19555 (I335512,I42587);
nand I_19556 (I335529,I335512,I42602);
not I_19557 (I335546,I335529);
nor I_19558 (I335563,I335546,I42590);
nor I_19559 (I335580,I335478,I335563);
DFFARX1 I_19560 (I335580,I3035,I335444,I335430,);
not I_19561 (I335611,I42590);
nand I_19562 (I335628,I335611,I335546);
and I_19563 (I335645,I335611,I42593);
nand I_19564 (I335662,I335645,I42608);
nor I_19565 (I335427,I335662,I335611);
and I_19566 (I335418,I335504,I335662);
not I_19567 (I335707,I335662);
nand I_19568 (I335421,I335504,I335707);
nor I_19569 (I335415,I335470,I335662);
not I_19570 (I335752,I42599);
nor I_19571 (I335769,I335752,I42593);
nand I_19572 (I335786,I335769,I335611);
nor I_19573 (I335424,I335529,I335786);
nor I_19574 (I335817,I335752,I42587);
and I_19575 (I335834,I335817,I42596);
or I_19576 (I335851,I335834,I42605);
DFFARX1 I_19577 (I335851,I3035,I335444,I335877,);
nor I_19578 (I335885,I335877,I335628);
DFFARX1 I_19579 (I335885,I3035,I335444,I335412,);
DFFARX1 I_19580 (I335877,I3035,I335444,I335436,);
not I_19581 (I335930,I335877);
nor I_19582 (I335947,I335930,I335504);
nor I_19583 (I335964,I335769,I335947);
DFFARX1 I_19584 (I335964,I3035,I335444,I335433,);
not I_19585 (I336022,I3042);
DFFARX1 I_19586 (I743633,I3035,I336022,I336048,);
not I_19587 (I336056,I336048);
DFFARX1 I_19588 (I743633,I3035,I336022,I336082,);
not I_19589 (I336090,I743657);
nand I_19590 (I336107,I336090,I743639);
not I_19591 (I336124,I336107);
nor I_19592 (I336141,I336124,I743654);
nor I_19593 (I336158,I336056,I336141);
DFFARX1 I_19594 (I336158,I3035,I336022,I336008,);
not I_19595 (I336189,I743654);
nand I_19596 (I336206,I336189,I336124);
and I_19597 (I336223,I336189,I743636);
nand I_19598 (I336240,I336223,I743645);
nor I_19599 (I336005,I336240,I336189);
and I_19600 (I335996,I336082,I336240);
not I_19601 (I336285,I336240);
nand I_19602 (I335999,I336082,I336285);
nor I_19603 (I335993,I336048,I336240);
not I_19604 (I336330,I743642);
nor I_19605 (I336347,I336330,I743636);
nand I_19606 (I336364,I336347,I336189);
nor I_19607 (I336002,I336107,I336364);
nor I_19608 (I336395,I336330,I743651);
and I_19609 (I336412,I336395,I743660);
or I_19610 (I336429,I336412,I743648);
DFFARX1 I_19611 (I336429,I3035,I336022,I336455,);
nor I_19612 (I336463,I336455,I336206);
DFFARX1 I_19613 (I336463,I3035,I336022,I335990,);
DFFARX1 I_19614 (I336455,I3035,I336022,I336014,);
not I_19615 (I336508,I336455);
nor I_19616 (I336525,I336508,I336082);
nor I_19617 (I336542,I336347,I336525);
DFFARX1 I_19618 (I336542,I3035,I336022,I336011,);
not I_19619 (I336600,I3042);
DFFARX1 I_19620 (I568384,I3035,I336600,I336626,);
not I_19621 (I336634,I336626);
DFFARX1 I_19622 (I568375,I3035,I336600,I336660,);
not I_19623 (I336668,I568369);
nand I_19624 (I336685,I336668,I568381);
not I_19625 (I336702,I336685);
nor I_19626 (I336719,I336702,I568372);
nor I_19627 (I336736,I336634,I336719);
DFFARX1 I_19628 (I336736,I3035,I336600,I336586,);
not I_19629 (I336767,I568372);
nand I_19630 (I336784,I336767,I336702);
and I_19631 (I336801,I336767,I568378);
nand I_19632 (I336818,I336801,I568363);
nor I_19633 (I336583,I336818,I336767);
and I_19634 (I336574,I336660,I336818);
not I_19635 (I336863,I336818);
nand I_19636 (I336577,I336660,I336863);
nor I_19637 (I336571,I336626,I336818);
not I_19638 (I336908,I568363);
nor I_19639 (I336925,I336908,I568378);
nand I_19640 (I336942,I336925,I336767);
nor I_19641 (I336580,I336685,I336942);
nor I_19642 (I336973,I336908,I568366);
and I_19643 (I336990,I336973,I568369);
or I_19644 (I337007,I336990,I568366);
DFFARX1 I_19645 (I337007,I3035,I336600,I337033,);
nor I_19646 (I337041,I337033,I336784);
DFFARX1 I_19647 (I337041,I3035,I336600,I336568,);
DFFARX1 I_19648 (I337033,I3035,I336600,I336592,);
not I_19649 (I337086,I337033);
nor I_19650 (I337103,I337086,I336660);
nor I_19651 (I337120,I336925,I337103);
DFFARX1 I_19652 (I337120,I3035,I336600,I336589,);
not I_19653 (I337178,I3042);
DFFARX1 I_19654 (I635870,I3035,I337178,I337204,);
not I_19655 (I337212,I337204);
DFFARX1 I_19656 (I635876,I3035,I337178,I337238,);
not I_19657 (I337246,I635870);
nand I_19658 (I337263,I337246,I635873);
not I_19659 (I337280,I337263);
nor I_19660 (I337297,I337280,I635891);
nor I_19661 (I337314,I337212,I337297);
DFFARX1 I_19662 (I337314,I3035,I337178,I337164,);
not I_19663 (I337345,I635891);
nand I_19664 (I337362,I337345,I337280);
and I_19665 (I337379,I337345,I635894);
nand I_19666 (I337396,I337379,I635873);
nor I_19667 (I337161,I337396,I337345);
and I_19668 (I337152,I337238,I337396);
not I_19669 (I337441,I337396);
nand I_19670 (I337155,I337238,I337441);
nor I_19671 (I337149,I337204,I337396);
not I_19672 (I337486,I635879);
nor I_19673 (I337503,I337486,I635894);
nand I_19674 (I337520,I337503,I337345);
nor I_19675 (I337158,I337263,I337520);
nor I_19676 (I337551,I337486,I635885);
and I_19677 (I337568,I337551,I635882);
or I_19678 (I337585,I337568,I635888);
DFFARX1 I_19679 (I337585,I3035,I337178,I337611,);
nor I_19680 (I337619,I337611,I337362);
DFFARX1 I_19681 (I337619,I3035,I337178,I337146,);
DFFARX1 I_19682 (I337611,I3035,I337178,I337170,);
not I_19683 (I337664,I337611);
nor I_19684 (I337681,I337664,I337238);
nor I_19685 (I337698,I337503,I337681);
DFFARX1 I_19686 (I337698,I3035,I337178,I337167,);
not I_19687 (I337756,I3042);
DFFARX1 I_19688 (I169277,I3035,I337756,I337782,);
not I_19689 (I337790,I337782);
DFFARX1 I_19690 (I169292,I3035,I337756,I337816,);
not I_19691 (I337824,I169295);
nand I_19692 (I337841,I337824,I169274);
not I_19693 (I337858,I337841);
nor I_19694 (I337875,I337858,I169298);
nor I_19695 (I337892,I337790,I337875);
DFFARX1 I_19696 (I337892,I3035,I337756,I337742,);
not I_19697 (I337923,I169298);
nand I_19698 (I337940,I337923,I337858);
and I_19699 (I337957,I337923,I169280);
nand I_19700 (I337974,I337957,I169271);
nor I_19701 (I337739,I337974,I337923);
and I_19702 (I337730,I337816,I337974);
not I_19703 (I338019,I337974);
nand I_19704 (I337733,I337816,I338019);
nor I_19705 (I337727,I337782,I337974);
not I_19706 (I338064,I169271);
nor I_19707 (I338081,I338064,I169280);
nand I_19708 (I338098,I338081,I337923);
nor I_19709 (I337736,I337841,I338098);
nor I_19710 (I338129,I338064,I169286);
and I_19711 (I338146,I338129,I169289);
or I_19712 (I338163,I338146,I169283);
DFFARX1 I_19713 (I338163,I3035,I337756,I338189,);
nor I_19714 (I338197,I338189,I337940);
DFFARX1 I_19715 (I338197,I3035,I337756,I337724,);
DFFARX1 I_19716 (I338189,I3035,I337756,I337748,);
not I_19717 (I338242,I338189);
nor I_19718 (I338259,I338242,I337816);
nor I_19719 (I338276,I338081,I338259);
DFFARX1 I_19720 (I338276,I3035,I337756,I337745,);
not I_19721 (I338334,I3042);
DFFARX1 I_19722 (I563881,I3035,I338334,I338360,);
not I_19723 (I338368,I338360);
nand I_19724 (I338385,I563878,I563896);
and I_19725 (I338402,I338385,I563893);
DFFARX1 I_19726 (I338402,I3035,I338334,I338428,);
not I_19727 (I338436,I563875);
DFFARX1 I_19728 (I563878,I3035,I338334,I338462,);
not I_19729 (I338470,I338462);
nor I_19730 (I338487,I338470,I338368);
and I_19731 (I338504,I338487,I563875);
nor I_19732 (I338521,I338470,I338436);
nor I_19733 (I338317,I338428,I338521);
DFFARX1 I_19734 (I563887,I3035,I338334,I338561,);
nor I_19735 (I338569,I338561,I338428);
not I_19736 (I338586,I338569);
not I_19737 (I338603,I338561);
nor I_19738 (I338620,I338603,I338504);
DFFARX1 I_19739 (I338620,I3035,I338334,I338320,);
nand I_19740 (I338651,I563890,I563875);
and I_19741 (I338668,I338651,I563881);
DFFARX1 I_19742 (I338668,I3035,I338334,I338694,);
nor I_19743 (I338702,I338694,I338561);
DFFARX1 I_19744 (I338702,I3035,I338334,I338302,);
nand I_19745 (I338733,I338694,I338603);
nand I_19746 (I338311,I338586,I338733);
not I_19747 (I338764,I338694);
nor I_19748 (I338781,I338764,I338504);
DFFARX1 I_19749 (I338781,I3035,I338334,I338323,);
nor I_19750 (I338812,I563884,I563875);
or I_19751 (I338314,I338561,I338812);
nor I_19752 (I338305,I338694,I338812);
or I_19753 (I338308,I338428,I338812);
DFFARX1 I_19754 (I338812,I3035,I338334,I338326,);
not I_19755 (I338912,I3042);
DFFARX1 I_19756 (I25735,I3035,I338912,I338938,);
not I_19757 (I338946,I338938);
nand I_19758 (I338963,I25732,I25723);
and I_19759 (I338980,I338963,I25723);
DFFARX1 I_19760 (I338980,I3035,I338912,I339006,);
not I_19761 (I339014,I25726);
DFFARX1 I_19762 (I25741,I3035,I338912,I339040,);
not I_19763 (I339048,I339040);
nor I_19764 (I339065,I339048,I338946);
and I_19765 (I339082,I339065,I25726);
nor I_19766 (I339099,I339048,I339014);
nor I_19767 (I338895,I339006,I339099);
DFFARX1 I_19768 (I25726,I3035,I338912,I339139,);
nor I_19769 (I339147,I339139,I339006);
not I_19770 (I339164,I339147);
not I_19771 (I339181,I339139);
nor I_19772 (I339198,I339181,I339082);
DFFARX1 I_19773 (I339198,I3035,I338912,I338898,);
nand I_19774 (I339229,I25744,I25729);
and I_19775 (I339246,I339229,I25747);
DFFARX1 I_19776 (I339246,I3035,I338912,I339272,);
nor I_19777 (I339280,I339272,I339139);
DFFARX1 I_19778 (I339280,I3035,I338912,I338880,);
nand I_19779 (I339311,I339272,I339181);
nand I_19780 (I338889,I339164,I339311);
not I_19781 (I339342,I339272);
nor I_19782 (I339359,I339342,I339082);
DFFARX1 I_19783 (I339359,I3035,I338912,I338901,);
nor I_19784 (I339390,I25738,I25729);
or I_19785 (I338892,I339139,I339390);
nor I_19786 (I338883,I339272,I339390);
or I_19787 (I338886,I339006,I339390);
DFFARX1 I_19788 (I339390,I3035,I338912,I338904,);
not I_19789 (I339490,I3042);
DFFARX1 I_19790 (I575198,I3035,I339490,I339516,);
not I_19791 (I339524,I339516);
nand I_19792 (I339541,I575180,I575192);
and I_19793 (I339558,I339541,I575195);
DFFARX1 I_19794 (I339558,I3035,I339490,I339584,);
not I_19795 (I339592,I575189);
DFFARX1 I_19796 (I575186,I3035,I339490,I339618,);
not I_19797 (I339626,I339618);
nor I_19798 (I339643,I339626,I339524);
and I_19799 (I339660,I339643,I575189);
nor I_19800 (I339677,I339626,I339592);
nor I_19801 (I339473,I339584,I339677);
DFFARX1 I_19802 (I575204,I3035,I339490,I339717,);
nor I_19803 (I339725,I339717,I339584);
not I_19804 (I339742,I339725);
not I_19805 (I339759,I339717);
nor I_19806 (I339776,I339759,I339660);
DFFARX1 I_19807 (I339776,I3035,I339490,I339476,);
nand I_19808 (I339807,I575183,I575183);
and I_19809 (I339824,I339807,I575180);
DFFARX1 I_19810 (I339824,I3035,I339490,I339850,);
nor I_19811 (I339858,I339850,I339717);
DFFARX1 I_19812 (I339858,I3035,I339490,I339458,);
nand I_19813 (I339889,I339850,I339759);
nand I_19814 (I339467,I339742,I339889);
not I_19815 (I339920,I339850);
nor I_19816 (I339937,I339920,I339660);
DFFARX1 I_19817 (I339937,I3035,I339490,I339479,);
nor I_19818 (I339968,I575201,I575183);
or I_19819 (I339470,I339717,I339968);
nor I_19820 (I339461,I339850,I339968);
or I_19821 (I339464,I339584,I339968);
DFFARX1 I_19822 (I339968,I3035,I339490,I339482,);
not I_19823 (I340068,I3042);
DFFARX1 I_19824 (I685782,I3035,I340068,I340094,);
not I_19825 (I340102,I340094);
nand I_19826 (I340119,I685806,I685788);
and I_19827 (I340136,I340119,I685794);
DFFARX1 I_19828 (I340136,I3035,I340068,I340162,);
not I_19829 (I340170,I685800);
DFFARX1 I_19830 (I685785,I3035,I340068,I340196,);
not I_19831 (I340204,I340196);
nor I_19832 (I340221,I340204,I340102);
and I_19833 (I340238,I340221,I685800);
nor I_19834 (I340255,I340204,I340170);
nor I_19835 (I340051,I340162,I340255);
DFFARX1 I_19836 (I685797,I3035,I340068,I340295,);
nor I_19837 (I340303,I340295,I340162);
not I_19838 (I340320,I340303);
not I_19839 (I340337,I340295);
nor I_19840 (I340354,I340337,I340238);
DFFARX1 I_19841 (I340354,I3035,I340068,I340054,);
nand I_19842 (I340385,I685803,I685791);
and I_19843 (I340402,I340385,I685785);
DFFARX1 I_19844 (I340402,I3035,I340068,I340428,);
nor I_19845 (I340436,I340428,I340295);
DFFARX1 I_19846 (I340436,I3035,I340068,I340036,);
nand I_19847 (I340467,I340428,I340337);
nand I_19848 (I340045,I340320,I340467);
not I_19849 (I340498,I340428);
nor I_19850 (I340515,I340498,I340238);
DFFARX1 I_19851 (I340515,I3035,I340068,I340057,);
nor I_19852 (I340546,I685782,I685791);
or I_19853 (I340048,I340295,I340546);
nor I_19854 (I340039,I340428,I340546);
or I_19855 (I340042,I340162,I340546);
DFFARX1 I_19856 (I340546,I3035,I340068,I340060,);
not I_19857 (I340646,I3042);
DFFARX1 I_19858 (I39428,I3035,I340646,I340672,);
not I_19859 (I340680,I340672);
nand I_19860 (I340697,I39437,I39446);
and I_19861 (I340714,I340697,I39425);
DFFARX1 I_19862 (I340714,I3035,I340646,I340740,);
not I_19863 (I340748,I39428);
DFFARX1 I_19864 (I39443,I3035,I340646,I340774,);
not I_19865 (I340782,I340774);
nor I_19866 (I340799,I340782,I340680);
and I_19867 (I340816,I340799,I39428);
nor I_19868 (I340833,I340782,I340748);
nor I_19869 (I340629,I340740,I340833);
DFFARX1 I_19870 (I39434,I3035,I340646,I340873,);
nor I_19871 (I340881,I340873,I340740);
not I_19872 (I340898,I340881);
not I_19873 (I340915,I340873);
nor I_19874 (I340932,I340915,I340816);
DFFARX1 I_19875 (I340932,I3035,I340646,I340632,);
nand I_19876 (I340963,I39449,I39425);
and I_19877 (I340980,I340963,I39431);
DFFARX1 I_19878 (I340980,I3035,I340646,I341006,);
nor I_19879 (I341014,I341006,I340873);
DFFARX1 I_19880 (I341014,I3035,I340646,I340614,);
nand I_19881 (I341045,I341006,I340915);
nand I_19882 (I340623,I340898,I341045);
not I_19883 (I341076,I341006);
nor I_19884 (I341093,I341076,I340816);
DFFARX1 I_19885 (I341093,I3035,I340646,I340635,);
nor I_19886 (I341124,I39440,I39425);
or I_19887 (I340626,I340873,I341124);
nor I_19888 (I340617,I341006,I341124);
or I_19889 (I340620,I340740,I341124);
DFFARX1 I_19890 (I341124,I3035,I340646,I340638,);
not I_19891 (I341224,I3042);
DFFARX1 I_19892 (I237518,I3035,I341224,I341250,);
not I_19893 (I341258,I341250);
nand I_19894 (I341275,I237509,I237527);
and I_19895 (I341292,I341275,I237530);
DFFARX1 I_19896 (I341292,I3035,I341224,I341318,);
not I_19897 (I341326,I237524);
DFFARX1 I_19898 (I237512,I3035,I341224,I341352,);
not I_19899 (I341360,I341352);
nor I_19900 (I341377,I341360,I341258);
and I_19901 (I341394,I341377,I237524);
nor I_19902 (I341411,I341360,I341326);
nor I_19903 (I341207,I341318,I341411);
DFFARX1 I_19904 (I237521,I3035,I341224,I341451,);
nor I_19905 (I341459,I341451,I341318);
not I_19906 (I341476,I341459);
not I_19907 (I341493,I341451);
nor I_19908 (I341510,I341493,I341394);
DFFARX1 I_19909 (I341510,I3035,I341224,I341210,);
nand I_19910 (I341541,I237536,I237533);
and I_19911 (I341558,I341541,I237515);
DFFARX1 I_19912 (I341558,I3035,I341224,I341584,);
nor I_19913 (I341592,I341584,I341451);
DFFARX1 I_19914 (I341592,I3035,I341224,I341192,);
nand I_19915 (I341623,I341584,I341493);
nand I_19916 (I341201,I341476,I341623);
not I_19917 (I341654,I341584);
nor I_19918 (I341671,I341654,I341394);
DFFARX1 I_19919 (I341671,I3035,I341224,I341213,);
nor I_19920 (I341702,I237509,I237533);
or I_19921 (I341204,I341451,I341702);
nor I_19922 (I341195,I341584,I341702);
or I_19923 (I341198,I341318,I341702);
DFFARX1 I_19924 (I341702,I3035,I341224,I341216,);
not I_19925 (I341802,I3042);
DFFARX1 I_19926 (I218833,I3035,I341802,I341828,);
not I_19927 (I341836,I341828);
nand I_19928 (I341853,I218836,I218812);
and I_19929 (I341870,I341853,I218809);
DFFARX1 I_19930 (I341870,I3035,I341802,I341896,);
not I_19931 (I341904,I218815);
DFFARX1 I_19932 (I218809,I3035,I341802,I341930,);
not I_19933 (I341938,I341930);
nor I_19934 (I341955,I341938,I341836);
and I_19935 (I341972,I341955,I218815);
nor I_19936 (I341989,I341938,I341904);
nor I_19937 (I341785,I341896,I341989);
DFFARX1 I_19938 (I218818,I3035,I341802,I342029,);
nor I_19939 (I342037,I342029,I341896);
not I_19940 (I342054,I342037);
not I_19941 (I342071,I342029);
nor I_19942 (I342088,I342071,I341972);
DFFARX1 I_19943 (I342088,I3035,I341802,I341788,);
nand I_19944 (I342119,I218821,I218830);
and I_19945 (I342136,I342119,I218827);
DFFARX1 I_19946 (I342136,I3035,I341802,I342162,);
nor I_19947 (I342170,I342162,I342029);
DFFARX1 I_19948 (I342170,I3035,I341802,I341770,);
nand I_19949 (I342201,I342162,I342071);
nand I_19950 (I341779,I342054,I342201);
not I_19951 (I342232,I342162);
nor I_19952 (I342249,I342232,I341972);
DFFARX1 I_19953 (I342249,I3035,I341802,I341791,);
nor I_19954 (I342280,I218824,I218830);
or I_19955 (I341782,I342029,I342280);
nor I_19956 (I341773,I342162,I342280);
or I_19957 (I341776,I341896,I342280);
DFFARX1 I_19958 (I342280,I3035,I341802,I341794,);
not I_19959 (I342380,I3042);
DFFARX1 I_19960 (I608144,I3035,I342380,I342406,);
not I_19961 (I342414,I342406);
nand I_19962 (I342431,I608126,I608138);
and I_19963 (I342448,I342431,I608141);
DFFARX1 I_19964 (I342448,I3035,I342380,I342474,);
not I_19965 (I342482,I608135);
DFFARX1 I_19966 (I608132,I3035,I342380,I342508,);
not I_19967 (I342516,I342508);
nor I_19968 (I342533,I342516,I342414);
and I_19969 (I342550,I342533,I608135);
nor I_19970 (I342567,I342516,I342482);
nor I_19971 (I342363,I342474,I342567);
DFFARX1 I_19972 (I608150,I3035,I342380,I342607,);
nor I_19973 (I342615,I342607,I342474);
not I_19974 (I342632,I342615);
not I_19975 (I342649,I342607);
nor I_19976 (I342666,I342649,I342550);
DFFARX1 I_19977 (I342666,I3035,I342380,I342366,);
nand I_19978 (I342697,I608129,I608129);
and I_19979 (I342714,I342697,I608126);
DFFARX1 I_19980 (I342714,I3035,I342380,I342740,);
nor I_19981 (I342748,I342740,I342607);
DFFARX1 I_19982 (I342748,I3035,I342380,I342348,);
nand I_19983 (I342779,I342740,I342649);
nand I_19984 (I342357,I342632,I342779);
not I_19985 (I342810,I342740);
nor I_19986 (I342827,I342810,I342550);
DFFARX1 I_19987 (I342827,I3035,I342380,I342369,);
nor I_19988 (I342858,I608147,I608129);
or I_19989 (I342360,I342607,I342858);
nor I_19990 (I342351,I342740,I342858);
or I_19991 (I342354,I342474,I342858);
DFFARX1 I_19992 (I342858,I3035,I342380,I342372,);
not I_19993 (I342958,I3042);
DFFARX1 I_19994 (I606410,I3035,I342958,I342984,);
not I_19995 (I342992,I342984);
nand I_19996 (I343009,I606392,I606404);
and I_19997 (I343026,I343009,I606407);
DFFARX1 I_19998 (I343026,I3035,I342958,I343052,);
not I_19999 (I343060,I606401);
DFFARX1 I_20000 (I606398,I3035,I342958,I343086,);
not I_20001 (I343094,I343086);
nor I_20002 (I343111,I343094,I342992);
and I_20003 (I343128,I343111,I606401);
nor I_20004 (I343145,I343094,I343060);
nor I_20005 (I342941,I343052,I343145);
DFFARX1 I_20006 (I606416,I3035,I342958,I343185,);
nor I_20007 (I343193,I343185,I343052);
not I_20008 (I343210,I343193);
not I_20009 (I343227,I343185);
nor I_20010 (I343244,I343227,I343128);
DFFARX1 I_20011 (I343244,I3035,I342958,I342944,);
nand I_20012 (I343275,I606395,I606395);
and I_20013 (I343292,I343275,I606392);
DFFARX1 I_20014 (I343292,I3035,I342958,I343318,);
nor I_20015 (I343326,I343318,I343185);
DFFARX1 I_20016 (I343326,I3035,I342958,I342926,);
nand I_20017 (I343357,I343318,I343227);
nand I_20018 (I342935,I343210,I343357);
not I_20019 (I343388,I343318);
nor I_20020 (I343405,I343388,I343128);
DFFARX1 I_20021 (I343405,I3035,I342958,I342947,);
nor I_20022 (I343436,I606413,I606395);
or I_20023 (I342938,I343185,I343436);
nor I_20024 (I342929,I343318,I343436);
or I_20025 (I342932,I343052,I343436);
DFFARX1 I_20026 (I343436,I3035,I342958,I342950,);
not I_20027 (I343536,I3042);
DFFARX1 I_20028 (I436679,I3035,I343536,I343562,);
not I_20029 (I343570,I343562);
nand I_20030 (I343587,I436667,I436685);
and I_20031 (I343604,I343587,I436682);
DFFARX1 I_20032 (I343604,I3035,I343536,I343630,);
not I_20033 (I343638,I436673);
DFFARX1 I_20034 (I436670,I3035,I343536,I343664,);
not I_20035 (I343672,I343664);
nor I_20036 (I343689,I343672,I343570);
and I_20037 (I343706,I343689,I436673);
nor I_20038 (I343723,I343672,I343638);
nor I_20039 (I343519,I343630,I343723);
DFFARX1 I_20040 (I436664,I3035,I343536,I343763,);
nor I_20041 (I343771,I343763,I343630);
not I_20042 (I343788,I343771);
not I_20043 (I343805,I343763);
nor I_20044 (I343822,I343805,I343706);
DFFARX1 I_20045 (I343822,I3035,I343536,I343522,);
nand I_20046 (I343853,I436664,I436667);
and I_20047 (I343870,I343853,I436670);
DFFARX1 I_20048 (I343870,I3035,I343536,I343896,);
nor I_20049 (I343904,I343896,I343763);
DFFARX1 I_20050 (I343904,I3035,I343536,I343504,);
nand I_20051 (I343935,I343896,I343805);
nand I_20052 (I343513,I343788,I343935);
not I_20053 (I343966,I343896);
nor I_20054 (I343983,I343966,I343706);
DFFARX1 I_20055 (I343983,I3035,I343536,I343525,);
nor I_20056 (I344014,I436676,I436667);
or I_20057 (I343516,I343763,I344014);
nor I_20058 (I343507,I343896,I344014);
or I_20059 (I343510,I343630,I344014);
DFFARX1 I_20060 (I344014,I3035,I343536,I343528,);
not I_20061 (I344114,I3042);
DFFARX1 I_20062 (I270158,I3035,I344114,I344140,);
not I_20063 (I344148,I344140);
nand I_20064 (I344165,I270149,I270167);
and I_20065 (I344182,I344165,I270170);
DFFARX1 I_20066 (I344182,I3035,I344114,I344208,);
not I_20067 (I344216,I270164);
DFFARX1 I_20068 (I270152,I3035,I344114,I344242,);
not I_20069 (I344250,I344242);
nor I_20070 (I344267,I344250,I344148);
and I_20071 (I344284,I344267,I270164);
nor I_20072 (I344301,I344250,I344216);
nor I_20073 (I344097,I344208,I344301);
DFFARX1 I_20074 (I270161,I3035,I344114,I344341,);
nor I_20075 (I344349,I344341,I344208);
not I_20076 (I344366,I344349);
not I_20077 (I344383,I344341);
nor I_20078 (I344400,I344383,I344284);
DFFARX1 I_20079 (I344400,I3035,I344114,I344100,);
nand I_20080 (I344431,I270176,I270173);
and I_20081 (I344448,I344431,I270155);
DFFARX1 I_20082 (I344448,I3035,I344114,I344474,);
nor I_20083 (I344482,I344474,I344341);
DFFARX1 I_20084 (I344482,I3035,I344114,I344082,);
nand I_20085 (I344513,I344474,I344383);
nand I_20086 (I344091,I344366,I344513);
not I_20087 (I344544,I344474);
nor I_20088 (I344561,I344544,I344284);
DFFARX1 I_20089 (I344561,I3035,I344114,I344103,);
nor I_20090 (I344592,I270149,I270173);
or I_20091 (I344094,I344341,I344592);
nor I_20092 (I344085,I344474,I344592);
or I_20093 (I344088,I344208,I344592);
DFFARX1 I_20094 (I344592,I3035,I344114,I344106,);
not I_20095 (I344692,I3042);
DFFARX1 I_20096 (I236974,I3035,I344692,I344718,);
not I_20097 (I344726,I344718);
nand I_20098 (I344743,I236965,I236983);
and I_20099 (I344760,I344743,I236986);
DFFARX1 I_20100 (I344760,I3035,I344692,I344786,);
not I_20101 (I344794,I236980);
DFFARX1 I_20102 (I236968,I3035,I344692,I344820,);
not I_20103 (I344828,I344820);
nor I_20104 (I344845,I344828,I344726);
and I_20105 (I344862,I344845,I236980);
nor I_20106 (I344879,I344828,I344794);
nor I_20107 (I344675,I344786,I344879);
DFFARX1 I_20108 (I236977,I3035,I344692,I344919,);
nor I_20109 (I344927,I344919,I344786);
not I_20110 (I344944,I344927);
not I_20111 (I344961,I344919);
nor I_20112 (I344978,I344961,I344862);
DFFARX1 I_20113 (I344978,I3035,I344692,I344678,);
nand I_20114 (I345009,I236992,I236989);
and I_20115 (I345026,I345009,I236971);
DFFARX1 I_20116 (I345026,I3035,I344692,I345052,);
nor I_20117 (I345060,I345052,I344919);
DFFARX1 I_20118 (I345060,I3035,I344692,I344660,);
nand I_20119 (I345091,I345052,I344961);
nand I_20120 (I344669,I344944,I345091);
not I_20121 (I345122,I345052);
nor I_20122 (I345139,I345122,I344862);
DFFARX1 I_20123 (I345139,I3035,I344692,I344681,);
nor I_20124 (I345170,I236965,I236989);
or I_20125 (I344672,I344919,I345170);
nor I_20126 (I344663,I345052,I345170);
or I_20127 (I344666,I344786,I345170);
DFFARX1 I_20128 (I345170,I3035,I344692,I344684,);
not I_20129 (I345270,I3042);
DFFARX1 I_20130 (I655046,I3035,I345270,I345296,);
not I_20131 (I345304,I345296);
nand I_20132 (I345321,I655049,I655058);
and I_20133 (I345338,I345321,I655061);
DFFARX1 I_20134 (I345338,I3035,I345270,I345364,);
not I_20135 (I345372,I655070);
DFFARX1 I_20136 (I655052,I3035,I345270,I345398,);
not I_20137 (I345406,I345398);
nor I_20138 (I345423,I345406,I345304);
and I_20139 (I345440,I345423,I655070);
nor I_20140 (I345457,I345406,I345372);
nor I_20141 (I345253,I345364,I345457);
DFFARX1 I_20142 (I655049,I3035,I345270,I345497,);
nor I_20143 (I345505,I345497,I345364);
not I_20144 (I345522,I345505);
not I_20145 (I345539,I345497);
nor I_20146 (I345556,I345539,I345440);
DFFARX1 I_20147 (I345556,I3035,I345270,I345256,);
nand I_20148 (I345587,I655067,I655046);
and I_20149 (I345604,I345587,I655064);
DFFARX1 I_20150 (I345604,I3035,I345270,I345630,);
nor I_20151 (I345638,I345630,I345497);
DFFARX1 I_20152 (I345638,I3035,I345270,I345238,);
nand I_20153 (I345669,I345630,I345539);
nand I_20154 (I345247,I345522,I345669);
not I_20155 (I345700,I345630);
nor I_20156 (I345717,I345700,I345440);
DFFARX1 I_20157 (I345717,I3035,I345270,I345259,);
nor I_20158 (I345748,I655055,I655046);
or I_20159 (I345250,I345497,I345748);
nor I_20160 (I345241,I345630,I345748);
or I_20161 (I345244,I345364,I345748);
DFFARX1 I_20162 (I345748,I3035,I345270,I345262,);
not I_20163 (I345848,I3042);
DFFARX1 I_20164 (I83659,I3035,I345848,I345874,);
not I_20165 (I345882,I345874);
nand I_20166 (I345899,I83662,I83683);
and I_20167 (I345916,I345899,I83671);
DFFARX1 I_20168 (I345916,I3035,I345848,I345942,);
not I_20169 (I345950,I83668);
DFFARX1 I_20170 (I83659,I3035,I345848,I345976,);
not I_20171 (I345984,I345976);
nor I_20172 (I346001,I345984,I345882);
and I_20173 (I346018,I346001,I83668);
nor I_20174 (I346035,I345984,I345950);
nor I_20175 (I345831,I345942,I346035);
DFFARX1 I_20176 (I83677,I3035,I345848,I346075,);
nor I_20177 (I346083,I346075,I345942);
not I_20178 (I346100,I346083);
not I_20179 (I346117,I346075);
nor I_20180 (I346134,I346117,I346018);
DFFARX1 I_20181 (I346134,I3035,I345848,I345834,);
nand I_20182 (I346165,I83662,I83665);
and I_20183 (I346182,I346165,I83674);
DFFARX1 I_20184 (I346182,I3035,I345848,I346208,);
nor I_20185 (I346216,I346208,I346075);
DFFARX1 I_20186 (I346216,I3035,I345848,I345816,);
nand I_20187 (I346247,I346208,I346117);
nand I_20188 (I345825,I346100,I346247);
not I_20189 (I346278,I346208);
nor I_20190 (I346295,I346278,I346018);
DFFARX1 I_20191 (I346295,I3035,I345848,I345837,);
nor I_20192 (I346326,I83680,I83665);
or I_20193 (I345828,I346075,I346326);
nor I_20194 (I345819,I346208,I346326);
or I_20195 (I345822,I345942,I346326);
DFFARX1 I_20196 (I346326,I3035,I345848,I345840,);
not I_20197 (I346426,I3042);
DFFARX1 I_20198 (I274510,I3035,I346426,I346452,);
not I_20199 (I346460,I346452);
nand I_20200 (I346477,I274501,I274519);
and I_20201 (I346494,I346477,I274522);
DFFARX1 I_20202 (I346494,I3035,I346426,I346520,);
not I_20203 (I346528,I274516);
DFFARX1 I_20204 (I274504,I3035,I346426,I346554,);
not I_20205 (I346562,I346554);
nor I_20206 (I346579,I346562,I346460);
and I_20207 (I346596,I346579,I274516);
nor I_20208 (I346613,I346562,I346528);
nor I_20209 (I346409,I346520,I346613);
DFFARX1 I_20210 (I274513,I3035,I346426,I346653,);
nor I_20211 (I346661,I346653,I346520);
not I_20212 (I346678,I346661);
not I_20213 (I346695,I346653);
nor I_20214 (I346712,I346695,I346596);
DFFARX1 I_20215 (I346712,I3035,I346426,I346412,);
nand I_20216 (I346743,I274528,I274525);
and I_20217 (I346760,I346743,I274507);
DFFARX1 I_20218 (I346760,I3035,I346426,I346786,);
nor I_20219 (I346794,I346786,I346653);
DFFARX1 I_20220 (I346794,I3035,I346426,I346394,);
nand I_20221 (I346825,I346786,I346695);
nand I_20222 (I346403,I346678,I346825);
not I_20223 (I346856,I346786);
nor I_20224 (I346873,I346856,I346596);
DFFARX1 I_20225 (I346873,I3035,I346426,I346415,);
nor I_20226 (I346904,I274501,I274525);
or I_20227 (I346406,I346653,I346904);
nor I_20228 (I346397,I346786,I346904);
or I_20229 (I346400,I346520,I346904);
DFFARX1 I_20230 (I346904,I3035,I346426,I346418,);
not I_20231 (I347004,I3042);
DFFARX1 I_20232 (I72629,I3035,I347004,I347030,);
not I_20233 (I347038,I347030);
nand I_20234 (I347055,I72638,I72647);
and I_20235 (I347072,I347055,I72626);
DFFARX1 I_20236 (I347072,I3035,I347004,I347098,);
not I_20237 (I347106,I72629);
DFFARX1 I_20238 (I72644,I3035,I347004,I347132,);
not I_20239 (I347140,I347132);
nor I_20240 (I347157,I347140,I347038);
and I_20241 (I347174,I347157,I72629);
nor I_20242 (I347191,I347140,I347106);
nor I_20243 (I346987,I347098,I347191);
DFFARX1 I_20244 (I72635,I3035,I347004,I347231,);
nor I_20245 (I347239,I347231,I347098);
not I_20246 (I347256,I347239);
not I_20247 (I347273,I347231);
nor I_20248 (I347290,I347273,I347174);
DFFARX1 I_20249 (I347290,I3035,I347004,I346990,);
nand I_20250 (I347321,I72650,I72626);
and I_20251 (I347338,I347321,I72632);
DFFARX1 I_20252 (I347338,I3035,I347004,I347364,);
nor I_20253 (I347372,I347364,I347231);
DFFARX1 I_20254 (I347372,I3035,I347004,I346972,);
nand I_20255 (I347403,I347364,I347273);
nand I_20256 (I346981,I347256,I347403);
not I_20257 (I347434,I347364);
nor I_20258 (I347451,I347434,I347174);
DFFARX1 I_20259 (I347451,I3035,I347004,I346993,);
nor I_20260 (I347482,I72641,I72626);
or I_20261 (I346984,I347231,I347482);
nor I_20262 (I346975,I347364,I347482);
or I_20263 (I346978,I347098,I347482);
DFFARX1 I_20264 (I347482,I3035,I347004,I346996,);
not I_20265 (I347582,I3042);
DFFARX1 I_20266 (I311714,I3035,I347582,I347608,);
not I_20267 (I347616,I347608);
nand I_20268 (I347633,I311723,I311732);
and I_20269 (I347650,I347633,I311738);
DFFARX1 I_20270 (I347650,I3035,I347582,I347676,);
not I_20271 (I347684,I311735);
DFFARX1 I_20272 (I311720,I3035,I347582,I347710,);
not I_20273 (I347718,I347710);
nor I_20274 (I347735,I347718,I347616);
and I_20275 (I347752,I347735,I311735);
nor I_20276 (I347769,I347718,I347684);
nor I_20277 (I347565,I347676,I347769);
DFFARX1 I_20278 (I311729,I3035,I347582,I347809,);
nor I_20279 (I347817,I347809,I347676);
not I_20280 (I347834,I347817);
not I_20281 (I347851,I347809);
nor I_20282 (I347868,I347851,I347752);
DFFARX1 I_20283 (I347868,I3035,I347582,I347568,);
nand I_20284 (I347899,I311726,I311717);
and I_20285 (I347916,I347899,I311714);
DFFARX1 I_20286 (I347916,I3035,I347582,I347942,);
nor I_20287 (I347950,I347942,I347809);
DFFARX1 I_20288 (I347950,I3035,I347582,I347550,);
nand I_20289 (I347981,I347942,I347851);
nand I_20290 (I347559,I347834,I347981);
not I_20291 (I348012,I347942);
nor I_20292 (I348029,I348012,I347752);
DFFARX1 I_20293 (I348029,I3035,I347582,I347571,);
nor I_20294 (I348060,I311717,I311717);
or I_20295 (I347562,I347809,I348060);
nor I_20296 (I347553,I347942,I348060);
or I_20297 (I347556,I347676,I348060);
DFFARX1 I_20298 (I348060,I3035,I347582,I347574,);
not I_20299 (I348160,I3042);
DFFARX1 I_20300 (I497412,I3035,I348160,I348186,);
not I_20301 (I348194,I348186);
nand I_20302 (I348211,I497388,I497403);
and I_20303 (I348228,I348211,I497415);
DFFARX1 I_20304 (I348228,I3035,I348160,I348254,);
not I_20305 (I348262,I497400);
DFFARX1 I_20306 (I497391,I3035,I348160,I348288,);
not I_20307 (I348296,I348288);
nor I_20308 (I348313,I348296,I348194);
and I_20309 (I348330,I348313,I497400);
nor I_20310 (I348347,I348296,I348262);
nor I_20311 (I348143,I348254,I348347);
DFFARX1 I_20312 (I497388,I3035,I348160,I348387,);
nor I_20313 (I348395,I348387,I348254);
not I_20314 (I348412,I348395);
not I_20315 (I348429,I348387);
nor I_20316 (I348446,I348429,I348330);
DFFARX1 I_20317 (I348446,I3035,I348160,I348146,);
nand I_20318 (I348477,I497406,I497397);
and I_20319 (I348494,I348477,I497409);
DFFARX1 I_20320 (I348494,I3035,I348160,I348520,);
nor I_20321 (I348528,I348520,I348387);
DFFARX1 I_20322 (I348528,I3035,I348160,I348128,);
nand I_20323 (I348559,I348520,I348429);
nand I_20324 (I348137,I348412,I348559);
not I_20325 (I348590,I348520);
nor I_20326 (I348607,I348590,I348330);
DFFARX1 I_20327 (I348607,I3035,I348160,I348149,);
nor I_20328 (I348638,I497394,I497397);
or I_20329 (I348140,I348387,I348638);
nor I_20330 (I348131,I348520,I348638);
or I_20331 (I348134,I348254,I348638);
DFFARX1 I_20332 (I348638,I3035,I348160,I348152,);
not I_20333 (I348738,I3042);
DFFARX1 I_20334 (I308246,I3035,I348738,I348764,);
not I_20335 (I348772,I348764);
nand I_20336 (I348789,I308255,I308264);
and I_20337 (I348806,I348789,I308270);
DFFARX1 I_20338 (I348806,I3035,I348738,I348832,);
not I_20339 (I348840,I308267);
DFFARX1 I_20340 (I308252,I3035,I348738,I348866,);
not I_20341 (I348874,I348866);
nor I_20342 (I348891,I348874,I348772);
and I_20343 (I348908,I348891,I308267);
nor I_20344 (I348925,I348874,I348840);
nor I_20345 (I348721,I348832,I348925);
DFFARX1 I_20346 (I308261,I3035,I348738,I348965,);
nor I_20347 (I348973,I348965,I348832);
not I_20348 (I348990,I348973);
not I_20349 (I349007,I348965);
nor I_20350 (I349024,I349007,I348908);
DFFARX1 I_20351 (I349024,I3035,I348738,I348724,);
nand I_20352 (I349055,I308258,I308249);
and I_20353 (I349072,I349055,I308246);
DFFARX1 I_20354 (I349072,I3035,I348738,I349098,);
nor I_20355 (I349106,I349098,I348965);
DFFARX1 I_20356 (I349106,I3035,I348738,I348706,);
nand I_20357 (I349137,I349098,I349007);
nand I_20358 (I348715,I348990,I349137);
not I_20359 (I349168,I349098);
nor I_20360 (I349185,I349168,I348908);
DFFARX1 I_20361 (I349185,I3035,I348738,I348727,);
nor I_20362 (I349216,I308249,I308249);
or I_20363 (I348718,I348965,I349216);
nor I_20364 (I348709,I349098,I349216);
or I_20365 (I348712,I348832,I349216);
DFFARX1 I_20366 (I349216,I3035,I348738,I348730,);
not I_20367 (I349316,I3042);
DFFARX1 I_20368 (I325586,I3035,I349316,I349342,);
not I_20369 (I349350,I349342);
nand I_20370 (I349367,I325595,I325604);
and I_20371 (I349384,I349367,I325610);
DFFARX1 I_20372 (I349384,I3035,I349316,I349410,);
not I_20373 (I349418,I325607);
DFFARX1 I_20374 (I325592,I3035,I349316,I349444,);
not I_20375 (I349452,I349444);
nor I_20376 (I349469,I349452,I349350);
and I_20377 (I349486,I349469,I325607);
nor I_20378 (I349503,I349452,I349418);
nor I_20379 (I349299,I349410,I349503);
DFFARX1 I_20380 (I325601,I3035,I349316,I349543,);
nor I_20381 (I349551,I349543,I349410);
not I_20382 (I349568,I349551);
not I_20383 (I349585,I349543);
nor I_20384 (I349602,I349585,I349486);
DFFARX1 I_20385 (I349602,I3035,I349316,I349302,);
nand I_20386 (I349633,I325598,I325589);
and I_20387 (I349650,I349633,I325586);
DFFARX1 I_20388 (I349650,I3035,I349316,I349676,);
nor I_20389 (I349684,I349676,I349543);
DFFARX1 I_20390 (I349684,I3035,I349316,I349284,);
nand I_20391 (I349715,I349676,I349585);
nand I_20392 (I349293,I349568,I349715);
not I_20393 (I349746,I349676);
nor I_20394 (I349763,I349746,I349486);
DFFARX1 I_20395 (I349763,I3035,I349316,I349305,);
nor I_20396 (I349794,I325589,I325589);
or I_20397 (I349296,I349543,I349794);
nor I_20398 (I349287,I349676,I349794);
or I_20399 (I349290,I349410,I349794);
DFFARX1 I_20400 (I349794,I3035,I349316,I349308,);
not I_20401 (I349894,I3042);
DFFARX1 I_20402 (I536172,I3035,I349894,I349920,);
not I_20403 (I349928,I349920);
nand I_20404 (I349945,I536148,I536163);
and I_20405 (I349962,I349945,I536175);
DFFARX1 I_20406 (I349962,I3035,I349894,I349988,);
not I_20407 (I349996,I536160);
DFFARX1 I_20408 (I536151,I3035,I349894,I350022,);
not I_20409 (I350030,I350022);
nor I_20410 (I350047,I350030,I349928);
and I_20411 (I350064,I350047,I536160);
nor I_20412 (I350081,I350030,I349996);
nor I_20413 (I349877,I349988,I350081);
DFFARX1 I_20414 (I536148,I3035,I349894,I350121,);
nor I_20415 (I350129,I350121,I349988);
not I_20416 (I350146,I350129);
not I_20417 (I350163,I350121);
nor I_20418 (I350180,I350163,I350064);
DFFARX1 I_20419 (I350180,I3035,I349894,I349880,);
nand I_20420 (I350211,I536166,I536157);
and I_20421 (I350228,I350211,I536169);
DFFARX1 I_20422 (I350228,I3035,I349894,I350254,);
nor I_20423 (I350262,I350254,I350121);
DFFARX1 I_20424 (I350262,I3035,I349894,I349862,);
nand I_20425 (I350293,I350254,I350163);
nand I_20426 (I349871,I350146,I350293);
not I_20427 (I350324,I350254);
nor I_20428 (I350341,I350324,I350064);
DFFARX1 I_20429 (I350341,I3035,I349894,I349883,);
nor I_20430 (I350372,I536154,I536157);
or I_20431 (I349874,I350121,I350372);
nor I_20432 (I349865,I350254,I350372);
or I_20433 (I349868,I349988,I350372);
DFFARX1 I_20434 (I350372,I3035,I349894,I349886,);
not I_20435 (I350472,I3042);
DFFARX1 I_20436 (I431409,I3035,I350472,I350498,);
not I_20437 (I350506,I350498);
nand I_20438 (I350523,I431397,I431415);
and I_20439 (I350540,I350523,I431412);
DFFARX1 I_20440 (I350540,I3035,I350472,I350566,);
not I_20441 (I350574,I431403);
DFFARX1 I_20442 (I431400,I3035,I350472,I350600,);
not I_20443 (I350608,I350600);
nor I_20444 (I350625,I350608,I350506);
and I_20445 (I350642,I350625,I431403);
nor I_20446 (I350659,I350608,I350574);
nor I_20447 (I350455,I350566,I350659);
DFFARX1 I_20448 (I431394,I3035,I350472,I350699,);
nor I_20449 (I350707,I350699,I350566);
not I_20450 (I350724,I350707);
not I_20451 (I350741,I350699);
nor I_20452 (I350758,I350741,I350642);
DFFARX1 I_20453 (I350758,I3035,I350472,I350458,);
nand I_20454 (I350789,I431394,I431397);
and I_20455 (I350806,I350789,I431400);
DFFARX1 I_20456 (I350806,I3035,I350472,I350832,);
nor I_20457 (I350840,I350832,I350699);
DFFARX1 I_20458 (I350840,I3035,I350472,I350440,);
nand I_20459 (I350871,I350832,I350741);
nand I_20460 (I350449,I350724,I350871);
not I_20461 (I350902,I350832);
nor I_20462 (I350919,I350902,I350642);
DFFARX1 I_20463 (I350919,I3035,I350472,I350461,);
nor I_20464 (I350950,I431406,I431397);
or I_20465 (I350452,I350699,I350950);
nor I_20466 (I350443,I350832,I350950);
or I_20467 (I350446,I350566,I350950);
DFFARX1 I_20468 (I350950,I3035,I350472,I350464,);
not I_20469 (I351050,I3042);
DFFARX1 I_20470 (I719860,I3035,I351050,I351076,);
not I_20471 (I351084,I351076);
nand I_20472 (I351101,I719845,I719833);
and I_20473 (I351118,I351101,I719848);
DFFARX1 I_20474 (I351118,I3035,I351050,I351144,);
not I_20475 (I351152,I719833);
DFFARX1 I_20476 (I719851,I3035,I351050,I351178,);
not I_20477 (I351186,I351178);
nor I_20478 (I351203,I351186,I351084);
and I_20479 (I351220,I351203,I719833);
nor I_20480 (I351237,I351186,I351152);
nor I_20481 (I351033,I351144,I351237);
DFFARX1 I_20482 (I719839,I3035,I351050,I351277,);
nor I_20483 (I351285,I351277,I351144);
not I_20484 (I351302,I351285);
not I_20485 (I351319,I351277);
nor I_20486 (I351336,I351319,I351220);
DFFARX1 I_20487 (I351336,I3035,I351050,I351036,);
nand I_20488 (I351367,I719836,I719842);
and I_20489 (I351384,I351367,I719857);
DFFARX1 I_20490 (I351384,I3035,I351050,I351410,);
nor I_20491 (I351418,I351410,I351277);
DFFARX1 I_20492 (I351418,I3035,I351050,I351018,);
nand I_20493 (I351449,I351410,I351319);
nand I_20494 (I351027,I351302,I351449);
not I_20495 (I351480,I351410);
nor I_20496 (I351497,I351480,I351220);
DFFARX1 I_20497 (I351497,I3035,I351050,I351039,);
nor I_20498 (I351528,I719854,I719842);
or I_20499 (I351030,I351277,I351528);
nor I_20500 (I351021,I351410,I351528);
or I_20501 (I351024,I351144,I351528);
DFFARX1 I_20502 (I351528,I3035,I351050,I351042,);
not I_20503 (I351628,I3042);
DFFARX1 I_20504 (I195645,I3035,I351628,I351654,);
not I_20505 (I351662,I351654);
nand I_20506 (I351679,I195648,I195624);
and I_20507 (I351696,I351679,I195621);
DFFARX1 I_20508 (I351696,I3035,I351628,I351722,);
not I_20509 (I351730,I195627);
DFFARX1 I_20510 (I195621,I3035,I351628,I351756,);
not I_20511 (I351764,I351756);
nor I_20512 (I351781,I351764,I351662);
and I_20513 (I351798,I351781,I195627);
nor I_20514 (I351815,I351764,I351730);
nor I_20515 (I351611,I351722,I351815);
DFFARX1 I_20516 (I195630,I3035,I351628,I351855,);
nor I_20517 (I351863,I351855,I351722);
not I_20518 (I351880,I351863);
not I_20519 (I351897,I351855);
nor I_20520 (I351914,I351897,I351798);
DFFARX1 I_20521 (I351914,I3035,I351628,I351614,);
nand I_20522 (I351945,I195633,I195642);
and I_20523 (I351962,I351945,I195639);
DFFARX1 I_20524 (I351962,I3035,I351628,I351988,);
nor I_20525 (I351996,I351988,I351855);
DFFARX1 I_20526 (I351996,I3035,I351628,I351596,);
nand I_20527 (I352027,I351988,I351897);
nand I_20528 (I351605,I351880,I352027);
not I_20529 (I352058,I351988);
nor I_20530 (I352075,I352058,I351798);
DFFARX1 I_20531 (I352075,I3035,I351628,I351617,);
nor I_20532 (I352106,I195636,I195642);
or I_20533 (I351608,I351855,I352106);
nor I_20534 (I351599,I351988,I352106);
or I_20535 (I351602,I351722,I352106);
DFFARX1 I_20536 (I352106,I3035,I351628,I351620,);
not I_20537 (I352206,I3042);
DFFARX1 I_20538 (I5431,I3035,I352206,I352232,);
not I_20539 (I352240,I352232);
nand I_20540 (I352257,I5434,I5446);
and I_20541 (I352274,I352257,I5425);
DFFARX1 I_20542 (I352274,I3035,I352206,I352300,);
not I_20543 (I352308,I5425);
DFFARX1 I_20544 (I5428,I3035,I352206,I352334,);
not I_20545 (I352342,I352334);
nor I_20546 (I352359,I352342,I352240);
and I_20547 (I352376,I352359,I5425);
nor I_20548 (I352393,I352342,I352308);
nor I_20549 (I352189,I352300,I352393);
DFFARX1 I_20550 (I5440,I3035,I352206,I352433,);
nor I_20551 (I352441,I352433,I352300);
not I_20552 (I352458,I352441);
not I_20553 (I352475,I352433);
nor I_20554 (I352492,I352475,I352376);
DFFARX1 I_20555 (I352492,I3035,I352206,I352192,);
nand I_20556 (I352523,I5443,I5428);
and I_20557 (I352540,I352523,I5437);
DFFARX1 I_20558 (I352540,I3035,I352206,I352566,);
nor I_20559 (I352574,I352566,I352433);
DFFARX1 I_20560 (I352574,I3035,I352206,I352174,);
nand I_20561 (I352605,I352566,I352475);
nand I_20562 (I352183,I352458,I352605);
not I_20563 (I352636,I352566);
nor I_20564 (I352653,I352636,I352376);
DFFARX1 I_20565 (I352653,I3035,I352206,I352195,);
nor I_20566 (I352684,I5431,I5428);
or I_20567 (I352186,I352433,I352684);
nor I_20568 (I352177,I352566,I352684);
or I_20569 (I352180,I352300,I352684);
DFFARX1 I_20570 (I352684,I3035,I352206,I352198,);
not I_20571 (I352784,I3042);
DFFARX1 I_20572 (I681736,I3035,I352784,I352810,);
not I_20573 (I352818,I352810);
nand I_20574 (I352835,I681760,I681742);
and I_20575 (I352852,I352835,I681748);
DFFARX1 I_20576 (I352852,I3035,I352784,I352878,);
not I_20577 (I352886,I681754);
DFFARX1 I_20578 (I681739,I3035,I352784,I352912,);
not I_20579 (I352920,I352912);
nor I_20580 (I352937,I352920,I352818);
and I_20581 (I352954,I352937,I681754);
nor I_20582 (I352971,I352920,I352886);
nor I_20583 (I352767,I352878,I352971);
DFFARX1 I_20584 (I681751,I3035,I352784,I353011,);
nor I_20585 (I353019,I353011,I352878);
not I_20586 (I353036,I353019);
not I_20587 (I353053,I353011);
nor I_20588 (I353070,I353053,I352954);
DFFARX1 I_20589 (I353070,I3035,I352784,I352770,);
nand I_20590 (I353101,I681757,I681745);
and I_20591 (I353118,I353101,I681739);
DFFARX1 I_20592 (I353118,I3035,I352784,I353144,);
nor I_20593 (I353152,I353144,I353011);
DFFARX1 I_20594 (I353152,I3035,I352784,I352752,);
nand I_20595 (I353183,I353144,I353053);
nand I_20596 (I352761,I353036,I353183);
not I_20597 (I353214,I353144);
nor I_20598 (I353231,I353214,I352954);
DFFARX1 I_20599 (I353231,I3035,I352784,I352773,);
nor I_20600 (I353262,I681736,I681745);
or I_20601 (I352764,I353011,I353262);
nor I_20602 (I352755,I353144,I353262);
or I_20603 (I352758,I352878,I353262);
DFFARX1 I_20604 (I353262,I3035,I352784,I352776,);
not I_20605 (I353362,I3042);
DFFARX1 I_20606 (I319228,I3035,I353362,I353388,);
not I_20607 (I353396,I353388);
nand I_20608 (I353413,I319237,I319246);
and I_20609 (I353430,I353413,I319252);
DFFARX1 I_20610 (I353430,I3035,I353362,I353456,);
not I_20611 (I353464,I319249);
DFFARX1 I_20612 (I319234,I3035,I353362,I353490,);
not I_20613 (I353498,I353490);
nor I_20614 (I353515,I353498,I353396);
and I_20615 (I353532,I353515,I319249);
nor I_20616 (I353549,I353498,I353464);
nor I_20617 (I353345,I353456,I353549);
DFFARX1 I_20618 (I319243,I3035,I353362,I353589,);
nor I_20619 (I353597,I353589,I353456);
not I_20620 (I353614,I353597);
not I_20621 (I353631,I353589);
nor I_20622 (I353648,I353631,I353532);
DFFARX1 I_20623 (I353648,I3035,I353362,I353348,);
nand I_20624 (I353679,I319240,I319231);
and I_20625 (I353696,I353679,I319228);
DFFARX1 I_20626 (I353696,I3035,I353362,I353722,);
nor I_20627 (I353730,I353722,I353589);
DFFARX1 I_20628 (I353730,I3035,I353362,I353330,);
nand I_20629 (I353761,I353722,I353631);
nand I_20630 (I353339,I353614,I353761);
not I_20631 (I353792,I353722);
nor I_20632 (I353809,I353792,I353532);
DFFARX1 I_20633 (I353809,I3035,I353362,I353351,);
nor I_20634 (I353840,I319231,I319231);
or I_20635 (I353342,I353589,I353840);
nor I_20636 (I353333,I353722,I353840);
or I_20637 (I353336,I353456,I353840);
DFFARX1 I_20638 (I353840,I3035,I353362,I353354,);
not I_20639 (I353940,I3042);
DFFARX1 I_20640 (I260910,I3035,I353940,I353966,);
not I_20641 (I353974,I353966);
nand I_20642 (I353991,I260901,I260919);
and I_20643 (I354008,I353991,I260922);
DFFARX1 I_20644 (I354008,I3035,I353940,I354034,);
not I_20645 (I354042,I260916);
DFFARX1 I_20646 (I260904,I3035,I353940,I354068,);
not I_20647 (I354076,I354068);
nor I_20648 (I354093,I354076,I353974);
and I_20649 (I354110,I354093,I260916);
nor I_20650 (I354127,I354076,I354042);
nor I_20651 (I353923,I354034,I354127);
DFFARX1 I_20652 (I260913,I3035,I353940,I354167,);
nor I_20653 (I354175,I354167,I354034);
not I_20654 (I354192,I354175);
not I_20655 (I354209,I354167);
nor I_20656 (I354226,I354209,I354110);
DFFARX1 I_20657 (I354226,I3035,I353940,I353926,);
nand I_20658 (I354257,I260928,I260925);
and I_20659 (I354274,I354257,I260907);
DFFARX1 I_20660 (I354274,I3035,I353940,I354300,);
nor I_20661 (I354308,I354300,I354167);
DFFARX1 I_20662 (I354308,I3035,I353940,I353908,);
nand I_20663 (I354339,I354300,I354209);
nand I_20664 (I353917,I354192,I354339);
not I_20665 (I354370,I354300);
nor I_20666 (I354387,I354370,I354110);
DFFARX1 I_20667 (I354387,I3035,I353940,I353929,);
nor I_20668 (I354418,I260901,I260925);
or I_20669 (I353920,I354167,I354418);
nor I_20670 (I353911,I354300,I354418);
or I_20671 (I353914,I354034,I354418);
DFFARX1 I_20672 (I354418,I3035,I353940,I353932,);
not I_20673 (I354518,I3042);
DFFARX1 I_20674 (I547051,I3035,I354518,I354544,);
not I_20675 (I354552,I354544);
nand I_20676 (I354569,I547048,I547066);
and I_20677 (I354586,I354569,I547063);
DFFARX1 I_20678 (I354586,I3035,I354518,I354612,);
not I_20679 (I354620,I547045);
DFFARX1 I_20680 (I547048,I3035,I354518,I354646,);
not I_20681 (I354654,I354646);
nor I_20682 (I354671,I354654,I354552);
and I_20683 (I354688,I354671,I547045);
nor I_20684 (I354705,I354654,I354620);
nor I_20685 (I354501,I354612,I354705);
DFFARX1 I_20686 (I547057,I3035,I354518,I354745,);
nor I_20687 (I354753,I354745,I354612);
not I_20688 (I354770,I354753);
not I_20689 (I354787,I354745);
nor I_20690 (I354804,I354787,I354688);
DFFARX1 I_20691 (I354804,I3035,I354518,I354504,);
nand I_20692 (I354835,I547060,I547045);
and I_20693 (I354852,I354835,I547051);
DFFARX1 I_20694 (I354852,I3035,I354518,I354878,);
nor I_20695 (I354886,I354878,I354745);
DFFARX1 I_20696 (I354886,I3035,I354518,I354486,);
nand I_20697 (I354917,I354878,I354787);
nand I_20698 (I354495,I354770,I354917);
not I_20699 (I354948,I354878);
nor I_20700 (I354965,I354948,I354688);
DFFARX1 I_20701 (I354965,I3035,I354518,I354507,);
nor I_20702 (I354996,I547054,I547045);
or I_20703 (I354498,I354745,I354996);
nor I_20704 (I354489,I354878,I354996);
or I_20705 (I354492,I354612,I354996);
DFFARX1 I_20706 (I354996,I3035,I354518,I354510,);
not I_20707 (I355096,I3042);
DFFARX1 I_20708 (I71575,I3035,I355096,I355122,);
not I_20709 (I355130,I355122);
nand I_20710 (I355147,I71584,I71593);
and I_20711 (I355164,I355147,I71572);
DFFARX1 I_20712 (I355164,I3035,I355096,I355190,);
not I_20713 (I355198,I71575);
DFFARX1 I_20714 (I71590,I3035,I355096,I355224,);
not I_20715 (I355232,I355224);
nor I_20716 (I355249,I355232,I355130);
and I_20717 (I355266,I355249,I71575);
nor I_20718 (I355283,I355232,I355198);
nor I_20719 (I355079,I355190,I355283);
DFFARX1 I_20720 (I71581,I3035,I355096,I355323,);
nor I_20721 (I355331,I355323,I355190);
not I_20722 (I355348,I355331);
not I_20723 (I355365,I355323);
nor I_20724 (I355382,I355365,I355266);
DFFARX1 I_20725 (I355382,I3035,I355096,I355082,);
nand I_20726 (I355413,I71596,I71572);
and I_20727 (I355430,I355413,I71578);
DFFARX1 I_20728 (I355430,I3035,I355096,I355456,);
nor I_20729 (I355464,I355456,I355323);
DFFARX1 I_20730 (I355464,I3035,I355096,I355064,);
nand I_20731 (I355495,I355456,I355365);
nand I_20732 (I355073,I355348,I355495);
not I_20733 (I355526,I355456);
nor I_20734 (I355543,I355526,I355266);
DFFARX1 I_20735 (I355543,I3035,I355096,I355085,);
nor I_20736 (I355574,I71587,I71572);
or I_20737 (I355076,I355323,I355574);
nor I_20738 (I355067,I355456,I355574);
or I_20739 (I355070,I355190,I355574);
DFFARX1 I_20740 (I355574,I3035,I355096,I355088,);
not I_20741 (I355674,I3042);
DFFARX1 I_20742 (I485138,I3035,I355674,I355700,);
not I_20743 (I355708,I355700);
nand I_20744 (I355725,I485114,I485129);
and I_20745 (I355742,I355725,I485141);
DFFARX1 I_20746 (I355742,I3035,I355674,I355768,);
not I_20747 (I355776,I485126);
DFFARX1 I_20748 (I485117,I3035,I355674,I355802,);
not I_20749 (I355810,I355802);
nor I_20750 (I355827,I355810,I355708);
and I_20751 (I355844,I355827,I485126);
nor I_20752 (I355861,I355810,I355776);
nor I_20753 (I355657,I355768,I355861);
DFFARX1 I_20754 (I485114,I3035,I355674,I355901,);
nor I_20755 (I355909,I355901,I355768);
not I_20756 (I355926,I355909);
not I_20757 (I355943,I355901);
nor I_20758 (I355960,I355943,I355844);
DFFARX1 I_20759 (I355960,I3035,I355674,I355660,);
nand I_20760 (I355991,I485132,I485123);
and I_20761 (I356008,I355991,I485135);
DFFARX1 I_20762 (I356008,I3035,I355674,I356034,);
nor I_20763 (I356042,I356034,I355901);
DFFARX1 I_20764 (I356042,I3035,I355674,I355642,);
nand I_20765 (I356073,I356034,I355943);
nand I_20766 (I355651,I355926,I356073);
not I_20767 (I356104,I356034);
nor I_20768 (I356121,I356104,I355844);
DFFARX1 I_20769 (I356121,I3035,I355674,I355663,);
nor I_20770 (I356152,I485120,I485123);
or I_20771 (I355654,I355901,I356152);
nor I_20772 (I355645,I356034,I356152);
or I_20773 (I355648,I355768,I356152);
DFFARX1 I_20774 (I356152,I3035,I355674,I355666,);
not I_20775 (I356252,I3042);
DFFARX1 I_20776 (I73156,I3035,I356252,I356278,);
not I_20777 (I356286,I356278);
nand I_20778 (I356303,I73165,I73174);
and I_20779 (I356320,I356303,I73153);
DFFARX1 I_20780 (I356320,I3035,I356252,I356346,);
not I_20781 (I356354,I73156);
DFFARX1 I_20782 (I73171,I3035,I356252,I356380,);
not I_20783 (I356388,I356380);
nor I_20784 (I356405,I356388,I356286);
and I_20785 (I356422,I356405,I73156);
nor I_20786 (I356439,I356388,I356354);
nor I_20787 (I356235,I356346,I356439);
DFFARX1 I_20788 (I73162,I3035,I356252,I356479,);
nor I_20789 (I356487,I356479,I356346);
not I_20790 (I356504,I356487);
not I_20791 (I356521,I356479);
nor I_20792 (I356538,I356521,I356422);
DFFARX1 I_20793 (I356538,I3035,I356252,I356238,);
nand I_20794 (I356569,I73177,I73153);
and I_20795 (I356586,I356569,I73159);
DFFARX1 I_20796 (I356586,I3035,I356252,I356612,);
nor I_20797 (I356620,I356612,I356479);
DFFARX1 I_20798 (I356620,I3035,I356252,I356220,);
nand I_20799 (I356651,I356612,I356521);
nand I_20800 (I356229,I356504,I356651);
not I_20801 (I356682,I356612);
nor I_20802 (I356699,I356682,I356422);
DFFARX1 I_20803 (I356699,I3035,I356252,I356241,);
nor I_20804 (I356730,I73168,I73153);
or I_20805 (I356232,I356479,I356730);
nor I_20806 (I356223,I356612,I356730);
or I_20807 (I356226,I356346,I356730);
DFFARX1 I_20808 (I356730,I3035,I356252,I356244,);
not I_20809 (I356830,I3042);
DFFARX1 I_20810 (I739495,I3035,I356830,I356856,);
not I_20811 (I356864,I356856);
nand I_20812 (I356881,I739480,I739468);
and I_20813 (I356898,I356881,I739483);
DFFARX1 I_20814 (I356898,I3035,I356830,I356924,);
not I_20815 (I356932,I739468);
DFFARX1 I_20816 (I739486,I3035,I356830,I356958,);
not I_20817 (I356966,I356958);
nor I_20818 (I356983,I356966,I356864);
and I_20819 (I357000,I356983,I739468);
nor I_20820 (I357017,I356966,I356932);
nor I_20821 (I356813,I356924,I357017);
DFFARX1 I_20822 (I739474,I3035,I356830,I357057,);
nor I_20823 (I357065,I357057,I356924);
not I_20824 (I357082,I357065);
not I_20825 (I357099,I357057);
nor I_20826 (I357116,I357099,I357000);
DFFARX1 I_20827 (I357116,I3035,I356830,I356816,);
nand I_20828 (I357147,I739471,I739477);
and I_20829 (I357164,I357147,I739492);
DFFARX1 I_20830 (I357164,I3035,I356830,I357190,);
nor I_20831 (I357198,I357190,I357057);
DFFARX1 I_20832 (I357198,I3035,I356830,I356798,);
nand I_20833 (I357229,I357190,I357099);
nand I_20834 (I356807,I357082,I357229);
not I_20835 (I357260,I357190);
nor I_20836 (I357277,I357260,I357000);
DFFARX1 I_20837 (I357277,I3035,I356830,I356819,);
nor I_20838 (I357308,I739489,I739477);
or I_20839 (I356810,I357057,I357308);
nor I_20840 (I356801,I357190,I357308);
or I_20841 (I356804,I356924,I357308);
DFFARX1 I_20842 (I357308,I3035,I356830,I356822,);
not I_20843 (I357408,I3042);
DFFARX1 I_20844 (I622016,I3035,I357408,I357434,);
not I_20845 (I357442,I357434);
nand I_20846 (I357459,I621998,I622010);
and I_20847 (I357476,I357459,I622013);
DFFARX1 I_20848 (I357476,I3035,I357408,I357502,);
not I_20849 (I357510,I622007);
DFFARX1 I_20850 (I622004,I3035,I357408,I357536,);
not I_20851 (I357544,I357536);
nor I_20852 (I357561,I357544,I357442);
and I_20853 (I357578,I357561,I622007);
nor I_20854 (I357595,I357544,I357510);
nor I_20855 (I357391,I357502,I357595);
DFFARX1 I_20856 (I622022,I3035,I357408,I357635,);
nor I_20857 (I357643,I357635,I357502);
not I_20858 (I357660,I357643);
not I_20859 (I357677,I357635);
nor I_20860 (I357694,I357677,I357578);
DFFARX1 I_20861 (I357694,I3035,I357408,I357394,);
nand I_20862 (I357725,I622001,I622001);
and I_20863 (I357742,I357725,I621998);
DFFARX1 I_20864 (I357742,I3035,I357408,I357768,);
nor I_20865 (I357776,I357768,I357635);
DFFARX1 I_20866 (I357776,I3035,I357408,I357376,);
nand I_20867 (I357807,I357768,I357677);
nand I_20868 (I357385,I357660,I357807);
not I_20869 (I357838,I357768);
nor I_20870 (I357855,I357838,I357578);
DFFARX1 I_20871 (I357855,I3035,I357408,I357397,);
nor I_20872 (I357886,I622019,I622001);
or I_20873 (I357388,I357635,I357886);
nor I_20874 (I357379,I357768,I357886);
or I_20875 (I357382,I357502,I357886);
DFFARX1 I_20876 (I357886,I3035,I357408,I357400,);
not I_20877 (I357986,I3042);
DFFARX1 I_20878 (I333678,I3035,I357986,I358012,);
not I_20879 (I358020,I358012);
nand I_20880 (I358037,I333687,I333696);
and I_20881 (I358054,I358037,I333702);
DFFARX1 I_20882 (I358054,I3035,I357986,I358080,);
not I_20883 (I358088,I333699);
DFFARX1 I_20884 (I333684,I3035,I357986,I358114,);
not I_20885 (I358122,I358114);
nor I_20886 (I358139,I358122,I358020);
and I_20887 (I358156,I358139,I333699);
nor I_20888 (I358173,I358122,I358088);
nor I_20889 (I357969,I358080,I358173);
DFFARX1 I_20890 (I333693,I3035,I357986,I358213,);
nor I_20891 (I358221,I358213,I358080);
not I_20892 (I358238,I358221);
not I_20893 (I358255,I358213);
nor I_20894 (I358272,I358255,I358156);
DFFARX1 I_20895 (I358272,I3035,I357986,I357972,);
nand I_20896 (I358303,I333690,I333681);
and I_20897 (I358320,I358303,I333678);
DFFARX1 I_20898 (I358320,I3035,I357986,I358346,);
nor I_20899 (I358354,I358346,I358213);
DFFARX1 I_20900 (I358354,I3035,I357986,I357954,);
nand I_20901 (I358385,I358346,I358255);
nand I_20902 (I357963,I358238,I358385);
not I_20903 (I358416,I358346);
nor I_20904 (I358433,I358416,I358156);
DFFARX1 I_20905 (I358433,I3035,I357986,I357975,);
nor I_20906 (I358464,I333681,I333681);
or I_20907 (I357966,I358213,I358464);
nor I_20908 (I357957,I358346,I358464);
or I_20909 (I357960,I358080,I358464);
DFFARX1 I_20910 (I358464,I3035,I357986,I357978,);
not I_20911 (I358564,I3042);
DFFARX1 I_20912 (I41536,I3035,I358564,I358590,);
not I_20913 (I358598,I358590);
nand I_20914 (I358615,I41545,I41554);
and I_20915 (I358632,I358615,I41533);
DFFARX1 I_20916 (I358632,I3035,I358564,I358658,);
not I_20917 (I358666,I41536);
DFFARX1 I_20918 (I41551,I3035,I358564,I358692,);
not I_20919 (I358700,I358692);
nor I_20920 (I358717,I358700,I358598);
and I_20921 (I358734,I358717,I41536);
nor I_20922 (I358751,I358700,I358666);
nor I_20923 (I358547,I358658,I358751);
DFFARX1 I_20924 (I41542,I3035,I358564,I358791,);
nor I_20925 (I358799,I358791,I358658);
not I_20926 (I358816,I358799);
not I_20927 (I358833,I358791);
nor I_20928 (I358850,I358833,I358734);
DFFARX1 I_20929 (I358850,I3035,I358564,I358550,);
nand I_20930 (I358881,I41557,I41533);
and I_20931 (I358898,I358881,I41539);
DFFARX1 I_20932 (I358898,I3035,I358564,I358924,);
nor I_20933 (I358932,I358924,I358791);
DFFARX1 I_20934 (I358932,I3035,I358564,I358532,);
nand I_20935 (I358963,I358924,I358833);
nand I_20936 (I358541,I358816,I358963);
not I_20937 (I358994,I358924);
nor I_20938 (I359011,I358994,I358734);
DFFARX1 I_20939 (I359011,I3035,I358564,I358553,);
nor I_20940 (I359042,I41548,I41533);
or I_20941 (I358544,I358791,I359042);
nor I_20942 (I358535,I358924,I359042);
or I_20943 (I358538,I358658,I359042);
DFFARX1 I_20944 (I359042,I3035,I358564,I358556,);
not I_20945 (I359142,I3042);
DFFARX1 I_20946 (I472515,I3035,I359142,I359168,);
not I_20947 (I359176,I359168);
nand I_20948 (I359193,I472503,I472521);
and I_20949 (I359210,I359193,I472518);
DFFARX1 I_20950 (I359210,I3035,I359142,I359236,);
not I_20951 (I359244,I472509);
DFFARX1 I_20952 (I472506,I3035,I359142,I359270,);
not I_20953 (I359278,I359270);
nor I_20954 (I359295,I359278,I359176);
and I_20955 (I359312,I359295,I472509);
nor I_20956 (I359329,I359278,I359244);
nor I_20957 (I359125,I359236,I359329);
DFFARX1 I_20958 (I472500,I3035,I359142,I359369,);
nor I_20959 (I359377,I359369,I359236);
not I_20960 (I359394,I359377);
not I_20961 (I359411,I359369);
nor I_20962 (I359428,I359411,I359312);
DFFARX1 I_20963 (I359428,I3035,I359142,I359128,);
nand I_20964 (I359459,I472500,I472503);
and I_20965 (I359476,I359459,I472506);
DFFARX1 I_20966 (I359476,I3035,I359142,I359502,);
nor I_20967 (I359510,I359502,I359369);
DFFARX1 I_20968 (I359510,I3035,I359142,I359110,);
nand I_20969 (I359541,I359502,I359411);
nand I_20970 (I359119,I359394,I359541);
not I_20971 (I359572,I359502);
nor I_20972 (I359589,I359572,I359312);
DFFARX1 I_20973 (I359589,I3035,I359142,I359131,);
nor I_20974 (I359620,I472512,I472503);
or I_20975 (I359122,I359369,I359620);
nor I_20976 (I359113,I359502,I359620);
or I_20977 (I359116,I359236,I359620);
DFFARX1 I_20978 (I359620,I3035,I359142,I359134,);
not I_20979 (I359720,I3042);
DFFARX1 I_20980 (I35739,I3035,I359720,I359746,);
not I_20981 (I359754,I359746);
nand I_20982 (I359771,I35748,I35757);
and I_20983 (I359788,I359771,I35736);
DFFARX1 I_20984 (I359788,I3035,I359720,I359814,);
not I_20985 (I359822,I35739);
DFFARX1 I_20986 (I35754,I3035,I359720,I359848,);
not I_20987 (I359856,I359848);
nor I_20988 (I359873,I359856,I359754);
and I_20989 (I359890,I359873,I35739);
nor I_20990 (I359907,I359856,I359822);
nor I_20991 (I359703,I359814,I359907);
DFFARX1 I_20992 (I35745,I3035,I359720,I359947,);
nor I_20993 (I359955,I359947,I359814);
not I_20994 (I359972,I359955);
not I_20995 (I359989,I359947);
nor I_20996 (I360006,I359989,I359890);
DFFARX1 I_20997 (I360006,I3035,I359720,I359706,);
nand I_20998 (I360037,I35760,I35736);
and I_20999 (I360054,I360037,I35742);
DFFARX1 I_21000 (I360054,I3035,I359720,I360080,);
nor I_21001 (I360088,I360080,I359947);
DFFARX1 I_21002 (I360088,I3035,I359720,I359688,);
nand I_21003 (I360119,I360080,I359989);
nand I_21004 (I359697,I359972,I360119);
not I_21005 (I360150,I360080);
nor I_21006 (I360167,I360150,I359890);
DFFARX1 I_21007 (I360167,I3035,I359720,I359709,);
nor I_21008 (I360198,I35751,I35736);
or I_21009 (I359700,I359947,I360198);
nor I_21010 (I359691,I360080,I360198);
or I_21011 (I359694,I359814,I360198);
DFFARX1 I_21012 (I360198,I3035,I359720,I359712,);
not I_21013 (I360298,I3042);
DFFARX1 I_21014 (I215671,I3035,I360298,I360324,);
not I_21015 (I360332,I360324);
nand I_21016 (I360349,I215674,I215650);
and I_21017 (I360366,I360349,I215647);
DFFARX1 I_21018 (I360366,I3035,I360298,I360392,);
not I_21019 (I360400,I215653);
DFFARX1 I_21020 (I215647,I3035,I360298,I360426,);
not I_21021 (I360434,I360426);
nor I_21022 (I360451,I360434,I360332);
and I_21023 (I360468,I360451,I215653);
nor I_21024 (I360485,I360434,I360400);
nor I_21025 (I360281,I360392,I360485);
DFFARX1 I_21026 (I215656,I3035,I360298,I360525,);
nor I_21027 (I360533,I360525,I360392);
not I_21028 (I360550,I360533);
not I_21029 (I360567,I360525);
nor I_21030 (I360584,I360567,I360468);
DFFARX1 I_21031 (I360584,I3035,I360298,I360284,);
nand I_21032 (I360615,I215659,I215668);
and I_21033 (I360632,I360615,I215665);
DFFARX1 I_21034 (I360632,I3035,I360298,I360658,);
nor I_21035 (I360666,I360658,I360525);
DFFARX1 I_21036 (I360666,I3035,I360298,I360266,);
nand I_21037 (I360697,I360658,I360567);
nand I_21038 (I360275,I360550,I360697);
not I_21039 (I360728,I360658);
nor I_21040 (I360745,I360728,I360468);
DFFARX1 I_21041 (I360745,I3035,I360298,I360287,);
nor I_21042 (I360776,I215662,I215668);
or I_21043 (I360278,I360525,I360776);
nor I_21044 (I360269,I360658,I360776);
or I_21045 (I360272,I360392,I360776);
DFFARX1 I_21046 (I360776,I3035,I360298,I360290,);
not I_21047 (I360876,I3042);
DFFARX1 I_21048 (I672488,I3035,I360876,I360902,);
not I_21049 (I360910,I360902);
nand I_21050 (I360927,I672512,I672494);
and I_21051 (I360944,I360927,I672500);
DFFARX1 I_21052 (I360944,I3035,I360876,I360970,);
not I_21053 (I360978,I672506);
DFFARX1 I_21054 (I672491,I3035,I360876,I361004,);
not I_21055 (I361012,I361004);
nor I_21056 (I361029,I361012,I360910);
and I_21057 (I361046,I361029,I672506);
nor I_21058 (I361063,I361012,I360978);
nor I_21059 (I360859,I360970,I361063);
DFFARX1 I_21060 (I672503,I3035,I360876,I361103,);
nor I_21061 (I361111,I361103,I360970);
not I_21062 (I361128,I361111);
not I_21063 (I361145,I361103);
nor I_21064 (I361162,I361145,I361046);
DFFARX1 I_21065 (I361162,I3035,I360876,I360862,);
nand I_21066 (I361193,I672509,I672497);
and I_21067 (I361210,I361193,I672491);
DFFARX1 I_21068 (I361210,I3035,I360876,I361236,);
nor I_21069 (I361244,I361236,I361103);
DFFARX1 I_21070 (I361244,I3035,I360876,I360844,);
nand I_21071 (I361275,I361236,I361145);
nand I_21072 (I360853,I361128,I361275);
not I_21073 (I361306,I361236);
nor I_21074 (I361323,I361306,I361046);
DFFARX1 I_21075 (I361323,I3035,I360876,I360865,);
nor I_21076 (I361354,I672488,I672497);
or I_21077 (I360856,I361103,I361354);
nor I_21078 (I360847,I361236,I361354);
or I_21079 (I360850,I360970,I361354);
DFFARX1 I_21080 (I361354,I3035,I360876,I360868,);
not I_21081 (I361454,I3042);
DFFARX1 I_21082 (I624906,I3035,I361454,I361480,);
not I_21083 (I361488,I361480);
nand I_21084 (I361505,I624888,I624900);
and I_21085 (I361522,I361505,I624903);
DFFARX1 I_21086 (I361522,I3035,I361454,I361548,);
not I_21087 (I361556,I624897);
DFFARX1 I_21088 (I624894,I3035,I361454,I361582,);
not I_21089 (I361590,I361582);
nor I_21090 (I361607,I361590,I361488);
and I_21091 (I361624,I361607,I624897);
nor I_21092 (I361641,I361590,I361556);
nor I_21093 (I361437,I361548,I361641);
DFFARX1 I_21094 (I624912,I3035,I361454,I361681,);
nor I_21095 (I361689,I361681,I361548);
not I_21096 (I361706,I361689);
not I_21097 (I361723,I361681);
nor I_21098 (I361740,I361723,I361624);
DFFARX1 I_21099 (I361740,I3035,I361454,I361440,);
nand I_21100 (I361771,I624891,I624891);
and I_21101 (I361788,I361771,I624888);
DFFARX1 I_21102 (I361788,I3035,I361454,I361814,);
nor I_21103 (I361822,I361814,I361681);
DFFARX1 I_21104 (I361822,I3035,I361454,I361422,);
nand I_21105 (I361853,I361814,I361723);
nand I_21106 (I361431,I361706,I361853);
not I_21107 (I361884,I361814);
nor I_21108 (I361901,I361884,I361624);
DFFARX1 I_21109 (I361901,I3035,I361454,I361443,);
nor I_21110 (I361932,I624909,I624891);
or I_21111 (I361434,I361681,I361932);
nor I_21112 (I361425,I361814,I361932);
or I_21113 (I361428,I361548,I361932);
DFFARX1 I_21114 (I361932,I3035,I361454,I361446,);
not I_21115 (I362032,I3042);
DFFARX1 I_21116 (I426139,I3035,I362032,I362058,);
not I_21117 (I362066,I362058);
nand I_21118 (I362083,I426127,I426145);
and I_21119 (I362100,I362083,I426142);
DFFARX1 I_21120 (I362100,I3035,I362032,I362126,);
not I_21121 (I362134,I426133);
DFFARX1 I_21122 (I426130,I3035,I362032,I362160,);
not I_21123 (I362168,I362160);
nor I_21124 (I362185,I362168,I362066);
and I_21125 (I362202,I362185,I426133);
nor I_21126 (I362219,I362168,I362134);
nor I_21127 (I362015,I362126,I362219);
DFFARX1 I_21128 (I426124,I3035,I362032,I362259,);
nor I_21129 (I362267,I362259,I362126);
not I_21130 (I362284,I362267);
not I_21131 (I362301,I362259);
nor I_21132 (I362318,I362301,I362202);
DFFARX1 I_21133 (I362318,I3035,I362032,I362018,);
nand I_21134 (I362349,I426124,I426127);
and I_21135 (I362366,I362349,I426130);
DFFARX1 I_21136 (I362366,I3035,I362032,I362392,);
nor I_21137 (I362400,I362392,I362259);
DFFARX1 I_21138 (I362400,I3035,I362032,I362000,);
nand I_21139 (I362431,I362392,I362301);
nand I_21140 (I362009,I362284,I362431);
not I_21141 (I362462,I362392);
nor I_21142 (I362479,I362462,I362202);
DFFARX1 I_21143 (I362479,I3035,I362032,I362021,);
nor I_21144 (I362510,I426136,I426127);
or I_21145 (I362012,I362259,I362510);
nor I_21146 (I362003,I362392,I362510);
or I_21147 (I362006,I362126,I362510);
DFFARX1 I_21148 (I362510,I3035,I362032,I362024,);
not I_21149 (I362610,I3042);
DFFARX1 I_21150 (I715100,I3035,I362610,I362636,);
not I_21151 (I362644,I362636);
nand I_21152 (I362661,I715085,I715073);
and I_21153 (I362678,I362661,I715088);
DFFARX1 I_21154 (I362678,I3035,I362610,I362704,);
not I_21155 (I362712,I715073);
DFFARX1 I_21156 (I715091,I3035,I362610,I362738,);
not I_21157 (I362746,I362738);
nor I_21158 (I362763,I362746,I362644);
and I_21159 (I362780,I362763,I715073);
nor I_21160 (I362797,I362746,I362712);
nor I_21161 (I362593,I362704,I362797);
DFFARX1 I_21162 (I715079,I3035,I362610,I362837,);
nor I_21163 (I362845,I362837,I362704);
not I_21164 (I362862,I362845);
not I_21165 (I362879,I362837);
nor I_21166 (I362896,I362879,I362780);
DFFARX1 I_21167 (I362896,I3035,I362610,I362596,);
nand I_21168 (I362927,I715076,I715082);
and I_21169 (I362944,I362927,I715097);
DFFARX1 I_21170 (I362944,I3035,I362610,I362970,);
nor I_21171 (I362978,I362970,I362837);
DFFARX1 I_21172 (I362978,I3035,I362610,I362578,);
nand I_21173 (I363009,I362970,I362879);
nand I_21174 (I362587,I362862,I363009);
not I_21175 (I363040,I362970);
nor I_21176 (I363057,I363040,I362780);
DFFARX1 I_21177 (I363057,I3035,I362610,I362599,);
nor I_21178 (I363088,I715094,I715082);
or I_21179 (I362590,I362837,I363088);
nor I_21180 (I362581,I362970,I363088);
or I_21181 (I362584,I362704,I363088);
DFFARX1 I_21182 (I363088,I3035,I362610,I362602,);
not I_21183 (I363188,I3042);
DFFARX1 I_21184 (I62616,I3035,I363188,I363214,);
not I_21185 (I363222,I363214);
nand I_21186 (I363239,I62625,I62634);
and I_21187 (I363256,I363239,I62613);
DFFARX1 I_21188 (I363256,I3035,I363188,I363282,);
not I_21189 (I363290,I62616);
DFFARX1 I_21190 (I62631,I3035,I363188,I363316,);
not I_21191 (I363324,I363316);
nor I_21192 (I363341,I363324,I363222);
and I_21193 (I363358,I363341,I62616);
nor I_21194 (I363375,I363324,I363290);
nor I_21195 (I363171,I363282,I363375);
DFFARX1 I_21196 (I62622,I3035,I363188,I363415,);
nor I_21197 (I363423,I363415,I363282);
not I_21198 (I363440,I363423);
not I_21199 (I363457,I363415);
nor I_21200 (I363474,I363457,I363358);
DFFARX1 I_21201 (I363474,I3035,I363188,I363174,);
nand I_21202 (I363505,I62637,I62613);
and I_21203 (I363522,I363505,I62619);
DFFARX1 I_21204 (I363522,I3035,I363188,I363548,);
nor I_21205 (I363556,I363548,I363415);
DFFARX1 I_21206 (I363556,I3035,I363188,I363156,);
nand I_21207 (I363587,I363548,I363457);
nand I_21208 (I363165,I363440,I363587);
not I_21209 (I363618,I363548);
nor I_21210 (I363635,I363618,I363358);
DFFARX1 I_21211 (I363635,I3035,I363188,I363177,);
nor I_21212 (I363666,I62628,I62613);
or I_21213 (I363168,I363415,I363666);
nor I_21214 (I363159,I363548,I363666);
or I_21215 (I363162,I363282,I363666);
DFFARX1 I_21216 (I363666,I3035,I363188,I363180,);
not I_21217 (I363766,I3042);
DFFARX1 I_21218 (I197226,I3035,I363766,I363792,);
not I_21219 (I363800,I363792);
nand I_21220 (I363817,I197229,I197205);
and I_21221 (I363834,I363817,I197202);
DFFARX1 I_21222 (I363834,I3035,I363766,I363860,);
not I_21223 (I363868,I197208);
DFFARX1 I_21224 (I197202,I3035,I363766,I363894,);
not I_21225 (I363902,I363894);
nor I_21226 (I363919,I363902,I363800);
and I_21227 (I363936,I363919,I197208);
nor I_21228 (I363953,I363902,I363868);
nor I_21229 (I363749,I363860,I363953);
DFFARX1 I_21230 (I197211,I3035,I363766,I363993,);
nor I_21231 (I364001,I363993,I363860);
not I_21232 (I364018,I364001);
not I_21233 (I364035,I363993);
nor I_21234 (I364052,I364035,I363936);
DFFARX1 I_21235 (I364052,I3035,I363766,I363752,);
nand I_21236 (I364083,I197214,I197223);
and I_21237 (I364100,I364083,I197220);
DFFARX1 I_21238 (I364100,I3035,I363766,I364126,);
nor I_21239 (I364134,I364126,I363993);
DFFARX1 I_21240 (I364134,I3035,I363766,I363734,);
nand I_21241 (I364165,I364126,I364035);
nand I_21242 (I363743,I364018,I364165);
not I_21243 (I364196,I364126);
nor I_21244 (I364213,I364196,I363936);
DFFARX1 I_21245 (I364213,I3035,I363766,I363755,);
nor I_21246 (I364244,I197217,I197223);
or I_21247 (I363746,I363993,I364244);
nor I_21248 (I363737,I364126,I364244);
or I_21249 (I363740,I363860,I364244);
DFFARX1 I_21250 (I364244,I3035,I363766,I363758,);
not I_21251 (I364344,I3042);
DFFARX1 I_21252 (I221995,I3035,I364344,I364370,);
not I_21253 (I364378,I364370);
nand I_21254 (I364395,I221998,I221974);
and I_21255 (I364412,I364395,I221971);
DFFARX1 I_21256 (I364412,I3035,I364344,I364438,);
not I_21257 (I364446,I221977);
DFFARX1 I_21258 (I221971,I3035,I364344,I364472,);
not I_21259 (I364480,I364472);
nor I_21260 (I364497,I364480,I364378);
and I_21261 (I364514,I364497,I221977);
nor I_21262 (I364531,I364480,I364446);
nor I_21263 (I364327,I364438,I364531);
DFFARX1 I_21264 (I221980,I3035,I364344,I364571,);
nor I_21265 (I364579,I364571,I364438);
not I_21266 (I364596,I364579);
not I_21267 (I364613,I364571);
nor I_21268 (I364630,I364613,I364514);
DFFARX1 I_21269 (I364630,I3035,I364344,I364330,);
nand I_21270 (I364661,I221983,I221992);
and I_21271 (I364678,I364661,I221989);
DFFARX1 I_21272 (I364678,I3035,I364344,I364704,);
nor I_21273 (I364712,I364704,I364571);
DFFARX1 I_21274 (I364712,I3035,I364344,I364312,);
nand I_21275 (I364743,I364704,I364613);
nand I_21276 (I364321,I364596,I364743);
not I_21277 (I364774,I364704);
nor I_21278 (I364791,I364774,I364514);
DFFARX1 I_21279 (I364791,I3035,I364344,I364333,);
nor I_21280 (I364822,I221986,I221992);
or I_21281 (I364324,I364571,I364822);
nor I_21282 (I364315,I364704,I364822);
or I_21283 (I364318,I364438,I364822);
DFFARX1 I_21284 (I364822,I3035,I364344,I364336,);
not I_21285 (I364922,I3042);
DFFARX1 I_21286 (I329054,I3035,I364922,I364948,);
not I_21287 (I364956,I364948);
nand I_21288 (I364973,I329063,I329072);
and I_21289 (I364990,I364973,I329078);
DFFARX1 I_21290 (I364990,I3035,I364922,I365016,);
not I_21291 (I365024,I329075);
DFFARX1 I_21292 (I329060,I3035,I364922,I365050,);
not I_21293 (I365058,I365050);
nor I_21294 (I365075,I365058,I364956);
and I_21295 (I365092,I365075,I329075);
nor I_21296 (I365109,I365058,I365024);
nor I_21297 (I364905,I365016,I365109);
DFFARX1 I_21298 (I329069,I3035,I364922,I365149,);
nor I_21299 (I365157,I365149,I365016);
not I_21300 (I365174,I365157);
not I_21301 (I365191,I365149);
nor I_21302 (I365208,I365191,I365092);
DFFARX1 I_21303 (I365208,I3035,I364922,I364908,);
nand I_21304 (I365239,I329066,I329057);
and I_21305 (I365256,I365239,I329054);
DFFARX1 I_21306 (I365256,I3035,I364922,I365282,);
nor I_21307 (I365290,I365282,I365149);
DFFARX1 I_21308 (I365290,I3035,I364922,I364890,);
nand I_21309 (I365321,I365282,I365191);
nand I_21310 (I364899,I365174,I365321);
not I_21311 (I365352,I365282);
nor I_21312 (I365369,I365352,I365092);
DFFARX1 I_21313 (I365369,I3035,I364922,I364911,);
nor I_21314 (I365400,I329057,I329057);
or I_21315 (I364902,I365149,I365400);
nor I_21316 (I364893,I365282,I365400);
or I_21317 (I364896,I365016,I365400);
DFFARX1 I_21318 (I365400,I3035,I364922,I364914,);
not I_21319 (I365500,I3042);
DFFARX1 I_21320 (I119954,I3035,I365500,I365526,);
not I_21321 (I365534,I365526);
nand I_21322 (I365551,I119957,I119978);
and I_21323 (I365568,I365551,I119966);
DFFARX1 I_21324 (I365568,I3035,I365500,I365594,);
not I_21325 (I365602,I119963);
DFFARX1 I_21326 (I119954,I3035,I365500,I365628,);
not I_21327 (I365636,I365628);
nor I_21328 (I365653,I365636,I365534);
and I_21329 (I365670,I365653,I119963);
nor I_21330 (I365687,I365636,I365602);
nor I_21331 (I365483,I365594,I365687);
DFFARX1 I_21332 (I119972,I3035,I365500,I365727,);
nor I_21333 (I365735,I365727,I365594);
not I_21334 (I365752,I365735);
not I_21335 (I365769,I365727);
nor I_21336 (I365786,I365769,I365670);
DFFARX1 I_21337 (I365786,I3035,I365500,I365486,);
nand I_21338 (I365817,I119957,I119960);
and I_21339 (I365834,I365817,I119969);
DFFARX1 I_21340 (I365834,I3035,I365500,I365860,);
nor I_21341 (I365868,I365860,I365727);
DFFARX1 I_21342 (I365868,I3035,I365500,I365468,);
nand I_21343 (I365899,I365860,I365769);
nand I_21344 (I365477,I365752,I365899);
not I_21345 (I365930,I365860);
nor I_21346 (I365947,I365930,I365670);
DFFARX1 I_21347 (I365947,I3035,I365500,I365489,);
nor I_21348 (I365978,I119975,I119960);
or I_21349 (I365480,I365727,I365978);
nor I_21350 (I365471,I365860,I365978);
or I_21351 (I365474,I365594,I365978);
DFFARX1 I_21352 (I365978,I3035,I365500,I365492,);
not I_21353 (I366078,I3042);
DFFARX1 I_21354 (I425085,I3035,I366078,I366104,);
not I_21355 (I366112,I366104);
nand I_21356 (I366129,I425073,I425091);
and I_21357 (I366146,I366129,I425088);
DFFARX1 I_21358 (I366146,I3035,I366078,I366172,);
not I_21359 (I366180,I425079);
DFFARX1 I_21360 (I425076,I3035,I366078,I366206,);
not I_21361 (I366214,I366206);
nor I_21362 (I366231,I366214,I366112);
and I_21363 (I366248,I366231,I425079);
nor I_21364 (I366265,I366214,I366180);
nor I_21365 (I366061,I366172,I366265);
DFFARX1 I_21366 (I425070,I3035,I366078,I366305,);
nor I_21367 (I366313,I366305,I366172);
not I_21368 (I366330,I366313);
not I_21369 (I366347,I366305);
nor I_21370 (I366364,I366347,I366248);
DFFARX1 I_21371 (I366364,I3035,I366078,I366064,);
nand I_21372 (I366395,I425070,I425073);
and I_21373 (I366412,I366395,I425076);
DFFARX1 I_21374 (I366412,I3035,I366078,I366438,);
nor I_21375 (I366446,I366438,I366305);
DFFARX1 I_21376 (I366446,I3035,I366078,I366046,);
nand I_21377 (I366477,I366438,I366347);
nand I_21378 (I366055,I366330,I366477);
not I_21379 (I366508,I366438);
nor I_21380 (I366525,I366508,I366248);
DFFARX1 I_21381 (I366525,I3035,I366078,I366067,);
nor I_21382 (I366556,I425082,I425073);
or I_21383 (I366058,I366305,I366556);
nor I_21384 (I366049,I366438,I366556);
or I_21385 (I366052,I366172,I366556);
DFFARX1 I_21386 (I366556,I3035,I366078,I366070,);
not I_21387 (I366656,I3042);
DFFARX1 I_21388 (I157701,I3035,I366656,I366682,);
not I_21389 (I366690,I366682);
nand I_21390 (I366707,I157704,I157680);
and I_21391 (I366724,I366707,I157677);
DFFARX1 I_21392 (I366724,I3035,I366656,I366750,);
not I_21393 (I366758,I157683);
DFFARX1 I_21394 (I157677,I3035,I366656,I366784,);
not I_21395 (I366792,I366784);
nor I_21396 (I366809,I366792,I366690);
and I_21397 (I366826,I366809,I157683);
nor I_21398 (I366843,I366792,I366758);
nor I_21399 (I366639,I366750,I366843);
DFFARX1 I_21400 (I157686,I3035,I366656,I366883,);
nor I_21401 (I366891,I366883,I366750);
not I_21402 (I366908,I366891);
not I_21403 (I366925,I366883);
nor I_21404 (I366942,I366925,I366826);
DFFARX1 I_21405 (I366942,I3035,I366656,I366642,);
nand I_21406 (I366973,I157689,I157698);
and I_21407 (I366990,I366973,I157695);
DFFARX1 I_21408 (I366990,I3035,I366656,I367016,);
nor I_21409 (I367024,I367016,I366883);
DFFARX1 I_21410 (I367024,I3035,I366656,I366624,);
nand I_21411 (I367055,I367016,I366925);
nand I_21412 (I366633,I366908,I367055);
not I_21413 (I367086,I367016);
nor I_21414 (I367103,I367086,I366826);
DFFARX1 I_21415 (I367103,I3035,I366656,I366645,);
nor I_21416 (I367134,I157692,I157698);
or I_21417 (I366636,I366883,I367134);
nor I_21418 (I366627,I367016,I367134);
or I_21419 (I366630,I366750,I367134);
DFFARX1 I_21420 (I367134,I3035,I366656,I366648,);
not I_21421 (I367234,I3042);
DFFARX1 I_21422 (I11506,I3035,I367234,I367260,);
not I_21423 (I367268,I367260);
nand I_21424 (I367285,I11503,I11494);
and I_21425 (I367302,I367285,I11494);
DFFARX1 I_21426 (I367302,I3035,I367234,I367328,);
not I_21427 (I367336,I11497);
DFFARX1 I_21428 (I11512,I3035,I367234,I367362,);
not I_21429 (I367370,I367362);
nor I_21430 (I367387,I367370,I367268);
and I_21431 (I367404,I367387,I11497);
nor I_21432 (I367421,I367370,I367336);
nor I_21433 (I367217,I367328,I367421);
DFFARX1 I_21434 (I11497,I3035,I367234,I367461,);
nor I_21435 (I367469,I367461,I367328);
not I_21436 (I367486,I367469);
not I_21437 (I367503,I367461);
nor I_21438 (I367520,I367503,I367404);
DFFARX1 I_21439 (I367520,I3035,I367234,I367220,);
nand I_21440 (I367551,I11515,I11500);
and I_21441 (I367568,I367551,I11518);
DFFARX1 I_21442 (I367568,I3035,I367234,I367594,);
nor I_21443 (I367602,I367594,I367461);
DFFARX1 I_21444 (I367602,I3035,I367234,I367202,);
nand I_21445 (I367633,I367594,I367503);
nand I_21446 (I367211,I367486,I367633);
not I_21447 (I367664,I367594);
nor I_21448 (I367681,I367664,I367404);
DFFARX1 I_21449 (I367681,I3035,I367234,I367223,);
nor I_21450 (I367712,I11509,I11500);
or I_21451 (I367214,I367461,I367712);
nor I_21452 (I367205,I367594,I367712);
or I_21453 (I367208,I367328,I367712);
DFFARX1 I_21454 (I367712,I3035,I367234,I367226,);
not I_21455 (I367812,I3042);
DFFARX1 I_21456 (I106864,I3035,I367812,I367838,);
not I_21457 (I367846,I367838);
nand I_21458 (I367863,I106867,I106888);
and I_21459 (I367880,I367863,I106876);
DFFARX1 I_21460 (I367880,I3035,I367812,I367906,);
not I_21461 (I367914,I106873);
DFFARX1 I_21462 (I106864,I3035,I367812,I367940,);
not I_21463 (I367948,I367940);
nor I_21464 (I367965,I367948,I367846);
and I_21465 (I367982,I367965,I106873);
nor I_21466 (I367999,I367948,I367914);
nor I_21467 (I367795,I367906,I367999);
DFFARX1 I_21468 (I106882,I3035,I367812,I368039,);
nor I_21469 (I368047,I368039,I367906);
not I_21470 (I368064,I368047);
not I_21471 (I368081,I368039);
nor I_21472 (I368098,I368081,I367982);
DFFARX1 I_21473 (I368098,I3035,I367812,I367798,);
nand I_21474 (I368129,I106867,I106870);
and I_21475 (I368146,I368129,I106879);
DFFARX1 I_21476 (I368146,I3035,I367812,I368172,);
nor I_21477 (I368180,I368172,I368039);
DFFARX1 I_21478 (I368180,I3035,I367812,I367780,);
nand I_21479 (I368211,I368172,I368081);
nand I_21480 (I367789,I368064,I368211);
not I_21481 (I368242,I368172);
nor I_21482 (I368259,I368242,I367982);
DFFARX1 I_21483 (I368259,I3035,I367812,I367801,);
nor I_21484 (I368290,I106885,I106870);
or I_21485 (I367792,I368039,I368290);
nor I_21486 (I367783,I368172,I368290);
or I_21487 (I367786,I367906,I368290);
DFFARX1 I_21488 (I368290,I3035,I367812,I367804,);
not I_21489 (I368390,I3042);
DFFARX1 I_21490 (I701415,I3035,I368390,I368416,);
not I_21491 (I368424,I368416);
nand I_21492 (I368441,I701400,I701388);
and I_21493 (I368458,I368441,I701403);
DFFARX1 I_21494 (I368458,I3035,I368390,I368484,);
not I_21495 (I368492,I701388);
DFFARX1 I_21496 (I701406,I3035,I368390,I368518,);
not I_21497 (I368526,I368518);
nor I_21498 (I368543,I368526,I368424);
and I_21499 (I368560,I368543,I701388);
nor I_21500 (I368577,I368526,I368492);
nor I_21501 (I368373,I368484,I368577);
DFFARX1 I_21502 (I701394,I3035,I368390,I368617,);
nor I_21503 (I368625,I368617,I368484);
not I_21504 (I368642,I368625);
not I_21505 (I368659,I368617);
nor I_21506 (I368676,I368659,I368560);
DFFARX1 I_21507 (I368676,I3035,I368390,I368376,);
nand I_21508 (I368707,I701391,I701397);
and I_21509 (I368724,I368707,I701412);
DFFARX1 I_21510 (I368724,I3035,I368390,I368750,);
nor I_21511 (I368758,I368750,I368617);
DFFARX1 I_21512 (I368758,I3035,I368390,I368358,);
nand I_21513 (I368789,I368750,I368659);
nand I_21514 (I368367,I368642,I368789);
not I_21515 (I368820,I368750);
nor I_21516 (I368837,I368820,I368560);
DFFARX1 I_21517 (I368837,I3035,I368390,I368379,);
nor I_21518 (I368868,I701409,I701397);
or I_21519 (I368370,I368617,I368868);
nor I_21520 (I368361,I368750,I368868);
or I_21521 (I368364,I368484,I368868);
DFFARX1 I_21522 (I368868,I3035,I368390,I368382,);
not I_21523 (I368968,I3042);
DFFARX1 I_21524 (I204077,I3035,I368968,I368994,);
not I_21525 (I369002,I368994);
nand I_21526 (I369019,I204080,I204056);
and I_21527 (I369036,I369019,I204053);
DFFARX1 I_21528 (I369036,I3035,I368968,I369062,);
not I_21529 (I369070,I204059);
DFFARX1 I_21530 (I204053,I3035,I368968,I369096,);
not I_21531 (I369104,I369096);
nor I_21532 (I369121,I369104,I369002);
and I_21533 (I369138,I369121,I204059);
nor I_21534 (I369155,I369104,I369070);
nor I_21535 (I368951,I369062,I369155);
DFFARX1 I_21536 (I204062,I3035,I368968,I369195,);
nor I_21537 (I369203,I369195,I369062);
not I_21538 (I369220,I369203);
not I_21539 (I369237,I369195);
nor I_21540 (I369254,I369237,I369138);
DFFARX1 I_21541 (I369254,I3035,I368968,I368954,);
nand I_21542 (I369285,I204065,I204074);
and I_21543 (I369302,I369285,I204071);
DFFARX1 I_21544 (I369302,I3035,I368968,I369328,);
nor I_21545 (I369336,I369328,I369195);
DFFARX1 I_21546 (I369336,I3035,I368968,I368936,);
nand I_21547 (I369367,I369328,I369237);
nand I_21548 (I368945,I369220,I369367);
not I_21549 (I369398,I369328);
nor I_21550 (I369415,I369398,I369138);
DFFARX1 I_21551 (I369415,I3035,I368968,I368957,);
nor I_21552 (I369446,I204068,I204074);
or I_21553 (I368948,I369195,I369446);
nor I_21554 (I368939,I369328,I369446);
or I_21555 (I368942,I369062,I369446);
DFFARX1 I_21556 (I369446,I3035,I368968,I368960,);
not I_21557 (I369546,I3042);
DFFARX1 I_21558 (I38901,I3035,I369546,I369572,);
not I_21559 (I369580,I369572);
nand I_21560 (I369597,I38910,I38919);
and I_21561 (I369614,I369597,I38898);
DFFARX1 I_21562 (I369614,I3035,I369546,I369640,);
not I_21563 (I369648,I38901);
DFFARX1 I_21564 (I38916,I3035,I369546,I369674,);
not I_21565 (I369682,I369674);
nor I_21566 (I369699,I369682,I369580);
and I_21567 (I369716,I369699,I38901);
nor I_21568 (I369733,I369682,I369648);
nor I_21569 (I369529,I369640,I369733);
DFFARX1 I_21570 (I38907,I3035,I369546,I369773,);
nor I_21571 (I369781,I369773,I369640);
not I_21572 (I369798,I369781);
not I_21573 (I369815,I369773);
nor I_21574 (I369832,I369815,I369716);
DFFARX1 I_21575 (I369832,I3035,I369546,I369532,);
nand I_21576 (I369863,I38922,I38898);
and I_21577 (I369880,I369863,I38904);
DFFARX1 I_21578 (I369880,I3035,I369546,I369906,);
nor I_21579 (I369914,I369906,I369773);
DFFARX1 I_21580 (I369914,I3035,I369546,I369514,);
nand I_21581 (I369945,I369906,I369815);
nand I_21582 (I369523,I369798,I369945);
not I_21583 (I369976,I369906);
nor I_21584 (I369993,I369976,I369716);
DFFARX1 I_21585 (I369993,I3035,I369546,I369535,);
nor I_21586 (I370024,I38913,I38898);
or I_21587 (I369526,I369773,I370024);
nor I_21588 (I369517,I369906,I370024);
or I_21589 (I369520,I369640,I370024);
DFFARX1 I_21590 (I370024,I3035,I369546,I369538,);
not I_21591 (I370124,I3042);
DFFARX1 I_21592 (I114004,I3035,I370124,I370150,);
not I_21593 (I370158,I370150);
nand I_21594 (I370175,I114007,I114028);
and I_21595 (I370192,I370175,I114016);
DFFARX1 I_21596 (I370192,I3035,I370124,I370218,);
not I_21597 (I370226,I114013);
DFFARX1 I_21598 (I114004,I3035,I370124,I370252,);
not I_21599 (I370260,I370252);
nor I_21600 (I370277,I370260,I370158);
and I_21601 (I370294,I370277,I114013);
nor I_21602 (I370311,I370260,I370226);
nor I_21603 (I370107,I370218,I370311);
DFFARX1 I_21604 (I114022,I3035,I370124,I370351,);
nor I_21605 (I370359,I370351,I370218);
not I_21606 (I370376,I370359);
not I_21607 (I370393,I370351);
nor I_21608 (I370410,I370393,I370294);
DFFARX1 I_21609 (I370410,I3035,I370124,I370110,);
nand I_21610 (I370441,I114007,I114010);
and I_21611 (I370458,I370441,I114019);
DFFARX1 I_21612 (I370458,I3035,I370124,I370484,);
nor I_21613 (I370492,I370484,I370351);
DFFARX1 I_21614 (I370492,I3035,I370124,I370092,);
nand I_21615 (I370523,I370484,I370393);
nand I_21616 (I370101,I370376,I370523);
not I_21617 (I370554,I370484);
nor I_21618 (I370571,I370554,I370294);
DFFARX1 I_21619 (I370571,I3035,I370124,I370113,);
nor I_21620 (I370602,I114025,I114010);
or I_21621 (I370104,I370351,I370602);
nor I_21622 (I370095,I370484,I370602);
or I_21623 (I370098,I370218,I370602);
DFFARX1 I_21624 (I370602,I3035,I370124,I370116,);
not I_21625 (I370702,I3042);
DFFARX1 I_21626 (I44171,I3035,I370702,I370728,);
not I_21627 (I370736,I370728);
nand I_21628 (I370753,I44180,I44189);
and I_21629 (I370770,I370753,I44168);
DFFARX1 I_21630 (I370770,I3035,I370702,I370796,);
not I_21631 (I370804,I44171);
DFFARX1 I_21632 (I44186,I3035,I370702,I370830,);
not I_21633 (I370838,I370830);
nor I_21634 (I370855,I370838,I370736);
and I_21635 (I370872,I370855,I44171);
nor I_21636 (I370889,I370838,I370804);
nor I_21637 (I370685,I370796,I370889);
DFFARX1 I_21638 (I44177,I3035,I370702,I370929,);
nor I_21639 (I370937,I370929,I370796);
not I_21640 (I370954,I370937);
not I_21641 (I370971,I370929);
nor I_21642 (I370988,I370971,I370872);
DFFARX1 I_21643 (I370988,I3035,I370702,I370688,);
nand I_21644 (I371019,I44192,I44168);
and I_21645 (I371036,I371019,I44174);
DFFARX1 I_21646 (I371036,I3035,I370702,I371062,);
nor I_21647 (I371070,I371062,I370929);
DFFARX1 I_21648 (I371070,I3035,I370702,I370670,);
nand I_21649 (I371101,I371062,I370971);
nand I_21650 (I370679,I370954,I371101);
not I_21651 (I371132,I371062);
nor I_21652 (I371149,I371132,I370872);
DFFARX1 I_21653 (I371149,I3035,I370702,I370691,);
nor I_21654 (I371180,I44183,I44168);
or I_21655 (I370682,I370929,I371180);
nor I_21656 (I370673,I371062,I371180);
or I_21657 (I370676,I370796,I371180);
DFFARX1 I_21658 (I371180,I3035,I370702,I370694,);
not I_21659 (I371280,I3042);
DFFARX1 I_21660 (I305934,I3035,I371280,I371306,);
not I_21661 (I371314,I371306);
nand I_21662 (I371331,I305943,I305952);
and I_21663 (I371348,I371331,I305958);
DFFARX1 I_21664 (I371348,I3035,I371280,I371374,);
not I_21665 (I371382,I305955);
DFFARX1 I_21666 (I305940,I3035,I371280,I371408,);
not I_21667 (I371416,I371408);
nor I_21668 (I371433,I371416,I371314);
and I_21669 (I371450,I371433,I305955);
nor I_21670 (I371467,I371416,I371382);
nor I_21671 (I371263,I371374,I371467);
DFFARX1 I_21672 (I305949,I3035,I371280,I371507,);
nor I_21673 (I371515,I371507,I371374);
not I_21674 (I371532,I371515);
not I_21675 (I371549,I371507);
nor I_21676 (I371566,I371549,I371450);
DFFARX1 I_21677 (I371566,I3035,I371280,I371266,);
nand I_21678 (I371597,I305946,I305937);
and I_21679 (I371614,I371597,I305934);
DFFARX1 I_21680 (I371614,I3035,I371280,I371640,);
nor I_21681 (I371648,I371640,I371507);
DFFARX1 I_21682 (I371648,I3035,I371280,I371248,);
nand I_21683 (I371679,I371640,I371549);
nand I_21684 (I371257,I371532,I371679);
not I_21685 (I371710,I371640);
nor I_21686 (I371727,I371710,I371450);
DFFARX1 I_21687 (I371727,I3035,I371280,I371269,);
nor I_21688 (I371758,I305937,I305937);
or I_21689 (I371260,I371507,I371758);
nor I_21690 (I371251,I371640,I371758);
or I_21691 (I371254,I371374,I371758);
DFFARX1 I_21692 (I371758,I3035,I371280,I371272,);
not I_21693 (I371858,I3042);
DFFARX1 I_21694 (I681158,I3035,I371858,I371884,);
not I_21695 (I371892,I371884);
nand I_21696 (I371909,I681182,I681164);
and I_21697 (I371926,I371909,I681170);
DFFARX1 I_21698 (I371926,I3035,I371858,I371952,);
not I_21699 (I371960,I681176);
DFFARX1 I_21700 (I681161,I3035,I371858,I371986,);
not I_21701 (I371994,I371986);
nor I_21702 (I372011,I371994,I371892);
and I_21703 (I372028,I372011,I681176);
nor I_21704 (I372045,I371994,I371960);
nor I_21705 (I371841,I371952,I372045);
DFFARX1 I_21706 (I681173,I3035,I371858,I372085,);
nor I_21707 (I372093,I372085,I371952);
not I_21708 (I372110,I372093);
not I_21709 (I372127,I372085);
nor I_21710 (I372144,I372127,I372028);
DFFARX1 I_21711 (I372144,I3035,I371858,I371844,);
nand I_21712 (I372175,I681179,I681167);
and I_21713 (I372192,I372175,I681161);
DFFARX1 I_21714 (I372192,I3035,I371858,I372218,);
nor I_21715 (I372226,I372218,I372085);
DFFARX1 I_21716 (I372226,I3035,I371858,I371826,);
nand I_21717 (I372257,I372218,I372127);
nand I_21718 (I371835,I372110,I372257);
not I_21719 (I372288,I372218);
nor I_21720 (I372305,I372288,I372028);
DFFARX1 I_21721 (I372305,I3035,I371858,I371847,);
nor I_21722 (I372336,I681158,I681167);
or I_21723 (I371838,I372085,I372336);
nor I_21724 (I371829,I372218,I372336);
or I_21725 (I371832,I371952,I372336);
DFFARX1 I_21726 (I372336,I3035,I371858,I371850,);
not I_21727 (I372436,I3042);
DFFARX1 I_21728 (I652870,I3035,I372436,I372462,);
not I_21729 (I372470,I372462);
nand I_21730 (I372487,I652873,I652882);
and I_21731 (I372504,I372487,I652885);
DFFARX1 I_21732 (I372504,I3035,I372436,I372530,);
not I_21733 (I372538,I652894);
DFFARX1 I_21734 (I652876,I3035,I372436,I372564,);
not I_21735 (I372572,I372564);
nor I_21736 (I372589,I372572,I372470);
and I_21737 (I372606,I372589,I652894);
nor I_21738 (I372623,I372572,I372538);
nor I_21739 (I372419,I372530,I372623);
DFFARX1 I_21740 (I652873,I3035,I372436,I372663,);
nor I_21741 (I372671,I372663,I372530);
not I_21742 (I372688,I372671);
not I_21743 (I372705,I372663);
nor I_21744 (I372722,I372705,I372606);
DFFARX1 I_21745 (I372722,I3035,I372436,I372422,);
nand I_21746 (I372753,I652891,I652870);
and I_21747 (I372770,I372753,I652888);
DFFARX1 I_21748 (I372770,I3035,I372436,I372796,);
nor I_21749 (I372804,I372796,I372663);
DFFARX1 I_21750 (I372804,I3035,I372436,I372404,);
nand I_21751 (I372835,I372796,I372705);
nand I_21752 (I372413,I372688,I372835);
not I_21753 (I372866,I372796);
nor I_21754 (I372883,I372866,I372606);
DFFARX1 I_21755 (I372883,I3035,I372436,I372425,);
nor I_21756 (I372914,I652879,I652870);
or I_21757 (I372416,I372663,I372914);
nor I_21758 (I372407,I372796,I372914);
or I_21759 (I372410,I372530,I372914);
DFFARX1 I_21760 (I372914,I3035,I372436,I372428,);
not I_21761 (I373014,I3042);
DFFARX1 I_21762 (I69467,I3035,I373014,I373040,);
not I_21763 (I373048,I373040);
nand I_21764 (I373065,I69476,I69485);
and I_21765 (I373082,I373065,I69464);
DFFARX1 I_21766 (I373082,I3035,I373014,I373108,);
not I_21767 (I373116,I69467);
DFFARX1 I_21768 (I69482,I3035,I373014,I373142,);
not I_21769 (I373150,I373142);
nor I_21770 (I373167,I373150,I373048);
and I_21771 (I373184,I373167,I69467);
nor I_21772 (I373201,I373150,I373116);
nor I_21773 (I372997,I373108,I373201);
DFFARX1 I_21774 (I69473,I3035,I373014,I373241,);
nor I_21775 (I373249,I373241,I373108);
not I_21776 (I373266,I373249);
not I_21777 (I373283,I373241);
nor I_21778 (I373300,I373283,I373184);
DFFARX1 I_21779 (I373300,I3035,I373014,I373000,);
nand I_21780 (I373331,I69488,I69464);
and I_21781 (I373348,I373331,I69470);
DFFARX1 I_21782 (I373348,I3035,I373014,I373374,);
nor I_21783 (I373382,I373374,I373241);
DFFARX1 I_21784 (I373382,I3035,I373014,I372982,);
nand I_21785 (I373413,I373374,I373283);
nand I_21786 (I372991,I373266,I373413);
not I_21787 (I373444,I373374);
nor I_21788 (I373461,I373444,I373184);
DFFARX1 I_21789 (I373461,I3035,I373014,I373003,);
nor I_21790 (I373492,I69479,I69464);
or I_21791 (I372994,I373241,I373492);
nor I_21792 (I372985,I373374,I373492);
or I_21793 (I372988,I373108,I373492);
DFFARX1 I_21794 (I373492,I3035,I373014,I373006,);
not I_21795 (I373592,I3042);
DFFARX1 I_21796 (I745445,I3035,I373592,I373618,);
not I_21797 (I373626,I373618);
nand I_21798 (I373643,I745430,I745418);
and I_21799 (I373660,I373643,I745433);
DFFARX1 I_21800 (I373660,I3035,I373592,I373686,);
not I_21801 (I373694,I745418);
DFFARX1 I_21802 (I745436,I3035,I373592,I373720,);
not I_21803 (I373728,I373720);
nor I_21804 (I373745,I373728,I373626);
and I_21805 (I373762,I373745,I745418);
nor I_21806 (I373779,I373728,I373694);
nor I_21807 (I373575,I373686,I373779);
DFFARX1 I_21808 (I745424,I3035,I373592,I373819,);
nor I_21809 (I373827,I373819,I373686);
not I_21810 (I373844,I373827);
not I_21811 (I373861,I373819);
nor I_21812 (I373878,I373861,I373762);
DFFARX1 I_21813 (I373878,I3035,I373592,I373578,);
nand I_21814 (I373909,I745421,I745427);
and I_21815 (I373926,I373909,I745442);
DFFARX1 I_21816 (I373926,I3035,I373592,I373952,);
nor I_21817 (I373960,I373952,I373819);
DFFARX1 I_21818 (I373960,I3035,I373592,I373560,);
nand I_21819 (I373991,I373952,I373861);
nand I_21820 (I373569,I373844,I373991);
not I_21821 (I374022,I373952);
nor I_21822 (I374039,I374022,I373762);
DFFARX1 I_21823 (I374039,I3035,I373592,I373581,);
nor I_21824 (I374070,I745439,I745427);
or I_21825 (I373572,I373819,I374070);
nor I_21826 (I373563,I373952,I374070);
or I_21827 (I373566,I373686,I374070);
DFFARX1 I_21828 (I374070,I3035,I373592,I373584,);
not I_21829 (I374170,I3042);
DFFARX1 I_21830 (I520668,I3035,I374170,I374196,);
not I_21831 (I374204,I374196);
nand I_21832 (I374221,I520644,I520659);
and I_21833 (I374238,I374221,I520671);
DFFARX1 I_21834 (I374238,I3035,I374170,I374264,);
not I_21835 (I374272,I520656);
DFFARX1 I_21836 (I520647,I3035,I374170,I374298,);
not I_21837 (I374306,I374298);
nor I_21838 (I374323,I374306,I374204);
and I_21839 (I374340,I374323,I520656);
nor I_21840 (I374357,I374306,I374272);
nor I_21841 (I374153,I374264,I374357);
DFFARX1 I_21842 (I520644,I3035,I374170,I374397,);
nor I_21843 (I374405,I374397,I374264);
not I_21844 (I374422,I374405);
not I_21845 (I374439,I374397);
nor I_21846 (I374456,I374439,I374340);
DFFARX1 I_21847 (I374456,I3035,I374170,I374156,);
nand I_21848 (I374487,I520662,I520653);
and I_21849 (I374504,I374487,I520665);
DFFARX1 I_21850 (I374504,I3035,I374170,I374530,);
nor I_21851 (I374538,I374530,I374397);
DFFARX1 I_21852 (I374538,I3035,I374170,I374138,);
nand I_21853 (I374569,I374530,I374439);
nand I_21854 (I374147,I374422,I374569);
not I_21855 (I374600,I374530);
nor I_21856 (I374617,I374600,I374340);
DFFARX1 I_21857 (I374617,I3035,I374170,I374159,);
nor I_21858 (I374648,I520650,I520653);
or I_21859 (I374150,I374397,I374648);
nor I_21860 (I374141,I374530,I374648);
or I_21861 (I374144,I374264,I374648);
DFFARX1 I_21862 (I374648,I3035,I374170,I374162,);
not I_21863 (I374748,I3042);
DFFARX1 I_21864 (I294816,I3035,I374748,I374774,);
not I_21865 (I374782,I374774);
nand I_21866 (I374799,I294831,I294816);
and I_21867 (I374816,I374799,I294819);
DFFARX1 I_21868 (I374816,I3035,I374748,I374842,);
not I_21869 (I374850,I294819);
DFFARX1 I_21870 (I294828,I3035,I374748,I374876,);
not I_21871 (I374884,I374876);
nor I_21872 (I374901,I374884,I374782);
and I_21873 (I374918,I374901,I294819);
nor I_21874 (I374935,I374884,I374850);
nor I_21875 (I374731,I374842,I374935);
DFFARX1 I_21876 (I294822,I3035,I374748,I374975,);
nor I_21877 (I374983,I374975,I374842);
not I_21878 (I375000,I374983);
not I_21879 (I375017,I374975);
nor I_21880 (I375034,I375017,I374918);
DFFARX1 I_21881 (I375034,I3035,I374748,I374734,);
nand I_21882 (I375065,I294825,I294834);
and I_21883 (I375082,I375065,I294840);
DFFARX1 I_21884 (I375082,I3035,I374748,I375108,);
nor I_21885 (I375116,I375108,I374975);
DFFARX1 I_21886 (I375116,I3035,I374748,I374716,);
nand I_21887 (I375147,I375108,I375017);
nand I_21888 (I374725,I375000,I375147);
not I_21889 (I375178,I375108);
nor I_21890 (I375195,I375178,I374918);
DFFARX1 I_21891 (I375195,I3035,I374748,I374737,);
nor I_21892 (I375226,I294837,I294834);
or I_21893 (I374728,I374975,I375226);
nor I_21894 (I374719,I375108,I375226);
or I_21895 (I374722,I374842,I375226);
DFFARX1 I_21896 (I375226,I3035,I374748,I374740,);
not I_21897 (I375326,I3042);
DFFARX1 I_21898 (I306512,I3035,I375326,I375352,);
not I_21899 (I375360,I375352);
nand I_21900 (I375377,I306521,I306530);
and I_21901 (I375394,I375377,I306536);
DFFARX1 I_21902 (I375394,I3035,I375326,I375420,);
not I_21903 (I375428,I306533);
DFFARX1 I_21904 (I306518,I3035,I375326,I375454,);
not I_21905 (I375462,I375454);
nor I_21906 (I375479,I375462,I375360);
and I_21907 (I375496,I375479,I306533);
nor I_21908 (I375513,I375462,I375428);
nor I_21909 (I375309,I375420,I375513);
DFFARX1 I_21910 (I306527,I3035,I375326,I375553,);
nor I_21911 (I375561,I375553,I375420);
not I_21912 (I375578,I375561);
not I_21913 (I375595,I375553);
nor I_21914 (I375612,I375595,I375496);
DFFARX1 I_21915 (I375612,I3035,I375326,I375312,);
nand I_21916 (I375643,I306524,I306515);
and I_21917 (I375660,I375643,I306512);
DFFARX1 I_21918 (I375660,I3035,I375326,I375686,);
nor I_21919 (I375694,I375686,I375553);
DFFARX1 I_21920 (I375694,I3035,I375326,I375294,);
nand I_21921 (I375725,I375686,I375595);
nand I_21922 (I375303,I375578,I375725);
not I_21923 (I375756,I375686);
nor I_21924 (I375773,I375756,I375496);
DFFARX1 I_21925 (I375773,I3035,I375326,I375315,);
nor I_21926 (I375804,I306515,I306515);
or I_21927 (I375306,I375553,I375804);
nor I_21928 (I375297,I375686,I375804);
or I_21929 (I375300,I375420,I375804);
DFFARX1 I_21930 (I375804,I3035,I375326,I375318,);
not I_21931 (I375904,I3042);
DFFARX1 I_21932 (I171930,I3035,I375904,I375930,);
not I_21933 (I375938,I375930);
nand I_21934 (I375955,I171933,I171909);
and I_21935 (I375972,I375955,I171906);
DFFARX1 I_21936 (I375972,I3035,I375904,I375998,);
not I_21937 (I376006,I171912);
DFFARX1 I_21938 (I171906,I3035,I375904,I376032,);
not I_21939 (I376040,I376032);
nor I_21940 (I376057,I376040,I375938);
and I_21941 (I376074,I376057,I171912);
nor I_21942 (I376091,I376040,I376006);
nor I_21943 (I375887,I375998,I376091);
DFFARX1 I_21944 (I171915,I3035,I375904,I376131,);
nor I_21945 (I376139,I376131,I375998);
not I_21946 (I376156,I376139);
not I_21947 (I376173,I376131);
nor I_21948 (I376190,I376173,I376074);
DFFARX1 I_21949 (I376190,I3035,I375904,I375890,);
nand I_21950 (I376221,I171918,I171927);
and I_21951 (I376238,I376221,I171924);
DFFARX1 I_21952 (I376238,I3035,I375904,I376264,);
nor I_21953 (I376272,I376264,I376131);
DFFARX1 I_21954 (I376272,I3035,I375904,I375872,);
nand I_21955 (I376303,I376264,I376173);
nand I_21956 (I375881,I376156,I376303);
not I_21957 (I376334,I376264);
nor I_21958 (I376351,I376334,I376074);
DFFARX1 I_21959 (I376351,I3035,I375904,I375893,);
nor I_21960 (I376382,I171921,I171927);
or I_21961 (I375884,I376131,I376382);
nor I_21962 (I375875,I376264,I376382);
or I_21963 (I375878,I375998,I376382);
DFFARX1 I_21964 (I376382,I3035,I375904,I375896,);
not I_21965 (I376482,I3042);
DFFARX1 I_21966 (I112219,I3035,I376482,I376508,);
not I_21967 (I376516,I376508);
nand I_21968 (I376533,I112222,I112243);
and I_21969 (I376550,I376533,I112231);
DFFARX1 I_21970 (I376550,I3035,I376482,I376576,);
not I_21971 (I376584,I112228);
DFFARX1 I_21972 (I112219,I3035,I376482,I376610,);
not I_21973 (I376618,I376610);
nor I_21974 (I376635,I376618,I376516);
and I_21975 (I376652,I376635,I112228);
nor I_21976 (I376669,I376618,I376584);
nor I_21977 (I376465,I376576,I376669);
DFFARX1 I_21978 (I112237,I3035,I376482,I376709,);
nor I_21979 (I376717,I376709,I376576);
not I_21980 (I376734,I376717);
not I_21981 (I376751,I376709);
nor I_21982 (I376768,I376751,I376652);
DFFARX1 I_21983 (I376768,I3035,I376482,I376468,);
nand I_21984 (I376799,I112222,I112225);
and I_21985 (I376816,I376799,I112234);
DFFARX1 I_21986 (I376816,I3035,I376482,I376842,);
nor I_21987 (I376850,I376842,I376709);
DFFARX1 I_21988 (I376850,I3035,I376482,I376450,);
nand I_21989 (I376881,I376842,I376751);
nand I_21990 (I376459,I376734,I376881);
not I_21991 (I376912,I376842);
nor I_21992 (I376929,I376912,I376652);
DFFARX1 I_21993 (I376929,I3035,I376482,I376471,);
nor I_21994 (I376960,I112240,I112225);
or I_21995 (I376462,I376709,I376960);
nor I_21996 (I376453,I376842,I376960);
or I_21997 (I376456,I376576,I376960);
DFFARX1 I_21998 (I376960,I3035,I376482,I376474,);
not I_21999 (I377060,I3042);
DFFARX1 I_22000 (I519376,I3035,I377060,I377086,);
not I_22001 (I377094,I377086);
nand I_22002 (I377111,I519352,I519367);
and I_22003 (I377128,I377111,I519379);
DFFARX1 I_22004 (I377128,I3035,I377060,I377154,);
not I_22005 (I377162,I519364);
DFFARX1 I_22006 (I519355,I3035,I377060,I377188,);
not I_22007 (I377196,I377188);
nor I_22008 (I377213,I377196,I377094);
and I_22009 (I377230,I377213,I519364);
nor I_22010 (I377247,I377196,I377162);
nor I_22011 (I377043,I377154,I377247);
DFFARX1 I_22012 (I519352,I3035,I377060,I377287,);
nor I_22013 (I377295,I377287,I377154);
not I_22014 (I377312,I377295);
not I_22015 (I377329,I377287);
nor I_22016 (I377346,I377329,I377230);
DFFARX1 I_22017 (I377346,I3035,I377060,I377046,);
nand I_22018 (I377377,I519370,I519361);
and I_22019 (I377394,I377377,I519373);
DFFARX1 I_22020 (I377394,I3035,I377060,I377420,);
nor I_22021 (I377428,I377420,I377287);
DFFARX1 I_22022 (I377428,I3035,I377060,I377028,);
nand I_22023 (I377459,I377420,I377329);
nand I_22024 (I377037,I377312,I377459);
not I_22025 (I377490,I377420);
nor I_22026 (I377507,I377490,I377230);
DFFARX1 I_22027 (I377507,I3035,I377060,I377049,);
nor I_22028 (I377538,I519358,I519361);
or I_22029 (I377040,I377287,I377538);
nor I_22030 (I377031,I377420,I377538);
or I_22031 (I377034,I377154,I377538);
DFFARX1 I_22032 (I377538,I3035,I377060,I377052,);
not I_22033 (I377638,I3042);
DFFARX1 I_22034 (I448273,I3035,I377638,I377664,);
not I_22035 (I377672,I377664);
nand I_22036 (I377689,I448261,I448279);
and I_22037 (I377706,I377689,I448276);
DFFARX1 I_22038 (I377706,I3035,I377638,I377732,);
not I_22039 (I377740,I448267);
DFFARX1 I_22040 (I448264,I3035,I377638,I377766,);
not I_22041 (I377774,I377766);
nor I_22042 (I377791,I377774,I377672);
and I_22043 (I377808,I377791,I448267);
nor I_22044 (I377825,I377774,I377740);
nor I_22045 (I377621,I377732,I377825);
DFFARX1 I_22046 (I448258,I3035,I377638,I377865,);
nor I_22047 (I377873,I377865,I377732);
not I_22048 (I377890,I377873);
not I_22049 (I377907,I377865);
nor I_22050 (I377924,I377907,I377808);
DFFARX1 I_22051 (I377924,I3035,I377638,I377624,);
nand I_22052 (I377955,I448258,I448261);
and I_22053 (I377972,I377955,I448264);
DFFARX1 I_22054 (I377972,I3035,I377638,I377998,);
nor I_22055 (I378006,I377998,I377865);
DFFARX1 I_22056 (I378006,I3035,I377638,I377606,);
nand I_22057 (I378037,I377998,I377907);
nand I_22058 (I377615,I377890,I378037);
not I_22059 (I378068,I377998);
nor I_22060 (I378085,I378068,I377808);
DFFARX1 I_22061 (I378085,I3035,I377638,I377627,);
nor I_22062 (I378116,I448270,I448261);
or I_22063 (I377618,I377865,I378116);
nor I_22064 (I377609,I377998,I378116);
or I_22065 (I377612,I377732,I378116);
DFFARX1 I_22066 (I378116,I3035,I377638,I377630,);
not I_22067 (I378216,I3042);
DFFARX1 I_22068 (I627218,I3035,I378216,I378242,);
not I_22069 (I378250,I378242);
nand I_22070 (I378267,I627200,I627212);
and I_22071 (I378284,I378267,I627215);
DFFARX1 I_22072 (I378284,I3035,I378216,I378310,);
not I_22073 (I378318,I627209);
DFFARX1 I_22074 (I627206,I3035,I378216,I378344,);
not I_22075 (I378352,I378344);
nor I_22076 (I378369,I378352,I378250);
and I_22077 (I378386,I378369,I627209);
nor I_22078 (I378403,I378352,I378318);
nor I_22079 (I378199,I378310,I378403);
DFFARX1 I_22080 (I627224,I3035,I378216,I378443,);
nor I_22081 (I378451,I378443,I378310);
not I_22082 (I378468,I378451);
not I_22083 (I378485,I378443);
nor I_22084 (I378502,I378485,I378386);
DFFARX1 I_22085 (I378502,I3035,I378216,I378202,);
nand I_22086 (I378533,I627203,I627203);
and I_22087 (I378550,I378533,I627200);
DFFARX1 I_22088 (I378550,I3035,I378216,I378576,);
nor I_22089 (I378584,I378576,I378443);
DFFARX1 I_22090 (I378584,I3035,I378216,I378184,);
nand I_22091 (I378615,I378576,I378485);
nand I_22092 (I378193,I378468,I378615);
not I_22093 (I378646,I378576);
nor I_22094 (I378663,I378646,I378386);
DFFARX1 I_22095 (I378663,I3035,I378216,I378205,);
nor I_22096 (I378694,I627221,I627203);
or I_22097 (I378196,I378443,I378694);
nor I_22098 (I378187,I378576,I378694);
or I_22099 (I378190,I378310,I378694);
DFFARX1 I_22100 (I378694,I3035,I378216,I378208,);
not I_22101 (I378794,I3042);
DFFARX1 I_22102 (I543924,I3035,I378794,I378820,);
not I_22103 (I378828,I378820);
nand I_22104 (I378845,I543900,I543915);
and I_22105 (I378862,I378845,I543927);
DFFARX1 I_22106 (I378862,I3035,I378794,I378888,);
not I_22107 (I378896,I543912);
DFFARX1 I_22108 (I543903,I3035,I378794,I378922,);
not I_22109 (I378930,I378922);
nor I_22110 (I378947,I378930,I378828);
and I_22111 (I378964,I378947,I543912);
nor I_22112 (I378981,I378930,I378896);
nor I_22113 (I378777,I378888,I378981);
DFFARX1 I_22114 (I543900,I3035,I378794,I379021,);
nor I_22115 (I379029,I379021,I378888);
not I_22116 (I379046,I379029);
not I_22117 (I379063,I379021);
nor I_22118 (I379080,I379063,I378964);
DFFARX1 I_22119 (I379080,I3035,I378794,I378780,);
nand I_22120 (I379111,I543918,I543909);
and I_22121 (I379128,I379111,I543921);
DFFARX1 I_22122 (I379128,I3035,I378794,I379154,);
nor I_22123 (I379162,I379154,I379021);
DFFARX1 I_22124 (I379162,I3035,I378794,I378762,);
nand I_22125 (I379193,I379154,I379063);
nand I_22126 (I378771,I379046,I379193);
not I_22127 (I379224,I379154);
nor I_22128 (I379241,I379224,I378964);
DFFARX1 I_22129 (I379241,I3035,I378794,I378783,);
nor I_22130 (I379272,I543906,I543909);
or I_22131 (I378774,I379021,I379272);
nor I_22132 (I378765,I379154,I379272);
or I_22133 (I378768,I378888,I379272);
DFFARX1 I_22134 (I379272,I3035,I378794,I378786,);
not I_22135 (I379372,I3042);
DFFARX1 I_22136 (I428774,I3035,I379372,I379398,);
not I_22137 (I379406,I379398);
nand I_22138 (I379423,I428762,I428780);
and I_22139 (I379440,I379423,I428777);
DFFARX1 I_22140 (I379440,I3035,I379372,I379466,);
not I_22141 (I379474,I428768);
DFFARX1 I_22142 (I428765,I3035,I379372,I379500,);
not I_22143 (I379508,I379500);
nor I_22144 (I379525,I379508,I379406);
and I_22145 (I379542,I379525,I428768);
nor I_22146 (I379559,I379508,I379474);
nor I_22147 (I379355,I379466,I379559);
DFFARX1 I_22148 (I428759,I3035,I379372,I379599,);
nor I_22149 (I379607,I379599,I379466);
not I_22150 (I379624,I379607);
not I_22151 (I379641,I379599);
nor I_22152 (I379658,I379641,I379542);
DFFARX1 I_22153 (I379658,I3035,I379372,I379358,);
nand I_22154 (I379689,I428759,I428762);
and I_22155 (I379706,I379689,I428765);
DFFARX1 I_22156 (I379706,I3035,I379372,I379732,);
nor I_22157 (I379740,I379732,I379599);
DFFARX1 I_22158 (I379740,I3035,I379372,I379340,);
nand I_22159 (I379771,I379732,I379641);
nand I_22160 (I379349,I379624,I379771);
not I_22161 (I379802,I379732);
nor I_22162 (I379819,I379802,I379542);
DFFARX1 I_22163 (I379819,I3035,I379372,I379361,);
nor I_22164 (I379850,I428771,I428762);
or I_22165 (I379352,I379599,I379850);
nor I_22166 (I379343,I379732,I379850);
or I_22167 (I379346,I379466,I379850);
DFFARX1 I_22168 (I379850,I3035,I379372,I379364,);
not I_22169 (I379950,I3042);
DFFARX1 I_22170 (I247310,I3035,I379950,I379976,);
not I_22171 (I379984,I379976);
nand I_22172 (I380001,I247301,I247319);
and I_22173 (I380018,I380001,I247322);
DFFARX1 I_22174 (I380018,I3035,I379950,I380044,);
not I_22175 (I380052,I247316);
DFFARX1 I_22176 (I247304,I3035,I379950,I380078,);
not I_22177 (I380086,I380078);
nor I_22178 (I380103,I380086,I379984);
and I_22179 (I380120,I380103,I247316);
nor I_22180 (I380137,I380086,I380052);
nor I_22181 (I379933,I380044,I380137);
DFFARX1 I_22182 (I247313,I3035,I379950,I380177,);
nor I_22183 (I380185,I380177,I380044);
not I_22184 (I380202,I380185);
not I_22185 (I380219,I380177);
nor I_22186 (I380236,I380219,I380120);
DFFARX1 I_22187 (I380236,I3035,I379950,I379936,);
nand I_22188 (I380267,I247328,I247325);
and I_22189 (I380284,I380267,I247307);
DFFARX1 I_22190 (I380284,I3035,I379950,I380310,);
nor I_22191 (I380318,I380310,I380177);
DFFARX1 I_22192 (I380318,I3035,I379950,I379918,);
nand I_22193 (I380349,I380310,I380219);
nand I_22194 (I379927,I380202,I380349);
not I_22195 (I380380,I380310);
nor I_22196 (I380397,I380380,I380120);
DFFARX1 I_22197 (I380397,I3035,I379950,I379939,);
nor I_22198 (I380428,I247301,I247325);
or I_22199 (I379930,I380177,I380428);
nor I_22200 (I379921,I380310,I380428);
or I_22201 (I379924,I380044,I380428);
DFFARX1 I_22202 (I380428,I3035,I379950,I379942,);
not I_22203 (I380528,I3042);
DFFARX1 I_22204 (I25208,I3035,I380528,I380554,);
not I_22205 (I380562,I380554);
nand I_22206 (I380579,I25205,I25196);
and I_22207 (I380596,I380579,I25196);
DFFARX1 I_22208 (I380596,I3035,I380528,I380622,);
not I_22209 (I380630,I25199);
DFFARX1 I_22210 (I25214,I3035,I380528,I380656,);
not I_22211 (I380664,I380656);
nor I_22212 (I380681,I380664,I380562);
and I_22213 (I380698,I380681,I25199);
nor I_22214 (I380715,I380664,I380630);
nor I_22215 (I380511,I380622,I380715);
DFFARX1 I_22216 (I25199,I3035,I380528,I380755,);
nor I_22217 (I380763,I380755,I380622);
not I_22218 (I380780,I380763);
not I_22219 (I380797,I380755);
nor I_22220 (I380814,I380797,I380698);
DFFARX1 I_22221 (I380814,I3035,I380528,I380514,);
nand I_22222 (I380845,I25217,I25202);
and I_22223 (I380862,I380845,I25220);
DFFARX1 I_22224 (I380862,I3035,I380528,I380888,);
nor I_22225 (I380896,I380888,I380755);
DFFARX1 I_22226 (I380896,I3035,I380528,I380496,);
nand I_22227 (I380927,I380888,I380797);
nand I_22228 (I380505,I380780,I380927);
not I_22229 (I380958,I380888);
nor I_22230 (I380975,I380958,I380698);
DFFARX1 I_22231 (I380975,I3035,I380528,I380517,);
nor I_22232 (I381006,I25211,I25202);
or I_22233 (I380508,I380755,I381006);
nor I_22234 (I380499,I380888,I381006);
or I_22235 (I380502,I380622,I381006);
DFFARX1 I_22236 (I381006,I3035,I380528,I380520,);
not I_22237 (I381106,I3042);
DFFARX1 I_22238 (I734140,I3035,I381106,I381132,);
not I_22239 (I381140,I381132);
nand I_22240 (I381157,I734125,I734113);
and I_22241 (I381174,I381157,I734128);
DFFARX1 I_22242 (I381174,I3035,I381106,I381200,);
not I_22243 (I381208,I734113);
DFFARX1 I_22244 (I734131,I3035,I381106,I381234,);
not I_22245 (I381242,I381234);
nor I_22246 (I381259,I381242,I381140);
and I_22247 (I381276,I381259,I734113);
nor I_22248 (I381293,I381242,I381208);
nor I_22249 (I381089,I381200,I381293);
DFFARX1 I_22250 (I734119,I3035,I381106,I381333,);
nor I_22251 (I381341,I381333,I381200);
not I_22252 (I381358,I381341);
not I_22253 (I381375,I381333);
nor I_22254 (I381392,I381375,I381276);
DFFARX1 I_22255 (I381392,I3035,I381106,I381092,);
nand I_22256 (I381423,I734116,I734122);
and I_22257 (I381440,I381423,I734137);
DFFARX1 I_22258 (I381440,I3035,I381106,I381466,);
nor I_22259 (I381474,I381466,I381333);
DFFARX1 I_22260 (I381474,I3035,I381106,I381074,);
nand I_22261 (I381505,I381466,I381375);
nand I_22262 (I381083,I381358,I381505);
not I_22263 (I381536,I381466);
nor I_22264 (I381553,I381536,I381276);
DFFARX1 I_22265 (I381553,I3035,I381106,I381095,);
nor I_22266 (I381584,I734134,I734122);
or I_22267 (I381086,I381333,I381584);
nor I_22268 (I381077,I381466,I381584);
or I_22269 (I381080,I381200,I381584);
DFFARX1 I_22270 (I381584,I3035,I381106,I381098,);
not I_22271 (I381684,I3042);
DFFARX1 I_22272 (I48387,I3035,I381684,I381710,);
not I_22273 (I381718,I381710);
nand I_22274 (I381735,I48396,I48405);
and I_22275 (I381752,I381735,I48384);
DFFARX1 I_22276 (I381752,I3035,I381684,I381778,);
not I_22277 (I381786,I48387);
DFFARX1 I_22278 (I48402,I3035,I381684,I381812,);
not I_22279 (I381820,I381812);
nor I_22280 (I381837,I381820,I381718);
and I_22281 (I381854,I381837,I48387);
nor I_22282 (I381871,I381820,I381786);
nor I_22283 (I381667,I381778,I381871);
DFFARX1 I_22284 (I48393,I3035,I381684,I381911,);
nor I_22285 (I381919,I381911,I381778);
not I_22286 (I381936,I381919);
not I_22287 (I381953,I381911);
nor I_22288 (I381970,I381953,I381854);
DFFARX1 I_22289 (I381970,I3035,I381684,I381670,);
nand I_22290 (I382001,I48408,I48384);
and I_22291 (I382018,I382001,I48390);
DFFARX1 I_22292 (I382018,I3035,I381684,I382044,);
nor I_22293 (I382052,I382044,I381911);
DFFARX1 I_22294 (I382052,I3035,I381684,I381652,);
nand I_22295 (I382083,I382044,I381953);
nand I_22296 (I381661,I381936,I382083);
not I_22297 (I382114,I382044);
nor I_22298 (I382131,I382114,I381854);
DFFARX1 I_22299 (I382131,I3035,I381684,I381673,);
nor I_22300 (I382162,I48399,I48384);
or I_22301 (I381664,I381911,I382162);
nor I_22302 (I381655,I382044,I382162);
or I_22303 (I381658,I381778,I382162);
DFFARX1 I_22304 (I382162,I3035,I381684,I381676,);
not I_22305 (I382262,I3042);
DFFARX1 I_22306 (I721050,I3035,I382262,I382288,);
not I_22307 (I382296,I382288);
nand I_22308 (I382313,I721035,I721023);
and I_22309 (I382330,I382313,I721038);
DFFARX1 I_22310 (I382330,I3035,I382262,I382356,);
not I_22311 (I382364,I721023);
DFFARX1 I_22312 (I721041,I3035,I382262,I382390,);
not I_22313 (I382398,I382390);
nor I_22314 (I382415,I382398,I382296);
and I_22315 (I382432,I382415,I721023);
nor I_22316 (I382449,I382398,I382364);
nor I_22317 (I382245,I382356,I382449);
DFFARX1 I_22318 (I721029,I3035,I382262,I382489,);
nor I_22319 (I382497,I382489,I382356);
not I_22320 (I382514,I382497);
not I_22321 (I382531,I382489);
nor I_22322 (I382548,I382531,I382432);
DFFARX1 I_22323 (I382548,I3035,I382262,I382248,);
nand I_22324 (I382579,I721026,I721032);
and I_22325 (I382596,I382579,I721047);
DFFARX1 I_22326 (I382596,I3035,I382262,I382622,);
nor I_22327 (I382630,I382622,I382489);
DFFARX1 I_22328 (I382630,I3035,I382262,I382230,);
nand I_22329 (I382661,I382622,I382531);
nand I_22330 (I382239,I382514,I382661);
not I_22331 (I382692,I382622);
nor I_22332 (I382709,I382692,I382432);
DFFARX1 I_22333 (I382709,I3035,I382262,I382251,);
nor I_22334 (I382740,I721044,I721032);
or I_22335 (I382242,I382489,I382740);
nor I_22336 (I382233,I382622,I382740);
or I_22337 (I382236,I382356,I382740);
DFFARX1 I_22338 (I382740,I3035,I382262,I382254,);
not I_22339 (I382840,I3042);
DFFARX1 I_22340 (I84254,I3035,I382840,I382866,);
not I_22341 (I382874,I382866);
nand I_22342 (I382891,I84257,I84278);
and I_22343 (I382908,I382891,I84266);
DFFARX1 I_22344 (I382908,I3035,I382840,I382934,);
not I_22345 (I382942,I84263);
DFFARX1 I_22346 (I84254,I3035,I382840,I382968,);
not I_22347 (I382976,I382968);
nor I_22348 (I382993,I382976,I382874);
and I_22349 (I383010,I382993,I84263);
nor I_22350 (I383027,I382976,I382942);
nor I_22351 (I382823,I382934,I383027);
DFFARX1 I_22352 (I84272,I3035,I382840,I383067,);
nor I_22353 (I383075,I383067,I382934);
not I_22354 (I383092,I383075);
not I_22355 (I383109,I383067);
nor I_22356 (I383126,I383109,I383010);
DFFARX1 I_22357 (I383126,I3035,I382840,I382826,);
nand I_22358 (I383157,I84257,I84260);
and I_22359 (I383174,I383157,I84269);
DFFARX1 I_22360 (I383174,I3035,I382840,I383200,);
nor I_22361 (I383208,I383200,I383067);
DFFARX1 I_22362 (I383208,I3035,I382840,I382808,);
nand I_22363 (I383239,I383200,I383109);
nand I_22364 (I382817,I383092,I383239);
not I_22365 (I383270,I383200);
nor I_22366 (I383287,I383270,I383010);
DFFARX1 I_22367 (I383287,I3035,I382840,I382829,);
nor I_22368 (I383318,I84275,I84260);
or I_22369 (I382820,I383067,I383318);
nor I_22370 (I382811,I383200,I383318);
or I_22371 (I382814,I382934,I383318);
DFFARX1 I_22372 (I383318,I3035,I382840,I382832,);
not I_22373 (I383418,I3042);
DFFARX1 I_22374 (I224103,I3035,I383418,I383444,);
not I_22375 (I383452,I383444);
nand I_22376 (I383469,I224106,I224082);
and I_22377 (I383486,I383469,I224079);
DFFARX1 I_22378 (I383486,I3035,I383418,I383512,);
not I_22379 (I383520,I224085);
DFFARX1 I_22380 (I224079,I3035,I383418,I383546,);
not I_22381 (I383554,I383546);
nor I_22382 (I383571,I383554,I383452);
and I_22383 (I383588,I383571,I224085);
nor I_22384 (I383605,I383554,I383520);
nor I_22385 (I383401,I383512,I383605);
DFFARX1 I_22386 (I224088,I3035,I383418,I383645,);
nor I_22387 (I383653,I383645,I383512);
not I_22388 (I383670,I383653);
not I_22389 (I383687,I383645);
nor I_22390 (I383704,I383687,I383588);
DFFARX1 I_22391 (I383704,I3035,I383418,I383404,);
nand I_22392 (I383735,I224091,I224100);
and I_22393 (I383752,I383735,I224097);
DFFARX1 I_22394 (I383752,I3035,I383418,I383778,);
nor I_22395 (I383786,I383778,I383645);
DFFARX1 I_22396 (I383786,I3035,I383418,I383386,);
nand I_22397 (I383817,I383778,I383687);
nand I_22398 (I383395,I383670,I383817);
not I_22399 (I383848,I383778);
nor I_22400 (I383865,I383848,I383588);
DFFARX1 I_22401 (I383865,I3035,I383418,I383407,);
nor I_22402 (I383896,I224094,I224100);
or I_22403 (I383398,I383645,I383896);
nor I_22404 (I383389,I383778,I383896);
or I_22405 (I383392,I383512,I383896);
DFFARX1 I_22406 (I383896,I3035,I383418,I383410,);
not I_22407 (I383996,I3042);
DFFARX1 I_22408 (I589070,I3035,I383996,I384022,);
not I_22409 (I384030,I384022);
nand I_22410 (I384047,I589052,I589064);
and I_22411 (I384064,I384047,I589067);
DFFARX1 I_22412 (I384064,I3035,I383996,I384090,);
not I_22413 (I384098,I589061);
DFFARX1 I_22414 (I589058,I3035,I383996,I384124,);
not I_22415 (I384132,I384124);
nor I_22416 (I384149,I384132,I384030);
and I_22417 (I384166,I384149,I589061);
nor I_22418 (I384183,I384132,I384098);
nor I_22419 (I383979,I384090,I384183);
DFFARX1 I_22420 (I589076,I3035,I383996,I384223,);
nor I_22421 (I384231,I384223,I384090);
not I_22422 (I384248,I384231);
not I_22423 (I384265,I384223);
nor I_22424 (I384282,I384265,I384166);
DFFARX1 I_22425 (I384282,I3035,I383996,I383982,);
nand I_22426 (I384313,I589055,I589055);
and I_22427 (I384330,I384313,I589052);
DFFARX1 I_22428 (I384330,I3035,I383996,I384356,);
nor I_22429 (I384364,I384356,I384223);
DFFARX1 I_22430 (I384364,I3035,I383996,I383964,);
nand I_22431 (I384395,I384356,I384265);
nand I_22432 (I383973,I384248,I384395);
not I_22433 (I384426,I384356);
nor I_22434 (I384443,I384426,I384166);
DFFARX1 I_22435 (I384443,I3035,I383996,I383985,);
nor I_22436 (I384474,I589073,I589055);
or I_22437 (I383976,I384223,I384474);
nor I_22438 (I383967,I384356,I384474);
or I_22439 (I383970,I384090,I384474);
DFFARX1 I_22440 (I384474,I3035,I383996,I383988,);
not I_22441 (I384574,I3042);
DFFARX1 I_22442 (I19938,I3035,I384574,I384600,);
not I_22443 (I384608,I384600);
nand I_22444 (I384625,I19935,I19926);
and I_22445 (I384642,I384625,I19926);
DFFARX1 I_22446 (I384642,I3035,I384574,I384668,);
not I_22447 (I384676,I19929);
DFFARX1 I_22448 (I19944,I3035,I384574,I384702,);
not I_22449 (I384710,I384702);
nor I_22450 (I384727,I384710,I384608);
and I_22451 (I384744,I384727,I19929);
nor I_22452 (I384761,I384710,I384676);
nor I_22453 (I384557,I384668,I384761);
DFFARX1 I_22454 (I19929,I3035,I384574,I384801,);
nor I_22455 (I384809,I384801,I384668);
not I_22456 (I384826,I384809);
not I_22457 (I384843,I384801);
nor I_22458 (I384860,I384843,I384744);
DFFARX1 I_22459 (I384860,I3035,I384574,I384560,);
nand I_22460 (I384891,I19947,I19932);
and I_22461 (I384908,I384891,I19950);
DFFARX1 I_22462 (I384908,I3035,I384574,I384934,);
nor I_22463 (I384942,I384934,I384801);
DFFARX1 I_22464 (I384942,I3035,I384574,I384542,);
nand I_22465 (I384973,I384934,I384843);
nand I_22466 (I384551,I384826,I384973);
not I_22467 (I385004,I384934);
nor I_22468 (I385021,I385004,I384744);
DFFARX1 I_22469 (I385021,I3035,I384574,I384563,);
nor I_22470 (I385052,I19941,I19932);
or I_22471 (I384554,I384801,I385052);
nor I_22472 (I384545,I384934,I385052);
or I_22473 (I384548,I384668,I385052);
DFFARX1 I_22474 (I385052,I3035,I384574,I384566,);
not I_22475 (I385152,I3042);
DFFARX1 I_22476 (I318650,I3035,I385152,I385178,);
not I_22477 (I385186,I385178);
nand I_22478 (I385203,I318659,I318668);
and I_22479 (I385220,I385203,I318674);
DFFARX1 I_22480 (I385220,I3035,I385152,I385246,);
not I_22481 (I385254,I318671);
DFFARX1 I_22482 (I318656,I3035,I385152,I385280,);
not I_22483 (I385288,I385280);
nor I_22484 (I385305,I385288,I385186);
and I_22485 (I385322,I385305,I318671);
nor I_22486 (I385339,I385288,I385254);
nor I_22487 (I385135,I385246,I385339);
DFFARX1 I_22488 (I318665,I3035,I385152,I385379,);
nor I_22489 (I385387,I385379,I385246);
not I_22490 (I385404,I385387);
not I_22491 (I385421,I385379);
nor I_22492 (I385438,I385421,I385322);
DFFARX1 I_22493 (I385438,I3035,I385152,I385138,);
nand I_22494 (I385469,I318662,I318653);
and I_22495 (I385486,I385469,I318650);
DFFARX1 I_22496 (I385486,I3035,I385152,I385512,);
nor I_22497 (I385520,I385512,I385379);
DFFARX1 I_22498 (I385520,I3035,I385152,I385120,);
nand I_22499 (I385551,I385512,I385421);
nand I_22500 (I385129,I385404,I385551);
not I_22501 (I385582,I385512);
nor I_22502 (I385599,I385582,I385322);
DFFARX1 I_22503 (I385599,I3035,I385152,I385141,);
nor I_22504 (I385630,I318653,I318653);
or I_22505 (I385132,I385379,I385630);
nor I_22506 (I385123,I385512,I385630);
or I_22507 (I385126,I385246,I385630);
DFFARX1 I_22508 (I385630,I3035,I385152,I385144,);
not I_22509 (I385730,I3042);
DFFARX1 I_22510 (I2116,I3035,I385730,I385756,);
not I_22511 (I385764,I385756);
nand I_22512 (I385781,I1428,I2012);
and I_22513 (I385798,I385781,I2076);
DFFARX1 I_22514 (I385798,I3035,I385730,I385824,);
not I_22515 (I385832,I1684);
DFFARX1 I_22516 (I2188,I3035,I385730,I385858,);
not I_22517 (I385866,I385858);
nor I_22518 (I385883,I385866,I385764);
and I_22519 (I385900,I385883,I1684);
nor I_22520 (I385917,I385866,I385832);
nor I_22521 (I385713,I385824,I385917);
DFFARX1 I_22522 (I1820,I3035,I385730,I385957,);
nor I_22523 (I385965,I385957,I385824);
not I_22524 (I385982,I385965);
not I_22525 (I385999,I385957);
nor I_22526 (I386016,I385999,I385900);
DFFARX1 I_22527 (I386016,I3035,I385730,I385716,);
nand I_22528 (I386047,I2988,I2140);
and I_22529 (I386064,I386047,I1564);
DFFARX1 I_22530 (I386064,I3035,I385730,I386090,);
nor I_22531 (I386098,I386090,I385957);
DFFARX1 I_22532 (I386098,I3035,I385730,I385698,);
nand I_22533 (I386129,I386090,I385999);
nand I_22534 (I385707,I385982,I386129);
not I_22535 (I386160,I386090);
nor I_22536 (I386177,I386160,I385900);
DFFARX1 I_22537 (I386177,I3035,I385730,I385719,);
nor I_22538 (I386208,I1972,I2140);
or I_22539 (I385710,I385957,I386208);
nor I_22540 (I385701,I386090,I386208);
or I_22541 (I385704,I385824,I386208);
DFFARX1 I_22542 (I386208,I3035,I385730,I385722,);
not I_22543 (I386308,I3042);
DFFARX1 I_22544 (I29415,I3035,I386308,I386334,);
not I_22545 (I386342,I386334);
nand I_22546 (I386359,I29424,I29433);
and I_22547 (I386376,I386359,I29412);
DFFARX1 I_22548 (I386376,I3035,I386308,I386402,);
not I_22549 (I386410,I29415);
DFFARX1 I_22550 (I29430,I3035,I386308,I386436,);
not I_22551 (I386444,I386436);
nor I_22552 (I386461,I386444,I386342);
and I_22553 (I386478,I386461,I29415);
nor I_22554 (I386495,I386444,I386410);
nor I_22555 (I386291,I386402,I386495);
DFFARX1 I_22556 (I29421,I3035,I386308,I386535,);
nor I_22557 (I386543,I386535,I386402);
not I_22558 (I386560,I386543);
not I_22559 (I386577,I386535);
nor I_22560 (I386594,I386577,I386478);
DFFARX1 I_22561 (I386594,I3035,I386308,I386294,);
nand I_22562 (I386625,I29436,I29412);
and I_22563 (I386642,I386625,I29418);
DFFARX1 I_22564 (I386642,I3035,I386308,I386668,);
nor I_22565 (I386676,I386668,I386535);
DFFARX1 I_22566 (I386676,I3035,I386308,I386276,);
nand I_22567 (I386707,I386668,I386577);
nand I_22568 (I386285,I386560,I386707);
not I_22569 (I386738,I386668);
nor I_22570 (I386755,I386738,I386478);
DFFARX1 I_22571 (I386755,I3035,I386308,I386297,);
nor I_22572 (I386786,I29427,I29412);
or I_22573 (I386288,I386535,I386786);
nor I_22574 (I386279,I386668,I386786);
or I_22575 (I386282,I386402,I386786);
DFFARX1 I_22576 (I386786,I3035,I386308,I386300,);
not I_22577 (I386886,I3042);
DFFARX1 I_22578 (I36793,I3035,I386886,I386912,);
not I_22579 (I386920,I386912);
nand I_22580 (I386937,I36802,I36811);
and I_22581 (I386954,I386937,I36790);
DFFARX1 I_22582 (I386954,I3035,I386886,I386980,);
not I_22583 (I386988,I36793);
DFFARX1 I_22584 (I36808,I3035,I386886,I387014,);
not I_22585 (I387022,I387014);
nor I_22586 (I387039,I387022,I386920);
and I_22587 (I387056,I387039,I36793);
nor I_22588 (I387073,I387022,I386988);
nor I_22589 (I386869,I386980,I387073);
DFFARX1 I_22590 (I36799,I3035,I386886,I387113,);
nor I_22591 (I387121,I387113,I386980);
not I_22592 (I387138,I387121);
not I_22593 (I387155,I387113);
nor I_22594 (I387172,I387155,I387056);
DFFARX1 I_22595 (I387172,I3035,I386886,I386872,);
nand I_22596 (I387203,I36814,I36790);
and I_22597 (I387220,I387203,I36796);
DFFARX1 I_22598 (I387220,I3035,I386886,I387246,);
nor I_22599 (I387254,I387246,I387113);
DFFARX1 I_22600 (I387254,I3035,I386886,I386854,);
nand I_22601 (I387285,I387246,I387155);
nand I_22602 (I386863,I387138,I387285);
not I_22603 (I387316,I387246);
nor I_22604 (I387333,I387316,I387056);
DFFARX1 I_22605 (I387333,I3035,I386886,I386875,);
nor I_22606 (I387364,I36805,I36790);
or I_22607 (I386866,I387113,I387364);
nor I_22608 (I386857,I387246,I387364);
or I_22609 (I386860,I386980,I387364);
DFFARX1 I_22610 (I387364,I3035,I386886,I386878,);
not I_22611 (I387464,I3042);
DFFARX1 I_22612 (I234254,I3035,I387464,I387490,);
not I_22613 (I387498,I387490);
nand I_22614 (I387515,I234245,I234263);
and I_22615 (I387532,I387515,I234266);
DFFARX1 I_22616 (I387532,I3035,I387464,I387558,);
not I_22617 (I387566,I234260);
DFFARX1 I_22618 (I234248,I3035,I387464,I387592,);
not I_22619 (I387600,I387592);
nor I_22620 (I387617,I387600,I387498);
and I_22621 (I387634,I387617,I234260);
nor I_22622 (I387651,I387600,I387566);
nor I_22623 (I387447,I387558,I387651);
DFFARX1 I_22624 (I234257,I3035,I387464,I387691,);
nor I_22625 (I387699,I387691,I387558);
not I_22626 (I387716,I387699);
not I_22627 (I387733,I387691);
nor I_22628 (I387750,I387733,I387634);
DFFARX1 I_22629 (I387750,I3035,I387464,I387450,);
nand I_22630 (I387781,I234272,I234269);
and I_22631 (I387798,I387781,I234251);
DFFARX1 I_22632 (I387798,I3035,I387464,I387824,);
nor I_22633 (I387832,I387824,I387691);
DFFARX1 I_22634 (I387832,I3035,I387464,I387432,);
nand I_22635 (I387863,I387824,I387733);
nand I_22636 (I387441,I387716,I387863);
not I_22637 (I387894,I387824);
nor I_22638 (I387911,I387894,I387634);
DFFARX1 I_22639 (I387911,I3035,I387464,I387453,);
nor I_22640 (I387942,I234245,I234269);
or I_22641 (I387444,I387691,I387942);
nor I_22642 (I387435,I387824,I387942);
or I_22643 (I387438,I387558,I387942);
DFFARX1 I_22644 (I387942,I3035,I387464,I387456,);
not I_22645 (I388042,I3042);
DFFARX1 I_22646 (I63670,I3035,I388042,I388068,);
not I_22647 (I388076,I388068);
nand I_22648 (I388093,I63679,I63688);
and I_22649 (I388110,I388093,I63667);
DFFARX1 I_22650 (I388110,I3035,I388042,I388136,);
not I_22651 (I388144,I63670);
DFFARX1 I_22652 (I63685,I3035,I388042,I388170,);
not I_22653 (I388178,I388170);
nor I_22654 (I388195,I388178,I388076);
and I_22655 (I388212,I388195,I63670);
nor I_22656 (I388229,I388178,I388144);
nor I_22657 (I388025,I388136,I388229);
DFFARX1 I_22658 (I63676,I3035,I388042,I388269,);
nor I_22659 (I388277,I388269,I388136);
not I_22660 (I388294,I388277);
not I_22661 (I388311,I388269);
nor I_22662 (I388328,I388311,I388212);
DFFARX1 I_22663 (I388328,I3035,I388042,I388028,);
nand I_22664 (I388359,I63691,I63667);
and I_22665 (I388376,I388359,I63673);
DFFARX1 I_22666 (I388376,I3035,I388042,I388402,);
nor I_22667 (I388410,I388402,I388269);
DFFARX1 I_22668 (I388410,I3035,I388042,I388010,);
nand I_22669 (I388441,I388402,I388311);
nand I_22670 (I388019,I388294,I388441);
not I_22671 (I388472,I388402);
nor I_22672 (I388489,I388472,I388212);
DFFARX1 I_22673 (I388489,I3035,I388042,I388031,);
nor I_22674 (I388520,I63682,I63667);
or I_22675 (I388022,I388269,I388520);
nor I_22676 (I388013,I388402,I388520);
or I_22677 (I388016,I388136,I388520);
DFFARX1 I_22678 (I388520,I3035,I388042,I388034,);
not I_22679 (I388620,I3042);
DFFARX1 I_22680 (I715695,I3035,I388620,I388646,);
not I_22681 (I388654,I388646);
nand I_22682 (I388671,I715680,I715668);
and I_22683 (I388688,I388671,I715683);
DFFARX1 I_22684 (I388688,I3035,I388620,I388714,);
not I_22685 (I388722,I715668);
DFFARX1 I_22686 (I715686,I3035,I388620,I388748,);
not I_22687 (I388756,I388748);
nor I_22688 (I388773,I388756,I388654);
and I_22689 (I388790,I388773,I715668);
nor I_22690 (I388807,I388756,I388722);
nor I_22691 (I388603,I388714,I388807);
DFFARX1 I_22692 (I715674,I3035,I388620,I388847,);
nor I_22693 (I388855,I388847,I388714);
not I_22694 (I388872,I388855);
not I_22695 (I388889,I388847);
nor I_22696 (I388906,I388889,I388790);
DFFARX1 I_22697 (I388906,I3035,I388620,I388606,);
nand I_22698 (I388937,I715671,I715677);
and I_22699 (I388954,I388937,I715692);
DFFARX1 I_22700 (I388954,I3035,I388620,I388980,);
nor I_22701 (I388988,I388980,I388847);
DFFARX1 I_22702 (I388988,I3035,I388620,I388588,);
nand I_22703 (I389019,I388980,I388889);
nand I_22704 (I388597,I388872,I389019);
not I_22705 (I389050,I388980);
nor I_22706 (I389067,I389050,I388790);
DFFARX1 I_22707 (I389067,I3035,I388620,I388609,);
nor I_22708 (I389098,I715689,I715677);
or I_22709 (I388600,I388847,I389098);
nor I_22710 (I388591,I388980,I389098);
or I_22711 (I388594,I388714,I389098);
DFFARX1 I_22712 (I389098,I3035,I388620,I388612,);
not I_22713 (I389198,I3042);
DFFARX1 I_22714 (I214617,I3035,I389198,I389224,);
not I_22715 (I389232,I389224);
nand I_22716 (I389249,I214620,I214596);
and I_22717 (I389266,I389249,I214593);
DFFARX1 I_22718 (I389266,I3035,I389198,I389292,);
not I_22719 (I389300,I214599);
DFFARX1 I_22720 (I214593,I3035,I389198,I389326,);
not I_22721 (I389334,I389326);
nor I_22722 (I389351,I389334,I389232);
and I_22723 (I389368,I389351,I214599);
nor I_22724 (I389385,I389334,I389300);
nor I_22725 (I389181,I389292,I389385);
DFFARX1 I_22726 (I214602,I3035,I389198,I389425,);
nor I_22727 (I389433,I389425,I389292);
not I_22728 (I389450,I389433);
not I_22729 (I389467,I389425);
nor I_22730 (I389484,I389467,I389368);
DFFARX1 I_22731 (I389484,I3035,I389198,I389184,);
nand I_22732 (I389515,I214605,I214614);
and I_22733 (I389532,I389515,I214611);
DFFARX1 I_22734 (I389532,I3035,I389198,I389558,);
nor I_22735 (I389566,I389558,I389425);
DFFARX1 I_22736 (I389566,I3035,I389198,I389166,);
nand I_22737 (I389597,I389558,I389467);
nand I_22738 (I389175,I389450,I389597);
not I_22739 (I389628,I389558);
nor I_22740 (I389645,I389628,I389368);
DFFARX1 I_22741 (I389645,I3035,I389198,I389187,);
nor I_22742 (I389676,I214608,I214614);
or I_22743 (I389178,I389425,I389676);
nor I_22744 (I389169,I389558,I389676);
or I_22745 (I389172,I389292,I389676);
DFFARX1 I_22746 (I389676,I3035,I389198,I389190,);
not I_22747 (I389776,I3042);
DFFARX1 I_22748 (I209347,I3035,I389776,I389802,);
not I_22749 (I389810,I389802);
nand I_22750 (I389827,I209350,I209326);
and I_22751 (I389844,I389827,I209323);
DFFARX1 I_22752 (I389844,I3035,I389776,I389870,);
not I_22753 (I389878,I209329);
DFFARX1 I_22754 (I209323,I3035,I389776,I389904,);
not I_22755 (I389912,I389904);
nor I_22756 (I389929,I389912,I389810);
and I_22757 (I389946,I389929,I209329);
nor I_22758 (I389963,I389912,I389878);
nor I_22759 (I389759,I389870,I389963);
DFFARX1 I_22760 (I209332,I3035,I389776,I390003,);
nor I_22761 (I390011,I390003,I389870);
not I_22762 (I390028,I390011);
not I_22763 (I390045,I390003);
nor I_22764 (I390062,I390045,I389946);
DFFARX1 I_22765 (I390062,I3035,I389776,I389762,);
nand I_22766 (I390093,I209335,I209344);
and I_22767 (I390110,I390093,I209341);
DFFARX1 I_22768 (I390110,I3035,I389776,I390136,);
nor I_22769 (I390144,I390136,I390003);
DFFARX1 I_22770 (I390144,I3035,I389776,I389744,);
nand I_22771 (I390175,I390136,I390045);
nand I_22772 (I389753,I390028,I390175);
not I_22773 (I390206,I390136);
nor I_22774 (I390223,I390206,I389946);
DFFARX1 I_22775 (I390223,I3035,I389776,I389765,);
nor I_22776 (I390254,I209338,I209344);
or I_22777 (I389756,I390003,I390254);
nor I_22778 (I389747,I390136,I390254);
or I_22779 (I389750,I389870,I390254);
DFFARX1 I_22780 (I390254,I3035,I389776,I389768,);
not I_22781 (I390354,I3042);
DFFARX1 I_22782 (I264174,I3035,I390354,I390380,);
not I_22783 (I390388,I390380);
nand I_22784 (I390405,I264165,I264183);
and I_22785 (I390422,I390405,I264186);
DFFARX1 I_22786 (I390422,I3035,I390354,I390448,);
not I_22787 (I390456,I264180);
DFFARX1 I_22788 (I264168,I3035,I390354,I390482,);
not I_22789 (I390490,I390482);
nor I_22790 (I390507,I390490,I390388);
and I_22791 (I390524,I390507,I264180);
nor I_22792 (I390541,I390490,I390456);
nor I_22793 (I390337,I390448,I390541);
DFFARX1 I_22794 (I264177,I3035,I390354,I390581,);
nor I_22795 (I390589,I390581,I390448);
not I_22796 (I390606,I390589);
not I_22797 (I390623,I390581);
nor I_22798 (I390640,I390623,I390524);
DFFARX1 I_22799 (I390640,I3035,I390354,I390340,);
nand I_22800 (I390671,I264192,I264189);
and I_22801 (I390688,I390671,I264171);
DFFARX1 I_22802 (I390688,I3035,I390354,I390714,);
nor I_22803 (I390722,I390714,I390581);
DFFARX1 I_22804 (I390722,I3035,I390354,I390322,);
nand I_22805 (I390753,I390714,I390623);
nand I_22806 (I390331,I390606,I390753);
not I_22807 (I390784,I390714);
nor I_22808 (I390801,I390784,I390524);
DFFARX1 I_22809 (I390801,I3035,I390354,I390343,);
nor I_22810 (I390832,I264165,I264189);
or I_22811 (I390334,I390581,I390832);
nor I_22812 (I390325,I390714,I390832);
or I_22813 (I390328,I390448,I390832);
DFFARX1 I_22814 (I390832,I3035,I390354,I390346,);
not I_22815 (I390932,I3042);
DFFARX1 I_22816 (I58927,I3035,I390932,I390958,);
not I_22817 (I390966,I390958);
nand I_22818 (I390983,I58936,I58945);
and I_22819 (I391000,I390983,I58924);
DFFARX1 I_22820 (I391000,I3035,I390932,I391026,);
not I_22821 (I391034,I58927);
DFFARX1 I_22822 (I58942,I3035,I390932,I391060,);
not I_22823 (I391068,I391060);
nor I_22824 (I391085,I391068,I390966);
and I_22825 (I391102,I391085,I58927);
nor I_22826 (I391119,I391068,I391034);
nor I_22827 (I390915,I391026,I391119);
DFFARX1 I_22828 (I58933,I3035,I390932,I391159,);
nor I_22829 (I391167,I391159,I391026);
not I_22830 (I391184,I391167);
not I_22831 (I391201,I391159);
nor I_22832 (I391218,I391201,I391102);
DFFARX1 I_22833 (I391218,I3035,I390932,I390918,);
nand I_22834 (I391249,I58948,I58924);
and I_22835 (I391266,I391249,I58930);
DFFARX1 I_22836 (I391266,I3035,I390932,I391292,);
nor I_22837 (I391300,I391292,I391159);
DFFARX1 I_22838 (I391300,I3035,I390932,I390900,);
nand I_22839 (I391331,I391292,I391201);
nand I_22840 (I390909,I391184,I391331);
not I_22841 (I391362,I391292);
nor I_22842 (I391379,I391362,I391102);
DFFARX1 I_22843 (I391379,I3035,I390932,I390921,);
nor I_22844 (I391410,I58939,I58924);
or I_22845 (I390912,I391159,I391410);
nor I_22846 (I390903,I391292,I391410);
or I_22847 (I390906,I391026,I391410);
DFFARX1 I_22848 (I391410,I3035,I390932,I390924,);
not I_22849 (I391510,I3042);
DFFARX1 I_22850 (I66832,I3035,I391510,I391536,);
not I_22851 (I391544,I391536);
nand I_22852 (I391561,I66841,I66850);
and I_22853 (I391578,I391561,I66829);
DFFARX1 I_22854 (I391578,I3035,I391510,I391604,);
not I_22855 (I391612,I66832);
DFFARX1 I_22856 (I66847,I3035,I391510,I391638,);
not I_22857 (I391646,I391638);
nor I_22858 (I391663,I391646,I391544);
and I_22859 (I391680,I391663,I66832);
nor I_22860 (I391697,I391646,I391612);
nor I_22861 (I391493,I391604,I391697);
DFFARX1 I_22862 (I66838,I3035,I391510,I391737,);
nor I_22863 (I391745,I391737,I391604);
not I_22864 (I391762,I391745);
not I_22865 (I391779,I391737);
nor I_22866 (I391796,I391779,I391680);
DFFARX1 I_22867 (I391796,I3035,I391510,I391496,);
nand I_22868 (I391827,I66853,I66829);
and I_22869 (I391844,I391827,I66835);
DFFARX1 I_22870 (I391844,I3035,I391510,I391870,);
nor I_22871 (I391878,I391870,I391737);
DFFARX1 I_22872 (I391878,I3035,I391510,I391478,);
nand I_22873 (I391909,I391870,I391779);
nand I_22874 (I391487,I391762,I391909);
not I_22875 (I391940,I391870);
nor I_22876 (I391957,I391940,I391680);
DFFARX1 I_22877 (I391957,I3035,I391510,I391499,);
nor I_22878 (I391988,I66844,I66829);
or I_22879 (I391490,I391737,I391988);
nor I_22880 (I391481,I391870,I391988);
or I_22881 (I391484,I391604,I391988);
DFFARX1 I_22882 (I391988,I3035,I391510,I391502,);
not I_22883 (I392088,I3042);
DFFARX1 I_22884 (I181943,I3035,I392088,I392114,);
not I_22885 (I392122,I392114);
nand I_22886 (I392139,I181946,I181922);
and I_22887 (I392156,I392139,I181919);
DFFARX1 I_22888 (I392156,I3035,I392088,I392182,);
not I_22889 (I392190,I181925);
DFFARX1 I_22890 (I181919,I3035,I392088,I392216,);
not I_22891 (I392224,I392216);
nor I_22892 (I392241,I392224,I392122);
and I_22893 (I392258,I392241,I181925);
nor I_22894 (I392275,I392224,I392190);
nor I_22895 (I392071,I392182,I392275);
DFFARX1 I_22896 (I181928,I3035,I392088,I392315,);
nor I_22897 (I392323,I392315,I392182);
not I_22898 (I392340,I392323);
not I_22899 (I392357,I392315);
nor I_22900 (I392374,I392357,I392258);
DFFARX1 I_22901 (I392374,I3035,I392088,I392074,);
nand I_22902 (I392405,I181931,I181940);
and I_22903 (I392422,I392405,I181937);
DFFARX1 I_22904 (I392422,I3035,I392088,I392448,);
nor I_22905 (I392456,I392448,I392315);
DFFARX1 I_22906 (I392456,I3035,I392088,I392056,);
nand I_22907 (I392487,I392448,I392357);
nand I_22908 (I392065,I392340,I392487);
not I_22909 (I392518,I392448);
nor I_22910 (I392535,I392518,I392258);
DFFARX1 I_22911 (I392535,I3035,I392088,I392077,);
nor I_22912 (I392566,I181934,I181940);
or I_22913 (I392068,I392315,I392566);
nor I_22914 (I392059,I392448,I392566);
or I_22915 (I392062,I392182,I392566);
DFFARX1 I_22916 (I392566,I3035,I392088,I392080,);
not I_22917 (I392666,I3042);
DFFARX1 I_22918 (I242414,I3035,I392666,I392692,);
not I_22919 (I392700,I392692);
nand I_22920 (I392717,I242405,I242423);
and I_22921 (I392734,I392717,I242426);
DFFARX1 I_22922 (I392734,I3035,I392666,I392760,);
not I_22923 (I392768,I242420);
DFFARX1 I_22924 (I242408,I3035,I392666,I392794,);
not I_22925 (I392802,I392794);
nor I_22926 (I392819,I392802,I392700);
and I_22927 (I392836,I392819,I242420);
nor I_22928 (I392853,I392802,I392768);
nor I_22929 (I392649,I392760,I392853);
DFFARX1 I_22930 (I242417,I3035,I392666,I392893,);
nor I_22931 (I392901,I392893,I392760);
not I_22932 (I392918,I392901);
not I_22933 (I392935,I392893);
nor I_22934 (I392952,I392935,I392836);
DFFARX1 I_22935 (I392952,I3035,I392666,I392652,);
nand I_22936 (I392983,I242432,I242429);
and I_22937 (I393000,I392983,I242411);
DFFARX1 I_22938 (I393000,I3035,I392666,I393026,);
nor I_22939 (I393034,I393026,I392893);
DFFARX1 I_22940 (I393034,I3035,I392666,I392634,);
nand I_22941 (I393065,I393026,I392935);
nand I_22942 (I392643,I392918,I393065);
not I_22943 (I393096,I393026);
nor I_22944 (I393113,I393096,I392836);
DFFARX1 I_22945 (I393113,I3035,I392666,I392655,);
nor I_22946 (I393144,I242405,I242429);
or I_22947 (I392646,I392893,I393144);
nor I_22948 (I392637,I393026,I393144);
or I_22949 (I392640,I392760,I393144);
DFFARX1 I_22950 (I393144,I3035,I392666,I392658,);
not I_22951 (I393244,I3042);
DFFARX1 I_22952 (I475150,I3035,I393244,I393270,);
not I_22953 (I393278,I393270);
nand I_22954 (I393295,I475138,I475156);
and I_22955 (I393312,I393295,I475153);
DFFARX1 I_22956 (I393312,I3035,I393244,I393338,);
not I_22957 (I393346,I475144);
DFFARX1 I_22958 (I475141,I3035,I393244,I393372,);
not I_22959 (I393380,I393372);
nor I_22960 (I393397,I393380,I393278);
and I_22961 (I393414,I393397,I475144);
nor I_22962 (I393431,I393380,I393346);
nor I_22963 (I393227,I393338,I393431);
DFFARX1 I_22964 (I475135,I3035,I393244,I393471,);
nor I_22965 (I393479,I393471,I393338);
not I_22966 (I393496,I393479);
not I_22967 (I393513,I393471);
nor I_22968 (I393530,I393513,I393414);
DFFARX1 I_22969 (I393530,I3035,I393244,I393230,);
nand I_22970 (I393561,I475135,I475138);
and I_22971 (I393578,I393561,I475141);
DFFARX1 I_22972 (I393578,I3035,I393244,I393604,);
nor I_22973 (I393612,I393604,I393471);
DFFARX1 I_22974 (I393612,I3035,I393244,I393212,);
nand I_22975 (I393643,I393604,I393513);
nand I_22976 (I393221,I393496,I393643);
not I_22977 (I393674,I393604);
nor I_22978 (I393691,I393674,I393414);
DFFARX1 I_22979 (I393691,I3035,I393244,I393233,);
nor I_22980 (I393722,I475147,I475138);
or I_22981 (I393224,I393471,I393722);
nor I_22982 (I393215,I393604,I393722);
or I_22983 (I393218,I393338,I393722);
DFFARX1 I_22984 (I393722,I3035,I393244,I393236,);
not I_22985 (I393822,I3042);
DFFARX1 I_22986 (I290651,I3035,I393822,I393848,);
not I_22987 (I393856,I393848);
nand I_22988 (I393873,I290666,I290651);
and I_22989 (I393890,I393873,I290654);
DFFARX1 I_22990 (I393890,I3035,I393822,I393916,);
not I_22991 (I393924,I290654);
DFFARX1 I_22992 (I290663,I3035,I393822,I393950,);
not I_22993 (I393958,I393950);
nor I_22994 (I393975,I393958,I393856);
and I_22995 (I393992,I393975,I290654);
nor I_22996 (I394009,I393958,I393924);
nor I_22997 (I393805,I393916,I394009);
DFFARX1 I_22998 (I290657,I3035,I393822,I394049,);
nor I_22999 (I394057,I394049,I393916);
not I_23000 (I394074,I394057);
not I_23001 (I394091,I394049);
nor I_23002 (I394108,I394091,I393992);
DFFARX1 I_23003 (I394108,I3035,I393822,I393808,);
nand I_23004 (I394139,I290660,I290669);
and I_23005 (I394156,I394139,I290675);
DFFARX1 I_23006 (I394156,I3035,I393822,I394182,);
nor I_23007 (I394190,I394182,I394049);
DFFARX1 I_23008 (I394190,I3035,I393822,I393790,);
nand I_23009 (I394221,I394182,I394091);
nand I_23010 (I393799,I394074,I394221);
not I_23011 (I394252,I394182);
nor I_23012 (I394269,I394252,I393992);
DFFARX1 I_23013 (I394269,I3035,I393822,I393811,);
nor I_23014 (I394300,I290672,I290669);
or I_23015 (I393802,I394049,I394300);
nor I_23016 (I393793,I394182,I394300);
or I_23017 (I393796,I393916,I394300);
DFFARX1 I_23018 (I394300,I3035,I393822,I393814,);
not I_23019 (I394400,I3042);
DFFARX1 I_23020 (I555466,I3035,I394400,I394426,);
not I_23021 (I394434,I394426);
nand I_23022 (I394451,I555463,I555481);
and I_23023 (I394468,I394451,I555478);
DFFARX1 I_23024 (I394468,I3035,I394400,I394494,);
not I_23025 (I394502,I555460);
DFFARX1 I_23026 (I555463,I3035,I394400,I394528,);
not I_23027 (I394536,I394528);
nor I_23028 (I394553,I394536,I394434);
and I_23029 (I394570,I394553,I555460);
nor I_23030 (I394587,I394536,I394502);
nor I_23031 (I394383,I394494,I394587);
DFFARX1 I_23032 (I555472,I3035,I394400,I394627,);
nor I_23033 (I394635,I394627,I394494);
not I_23034 (I394652,I394635);
not I_23035 (I394669,I394627);
nor I_23036 (I394686,I394669,I394570);
DFFARX1 I_23037 (I394686,I3035,I394400,I394386,);
nand I_23038 (I394717,I555475,I555460);
and I_23039 (I394734,I394717,I555466);
DFFARX1 I_23040 (I394734,I3035,I394400,I394760,);
nor I_23041 (I394768,I394760,I394627);
DFFARX1 I_23042 (I394768,I3035,I394400,I394368,);
nand I_23043 (I394799,I394760,I394669);
nand I_23044 (I394377,I394652,I394799);
not I_23045 (I394830,I394760);
nor I_23046 (I394847,I394830,I394570);
DFFARX1 I_23047 (I394847,I3035,I394400,I394389,);
nor I_23048 (I394878,I555469,I555460);
or I_23049 (I394380,I394627,I394878);
nor I_23050 (I394371,I394760,I394878);
or I_23051 (I394374,I394494,I394878);
DFFARX1 I_23052 (I394878,I3035,I394400,I394392,);
not I_23053 (I394978,I3042);
DFFARX1 I_23054 (I44698,I3035,I394978,I395004,);
not I_23055 (I395012,I395004);
nand I_23056 (I395029,I44707,I44716);
and I_23057 (I395046,I395029,I44695);
DFFARX1 I_23058 (I395046,I3035,I394978,I395072,);
not I_23059 (I395080,I44698);
DFFARX1 I_23060 (I44713,I3035,I394978,I395106,);
not I_23061 (I395114,I395106);
nor I_23062 (I395131,I395114,I395012);
and I_23063 (I395148,I395131,I44698);
nor I_23064 (I395165,I395114,I395080);
nor I_23065 (I394961,I395072,I395165);
DFFARX1 I_23066 (I44704,I3035,I394978,I395205,);
nor I_23067 (I395213,I395205,I395072);
not I_23068 (I395230,I395213);
not I_23069 (I395247,I395205);
nor I_23070 (I395264,I395247,I395148);
DFFARX1 I_23071 (I395264,I3035,I394978,I394964,);
nand I_23072 (I395295,I44719,I44695);
and I_23073 (I395312,I395295,I44701);
DFFARX1 I_23074 (I395312,I3035,I394978,I395338,);
nor I_23075 (I395346,I395338,I395205);
DFFARX1 I_23076 (I395346,I3035,I394978,I394946,);
nand I_23077 (I395377,I395338,I395247);
nand I_23078 (I394955,I395230,I395377);
not I_23079 (I395408,I395338);
nor I_23080 (I395425,I395408,I395148);
DFFARX1 I_23081 (I395425,I3035,I394978,I394967,);
nor I_23082 (I395456,I44710,I44695);
or I_23083 (I394958,I395205,I395456);
nor I_23084 (I394949,I395338,I395456);
or I_23085 (I394952,I395072,I395456);
DFFARX1 I_23086 (I395456,I3035,I394978,I394970,);
not I_23087 (I395556,I3042);
DFFARX1 I_23088 (I135424,I3035,I395556,I395582,);
not I_23089 (I395590,I395582);
nand I_23090 (I395607,I135427,I135448);
and I_23091 (I395624,I395607,I135436);
DFFARX1 I_23092 (I395624,I3035,I395556,I395650,);
not I_23093 (I395658,I135433);
DFFARX1 I_23094 (I135424,I3035,I395556,I395684,);
not I_23095 (I395692,I395684);
nor I_23096 (I395709,I395692,I395590);
and I_23097 (I395726,I395709,I135433);
nor I_23098 (I395743,I395692,I395658);
nor I_23099 (I395539,I395650,I395743);
DFFARX1 I_23100 (I135442,I3035,I395556,I395783,);
nor I_23101 (I395791,I395783,I395650);
not I_23102 (I395808,I395791);
not I_23103 (I395825,I395783);
nor I_23104 (I395842,I395825,I395726);
DFFARX1 I_23105 (I395842,I3035,I395556,I395542,);
nand I_23106 (I395873,I135427,I135430);
and I_23107 (I395890,I395873,I135439);
DFFARX1 I_23108 (I395890,I3035,I395556,I395916,);
nor I_23109 (I395924,I395916,I395783);
DFFARX1 I_23110 (I395924,I3035,I395556,I395524,);
nand I_23111 (I395955,I395916,I395825);
nand I_23112 (I395533,I395808,I395955);
not I_23113 (I395986,I395916);
nor I_23114 (I396003,I395986,I395726);
DFFARX1 I_23115 (I396003,I3035,I395556,I395545,);
nor I_23116 (I396034,I135445,I135430);
or I_23117 (I395536,I395783,I396034);
nor I_23118 (I395527,I395916,I396034);
or I_23119 (I395530,I395650,I396034);
DFFARX1 I_23120 (I396034,I3035,I395556,I395548,);
not I_23121 (I396134,I3042);
DFFARX1 I_23122 (I168241,I3035,I396134,I396160,);
not I_23123 (I396168,I396160);
nand I_23124 (I396185,I168244,I168220);
and I_23125 (I396202,I396185,I168217);
DFFARX1 I_23126 (I396202,I3035,I396134,I396228,);
not I_23127 (I396236,I168223);
DFFARX1 I_23128 (I168217,I3035,I396134,I396262,);
not I_23129 (I396270,I396262);
nor I_23130 (I396287,I396270,I396168);
and I_23131 (I396304,I396287,I168223);
nor I_23132 (I396321,I396270,I396236);
nor I_23133 (I396117,I396228,I396321);
DFFARX1 I_23134 (I168226,I3035,I396134,I396361,);
nor I_23135 (I396369,I396361,I396228);
not I_23136 (I396386,I396369);
not I_23137 (I396403,I396361);
nor I_23138 (I396420,I396403,I396304);
DFFARX1 I_23139 (I396420,I3035,I396134,I396120,);
nand I_23140 (I396451,I168229,I168238);
and I_23141 (I396468,I396451,I168235);
DFFARX1 I_23142 (I396468,I3035,I396134,I396494,);
nor I_23143 (I396502,I396494,I396361);
DFFARX1 I_23144 (I396502,I3035,I396134,I396102,);
nand I_23145 (I396533,I396494,I396403);
nand I_23146 (I396111,I396386,I396533);
not I_23147 (I396564,I396494);
nor I_23148 (I396581,I396564,I396304);
DFFARX1 I_23149 (I396581,I3035,I396134,I396123,);
nor I_23150 (I396612,I168232,I168238);
or I_23151 (I396114,I396361,I396612);
nor I_23152 (I396105,I396494,I396612);
or I_23153 (I396108,I396228,I396612);
DFFARX1 I_23154 (I396612,I3035,I396134,I396126,);
not I_23155 (I396712,I3042);
DFFARX1 I_23156 (I686360,I3035,I396712,I396738,);
not I_23157 (I396746,I396738);
nand I_23158 (I396763,I686384,I686366);
and I_23159 (I396780,I396763,I686372);
DFFARX1 I_23160 (I396780,I3035,I396712,I396806,);
not I_23161 (I396814,I686378);
DFFARX1 I_23162 (I686363,I3035,I396712,I396840,);
not I_23163 (I396848,I396840);
nor I_23164 (I396865,I396848,I396746);
and I_23165 (I396882,I396865,I686378);
nor I_23166 (I396899,I396848,I396814);
nor I_23167 (I396695,I396806,I396899);
DFFARX1 I_23168 (I686375,I3035,I396712,I396939,);
nor I_23169 (I396947,I396939,I396806);
not I_23170 (I396964,I396947);
not I_23171 (I396981,I396939);
nor I_23172 (I396998,I396981,I396882);
DFFARX1 I_23173 (I396998,I3035,I396712,I396698,);
nand I_23174 (I397029,I686381,I686369);
and I_23175 (I397046,I397029,I686363);
DFFARX1 I_23176 (I397046,I3035,I396712,I397072,);
nor I_23177 (I397080,I397072,I396939);
DFFARX1 I_23178 (I397080,I3035,I396712,I396680,);
nand I_23179 (I397111,I397072,I396981);
nand I_23180 (I396689,I396964,I397111);
not I_23181 (I397142,I397072);
nor I_23182 (I397159,I397142,I396882);
DFFARX1 I_23183 (I397159,I3035,I396712,I396701,);
nor I_23184 (I397190,I686360,I686369);
or I_23185 (I396692,I396939,I397190);
nor I_23186 (I396683,I397072,I397190);
or I_23187 (I396686,I396806,I397190);
DFFARX1 I_23188 (I397190,I3035,I396712,I396704,);
not I_23189 (I397290,I3042);
DFFARX1 I_23190 (I313448,I3035,I397290,I397316,);
not I_23191 (I397324,I397316);
nand I_23192 (I397341,I313457,I313466);
and I_23193 (I397358,I397341,I313472);
DFFARX1 I_23194 (I397358,I3035,I397290,I397384,);
not I_23195 (I397392,I313469);
DFFARX1 I_23196 (I313454,I3035,I397290,I397418,);
not I_23197 (I397426,I397418);
nor I_23198 (I397443,I397426,I397324);
and I_23199 (I397460,I397443,I313469);
nor I_23200 (I397477,I397426,I397392);
nor I_23201 (I397273,I397384,I397477);
DFFARX1 I_23202 (I313463,I3035,I397290,I397517,);
nor I_23203 (I397525,I397517,I397384);
not I_23204 (I397542,I397525);
not I_23205 (I397559,I397517);
nor I_23206 (I397576,I397559,I397460);
DFFARX1 I_23207 (I397576,I3035,I397290,I397276,);
nand I_23208 (I397607,I313460,I313451);
and I_23209 (I397624,I397607,I313448);
DFFARX1 I_23210 (I397624,I3035,I397290,I397650,);
nor I_23211 (I397658,I397650,I397517);
DFFARX1 I_23212 (I397658,I3035,I397290,I397258,);
nand I_23213 (I397689,I397650,I397559);
nand I_23214 (I397267,I397542,I397689);
not I_23215 (I397720,I397650);
nor I_23216 (I397737,I397720,I397460);
DFFARX1 I_23217 (I397737,I3035,I397290,I397279,);
nor I_23218 (I397768,I313451,I313451);
or I_23219 (I397270,I397517,I397768);
nor I_23220 (I397261,I397650,I397768);
or I_23221 (I397264,I397384,I397768);
DFFARX1 I_23222 (I397768,I3035,I397290,I397282,);
not I_23223 (I397868,I3042);
DFFARX1 I_23224 (I454597,I3035,I397868,I397894,);
not I_23225 (I397902,I397894);
nand I_23226 (I397919,I454585,I454603);
and I_23227 (I397936,I397919,I454600);
DFFARX1 I_23228 (I397936,I3035,I397868,I397962,);
not I_23229 (I397970,I454591);
DFFARX1 I_23230 (I454588,I3035,I397868,I397996,);
not I_23231 (I398004,I397996);
nor I_23232 (I398021,I398004,I397902);
and I_23233 (I398038,I398021,I454591);
nor I_23234 (I398055,I398004,I397970);
nor I_23235 (I397851,I397962,I398055);
DFFARX1 I_23236 (I454582,I3035,I397868,I398095,);
nor I_23237 (I398103,I398095,I397962);
not I_23238 (I398120,I398103);
not I_23239 (I398137,I398095);
nor I_23240 (I398154,I398137,I398038);
DFFARX1 I_23241 (I398154,I3035,I397868,I397854,);
nand I_23242 (I398185,I454582,I454585);
and I_23243 (I398202,I398185,I454588);
DFFARX1 I_23244 (I398202,I3035,I397868,I398228,);
nor I_23245 (I398236,I398228,I398095);
DFFARX1 I_23246 (I398236,I3035,I397868,I397836,);
nand I_23247 (I398267,I398228,I398137);
nand I_23248 (I397845,I398120,I398267);
not I_23249 (I398298,I398228);
nor I_23250 (I398315,I398298,I398038);
DFFARX1 I_23251 (I398315,I3035,I397868,I397857,);
nor I_23252 (I398346,I454594,I454585);
or I_23253 (I397848,I398095,I398346);
nor I_23254 (I397839,I398228,I398346);
or I_23255 (I397842,I397962,I398346);
DFFARX1 I_23256 (I398346,I3035,I397868,I397860,);
not I_23257 (I398446,I3042);
DFFARX1 I_23258 (I669190,I3035,I398446,I398472,);
not I_23259 (I398480,I398472);
nand I_23260 (I398497,I669193,I669202);
and I_23261 (I398514,I398497,I669205);
DFFARX1 I_23262 (I398514,I3035,I398446,I398540,);
not I_23263 (I398548,I669214);
DFFARX1 I_23264 (I669196,I3035,I398446,I398574,);
not I_23265 (I398582,I398574);
nor I_23266 (I398599,I398582,I398480);
and I_23267 (I398616,I398599,I669214);
nor I_23268 (I398633,I398582,I398548);
nor I_23269 (I398429,I398540,I398633);
DFFARX1 I_23270 (I669193,I3035,I398446,I398673,);
nor I_23271 (I398681,I398673,I398540);
not I_23272 (I398698,I398681);
not I_23273 (I398715,I398673);
nor I_23274 (I398732,I398715,I398616);
DFFARX1 I_23275 (I398732,I3035,I398446,I398432,);
nand I_23276 (I398763,I669211,I669190);
and I_23277 (I398780,I398763,I669208);
DFFARX1 I_23278 (I398780,I3035,I398446,I398806,);
nor I_23279 (I398814,I398806,I398673);
DFFARX1 I_23280 (I398814,I3035,I398446,I398414,);
nand I_23281 (I398845,I398806,I398715);
nand I_23282 (I398423,I398698,I398845);
not I_23283 (I398876,I398806);
nor I_23284 (I398893,I398876,I398616);
DFFARX1 I_23285 (I398893,I3035,I398446,I398435,);
nor I_23286 (I398924,I669199,I669190);
or I_23287 (I398426,I398673,I398924);
nor I_23288 (I398417,I398806,I398924);
or I_23289 (I398420,I398540,I398924);
DFFARX1 I_23290 (I398924,I3035,I398446,I398438,);
not I_23291 (I399024,I3042);
DFFARX1 I_23292 (I22046,I3035,I399024,I399050,);
not I_23293 (I399058,I399050);
nand I_23294 (I399075,I22043,I22034);
and I_23295 (I399092,I399075,I22034);
DFFARX1 I_23296 (I399092,I3035,I399024,I399118,);
not I_23297 (I399126,I22037);
DFFARX1 I_23298 (I22052,I3035,I399024,I399152,);
not I_23299 (I399160,I399152);
nor I_23300 (I399177,I399160,I399058);
and I_23301 (I399194,I399177,I22037);
nor I_23302 (I399211,I399160,I399126);
nor I_23303 (I399007,I399118,I399211);
DFFARX1 I_23304 (I22037,I3035,I399024,I399251,);
nor I_23305 (I399259,I399251,I399118);
not I_23306 (I399276,I399259);
not I_23307 (I399293,I399251);
nor I_23308 (I399310,I399293,I399194);
DFFARX1 I_23309 (I399310,I3035,I399024,I399010,);
nand I_23310 (I399341,I22055,I22040);
and I_23311 (I399358,I399341,I22058);
DFFARX1 I_23312 (I399358,I3035,I399024,I399384,);
nor I_23313 (I399392,I399384,I399251);
DFFARX1 I_23314 (I399392,I3035,I399024,I398992,);
nand I_23315 (I399423,I399384,I399293);
nand I_23316 (I399001,I399276,I399423);
not I_23317 (I399454,I399384);
nor I_23318 (I399471,I399454,I399194);
DFFARX1 I_23319 (I399471,I3035,I399024,I399013,);
nor I_23320 (I399502,I22049,I22040);
or I_23321 (I399004,I399251,I399502);
nor I_23322 (I398995,I399384,I399502);
or I_23323 (I398998,I399118,I399502);
DFFARX1 I_23324 (I399502,I3035,I399024,I399016,);
not I_23325 (I399602,I3042);
DFFARX1 I_23326 (I150850,I3035,I399602,I399628,);
not I_23327 (I399636,I399628);
nand I_23328 (I399653,I150853,I150829);
and I_23329 (I399670,I399653,I150826);
DFFARX1 I_23330 (I399670,I3035,I399602,I399696,);
not I_23331 (I399704,I150832);
DFFARX1 I_23332 (I150826,I3035,I399602,I399730,);
not I_23333 (I399738,I399730);
nor I_23334 (I399755,I399738,I399636);
and I_23335 (I399772,I399755,I150832);
nor I_23336 (I399789,I399738,I399704);
nor I_23337 (I399585,I399696,I399789);
DFFARX1 I_23338 (I150835,I3035,I399602,I399829,);
nor I_23339 (I399837,I399829,I399696);
not I_23340 (I399854,I399837);
not I_23341 (I399871,I399829);
nor I_23342 (I399888,I399871,I399772);
DFFARX1 I_23343 (I399888,I3035,I399602,I399588,);
nand I_23344 (I399919,I150838,I150847);
and I_23345 (I399936,I399919,I150844);
DFFARX1 I_23346 (I399936,I3035,I399602,I399962,);
nor I_23347 (I399970,I399962,I399829);
DFFARX1 I_23348 (I399970,I3035,I399602,I399570,);
nand I_23349 (I400001,I399962,I399871);
nand I_23350 (I399579,I399854,I400001);
not I_23351 (I400032,I399962);
nor I_23352 (I400049,I400032,I399772);
DFFARX1 I_23353 (I400049,I3035,I399602,I399591,);
nor I_23354 (I400080,I150841,I150847);
or I_23355 (I399582,I399829,I400080);
nor I_23356 (I399573,I399962,I400080);
or I_23357 (I399576,I399696,I400080);
DFFARX1 I_23358 (I400080,I3035,I399602,I399594,);
not I_23359 (I400180,I3042);
DFFARX1 I_23360 (I670822,I3035,I400180,I400206,);
not I_23361 (I400214,I400206);
nand I_23362 (I400231,I670825,I670834);
and I_23363 (I400248,I400231,I670837);
DFFARX1 I_23364 (I400248,I3035,I400180,I400274,);
not I_23365 (I400282,I670846);
DFFARX1 I_23366 (I670828,I3035,I400180,I400308,);
not I_23367 (I400316,I400308);
nor I_23368 (I400333,I400316,I400214);
and I_23369 (I400350,I400333,I670846);
nor I_23370 (I400367,I400316,I400282);
nor I_23371 (I400163,I400274,I400367);
DFFARX1 I_23372 (I670825,I3035,I400180,I400407,);
nor I_23373 (I400415,I400407,I400274);
not I_23374 (I400432,I400415);
not I_23375 (I400449,I400407);
nor I_23376 (I400466,I400449,I400350);
DFFARX1 I_23377 (I400466,I3035,I400180,I400166,);
nand I_23378 (I400497,I670843,I670822);
and I_23379 (I400514,I400497,I670840);
DFFARX1 I_23380 (I400514,I3035,I400180,I400540,);
nor I_23381 (I400548,I400540,I400407);
DFFARX1 I_23382 (I400548,I3035,I400180,I400148,);
nand I_23383 (I400579,I400540,I400449);
nand I_23384 (I400157,I400432,I400579);
not I_23385 (I400610,I400540);
nor I_23386 (I400627,I400610,I400350);
DFFARX1 I_23387 (I400627,I3035,I400180,I400169,);
nor I_23388 (I400658,I670831,I670822);
or I_23389 (I400160,I400407,I400658);
nor I_23390 (I400151,I400540,I400658);
or I_23391 (I400154,I400274,I400658);
DFFARX1 I_23392 (I400658,I3035,I400180,I400172,);
not I_23393 (I400758,I3042);
DFFARX1 I_23394 (I545862,I3035,I400758,I400784,);
not I_23395 (I400792,I400784);
nand I_23396 (I400809,I545838,I545853);
and I_23397 (I400826,I400809,I545865);
DFFARX1 I_23398 (I400826,I3035,I400758,I400852,);
not I_23399 (I400860,I545850);
DFFARX1 I_23400 (I545841,I3035,I400758,I400886,);
not I_23401 (I400894,I400886);
nor I_23402 (I400911,I400894,I400792);
and I_23403 (I400928,I400911,I545850);
nor I_23404 (I400945,I400894,I400860);
nor I_23405 (I400741,I400852,I400945);
DFFARX1 I_23406 (I545838,I3035,I400758,I400985,);
nor I_23407 (I400993,I400985,I400852);
not I_23408 (I401010,I400993);
not I_23409 (I401027,I400985);
nor I_23410 (I401044,I401027,I400928);
DFFARX1 I_23411 (I401044,I3035,I400758,I400744,);
nand I_23412 (I401075,I545856,I545847);
and I_23413 (I401092,I401075,I545859);
DFFARX1 I_23414 (I401092,I3035,I400758,I401118,);
nor I_23415 (I401126,I401118,I400985);
DFFARX1 I_23416 (I401126,I3035,I400758,I400726,);
nand I_23417 (I401157,I401118,I401027);
nand I_23418 (I400735,I401010,I401157);
not I_23419 (I401188,I401118);
nor I_23420 (I401205,I401188,I400928);
DFFARX1 I_23421 (I401205,I3035,I400758,I400747,);
nor I_23422 (I401236,I545844,I545847);
or I_23423 (I400738,I400985,I401236);
nor I_23424 (I400729,I401118,I401236);
or I_23425 (I400732,I400852,I401236);
DFFARX1 I_23426 (I401236,I3035,I400758,I400750,);
not I_23427 (I401336,I3042);
DFFARX1 I_23428 (I7817,I3035,I401336,I401362,);
not I_23429 (I401370,I401362);
nand I_23430 (I401387,I7814,I7805);
and I_23431 (I401404,I401387,I7805);
DFFARX1 I_23432 (I401404,I3035,I401336,I401430,);
not I_23433 (I401438,I7808);
DFFARX1 I_23434 (I7823,I3035,I401336,I401464,);
not I_23435 (I401472,I401464);
nor I_23436 (I401489,I401472,I401370);
and I_23437 (I401506,I401489,I7808);
nor I_23438 (I401523,I401472,I401438);
nor I_23439 (I401319,I401430,I401523);
DFFARX1 I_23440 (I7808,I3035,I401336,I401563,);
nor I_23441 (I401571,I401563,I401430);
not I_23442 (I401588,I401571);
not I_23443 (I401605,I401563);
nor I_23444 (I401622,I401605,I401506);
DFFARX1 I_23445 (I401622,I3035,I401336,I401322,);
nand I_23446 (I401653,I7826,I7811);
and I_23447 (I401670,I401653,I7829);
DFFARX1 I_23448 (I401670,I3035,I401336,I401696,);
nor I_23449 (I401704,I401696,I401563);
DFFARX1 I_23450 (I401704,I3035,I401336,I401304,);
nand I_23451 (I401735,I401696,I401605);
nand I_23452 (I401313,I401588,I401735);
not I_23453 (I401766,I401696);
nor I_23454 (I401783,I401766,I401506);
DFFARX1 I_23455 (I401783,I3035,I401336,I401325,);
nor I_23456 (I401814,I7820,I7811);
or I_23457 (I401316,I401563,I401814);
nor I_23458 (I401307,I401696,I401814);
or I_23459 (I401310,I401430,I401814);
DFFARX1 I_23460 (I401814,I3035,I401336,I401328,);
not I_23461 (I401914,I3042);
DFFARX1 I_23462 (I706770,I3035,I401914,I401940,);
not I_23463 (I401948,I401940);
nand I_23464 (I401965,I706755,I706743);
and I_23465 (I401982,I401965,I706758);
DFFARX1 I_23466 (I401982,I3035,I401914,I402008,);
not I_23467 (I402016,I706743);
DFFARX1 I_23468 (I706761,I3035,I401914,I402042,);
not I_23469 (I402050,I402042);
nor I_23470 (I402067,I402050,I401948);
and I_23471 (I402084,I402067,I706743);
nor I_23472 (I402101,I402050,I402016);
nor I_23473 (I401897,I402008,I402101);
DFFARX1 I_23474 (I706749,I3035,I401914,I402141,);
nor I_23475 (I402149,I402141,I402008);
not I_23476 (I402166,I402149);
not I_23477 (I402183,I402141);
nor I_23478 (I402200,I402183,I402084);
DFFARX1 I_23479 (I402200,I3035,I401914,I401900,);
nand I_23480 (I402231,I706746,I706752);
and I_23481 (I402248,I402231,I706767);
DFFARX1 I_23482 (I402248,I3035,I401914,I402274,);
nor I_23483 (I402282,I402274,I402141);
DFFARX1 I_23484 (I402282,I3035,I401914,I401882,);
nand I_23485 (I402313,I402274,I402183);
nand I_23486 (I401891,I402166,I402313);
not I_23487 (I402344,I402274);
nor I_23488 (I402361,I402344,I402084);
DFFARX1 I_23489 (I402361,I3035,I401914,I401903,);
nor I_23490 (I402392,I706764,I706752);
or I_23491 (I401894,I402141,I402392);
nor I_23492 (I401885,I402274,I402392);
or I_23493 (I401888,I402008,I402392);
DFFARX1 I_23494 (I402392,I3035,I401914,I401906,);
not I_23495 (I402492,I3042);
DFFARX1 I_23496 (I268526,I3035,I402492,I402518,);
not I_23497 (I402526,I402518);
nand I_23498 (I402543,I268517,I268535);
and I_23499 (I402560,I402543,I268538);
DFFARX1 I_23500 (I402560,I3035,I402492,I402586,);
not I_23501 (I402594,I268532);
DFFARX1 I_23502 (I268520,I3035,I402492,I402620,);
not I_23503 (I402628,I402620);
nor I_23504 (I402645,I402628,I402526);
and I_23505 (I402662,I402645,I268532);
nor I_23506 (I402679,I402628,I402594);
nor I_23507 (I402475,I402586,I402679);
DFFARX1 I_23508 (I268529,I3035,I402492,I402719,);
nor I_23509 (I402727,I402719,I402586);
not I_23510 (I402744,I402727);
not I_23511 (I402761,I402719);
nor I_23512 (I402778,I402761,I402662);
DFFARX1 I_23513 (I402778,I3035,I402492,I402478,);
nand I_23514 (I402809,I268544,I268541);
and I_23515 (I402826,I402809,I268523);
DFFARX1 I_23516 (I402826,I3035,I402492,I402852,);
nor I_23517 (I402860,I402852,I402719);
DFFARX1 I_23518 (I402860,I3035,I402492,I402460,);
nand I_23519 (I402891,I402852,I402761);
nand I_23520 (I402469,I402744,I402891);
not I_23521 (I402922,I402852);
nor I_23522 (I402939,I402922,I402662);
DFFARX1 I_23523 (I402939,I3035,I402492,I402481,);
nor I_23524 (I402970,I268517,I268541);
or I_23525 (I402472,I402719,I402970);
nor I_23526 (I402463,I402852,I402970);
or I_23527 (I402466,I402586,I402970);
DFFARX1 I_23528 (I402970,I3035,I402492,I402484,);
not I_23529 (I403070,I3042);
DFFARX1 I_23530 (I207239,I3035,I403070,I403096,);
not I_23531 (I403104,I403096);
nand I_23532 (I403121,I207242,I207218);
and I_23533 (I403138,I403121,I207215);
DFFARX1 I_23534 (I403138,I3035,I403070,I403164,);
not I_23535 (I403172,I207221);
DFFARX1 I_23536 (I207215,I3035,I403070,I403198,);
not I_23537 (I403206,I403198);
nor I_23538 (I403223,I403206,I403104);
and I_23539 (I403240,I403223,I207221);
nor I_23540 (I403257,I403206,I403172);
nor I_23541 (I403053,I403164,I403257);
DFFARX1 I_23542 (I207224,I3035,I403070,I403297,);
nor I_23543 (I403305,I403297,I403164);
not I_23544 (I403322,I403305);
not I_23545 (I403339,I403297);
nor I_23546 (I403356,I403339,I403240);
DFFARX1 I_23547 (I403356,I3035,I403070,I403056,);
nand I_23548 (I403387,I207227,I207236);
and I_23549 (I403404,I403387,I207233);
DFFARX1 I_23550 (I403404,I3035,I403070,I403430,);
nor I_23551 (I403438,I403430,I403297);
DFFARX1 I_23552 (I403438,I3035,I403070,I403038,);
nand I_23553 (I403469,I403430,I403339);
nand I_23554 (I403047,I403322,I403469);
not I_23555 (I403500,I403430);
nor I_23556 (I403517,I403500,I403240);
DFFARX1 I_23557 (I403517,I3035,I403070,I403059,);
nor I_23558 (I403548,I207230,I207236);
or I_23559 (I403050,I403297,I403548);
nor I_23560 (I403041,I403430,I403548);
or I_23561 (I403044,I403164,I403548);
DFFARX1 I_23562 (I403548,I3035,I403070,I403062,);
not I_23563 (I403648,I3042);
DFFARX1 I_23564 (I62089,I3035,I403648,I403674,);
not I_23565 (I403682,I403674);
nand I_23566 (I403699,I62098,I62107);
and I_23567 (I403716,I403699,I62086);
DFFARX1 I_23568 (I403716,I3035,I403648,I403742,);
not I_23569 (I403750,I62089);
DFFARX1 I_23570 (I62104,I3035,I403648,I403776,);
not I_23571 (I403784,I403776);
nor I_23572 (I403801,I403784,I403682);
and I_23573 (I403818,I403801,I62089);
nor I_23574 (I403835,I403784,I403750);
nor I_23575 (I403631,I403742,I403835);
DFFARX1 I_23576 (I62095,I3035,I403648,I403875,);
nor I_23577 (I403883,I403875,I403742);
not I_23578 (I403900,I403883);
not I_23579 (I403917,I403875);
nor I_23580 (I403934,I403917,I403818);
DFFARX1 I_23581 (I403934,I3035,I403648,I403634,);
nand I_23582 (I403965,I62110,I62086);
and I_23583 (I403982,I403965,I62092);
DFFARX1 I_23584 (I403982,I3035,I403648,I404008,);
nor I_23585 (I404016,I404008,I403875);
DFFARX1 I_23586 (I404016,I3035,I403648,I403616,);
nand I_23587 (I404047,I404008,I403917);
nand I_23588 (I403625,I403900,I404047);
not I_23589 (I404078,I404008);
nor I_23590 (I404095,I404078,I403818);
DFFARX1 I_23591 (I404095,I3035,I403648,I403637,);
nor I_23592 (I404126,I62101,I62086);
or I_23593 (I403628,I403875,I404126);
nor I_23594 (I403619,I404008,I404126);
or I_23595 (I403622,I403742,I404126);
DFFARX1 I_23596 (I404126,I3035,I403648,I403640,);
not I_23597 (I404226,I3042);
DFFARX1 I_23598 (I550978,I3035,I404226,I404252,);
not I_23599 (I404260,I404252);
nand I_23600 (I404277,I550975,I550993);
and I_23601 (I404294,I404277,I550990);
DFFARX1 I_23602 (I404294,I3035,I404226,I404320,);
not I_23603 (I404328,I550972);
DFFARX1 I_23604 (I550975,I3035,I404226,I404354,);
not I_23605 (I404362,I404354);
nor I_23606 (I404379,I404362,I404260);
and I_23607 (I404396,I404379,I550972);
nor I_23608 (I404413,I404362,I404328);
nor I_23609 (I404209,I404320,I404413);
DFFARX1 I_23610 (I550984,I3035,I404226,I404453,);
nor I_23611 (I404461,I404453,I404320);
not I_23612 (I404478,I404461);
not I_23613 (I404495,I404453);
nor I_23614 (I404512,I404495,I404396);
DFFARX1 I_23615 (I404512,I3035,I404226,I404212,);
nand I_23616 (I404543,I550987,I550972);
and I_23617 (I404560,I404543,I550978);
DFFARX1 I_23618 (I404560,I3035,I404226,I404586,);
nor I_23619 (I404594,I404586,I404453);
DFFARX1 I_23620 (I404594,I3035,I404226,I404194,);
nand I_23621 (I404625,I404586,I404495);
nand I_23622 (I404203,I404478,I404625);
not I_23623 (I404656,I404586);
nor I_23624 (I404673,I404656,I404396);
DFFARX1 I_23625 (I404673,I3035,I404226,I404215,);
nor I_23626 (I404704,I550981,I550972);
or I_23627 (I404206,I404453,I404704);
nor I_23628 (I404197,I404586,I404704);
or I_23629 (I404200,I404320,I404704);
DFFARX1 I_23630 (I404704,I3035,I404226,I404218,);
not I_23631 (I404804,I3042);
DFFARX1 I_23632 (I102699,I3035,I404804,I404830,);
not I_23633 (I404838,I404830);
nand I_23634 (I404855,I102702,I102723);
and I_23635 (I404872,I404855,I102711);
DFFARX1 I_23636 (I404872,I3035,I404804,I404898,);
not I_23637 (I404906,I102708);
DFFARX1 I_23638 (I102699,I3035,I404804,I404932,);
not I_23639 (I404940,I404932);
nor I_23640 (I404957,I404940,I404838);
and I_23641 (I404974,I404957,I102708);
nor I_23642 (I404991,I404940,I404906);
nor I_23643 (I404787,I404898,I404991);
DFFARX1 I_23644 (I102717,I3035,I404804,I405031,);
nor I_23645 (I405039,I405031,I404898);
not I_23646 (I405056,I405039);
not I_23647 (I405073,I405031);
nor I_23648 (I405090,I405073,I404974);
DFFARX1 I_23649 (I405090,I3035,I404804,I404790,);
nand I_23650 (I405121,I102702,I102705);
and I_23651 (I405138,I405121,I102714);
DFFARX1 I_23652 (I405138,I3035,I404804,I405164,);
nor I_23653 (I405172,I405164,I405031);
DFFARX1 I_23654 (I405172,I3035,I404804,I404772,);
nand I_23655 (I405203,I405164,I405073);
nand I_23656 (I404781,I405056,I405203);
not I_23657 (I405234,I405164);
nor I_23658 (I405251,I405234,I404974);
DFFARX1 I_23659 (I405251,I3035,I404804,I404793,);
nor I_23660 (I405282,I102720,I102705);
or I_23661 (I404784,I405031,I405282);
nor I_23662 (I404775,I405164,I405282);
or I_23663 (I404778,I404898,I405282);
DFFARX1 I_23664 (I405282,I3035,I404804,I404796,);
not I_23665 (I405382,I3042);
DFFARX1 I_23666 (I480616,I3035,I405382,I405408,);
not I_23667 (I405416,I405408);
nand I_23668 (I405433,I480592,I480607);
and I_23669 (I405450,I405433,I480619);
DFFARX1 I_23670 (I405450,I3035,I405382,I405476,);
not I_23671 (I405484,I480604);
DFFARX1 I_23672 (I480595,I3035,I405382,I405510,);
not I_23673 (I405518,I405510);
nor I_23674 (I405535,I405518,I405416);
and I_23675 (I405552,I405535,I480604);
nor I_23676 (I405569,I405518,I405484);
nor I_23677 (I405365,I405476,I405569);
DFFARX1 I_23678 (I480592,I3035,I405382,I405609,);
nor I_23679 (I405617,I405609,I405476);
not I_23680 (I405634,I405617);
not I_23681 (I405651,I405609);
nor I_23682 (I405668,I405651,I405552);
DFFARX1 I_23683 (I405668,I3035,I405382,I405368,);
nand I_23684 (I405699,I480610,I480601);
and I_23685 (I405716,I405699,I480613);
DFFARX1 I_23686 (I405716,I3035,I405382,I405742,);
nor I_23687 (I405750,I405742,I405609);
DFFARX1 I_23688 (I405750,I3035,I405382,I405350,);
nand I_23689 (I405781,I405742,I405651);
nand I_23690 (I405359,I405634,I405781);
not I_23691 (I405812,I405742);
nor I_23692 (I405829,I405812,I405552);
DFFARX1 I_23693 (I405829,I3035,I405382,I405371,);
nor I_23694 (I405860,I480598,I480601);
or I_23695 (I405362,I405609,I405860);
nor I_23696 (I405353,I405742,I405860);
or I_23697 (I405356,I405476,I405860);
DFFARX1 I_23698 (I405860,I3035,I405382,I405374,);
not I_23699 (I405960,I3042);
DFFARX1 I_23700 (I75341,I3035,I405960,I405986,);
not I_23701 (I405994,I405986);
nand I_23702 (I406011,I75356,I75329);
and I_23703 (I406028,I406011,I75344);
DFFARX1 I_23704 (I406028,I3035,I405960,I406054,);
not I_23705 (I406062,I75347);
DFFARX1 I_23706 (I75332,I3035,I405960,I406088,);
not I_23707 (I406096,I406088);
nor I_23708 (I406113,I406096,I405994);
and I_23709 (I406130,I406113,I75347);
nor I_23710 (I406147,I406096,I406062);
nor I_23711 (I405943,I406054,I406147);
DFFARX1 I_23712 (I75338,I3035,I405960,I406187,);
nor I_23713 (I406195,I406187,I406054);
not I_23714 (I406212,I406195);
not I_23715 (I406229,I406187);
nor I_23716 (I406246,I406229,I406130);
DFFARX1 I_23717 (I406246,I3035,I405960,I405946,);
nand I_23718 (I406277,I75353,I75335);
and I_23719 (I406294,I406277,I75350);
DFFARX1 I_23720 (I406294,I3035,I405960,I406320,);
nor I_23721 (I406328,I406320,I406187);
DFFARX1 I_23722 (I406328,I3035,I405960,I405928,);
nand I_23723 (I406359,I406320,I406229);
nand I_23724 (I405937,I406212,I406359);
not I_23725 (I406390,I406320);
nor I_23726 (I406407,I406390,I406130);
DFFARX1 I_23727 (I406407,I3035,I405960,I405949,);
nor I_23728 (I406438,I75329,I75335);
or I_23729 (I405940,I406187,I406438);
nor I_23730 (I405931,I406320,I406438);
or I_23731 (I405934,I406054,I406438);
DFFARX1 I_23732 (I406438,I3035,I405960,I405952,);
not I_23733 (I406538,I3042);
DFFARX1 I_23734 (I3051,I3035,I406538,I406564,);
not I_23735 (I406572,I406564);
nand I_23736 (I406589,I3054,I3066);
and I_23737 (I406606,I406589,I3045);
DFFARX1 I_23738 (I406606,I3035,I406538,I406632,);
not I_23739 (I406640,I3045);
DFFARX1 I_23740 (I3048,I3035,I406538,I406666,);
not I_23741 (I406674,I406666);
nor I_23742 (I406691,I406674,I406572);
and I_23743 (I406708,I406691,I3045);
nor I_23744 (I406725,I406674,I406640);
nor I_23745 (I406521,I406632,I406725);
DFFARX1 I_23746 (I3060,I3035,I406538,I406765,);
nor I_23747 (I406773,I406765,I406632);
not I_23748 (I406790,I406773);
not I_23749 (I406807,I406765);
nor I_23750 (I406824,I406807,I406708);
DFFARX1 I_23751 (I406824,I3035,I406538,I406524,);
nand I_23752 (I406855,I3063,I3048);
and I_23753 (I406872,I406855,I3057);
DFFARX1 I_23754 (I406872,I3035,I406538,I406898,);
nor I_23755 (I406906,I406898,I406765);
DFFARX1 I_23756 (I406906,I3035,I406538,I406506,);
nand I_23757 (I406937,I406898,I406807);
nand I_23758 (I406515,I406790,I406937);
not I_23759 (I406968,I406898);
nor I_23760 (I406985,I406968,I406708);
DFFARX1 I_23761 (I406985,I3035,I406538,I406527,);
nor I_23762 (I407016,I3051,I3048);
or I_23763 (I406518,I406765,I407016);
nor I_23764 (I406509,I406898,I407016);
or I_23765 (I406512,I406632,I407016);
DFFARX1 I_23766 (I407016,I3035,I406538,I406530,);
not I_23767 (I407116,I3042);
DFFARX1 I_23768 (I272334,I3035,I407116,I407142,);
not I_23769 (I407150,I407142);
nand I_23770 (I407167,I272325,I272343);
and I_23771 (I407184,I407167,I272346);
DFFARX1 I_23772 (I407184,I3035,I407116,I407210,);
not I_23773 (I407218,I272340);
DFFARX1 I_23774 (I272328,I3035,I407116,I407244,);
not I_23775 (I407252,I407244);
nor I_23776 (I407269,I407252,I407150);
and I_23777 (I407286,I407269,I272340);
nor I_23778 (I407303,I407252,I407218);
nor I_23779 (I407099,I407210,I407303);
DFFARX1 I_23780 (I272337,I3035,I407116,I407343,);
nor I_23781 (I407351,I407343,I407210);
not I_23782 (I407368,I407351);
not I_23783 (I407385,I407343);
nor I_23784 (I407402,I407385,I407286);
DFFARX1 I_23785 (I407402,I3035,I407116,I407102,);
nand I_23786 (I407433,I272352,I272349);
and I_23787 (I407450,I407433,I272331);
DFFARX1 I_23788 (I407450,I3035,I407116,I407476,);
nor I_23789 (I407484,I407476,I407343);
DFFARX1 I_23790 (I407484,I3035,I407116,I407084,);
nand I_23791 (I407515,I407476,I407385);
nand I_23792 (I407093,I407368,I407515);
not I_23793 (I407546,I407476);
nor I_23794 (I407563,I407546,I407286);
DFFARX1 I_23795 (I407563,I3035,I407116,I407105,);
nor I_23796 (I407594,I272325,I272349);
or I_23797 (I407096,I407343,I407594);
nor I_23798 (I407087,I407476,I407594);
or I_23799 (I407090,I407210,I407594);
DFFARX1 I_23800 (I407594,I3035,I407116,I407108,);
not I_23801 (I407694,I3042);
DFFARX1 I_23802 (I118169,I3035,I407694,I407720,);
not I_23803 (I407728,I407720);
nand I_23804 (I407745,I118172,I118193);
and I_23805 (I407762,I407745,I118181);
DFFARX1 I_23806 (I407762,I3035,I407694,I407788,);
not I_23807 (I407796,I118178);
DFFARX1 I_23808 (I118169,I3035,I407694,I407822,);
not I_23809 (I407830,I407822);
nor I_23810 (I407847,I407830,I407728);
and I_23811 (I407864,I407847,I118178);
nor I_23812 (I407881,I407830,I407796);
nor I_23813 (I407677,I407788,I407881);
DFFARX1 I_23814 (I118187,I3035,I407694,I407921,);
nor I_23815 (I407929,I407921,I407788);
not I_23816 (I407946,I407929);
not I_23817 (I407963,I407921);
nor I_23818 (I407980,I407963,I407864);
DFFARX1 I_23819 (I407980,I3035,I407694,I407680,);
nand I_23820 (I408011,I118172,I118175);
and I_23821 (I408028,I408011,I118184);
DFFARX1 I_23822 (I408028,I3035,I407694,I408054,);
nor I_23823 (I408062,I408054,I407921);
DFFARX1 I_23824 (I408062,I3035,I407694,I407662,);
nand I_23825 (I408093,I408054,I407963);
nand I_23826 (I407671,I407946,I408093);
not I_23827 (I408124,I408054);
nor I_23828 (I408141,I408124,I407864);
DFFARX1 I_23829 (I408141,I3035,I407694,I407683,);
nor I_23830 (I408172,I118190,I118175);
or I_23831 (I407674,I407921,I408172);
nor I_23832 (I407665,I408054,I408172);
or I_23833 (I407668,I407788,I408172);
DFFARX1 I_23834 (I408172,I3035,I407694,I407686,);
not I_23835 (I408272,I3042);
DFFARX1 I_23836 (I740685,I3035,I408272,I408298,);
not I_23837 (I408306,I408298);
nand I_23838 (I408323,I740670,I740658);
and I_23839 (I408340,I408323,I740673);
DFFARX1 I_23840 (I408340,I3035,I408272,I408366,);
not I_23841 (I408374,I740658);
DFFARX1 I_23842 (I740676,I3035,I408272,I408400,);
not I_23843 (I408408,I408400);
nor I_23844 (I408425,I408408,I408306);
and I_23845 (I408442,I408425,I740658);
nor I_23846 (I408459,I408408,I408374);
nor I_23847 (I408255,I408366,I408459);
DFFARX1 I_23848 (I740664,I3035,I408272,I408499,);
nor I_23849 (I408507,I408499,I408366);
not I_23850 (I408524,I408507);
not I_23851 (I408541,I408499);
nor I_23852 (I408558,I408541,I408442);
DFFARX1 I_23853 (I408558,I3035,I408272,I408258,);
nand I_23854 (I408589,I740661,I740667);
and I_23855 (I408606,I408589,I740682);
DFFARX1 I_23856 (I408606,I3035,I408272,I408632,);
nor I_23857 (I408640,I408632,I408499);
DFFARX1 I_23858 (I408640,I3035,I408272,I408240,);
nand I_23859 (I408671,I408632,I408541);
nand I_23860 (I408249,I408524,I408671);
not I_23861 (I408702,I408632);
nor I_23862 (I408719,I408702,I408442);
DFFARX1 I_23863 (I408719,I3035,I408272,I408261,);
nor I_23864 (I408750,I740679,I740667);
or I_23865 (I408252,I408499,I408750);
nor I_23866 (I408243,I408632,I408750);
or I_23867 (I408246,I408366,I408750);
DFFARX1 I_23868 (I408750,I3035,I408272,I408264,);
not I_23869 (I408850,I3042);
DFFARX1 I_23870 (I193010,I3035,I408850,I408876,);
not I_23871 (I408884,I408876);
nand I_23872 (I408901,I193013,I192989);
and I_23873 (I408918,I408901,I192986);
DFFARX1 I_23874 (I408918,I3035,I408850,I408944,);
not I_23875 (I408952,I192992);
DFFARX1 I_23876 (I192986,I3035,I408850,I408978,);
not I_23877 (I408986,I408978);
nor I_23878 (I409003,I408986,I408884);
and I_23879 (I409020,I409003,I192992);
nor I_23880 (I409037,I408986,I408952);
nor I_23881 (I408833,I408944,I409037);
DFFARX1 I_23882 (I192995,I3035,I408850,I409077,);
nor I_23883 (I409085,I409077,I408944);
not I_23884 (I409102,I409085);
not I_23885 (I409119,I409077);
nor I_23886 (I409136,I409119,I409020);
DFFARX1 I_23887 (I409136,I3035,I408850,I408836,);
nand I_23888 (I409167,I192998,I193007);
and I_23889 (I409184,I409167,I193004);
DFFARX1 I_23890 (I409184,I3035,I408850,I409210,);
nor I_23891 (I409218,I409210,I409077);
DFFARX1 I_23892 (I409218,I3035,I408850,I408818,);
nand I_23893 (I409249,I409210,I409119);
nand I_23894 (I408827,I409102,I409249);
not I_23895 (I409280,I409210);
nor I_23896 (I409297,I409280,I409020);
DFFARX1 I_23897 (I409297,I3035,I408850,I408839,);
nor I_23898 (I409328,I193001,I193007);
or I_23899 (I408830,I409077,I409328);
nor I_23900 (I408821,I409210,I409328);
or I_23901 (I408824,I408944,I409328);
DFFARX1 I_23902 (I409328,I3035,I408850,I408842,);
not I_23903 (I409428,I3042);
DFFARX1 I_23904 (I322696,I3035,I409428,I409454,);
not I_23905 (I409462,I409454);
nand I_23906 (I409479,I322705,I322714);
and I_23907 (I409496,I409479,I322720);
DFFARX1 I_23908 (I409496,I3035,I409428,I409522,);
not I_23909 (I409530,I322717);
DFFARX1 I_23910 (I322702,I3035,I409428,I409556,);
not I_23911 (I409564,I409556);
nor I_23912 (I409581,I409564,I409462);
and I_23913 (I409598,I409581,I322717);
nor I_23914 (I409615,I409564,I409530);
nor I_23915 (I409411,I409522,I409615);
DFFARX1 I_23916 (I322711,I3035,I409428,I409655,);
nor I_23917 (I409663,I409655,I409522);
not I_23918 (I409680,I409663);
not I_23919 (I409697,I409655);
nor I_23920 (I409714,I409697,I409598);
DFFARX1 I_23921 (I409714,I3035,I409428,I409414,);
nand I_23922 (I409745,I322708,I322699);
and I_23923 (I409762,I409745,I322696);
DFFARX1 I_23924 (I409762,I3035,I409428,I409788,);
nor I_23925 (I409796,I409788,I409655);
DFFARX1 I_23926 (I409796,I3035,I409428,I409396,);
nand I_23927 (I409827,I409788,I409697);
nand I_23928 (I409405,I409680,I409827);
not I_23929 (I409858,I409788);
nor I_23930 (I409875,I409858,I409598);
DFFARX1 I_23931 (I409875,I3035,I409428,I409417,);
nor I_23932 (I409906,I322699,I322699);
or I_23933 (I409408,I409655,I409906);
nor I_23934 (I409399,I409788,I409906);
or I_23935 (I409402,I409522,I409906);
DFFARX1 I_23936 (I409906,I3035,I409428,I409420,);
not I_23937 (I410006,I3042);
DFFARX1 I_23938 (I104484,I3035,I410006,I410032,);
not I_23939 (I410040,I410032);
nand I_23940 (I410057,I104487,I104508);
and I_23941 (I410074,I410057,I104496);
DFFARX1 I_23942 (I410074,I3035,I410006,I410100,);
not I_23943 (I410108,I104493);
DFFARX1 I_23944 (I104484,I3035,I410006,I410134,);
not I_23945 (I410142,I410134);
nor I_23946 (I410159,I410142,I410040);
and I_23947 (I410176,I410159,I104493);
nor I_23948 (I410193,I410142,I410108);
nor I_23949 (I409989,I410100,I410193);
DFFARX1 I_23950 (I104502,I3035,I410006,I410233,);
nor I_23951 (I410241,I410233,I410100);
not I_23952 (I410258,I410241);
not I_23953 (I410275,I410233);
nor I_23954 (I410292,I410275,I410176);
DFFARX1 I_23955 (I410292,I3035,I410006,I409992,);
nand I_23956 (I410323,I104487,I104490);
and I_23957 (I410340,I410323,I104499);
DFFARX1 I_23958 (I410340,I3035,I410006,I410366,);
nor I_23959 (I410374,I410366,I410233);
DFFARX1 I_23960 (I410374,I3035,I410006,I409974,);
nand I_23961 (I410405,I410366,I410275);
nand I_23962 (I409983,I410258,I410405);
not I_23963 (I410436,I410366);
nor I_23964 (I410453,I410436,I410176);
DFFARX1 I_23965 (I410453,I3035,I410006,I409995,);
nor I_23966 (I410484,I104505,I104490);
or I_23967 (I409986,I410233,I410484);
nor I_23968 (I409977,I410366,I410484);
or I_23969 (I409980,I410100,I410484);
DFFARX1 I_23970 (I410484,I3035,I410006,I409998,);
not I_23971 (I410584,I3042);
DFFARX1 I_23972 (I598318,I3035,I410584,I410610,);
not I_23973 (I410618,I410610);
nand I_23974 (I410635,I598300,I598312);
and I_23975 (I410652,I410635,I598315);
DFFARX1 I_23976 (I410652,I3035,I410584,I410678,);
not I_23977 (I410686,I598309);
DFFARX1 I_23978 (I598306,I3035,I410584,I410712,);
not I_23979 (I410720,I410712);
nor I_23980 (I410737,I410720,I410618);
and I_23981 (I410754,I410737,I598309);
nor I_23982 (I410771,I410720,I410686);
nor I_23983 (I410567,I410678,I410771);
DFFARX1 I_23984 (I598324,I3035,I410584,I410811,);
nor I_23985 (I410819,I410811,I410678);
not I_23986 (I410836,I410819);
not I_23987 (I410853,I410811);
nor I_23988 (I410870,I410853,I410754);
DFFARX1 I_23989 (I410870,I3035,I410584,I410570,);
nand I_23990 (I410901,I598303,I598303);
and I_23991 (I410918,I410901,I598300);
DFFARX1 I_23992 (I410918,I3035,I410584,I410944,);
nor I_23993 (I410952,I410944,I410811);
DFFARX1 I_23994 (I410952,I3035,I410584,I410552,);
nand I_23995 (I410983,I410944,I410853);
nand I_23996 (I410561,I410836,I410983);
not I_23997 (I411014,I410944);
nor I_23998 (I411031,I411014,I410754);
DFFARX1 I_23999 (I411031,I3035,I410584,I410573,);
nor I_24000 (I411062,I598321,I598303);
or I_24001 (I410564,I410811,I411062);
nor I_24002 (I410555,I410944,I411062);
or I_24003 (I410558,I410678,I411062);
DFFARX1 I_24004 (I411062,I3035,I410584,I410576,);
not I_24005 (I411162,I3042);
DFFARX1 I_24006 (I188794,I3035,I411162,I411188,);
not I_24007 (I411196,I411188);
nand I_24008 (I411213,I188797,I188773);
and I_24009 (I411230,I411213,I188770);
DFFARX1 I_24010 (I411230,I3035,I411162,I411256,);
not I_24011 (I411264,I188776);
DFFARX1 I_24012 (I188770,I3035,I411162,I411290,);
not I_24013 (I411298,I411290);
nor I_24014 (I411315,I411298,I411196);
and I_24015 (I411332,I411315,I188776);
nor I_24016 (I411349,I411298,I411264);
nor I_24017 (I411145,I411256,I411349);
DFFARX1 I_24018 (I188779,I3035,I411162,I411389,);
nor I_24019 (I411397,I411389,I411256);
not I_24020 (I411414,I411397);
not I_24021 (I411431,I411389);
nor I_24022 (I411448,I411431,I411332);
DFFARX1 I_24023 (I411448,I3035,I411162,I411148,);
nand I_24024 (I411479,I188782,I188791);
and I_24025 (I411496,I411479,I188788);
DFFARX1 I_24026 (I411496,I3035,I411162,I411522,);
nor I_24027 (I411530,I411522,I411389);
DFFARX1 I_24028 (I411530,I3035,I411162,I411130,);
nand I_24029 (I411561,I411522,I411431);
nand I_24030 (I411139,I411414,I411561);
not I_24031 (I411592,I411522);
nor I_24032 (I411609,I411592,I411332);
DFFARX1 I_24033 (I411609,I3035,I411162,I411151,);
nor I_24034 (I411640,I188785,I188791);
or I_24035 (I411142,I411389,I411640);
nor I_24036 (I411133,I411522,I411640);
or I_24037 (I411136,I411256,I411640);
DFFARX1 I_24038 (I411640,I3035,I411162,I411154,);
not I_24039 (I411740,I3042);
DFFARX1 I_24040 (I96154,I3035,I411740,I411766,);
not I_24041 (I411774,I411766);
nand I_24042 (I411791,I96157,I96178);
and I_24043 (I411808,I411791,I96166);
DFFARX1 I_24044 (I411808,I3035,I411740,I411834,);
not I_24045 (I411842,I96163);
DFFARX1 I_24046 (I96154,I3035,I411740,I411868,);
not I_24047 (I411876,I411868);
nor I_24048 (I411893,I411876,I411774);
and I_24049 (I411910,I411893,I96163);
nor I_24050 (I411927,I411876,I411842);
nor I_24051 (I411723,I411834,I411927);
DFFARX1 I_24052 (I96172,I3035,I411740,I411967,);
nor I_24053 (I411975,I411967,I411834);
not I_24054 (I411992,I411975);
not I_24055 (I412009,I411967);
nor I_24056 (I412026,I412009,I411910);
DFFARX1 I_24057 (I412026,I3035,I411740,I411726,);
nand I_24058 (I412057,I96157,I96160);
and I_24059 (I412074,I412057,I96169);
DFFARX1 I_24060 (I412074,I3035,I411740,I412100,);
nor I_24061 (I412108,I412100,I411967);
DFFARX1 I_24062 (I412108,I3035,I411740,I411708,);
nand I_24063 (I412139,I412100,I412009);
nand I_24064 (I411717,I411992,I412139);
not I_24065 (I412170,I412100);
nor I_24066 (I412187,I412170,I411910);
DFFARX1 I_24067 (I412187,I3035,I411740,I411729,);
nor I_24068 (I412218,I96175,I96160);
or I_24069 (I411720,I411967,I412218);
nor I_24070 (I411711,I412100,I412218);
or I_24071 (I411714,I411834,I412218);
DFFARX1 I_24072 (I412218,I3035,I411740,I411732,);
not I_24073 (I412318,I3042);
DFFARX1 I_24074 (I134829,I3035,I412318,I412344,);
not I_24075 (I412352,I412344);
nand I_24076 (I412369,I134832,I134853);
and I_24077 (I412386,I412369,I134841);
DFFARX1 I_24078 (I412386,I3035,I412318,I412412,);
not I_24079 (I412420,I134838);
DFFARX1 I_24080 (I134829,I3035,I412318,I412446,);
not I_24081 (I412454,I412446);
nor I_24082 (I412471,I412454,I412352);
and I_24083 (I412488,I412471,I134838);
nor I_24084 (I412505,I412454,I412420);
nor I_24085 (I412301,I412412,I412505);
DFFARX1 I_24086 (I134847,I3035,I412318,I412545,);
nor I_24087 (I412553,I412545,I412412);
not I_24088 (I412570,I412553);
not I_24089 (I412587,I412545);
nor I_24090 (I412604,I412587,I412488);
DFFARX1 I_24091 (I412604,I3035,I412318,I412304,);
nand I_24092 (I412635,I134832,I134835);
and I_24093 (I412652,I412635,I134844);
DFFARX1 I_24094 (I412652,I3035,I412318,I412678,);
nor I_24095 (I412686,I412678,I412545);
DFFARX1 I_24096 (I412686,I3035,I412318,I412286,);
nand I_24097 (I412717,I412678,I412587);
nand I_24098 (I412295,I412570,I412717);
not I_24099 (I412748,I412678);
nor I_24100 (I412765,I412748,I412488);
DFFARX1 I_24101 (I412765,I3035,I412318,I412307,);
nor I_24102 (I412796,I134850,I134835);
or I_24103 (I412298,I412545,I412796);
nor I_24104 (I412289,I412678,I412796);
or I_24105 (I412292,I412412,I412796);
DFFARX1 I_24106 (I412796,I3035,I412318,I412310,);
not I_24107 (I412896,I3042);
DFFARX1 I_24108 (I9398,I3035,I412896,I412922,);
not I_24109 (I412930,I412922);
nand I_24110 (I412947,I9395,I9386);
and I_24111 (I412964,I412947,I9386);
DFFARX1 I_24112 (I412964,I3035,I412896,I412990,);
not I_24113 (I412998,I9389);
DFFARX1 I_24114 (I9404,I3035,I412896,I413024,);
not I_24115 (I413032,I413024);
nor I_24116 (I413049,I413032,I412930);
and I_24117 (I413066,I413049,I9389);
nor I_24118 (I413083,I413032,I412998);
nor I_24119 (I412879,I412990,I413083);
DFFARX1 I_24120 (I9389,I3035,I412896,I413123,);
nor I_24121 (I413131,I413123,I412990);
not I_24122 (I413148,I413131);
not I_24123 (I413165,I413123);
nor I_24124 (I413182,I413165,I413066);
DFFARX1 I_24125 (I413182,I3035,I412896,I412882,);
nand I_24126 (I413213,I9407,I9392);
and I_24127 (I413230,I413213,I9410);
DFFARX1 I_24128 (I413230,I3035,I412896,I413256,);
nor I_24129 (I413264,I413256,I413123);
DFFARX1 I_24130 (I413264,I3035,I412896,I412864,);
nand I_24131 (I413295,I413256,I413165);
nand I_24132 (I412873,I413148,I413295);
not I_24133 (I413326,I413256);
nor I_24134 (I413343,I413326,I413066);
DFFARX1 I_24135 (I413343,I3035,I412896,I412885,);
nor I_24136 (I413374,I9401,I9392);
or I_24137 (I412876,I413123,I413374);
nor I_24138 (I412867,I413256,I413374);
or I_24139 (I412870,I412990,I413374);
DFFARX1 I_24140 (I413374,I3035,I412896,I412888,);
not I_24141 (I413474,I3042);
DFFARX1 I_24142 (I148514,I3035,I413474,I413500,);
not I_24143 (I413508,I413500);
nand I_24144 (I413525,I148517,I148538);
and I_24145 (I413542,I413525,I148526);
DFFARX1 I_24146 (I413542,I3035,I413474,I413568,);
not I_24147 (I413576,I148523);
DFFARX1 I_24148 (I148514,I3035,I413474,I413602,);
not I_24149 (I413610,I413602);
nor I_24150 (I413627,I413610,I413508);
and I_24151 (I413644,I413627,I148523);
nor I_24152 (I413661,I413610,I413576);
nor I_24153 (I413457,I413568,I413661);
DFFARX1 I_24154 (I148532,I3035,I413474,I413701,);
nor I_24155 (I413709,I413701,I413568);
not I_24156 (I413726,I413709);
not I_24157 (I413743,I413701);
nor I_24158 (I413760,I413743,I413644);
DFFARX1 I_24159 (I413760,I3035,I413474,I413460,);
nand I_24160 (I413791,I148517,I148520);
and I_24161 (I413808,I413791,I148529);
DFFARX1 I_24162 (I413808,I3035,I413474,I413834,);
nor I_24163 (I413842,I413834,I413701);
DFFARX1 I_24164 (I413842,I3035,I413474,I413442,);
nand I_24165 (I413873,I413834,I413743);
nand I_24166 (I413451,I413726,I413873);
not I_24167 (I413904,I413834);
nor I_24168 (I413921,I413904,I413644);
DFFARX1 I_24169 (I413921,I3035,I413474,I413463,);
nor I_24170 (I413952,I148535,I148520);
or I_24171 (I413454,I413701,I413952);
nor I_24172 (I413445,I413834,I413952);
or I_24173 (I413448,I413568,I413952);
DFFARX1 I_24174 (I413952,I3035,I413474,I413466,);
not I_24175 (I414052,I3042);
DFFARX1 I_24176 (I553783,I3035,I414052,I414078,);
not I_24177 (I414086,I414078);
nand I_24178 (I414103,I553780,I553798);
and I_24179 (I414120,I414103,I553795);
DFFARX1 I_24180 (I414120,I3035,I414052,I414146,);
not I_24181 (I414154,I553777);
DFFARX1 I_24182 (I553780,I3035,I414052,I414180,);
not I_24183 (I414188,I414180);
nor I_24184 (I414205,I414188,I414086);
and I_24185 (I414222,I414205,I553777);
nor I_24186 (I414239,I414188,I414154);
nor I_24187 (I414035,I414146,I414239);
DFFARX1 I_24188 (I553789,I3035,I414052,I414279,);
nor I_24189 (I414287,I414279,I414146);
not I_24190 (I414304,I414287);
not I_24191 (I414321,I414279);
nor I_24192 (I414338,I414321,I414222);
DFFARX1 I_24193 (I414338,I3035,I414052,I414038,);
nand I_24194 (I414369,I553792,I553777);
and I_24195 (I414386,I414369,I553783);
DFFARX1 I_24196 (I414386,I3035,I414052,I414412,);
nor I_24197 (I414420,I414412,I414279);
DFFARX1 I_24198 (I414420,I3035,I414052,I414020,);
nand I_24199 (I414451,I414412,I414321);
nand I_24200 (I414029,I414304,I414451);
not I_24201 (I414482,I414412);
nor I_24202 (I414499,I414482,I414222);
DFFARX1 I_24203 (I414499,I3035,I414052,I414041,);
nor I_24204 (I414530,I553786,I553777);
or I_24205 (I414032,I414279,I414530);
nor I_24206 (I414023,I414412,I414530);
or I_24207 (I414026,I414146,I414530);
DFFARX1 I_24208 (I414530,I3035,I414052,I414044,);
not I_24209 (I414630,I3042);
DFFARX1 I_24210 (I544570,I3035,I414630,I414656,);
not I_24211 (I414664,I414656);
nand I_24212 (I414681,I544546,I544561);
and I_24213 (I414698,I414681,I544573);
DFFARX1 I_24214 (I414698,I3035,I414630,I414724,);
not I_24215 (I414732,I544558);
DFFARX1 I_24216 (I544549,I3035,I414630,I414758,);
not I_24217 (I414766,I414758);
nor I_24218 (I414783,I414766,I414664);
and I_24219 (I414800,I414783,I544558);
nor I_24220 (I414817,I414766,I414732);
nor I_24221 (I414613,I414724,I414817);
DFFARX1 I_24222 (I544546,I3035,I414630,I414857,);
nor I_24223 (I414865,I414857,I414724);
not I_24224 (I414882,I414865);
not I_24225 (I414899,I414857);
nor I_24226 (I414916,I414899,I414800);
DFFARX1 I_24227 (I414916,I3035,I414630,I414616,);
nand I_24228 (I414947,I544564,I544555);
and I_24229 (I414964,I414947,I544567);
DFFARX1 I_24230 (I414964,I3035,I414630,I414990,);
nor I_24231 (I414998,I414990,I414857);
DFFARX1 I_24232 (I414998,I3035,I414630,I414598,);
nand I_24233 (I415029,I414990,I414899);
nand I_24234 (I414607,I414882,I415029);
not I_24235 (I415060,I414990);
nor I_24236 (I415077,I415060,I414800);
DFFARX1 I_24237 (I415077,I3035,I414630,I414619,);
nor I_24238 (I415108,I544552,I544555);
or I_24239 (I414610,I414857,I415108);
nor I_24240 (I414601,I414990,I415108);
or I_24241 (I414604,I414724,I415108);
DFFARX1 I_24242 (I415108,I3035,I414630,I414622,);
not I_24243 (I415208,I3042);
DFFARX1 I_24244 (I473569,I3035,I415208,I415234,);
not I_24245 (I415242,I415234);
nand I_24246 (I415259,I473557,I473575);
and I_24247 (I415276,I415259,I473572);
DFFARX1 I_24248 (I415276,I3035,I415208,I415302,);
not I_24249 (I415310,I473563);
DFFARX1 I_24250 (I473560,I3035,I415208,I415336,);
not I_24251 (I415344,I415336);
nor I_24252 (I415361,I415344,I415242);
and I_24253 (I415378,I415361,I473563);
nor I_24254 (I415395,I415344,I415310);
nor I_24255 (I415191,I415302,I415395);
DFFARX1 I_24256 (I473554,I3035,I415208,I415435,);
nor I_24257 (I415443,I415435,I415302);
not I_24258 (I415460,I415443);
not I_24259 (I415477,I415435);
nor I_24260 (I415494,I415477,I415378);
DFFARX1 I_24261 (I415494,I3035,I415208,I415194,);
nand I_24262 (I415525,I473554,I473557);
and I_24263 (I415542,I415525,I473560);
DFFARX1 I_24264 (I415542,I3035,I415208,I415568,);
nor I_24265 (I415576,I415568,I415435);
DFFARX1 I_24266 (I415576,I3035,I415208,I415176,);
nand I_24267 (I415607,I415568,I415477);
nand I_24268 (I415185,I415460,I415607);
not I_24269 (I415638,I415568);
nor I_24270 (I415655,I415638,I415378);
DFFARX1 I_24271 (I415655,I3035,I415208,I415197,);
nor I_24272 (I415686,I473566,I473557);
or I_24273 (I415188,I415435,I415686);
nor I_24274 (I415179,I415568,I415686);
or I_24275 (I415182,I415302,I415686);
DFFARX1 I_24276 (I415686,I3035,I415208,I415200,);
not I_24277 (I415786,I3042);
DFFARX1 I_24278 (I95559,I3035,I415786,I415812,);
not I_24279 (I415820,I415812);
nand I_24280 (I415837,I95562,I95583);
and I_24281 (I415854,I415837,I95571);
DFFARX1 I_24282 (I415854,I3035,I415786,I415880,);
not I_24283 (I415888,I95568);
DFFARX1 I_24284 (I95559,I3035,I415786,I415914,);
not I_24285 (I415922,I415914);
nor I_24286 (I415939,I415922,I415820);
and I_24287 (I415956,I415939,I95568);
nor I_24288 (I415973,I415922,I415888);
nor I_24289 (I415769,I415880,I415973);
DFFARX1 I_24290 (I95577,I3035,I415786,I416013,);
nor I_24291 (I416021,I416013,I415880);
not I_24292 (I416038,I416021);
not I_24293 (I416055,I416013);
nor I_24294 (I416072,I416055,I415956);
DFFARX1 I_24295 (I416072,I3035,I415786,I415772,);
nand I_24296 (I416103,I95562,I95565);
and I_24297 (I416120,I416103,I95574);
DFFARX1 I_24298 (I416120,I3035,I415786,I416146,);
nor I_24299 (I416154,I416146,I416013);
DFFARX1 I_24300 (I416154,I3035,I415786,I415754,);
nand I_24301 (I416185,I416146,I416055);
nand I_24302 (I415763,I416038,I416185);
not I_24303 (I416216,I416146);
nor I_24304 (I416233,I416216,I415956);
DFFARX1 I_24305 (I416233,I3035,I415786,I415775,);
nor I_24306 (I416264,I95580,I95565);
or I_24307 (I415766,I416013,I416264);
nor I_24308 (I415757,I416146,I416264);
or I_24309 (I415760,I415880,I416264);
DFFARX1 I_24310 (I416264,I3035,I415786,I415778,);
not I_24311 (I416364,I3042);
DFFARX1 I_24312 (I150323,I3035,I416364,I416390,);
not I_24313 (I416398,I416390);
nand I_24314 (I416415,I150326,I150302);
and I_24315 (I416432,I416415,I150299);
DFFARX1 I_24316 (I416432,I3035,I416364,I416458,);
not I_24317 (I416466,I150305);
DFFARX1 I_24318 (I150299,I3035,I416364,I416492,);
not I_24319 (I416500,I416492);
nor I_24320 (I416517,I416500,I416398);
and I_24321 (I416534,I416517,I150305);
nor I_24322 (I416551,I416500,I416466);
nor I_24323 (I416347,I416458,I416551);
DFFARX1 I_24324 (I150308,I3035,I416364,I416591,);
nor I_24325 (I416599,I416591,I416458);
not I_24326 (I416616,I416599);
not I_24327 (I416633,I416591);
nor I_24328 (I416650,I416633,I416534);
DFFARX1 I_24329 (I416650,I3035,I416364,I416350,);
nand I_24330 (I416681,I150311,I150320);
and I_24331 (I416698,I416681,I150317);
DFFARX1 I_24332 (I416698,I3035,I416364,I416724,);
nor I_24333 (I416732,I416724,I416591);
DFFARX1 I_24334 (I416732,I3035,I416364,I416332,);
nand I_24335 (I416763,I416724,I416633);
nand I_24336 (I416341,I416616,I416763);
not I_24337 (I416794,I416724);
nor I_24338 (I416811,I416794,I416534);
DFFARX1 I_24339 (I416811,I3035,I416364,I416353,);
nor I_24340 (I416842,I150314,I150320);
or I_24341 (I416344,I416591,I416842);
nor I_24342 (I416335,I416724,I416842);
or I_24343 (I416338,I416458,I416842);
DFFARX1 I_24344 (I416842,I3035,I416364,I416356,);
not I_24345 (I416942,I3042);
DFFARX1 I_24346 (I329632,I3035,I416942,I416968,);
not I_24347 (I416976,I416968);
nand I_24348 (I416993,I329641,I329650);
and I_24349 (I417010,I416993,I329656);
DFFARX1 I_24350 (I417010,I3035,I416942,I417036,);
not I_24351 (I417044,I329653);
DFFARX1 I_24352 (I329638,I3035,I416942,I417070,);
not I_24353 (I417078,I417070);
nor I_24354 (I417095,I417078,I416976);
and I_24355 (I417112,I417095,I329653);
nor I_24356 (I417129,I417078,I417044);
nor I_24357 (I416925,I417036,I417129);
DFFARX1 I_24358 (I329647,I3035,I416942,I417169,);
nor I_24359 (I417177,I417169,I417036);
not I_24360 (I417194,I417177);
not I_24361 (I417211,I417169);
nor I_24362 (I417228,I417211,I417112);
DFFARX1 I_24363 (I417228,I3035,I416942,I416928,);
nand I_24364 (I417259,I329644,I329635);
and I_24365 (I417276,I417259,I329632);
DFFARX1 I_24366 (I417276,I3035,I416942,I417302,);
nor I_24367 (I417310,I417302,I417169);
DFFARX1 I_24368 (I417310,I3035,I416942,I416910,);
nand I_24369 (I417341,I417302,I417211);
nand I_24370 (I416919,I417194,I417341);
not I_24371 (I417372,I417302);
nor I_24372 (I417389,I417372,I417112);
DFFARX1 I_24373 (I417389,I3035,I416942,I416931,);
nor I_24374 (I417420,I329635,I329635);
or I_24375 (I416922,I417169,I417420);
nor I_24376 (I416913,I417302,I417420);
or I_24377 (I416916,I417036,I417420);
DFFARX1 I_24378 (I417420,I3035,I416942,I416934,);
not I_24379 (I417520,I3042);
DFFARX1 I_24380 (I315760,I3035,I417520,I417546,);
not I_24381 (I417554,I417546);
nand I_24382 (I417571,I315769,I315778);
and I_24383 (I417588,I417571,I315784);
DFFARX1 I_24384 (I417588,I3035,I417520,I417614,);
not I_24385 (I417622,I315781);
DFFARX1 I_24386 (I315766,I3035,I417520,I417648,);
not I_24387 (I417656,I417648);
nor I_24388 (I417673,I417656,I417554);
and I_24389 (I417690,I417673,I315781);
nor I_24390 (I417707,I417656,I417622);
nor I_24391 (I417503,I417614,I417707);
DFFARX1 I_24392 (I315775,I3035,I417520,I417747,);
nor I_24393 (I417755,I417747,I417614);
not I_24394 (I417772,I417755);
not I_24395 (I417789,I417747);
nor I_24396 (I417806,I417789,I417690);
DFFARX1 I_24397 (I417806,I3035,I417520,I417506,);
nand I_24398 (I417837,I315772,I315763);
and I_24399 (I417854,I417837,I315760);
DFFARX1 I_24400 (I417854,I3035,I417520,I417880,);
nor I_24401 (I417888,I417880,I417747);
DFFARX1 I_24402 (I417888,I3035,I417520,I417488,);
nand I_24403 (I417919,I417880,I417789);
nand I_24404 (I417497,I417772,I417919);
not I_24405 (I417950,I417880);
nor I_24406 (I417967,I417950,I417690);
DFFARX1 I_24407 (I417967,I3035,I417520,I417509,);
nor I_24408 (I417998,I315763,I315763);
or I_24409 (I417500,I417747,I417998);
nor I_24410 (I417491,I417880,I417998);
or I_24411 (I417494,I417614,I417998);
DFFARX1 I_24412 (I417998,I3035,I417520,I417512,);
not I_24413 (I418098,I3042);
DFFARX1 I_24414 (I4836,I3035,I418098,I418124,);
not I_24415 (I418132,I418124);
nand I_24416 (I418149,I4839,I4851);
and I_24417 (I418166,I418149,I4830);
DFFARX1 I_24418 (I418166,I3035,I418098,I418192,);
not I_24419 (I418200,I4830);
DFFARX1 I_24420 (I4833,I3035,I418098,I418226,);
not I_24421 (I418234,I418226);
nor I_24422 (I418251,I418234,I418132);
and I_24423 (I418268,I418251,I4830);
nor I_24424 (I418285,I418234,I418200);
nor I_24425 (I418081,I418192,I418285);
DFFARX1 I_24426 (I4845,I3035,I418098,I418325,);
nor I_24427 (I418333,I418325,I418192);
not I_24428 (I418350,I418333);
not I_24429 (I418367,I418325);
nor I_24430 (I418384,I418367,I418268);
DFFARX1 I_24431 (I418384,I3035,I418098,I418084,);
nand I_24432 (I418415,I4848,I4833);
and I_24433 (I418432,I418415,I4842);
DFFARX1 I_24434 (I418432,I3035,I418098,I418458,);
nor I_24435 (I418466,I418458,I418325);
DFFARX1 I_24436 (I418466,I3035,I418098,I418066,);
nand I_24437 (I418497,I418458,I418367);
nand I_24438 (I418075,I418350,I418497);
not I_24439 (I418528,I418458);
nor I_24440 (I418545,I418528,I418268);
DFFARX1 I_24441 (I418545,I3035,I418098,I418087,);
nor I_24442 (I418576,I4836,I4833);
or I_24443 (I418078,I418325,I418576);
nor I_24444 (I418069,I418458,I418576);
or I_24445 (I418072,I418192,I418576);
DFFARX1 I_24446 (I418576,I3035,I418098,I418090,);
not I_24447 (I418676,I3042);
DFFARX1 I_24448 (I42063,I3035,I418676,I418702,);
not I_24449 (I418710,I418702);
nand I_24450 (I418727,I42072,I42081);
and I_24451 (I418744,I418727,I42060);
DFFARX1 I_24452 (I418744,I3035,I418676,I418770,);
not I_24453 (I418778,I42063);
DFFARX1 I_24454 (I42078,I3035,I418676,I418804,);
not I_24455 (I418812,I418804);
nor I_24456 (I418829,I418812,I418710);
and I_24457 (I418846,I418829,I42063);
nor I_24458 (I418863,I418812,I418778);
nor I_24459 (I418659,I418770,I418863);
DFFARX1 I_24460 (I42069,I3035,I418676,I418903,);
nor I_24461 (I418911,I418903,I418770);
not I_24462 (I418928,I418911);
not I_24463 (I418945,I418903);
nor I_24464 (I418962,I418945,I418846);
DFFARX1 I_24465 (I418962,I3035,I418676,I418662,);
nand I_24466 (I418993,I42084,I42060);
and I_24467 (I419010,I418993,I42066);
DFFARX1 I_24468 (I419010,I3035,I418676,I419036,);
nor I_24469 (I419044,I419036,I418903);
DFFARX1 I_24470 (I419044,I3035,I418676,I418644,);
nand I_24471 (I419075,I419036,I418945);
nand I_24472 (I418653,I418928,I419075);
not I_24473 (I419106,I419036);
nor I_24474 (I419123,I419106,I418846);
DFFARX1 I_24475 (I419123,I3035,I418676,I418665,);
nor I_24476 (I419154,I42075,I42060);
or I_24477 (I418656,I418903,I419154);
nor I_24478 (I418647,I419036,I419154);
or I_24479 (I418650,I418770,I419154);
DFFARX1 I_24480 (I419154,I3035,I418676,I418668,);
not I_24481 (I419254,I3042);
DFFARX1 I_24482 (I636466,I3035,I419254,I419280,);
not I_24483 (I419288,I419280);
nand I_24484 (I419305,I636448,I636460);
and I_24485 (I419322,I419305,I636463);
DFFARX1 I_24486 (I419322,I3035,I419254,I419348,);
not I_24487 (I419356,I636457);
DFFARX1 I_24488 (I636454,I3035,I419254,I419382,);
not I_24489 (I419390,I419382);
nor I_24490 (I419407,I419390,I419288);
and I_24491 (I419424,I419407,I636457);
nor I_24492 (I419441,I419390,I419356);
nor I_24493 (I419237,I419348,I419441);
DFFARX1 I_24494 (I636472,I3035,I419254,I419481,);
nor I_24495 (I419489,I419481,I419348);
not I_24496 (I419506,I419489);
not I_24497 (I419523,I419481);
nor I_24498 (I419540,I419523,I419424);
DFFARX1 I_24499 (I419540,I3035,I419254,I419240,);
nand I_24500 (I419571,I636451,I636451);
and I_24501 (I419588,I419571,I636448);
DFFARX1 I_24502 (I419588,I3035,I419254,I419614,);
nor I_24503 (I419622,I419614,I419481);
DFFARX1 I_24504 (I419622,I3035,I419254,I419222,);
nand I_24505 (I419653,I419614,I419523);
nand I_24506 (I419231,I419506,I419653);
not I_24507 (I419684,I419614);
nor I_24508 (I419701,I419684,I419424);
DFFARX1 I_24509 (I419701,I3035,I419254,I419243,);
nor I_24510 (I419732,I636469,I636451);
or I_24511 (I419234,I419481,I419732);
nor I_24512 (I419225,I419614,I419732);
or I_24513 (I419228,I419348,I419732);
DFFARX1 I_24514 (I419732,I3035,I419254,I419246,);
not I_24515 (I419829,I3042);
DFFARX1 I_24516 (I101515,I3035,I419829,I419855,);
not I_24517 (I419863,I419855);
nand I_24518 (I419880,I101512,I101530);
and I_24519 (I419897,I419880,I101521);
DFFARX1 I_24520 (I419897,I3035,I419829,I419923,);
DFFARX1 I_24521 (I419923,I3035,I419829,I419818,);
DFFARX1 I_24522 (I101527,I3035,I419829,I419954,);
nand I_24523 (I419962,I419954,I101524);
not I_24524 (I419979,I419962);
DFFARX1 I_24525 (I419979,I3035,I419829,I420005,);
not I_24526 (I420013,I420005);
nor I_24527 (I419821,I419863,I420013);
DFFARX1 I_24528 (I101518,I3035,I419829,I420053,);
nor I_24529 (I419812,I420053,I419923);
nor I_24530 (I419803,I420053,I419979);
nand I_24531 (I420089,I101509,I101533);
and I_24532 (I420106,I420089,I101512);
DFFARX1 I_24533 (I420106,I3035,I419829,I420132,);
not I_24534 (I420140,I420132);
nand I_24535 (I420157,I420140,I420053);
nand I_24536 (I419806,I420140,I419962);
nor I_24537 (I420188,I101509,I101533);
and I_24538 (I420205,I420053,I420188);
nor I_24539 (I420222,I420140,I420205);
DFFARX1 I_24540 (I420222,I3035,I419829,I419815,);
nor I_24541 (I420253,I419855,I420188);
DFFARX1 I_24542 (I420253,I3035,I419829,I419800,);
nor I_24543 (I420284,I420132,I420188);
not I_24544 (I420301,I420284);
nand I_24545 (I419809,I420301,I420157);
not I_24546 (I420356,I3042);
DFFARX1 I_24547 (I586180,I3035,I420356,I420382,);
not I_24548 (I420390,I420382);
nand I_24549 (I420407,I586162,I586162);
and I_24550 (I420424,I420407,I586168);
DFFARX1 I_24551 (I420424,I3035,I420356,I420450,);
DFFARX1 I_24552 (I420450,I3035,I420356,I420345,);
DFFARX1 I_24553 (I586165,I3035,I420356,I420481,);
nand I_24554 (I420489,I420481,I586174);
not I_24555 (I420506,I420489);
DFFARX1 I_24556 (I420506,I3035,I420356,I420532,);
not I_24557 (I420540,I420532);
nor I_24558 (I420348,I420390,I420540);
DFFARX1 I_24559 (I586186,I3035,I420356,I420580,);
nor I_24560 (I420339,I420580,I420450);
nor I_24561 (I420330,I420580,I420506);
nand I_24562 (I420616,I586177,I586171);
and I_24563 (I420633,I420616,I586165);
DFFARX1 I_24564 (I420633,I3035,I420356,I420659,);
not I_24565 (I420667,I420659);
nand I_24566 (I420684,I420667,I420580);
nand I_24567 (I420333,I420667,I420489);
nor I_24568 (I420715,I586183,I586171);
and I_24569 (I420732,I420580,I420715);
nor I_24570 (I420749,I420667,I420732);
DFFARX1 I_24571 (I420749,I3035,I420356,I420342,);
nor I_24572 (I420780,I420382,I420715);
DFFARX1 I_24573 (I420780,I3035,I420356,I420327,);
nor I_24574 (I420811,I420659,I420715);
not I_24575 (I420828,I420811);
nand I_24576 (I420336,I420828,I420684);
not I_24577 (I420883,I3042);
DFFARX1 I_24578 (I94375,I3035,I420883,I420909,);
not I_24579 (I420917,I420909);
nand I_24580 (I420934,I94372,I94390);
and I_24581 (I420951,I420934,I94381);
DFFARX1 I_24582 (I420951,I3035,I420883,I420977,);
DFFARX1 I_24583 (I420977,I3035,I420883,I420872,);
DFFARX1 I_24584 (I94387,I3035,I420883,I421008,);
nand I_24585 (I421016,I421008,I94384);
not I_24586 (I421033,I421016);
DFFARX1 I_24587 (I421033,I3035,I420883,I421059,);
not I_24588 (I421067,I421059);
nor I_24589 (I420875,I420917,I421067);
DFFARX1 I_24590 (I94378,I3035,I420883,I421107,);
nor I_24591 (I420866,I421107,I420977);
nor I_24592 (I420857,I421107,I421033);
nand I_24593 (I421143,I94369,I94393);
and I_24594 (I421160,I421143,I94372);
DFFARX1 I_24595 (I421160,I3035,I420883,I421186,);
not I_24596 (I421194,I421186);
nand I_24597 (I421211,I421194,I421107);
nand I_24598 (I420860,I421194,I421016);
nor I_24599 (I421242,I94369,I94393);
and I_24600 (I421259,I421107,I421242);
nor I_24601 (I421276,I421194,I421259);
DFFARX1 I_24602 (I421276,I3035,I420883,I420869,);
nor I_24603 (I421307,I420909,I421242);
DFFARX1 I_24604 (I421307,I3035,I420883,I420854,);
nor I_24605 (I421338,I421186,I421242);
not I_24606 (I421355,I421338);
nand I_24607 (I420863,I421355,I421211);
not I_24608 (I421410,I3042);
DFFARX1 I_24609 (I486409,I3035,I421410,I421436,);
not I_24610 (I421444,I421436);
nand I_24611 (I421461,I486424,I486406);
and I_24612 (I421478,I421461,I486406);
DFFARX1 I_24613 (I421478,I3035,I421410,I421504,);
DFFARX1 I_24614 (I421504,I3035,I421410,I421399,);
DFFARX1 I_24615 (I486415,I3035,I421410,I421535,);
nand I_24616 (I421543,I421535,I486433);
not I_24617 (I421560,I421543);
DFFARX1 I_24618 (I421560,I3035,I421410,I421586,);
not I_24619 (I421594,I421586);
nor I_24620 (I421402,I421444,I421594);
DFFARX1 I_24621 (I486430,I3035,I421410,I421634,);
nor I_24622 (I421393,I421634,I421504);
nor I_24623 (I421384,I421634,I421560);
nand I_24624 (I421670,I486427,I486418);
and I_24625 (I421687,I421670,I486412);
DFFARX1 I_24626 (I421687,I3035,I421410,I421713,);
not I_24627 (I421721,I421713);
nand I_24628 (I421738,I421721,I421634);
nand I_24629 (I421387,I421721,I421543);
nor I_24630 (I421769,I486421,I486418);
and I_24631 (I421786,I421634,I421769);
nor I_24632 (I421803,I421721,I421786);
DFFARX1 I_24633 (I421803,I3035,I421410,I421396,);
nor I_24634 (I421834,I421436,I421769);
DFFARX1 I_24635 (I421834,I3035,I421410,I421381,);
nor I_24636 (I421865,I421713,I421769);
not I_24637 (I421882,I421865);
nand I_24638 (I421390,I421882,I421738);
not I_24639 (I421937,I3042);
DFFARX1 I_24640 (I304793,I3035,I421937,I421963,);
not I_24641 (I421971,I421963);
nand I_24642 (I421988,I304778,I304799);
and I_24643 (I422005,I421988,I304787);
DFFARX1 I_24644 (I422005,I3035,I421937,I422031,);
DFFARX1 I_24645 (I422031,I3035,I421937,I421926,);
DFFARX1 I_24646 (I304781,I3035,I421937,I422062,);
nand I_24647 (I422070,I422062,I304790);
not I_24648 (I422087,I422070);
DFFARX1 I_24649 (I422087,I3035,I421937,I422113,);
not I_24650 (I422121,I422113);
nor I_24651 (I421929,I421971,I422121);
DFFARX1 I_24652 (I304796,I3035,I421937,I422161,);
nor I_24653 (I421920,I422161,I422031);
nor I_24654 (I421911,I422161,I422087);
nand I_24655 (I422197,I304778,I304781);
and I_24656 (I422214,I422197,I304802);
DFFARX1 I_24657 (I422214,I3035,I421937,I422240,);
not I_24658 (I422248,I422240);
nand I_24659 (I422265,I422248,I422161);
nand I_24660 (I421914,I422248,I422070);
nor I_24661 (I422296,I304784,I304781);
and I_24662 (I422313,I422161,I422296);
nor I_24663 (I422330,I422248,I422313);
DFFARX1 I_24664 (I422330,I3035,I421937,I421923,);
nor I_24665 (I422361,I421963,I422296);
DFFARX1 I_24666 (I422361,I3035,I421937,I421908,);
nor I_24667 (I422392,I422240,I422296);
not I_24668 (I422409,I422392);
nand I_24669 (I421917,I422409,I422265);
not I_24670 (I422464,I3042);
DFFARX1 I_24671 (I308839,I3035,I422464,I422490,);
not I_24672 (I422498,I422490);
nand I_24673 (I422515,I308824,I308845);
and I_24674 (I422532,I422515,I308833);
DFFARX1 I_24675 (I422532,I3035,I422464,I422558,);
DFFARX1 I_24676 (I422558,I3035,I422464,I422453,);
DFFARX1 I_24677 (I308827,I3035,I422464,I422589,);
nand I_24678 (I422597,I422589,I308836);
not I_24679 (I422614,I422597);
DFFARX1 I_24680 (I422614,I3035,I422464,I422640,);
not I_24681 (I422648,I422640);
nor I_24682 (I422456,I422498,I422648);
DFFARX1 I_24683 (I308842,I3035,I422464,I422688,);
nor I_24684 (I422447,I422688,I422558);
nor I_24685 (I422438,I422688,I422614);
nand I_24686 (I422724,I308824,I308827);
and I_24687 (I422741,I422724,I308848);
DFFARX1 I_24688 (I422741,I3035,I422464,I422767,);
not I_24689 (I422775,I422767);
nand I_24690 (I422792,I422775,I422688);
nand I_24691 (I422441,I422775,I422597);
nor I_24692 (I422823,I308830,I308827);
and I_24693 (I422840,I422688,I422823);
nor I_24694 (I422857,I422775,I422840);
DFFARX1 I_24695 (I422857,I3035,I422464,I422450,);
nor I_24696 (I422888,I422490,I422823);
DFFARX1 I_24697 (I422888,I3035,I422464,I422435,);
nor I_24698 (I422919,I422767,I422823);
not I_24699 (I422936,I422919);
nand I_24700 (I422444,I422936,I422792);
not I_24701 (I422991,I3042);
DFFARX1 I_24702 (I165591,I3035,I422991,I423017,);
not I_24703 (I423025,I423017);
nand I_24704 (I423042,I165582,I165582);
and I_24705 (I423059,I423042,I165600);
DFFARX1 I_24706 (I423059,I3035,I422991,I423085,);
DFFARX1 I_24707 (I423085,I3035,I422991,I422980,);
DFFARX1 I_24708 (I165603,I3035,I422991,I423116,);
nand I_24709 (I423124,I423116,I165585);
not I_24710 (I423141,I423124);
DFFARX1 I_24711 (I423141,I3035,I422991,I423167,);
not I_24712 (I423175,I423167);
nor I_24713 (I422983,I423025,I423175);
DFFARX1 I_24714 (I165597,I3035,I422991,I423215,);
nor I_24715 (I422974,I423215,I423085);
nor I_24716 (I422965,I423215,I423141);
nand I_24717 (I423251,I165609,I165588);
and I_24718 (I423268,I423251,I165594);
DFFARX1 I_24719 (I423268,I3035,I422991,I423294,);
not I_24720 (I423302,I423294);
nand I_24721 (I423319,I423302,I423215);
nand I_24722 (I422968,I423302,I423124);
nor I_24723 (I423350,I165606,I165588);
and I_24724 (I423367,I423215,I423350);
nor I_24725 (I423384,I423302,I423367);
DFFARX1 I_24726 (I423384,I3035,I422991,I422977,);
nor I_24727 (I423415,I423017,I423350);
DFFARX1 I_24728 (I423415,I3035,I422991,I422962,);
nor I_24729 (I423446,I423294,I423350);
not I_24730 (I423463,I423446);
nand I_24731 (I422971,I423463,I423319);
not I_24732 (I423518,I3042);
DFFARX1 I_24733 (I710328,I3035,I423518,I423544,);
not I_24734 (I423552,I423544);
nand I_24735 (I423569,I710325,I710334);
and I_24736 (I423586,I423569,I710313);
DFFARX1 I_24737 (I423586,I3035,I423518,I423612,);
DFFARX1 I_24738 (I423612,I3035,I423518,I423507,);
DFFARX1 I_24739 (I710316,I3035,I423518,I423643,);
nand I_24740 (I423651,I423643,I710331);
not I_24741 (I423668,I423651);
DFFARX1 I_24742 (I423668,I3035,I423518,I423694,);
not I_24743 (I423702,I423694);
nor I_24744 (I423510,I423552,I423702);
DFFARX1 I_24745 (I710337,I3035,I423518,I423742,);
nor I_24746 (I423501,I423742,I423612);
nor I_24747 (I423492,I423742,I423668);
nand I_24748 (I423778,I710319,I710340);
and I_24749 (I423795,I423778,I710322);
DFFARX1 I_24750 (I423795,I3035,I423518,I423821,);
not I_24751 (I423829,I423821);
nand I_24752 (I423846,I423829,I423742);
nand I_24753 (I423495,I423829,I423651);
nor I_24754 (I423877,I710313,I710340);
and I_24755 (I423894,I423742,I423877);
nor I_24756 (I423911,I423829,I423894);
DFFARX1 I_24757 (I423911,I3035,I423518,I423504,);
nor I_24758 (I423942,I423544,I423877);
DFFARX1 I_24759 (I423942,I3035,I423518,I423489,);
nor I_24760 (I423973,I423821,I423877);
not I_24761 (I423990,I423973);
nand I_24762 (I423498,I423990,I423846);
not I_24763 (I424045,I3042);
DFFARX1 I_24764 (I109250,I3035,I424045,I424071,);
not I_24765 (I424079,I424071);
nand I_24766 (I424096,I109247,I109265);
and I_24767 (I424113,I424096,I109256);
DFFARX1 I_24768 (I424113,I3035,I424045,I424139,);
DFFARX1 I_24769 (I424139,I3035,I424045,I424034,);
DFFARX1 I_24770 (I109262,I3035,I424045,I424170,);
nand I_24771 (I424178,I424170,I109259);
not I_24772 (I424195,I424178);
DFFARX1 I_24773 (I424195,I3035,I424045,I424221,);
not I_24774 (I424229,I424221);
nor I_24775 (I424037,I424079,I424229);
DFFARX1 I_24776 (I109253,I3035,I424045,I424269,);
nor I_24777 (I424028,I424269,I424139);
nor I_24778 (I424019,I424269,I424195);
nand I_24779 (I424305,I109244,I109268);
and I_24780 (I424322,I424305,I109247);
DFFARX1 I_24781 (I424322,I3035,I424045,I424348,);
not I_24782 (I424356,I424348);
nand I_24783 (I424373,I424356,I424269);
nand I_24784 (I424022,I424356,I424178);
nor I_24785 (I424404,I109244,I109268);
and I_24786 (I424421,I424269,I424404);
nor I_24787 (I424438,I424356,I424421);
DFFARX1 I_24788 (I424438,I3035,I424045,I424031,);
nor I_24789 (I424469,I424071,I424404);
DFFARX1 I_24790 (I424469,I3035,I424045,I424016,);
nor I_24791 (I424500,I424348,I424404);
not I_24792 (I424517,I424500);
nand I_24793 (I424025,I424517,I424373);
not I_24794 (I424572,I3042);
DFFARX1 I_24795 (I113415,I3035,I424572,I424598,);
not I_24796 (I424606,I424598);
nand I_24797 (I424623,I113412,I113430);
and I_24798 (I424640,I424623,I113421);
DFFARX1 I_24799 (I424640,I3035,I424572,I424666,);
DFFARX1 I_24800 (I424666,I3035,I424572,I424561,);
DFFARX1 I_24801 (I113427,I3035,I424572,I424697,);
nand I_24802 (I424705,I424697,I113424);
not I_24803 (I424722,I424705);
DFFARX1 I_24804 (I424722,I3035,I424572,I424748,);
not I_24805 (I424756,I424748);
nor I_24806 (I424564,I424606,I424756);
DFFARX1 I_24807 (I113418,I3035,I424572,I424796,);
nor I_24808 (I424555,I424796,I424666);
nor I_24809 (I424546,I424796,I424722);
nand I_24810 (I424832,I113409,I113433);
and I_24811 (I424849,I424832,I113412);
DFFARX1 I_24812 (I424849,I3035,I424572,I424875,);
not I_24813 (I424883,I424875);
nand I_24814 (I424900,I424883,I424796);
nand I_24815 (I424549,I424883,I424705);
nor I_24816 (I424931,I113409,I113433);
and I_24817 (I424948,I424796,I424931);
nor I_24818 (I424965,I424883,I424948);
DFFARX1 I_24819 (I424965,I3035,I424572,I424558,);
nor I_24820 (I424996,I424598,I424931);
DFFARX1 I_24821 (I424996,I3035,I424572,I424543,);
nor I_24822 (I425027,I424875,I424931);
not I_24823 (I425044,I425027);
nand I_24824 (I424552,I425044,I424900);
not I_24825 (I425099,I3042);
DFFARX1 I_24826 (I243499,I3035,I425099,I425125,);
not I_24827 (I425133,I425125);
nand I_24828 (I425150,I243496,I243505);
and I_24829 (I425167,I425150,I243514);
DFFARX1 I_24830 (I425167,I3035,I425099,I425193,);
DFFARX1 I_24831 (I425193,I3035,I425099,I425088,);
DFFARX1 I_24832 (I243517,I3035,I425099,I425224,);
nand I_24833 (I425232,I425224,I243520);
not I_24834 (I425249,I425232);
DFFARX1 I_24835 (I425249,I3035,I425099,I425275,);
not I_24836 (I425283,I425275);
nor I_24837 (I425091,I425133,I425283);
DFFARX1 I_24838 (I243493,I3035,I425099,I425323,);
nor I_24839 (I425082,I425323,I425193);
nor I_24840 (I425073,I425323,I425249);
nand I_24841 (I425359,I243508,I243511);
and I_24842 (I425376,I425359,I243502);
DFFARX1 I_24843 (I425376,I3035,I425099,I425402,);
not I_24844 (I425410,I425402);
nand I_24845 (I425427,I425410,I425323);
nand I_24846 (I425076,I425410,I425232);
nor I_24847 (I425458,I243493,I243511);
and I_24848 (I425475,I425323,I425458);
nor I_24849 (I425492,I425410,I425475);
DFFARX1 I_24850 (I425492,I3035,I425099,I425085,);
nor I_24851 (I425523,I425125,I425458);
DFFARX1 I_24852 (I425523,I3035,I425099,I425070,);
nor I_24853 (I425554,I425402,I425458);
not I_24854 (I425571,I425554);
nand I_24855 (I425079,I425571,I425427);
not I_24856 (I425626,I3042);
DFFARX1 I_24857 (I88425,I3035,I425626,I425652,);
not I_24858 (I425660,I425652);
nand I_24859 (I425677,I88422,I88440);
and I_24860 (I425694,I425677,I88431);
DFFARX1 I_24861 (I425694,I3035,I425626,I425720,);
DFFARX1 I_24862 (I425720,I3035,I425626,I425615,);
DFFARX1 I_24863 (I88437,I3035,I425626,I425751,);
nand I_24864 (I425759,I425751,I88434);
not I_24865 (I425776,I425759);
DFFARX1 I_24866 (I425776,I3035,I425626,I425802,);
not I_24867 (I425810,I425802);
nor I_24868 (I425618,I425660,I425810);
DFFARX1 I_24869 (I88428,I3035,I425626,I425850,);
nor I_24870 (I425609,I425850,I425720);
nor I_24871 (I425600,I425850,I425776);
nand I_24872 (I425886,I88419,I88443);
and I_24873 (I425903,I425886,I88422);
DFFARX1 I_24874 (I425903,I3035,I425626,I425929,);
not I_24875 (I425937,I425929);
nand I_24876 (I425954,I425937,I425850);
nand I_24877 (I425603,I425937,I425759);
nor I_24878 (I425985,I88419,I88443);
and I_24879 (I426002,I425850,I425985);
nor I_24880 (I426019,I425937,I426002);
DFFARX1 I_24881 (I426019,I3035,I425626,I425612,);
nor I_24882 (I426050,I425652,I425985);
DFFARX1 I_24883 (I426050,I3035,I425626,I425597,);
nor I_24884 (I426081,I425929,I425985);
not I_24885 (I426098,I426081);
nand I_24886 (I425606,I426098,I425954);
not I_24887 (I426153,I3042);
DFFARX1 I_24888 (I397836,I3035,I426153,I426179,);
not I_24889 (I426187,I426179);
nand I_24890 (I426204,I397839,I397836);
and I_24891 (I426221,I426204,I397848);
DFFARX1 I_24892 (I426221,I3035,I426153,I426247,);
DFFARX1 I_24893 (I426247,I3035,I426153,I426142,);
DFFARX1 I_24894 (I397845,I3035,I426153,I426278,);
nand I_24895 (I426286,I426278,I397851);
not I_24896 (I426303,I426286);
DFFARX1 I_24897 (I426303,I3035,I426153,I426329,);
not I_24898 (I426337,I426329);
nor I_24899 (I426145,I426187,I426337);
DFFARX1 I_24900 (I397860,I3035,I426153,I426377,);
nor I_24901 (I426136,I426377,I426247);
nor I_24902 (I426127,I426377,I426303);
nand I_24903 (I426413,I397854,I397842);
and I_24904 (I426430,I426413,I397839);
DFFARX1 I_24905 (I426430,I3035,I426153,I426456,);
not I_24906 (I426464,I426456);
nand I_24907 (I426481,I426464,I426377);
nand I_24908 (I426130,I426464,I426286);
nor I_24909 (I426512,I397857,I397842);
and I_24910 (I426529,I426377,I426512);
nor I_24911 (I426546,I426464,I426529);
DFFARX1 I_24912 (I426546,I3035,I426153,I426139,);
nor I_24913 (I426577,I426179,I426512);
DFFARX1 I_24914 (I426577,I3035,I426153,I426124,);
nor I_24915 (I426608,I426456,I426512);
not I_24916 (I426625,I426608);
nand I_24917 (I426133,I426625,I426481);
not I_24918 (I426680,I3042);
DFFARX1 I_24919 (I89020,I3035,I426680,I426706,);
not I_24920 (I426714,I426706);
nand I_24921 (I426731,I89017,I89035);
and I_24922 (I426748,I426731,I89026);
DFFARX1 I_24923 (I426748,I3035,I426680,I426774,);
DFFARX1 I_24924 (I426774,I3035,I426680,I426669,);
DFFARX1 I_24925 (I89032,I3035,I426680,I426805,);
nand I_24926 (I426813,I426805,I89029);
not I_24927 (I426830,I426813);
DFFARX1 I_24928 (I426830,I3035,I426680,I426856,);
not I_24929 (I426864,I426856);
nor I_24930 (I426672,I426714,I426864);
DFFARX1 I_24931 (I89023,I3035,I426680,I426904,);
nor I_24932 (I426663,I426904,I426774);
nor I_24933 (I426654,I426904,I426830);
nand I_24934 (I426940,I89014,I89038);
and I_24935 (I426957,I426940,I89017);
DFFARX1 I_24936 (I426957,I3035,I426680,I426983,);
not I_24937 (I426991,I426983);
nand I_24938 (I427008,I426991,I426904);
nand I_24939 (I426657,I426991,I426813);
nor I_24940 (I427039,I89014,I89038);
and I_24941 (I427056,I426904,I427039);
nor I_24942 (I427073,I426991,I427056);
DFFARX1 I_24943 (I427073,I3035,I426680,I426666,);
nor I_24944 (I427104,I426706,I427039);
DFFARX1 I_24945 (I427104,I3035,I426680,I426651,);
nor I_24946 (I427135,I426983,I427039);
not I_24947 (I427152,I427135);
nand I_24948 (I426660,I427152,I427008);
not I_24949 (I427207,I3042);
DFFARX1 I_24950 (I580400,I3035,I427207,I427233,);
not I_24951 (I427241,I427233);
nand I_24952 (I427258,I580382,I580382);
and I_24953 (I427275,I427258,I580388);
DFFARX1 I_24954 (I427275,I3035,I427207,I427301,);
DFFARX1 I_24955 (I427301,I3035,I427207,I427196,);
DFFARX1 I_24956 (I580385,I3035,I427207,I427332,);
nand I_24957 (I427340,I427332,I580394);
not I_24958 (I427357,I427340);
DFFARX1 I_24959 (I427357,I3035,I427207,I427383,);
not I_24960 (I427391,I427383);
nor I_24961 (I427199,I427241,I427391);
DFFARX1 I_24962 (I580406,I3035,I427207,I427431,);
nor I_24963 (I427190,I427431,I427301);
nor I_24964 (I427181,I427431,I427357);
nand I_24965 (I427467,I580397,I580391);
and I_24966 (I427484,I427467,I580385);
DFFARX1 I_24967 (I427484,I3035,I427207,I427510,);
not I_24968 (I427518,I427510);
nand I_24969 (I427535,I427518,I427431);
nand I_24970 (I427184,I427518,I427340);
nor I_24971 (I427566,I580403,I580391);
and I_24972 (I427583,I427431,I427566);
nor I_24973 (I427600,I427518,I427583);
DFFARX1 I_24974 (I427600,I3035,I427207,I427193,);
nor I_24975 (I427631,I427233,I427566);
DFFARX1 I_24976 (I427631,I3035,I427207,I427178,);
nor I_24977 (I427662,I427510,I427566);
not I_24978 (I427679,I427662);
nand I_24979 (I427187,I427679,I427535);
not I_24980 (I427734,I3042);
DFFARX1 I_24981 (I85450,I3035,I427734,I427760,);
not I_24982 (I427768,I427760);
nand I_24983 (I427785,I85447,I85465);
and I_24984 (I427802,I427785,I85456);
DFFARX1 I_24985 (I427802,I3035,I427734,I427828,);
DFFARX1 I_24986 (I427828,I3035,I427734,I427723,);
DFFARX1 I_24987 (I85462,I3035,I427734,I427859,);
nand I_24988 (I427867,I427859,I85459);
not I_24989 (I427884,I427867);
DFFARX1 I_24990 (I427884,I3035,I427734,I427910,);
not I_24991 (I427918,I427910);
nor I_24992 (I427726,I427768,I427918);
DFFARX1 I_24993 (I85453,I3035,I427734,I427958,);
nor I_24994 (I427717,I427958,I427828);
nor I_24995 (I427708,I427958,I427884);
nand I_24996 (I427994,I85444,I85468);
and I_24997 (I428011,I427994,I85447);
DFFARX1 I_24998 (I428011,I3035,I427734,I428037,);
not I_24999 (I428045,I428037);
nand I_25000 (I428062,I428045,I427958);
nand I_25001 (I427711,I428045,I427867);
nor I_25002 (I428093,I85444,I85468);
and I_25003 (I428110,I427958,I428093);
nor I_25004 (I428127,I428045,I428110);
DFFARX1 I_25005 (I428127,I3035,I427734,I427720,);
nor I_25006 (I428158,I427760,I428093);
DFFARX1 I_25007 (I428158,I3035,I427734,I427705,);
nor I_25008 (I428189,I428037,I428093);
not I_25009 (I428206,I428189);
nand I_25010 (I427714,I428206,I428062);
not I_25011 (I428261,I3042);
DFFARX1 I_25012 (I262539,I3035,I428261,I428287,);
not I_25013 (I428295,I428287);
nand I_25014 (I428312,I262536,I262545);
and I_25015 (I428329,I428312,I262554);
DFFARX1 I_25016 (I428329,I3035,I428261,I428355,);
DFFARX1 I_25017 (I428355,I3035,I428261,I428250,);
DFFARX1 I_25018 (I262557,I3035,I428261,I428386,);
nand I_25019 (I428394,I428386,I262560);
not I_25020 (I428411,I428394);
DFFARX1 I_25021 (I428411,I3035,I428261,I428437,);
not I_25022 (I428445,I428437);
nor I_25023 (I428253,I428295,I428445);
DFFARX1 I_25024 (I262533,I3035,I428261,I428485,);
nor I_25025 (I428244,I428485,I428355);
nor I_25026 (I428235,I428485,I428411);
nand I_25027 (I428521,I262548,I262551);
and I_25028 (I428538,I428521,I262542);
DFFARX1 I_25029 (I428538,I3035,I428261,I428564,);
not I_25030 (I428572,I428564);
nand I_25031 (I428589,I428572,I428485);
nand I_25032 (I428238,I428572,I428394);
nor I_25033 (I428620,I262533,I262551);
and I_25034 (I428637,I428485,I428620);
nor I_25035 (I428654,I428572,I428637);
DFFARX1 I_25036 (I428654,I3035,I428261,I428247,);
nor I_25037 (I428685,I428287,I428620);
DFFARX1 I_25038 (I428685,I3035,I428261,I428232,);
nor I_25039 (I428716,I428564,I428620);
not I_25040 (I428733,I428716);
nand I_25041 (I428241,I428733,I428589);
not I_25042 (I428788,I3042);
DFFARX1 I_25043 (I595428,I3035,I428788,I428814,);
not I_25044 (I428822,I428814);
nand I_25045 (I428839,I595410,I595410);
and I_25046 (I428856,I428839,I595416);
DFFARX1 I_25047 (I428856,I3035,I428788,I428882,);
DFFARX1 I_25048 (I428882,I3035,I428788,I428777,);
DFFARX1 I_25049 (I595413,I3035,I428788,I428913,);
nand I_25050 (I428921,I428913,I595422);
not I_25051 (I428938,I428921);
DFFARX1 I_25052 (I428938,I3035,I428788,I428964,);
not I_25053 (I428972,I428964);
nor I_25054 (I428780,I428822,I428972);
DFFARX1 I_25055 (I595434,I3035,I428788,I429012,);
nor I_25056 (I428771,I429012,I428882);
nor I_25057 (I428762,I429012,I428938);
nand I_25058 (I429048,I595425,I595419);
and I_25059 (I429065,I429048,I595413);
DFFARX1 I_25060 (I429065,I3035,I428788,I429091,);
not I_25061 (I429099,I429091);
nand I_25062 (I429116,I429099,I429012);
nand I_25063 (I428765,I429099,I428921);
nor I_25064 (I429147,I595431,I595419);
and I_25065 (I429164,I429012,I429147);
nor I_25066 (I429181,I429099,I429164);
DFFARX1 I_25067 (I429181,I3035,I428788,I428774,);
nor I_25068 (I429212,I428814,I429147);
DFFARX1 I_25069 (I429212,I3035,I428788,I428759,);
nor I_25070 (I429243,I429091,I429147);
not I_25071 (I429260,I429243);
nand I_25072 (I428768,I429260,I429116);
not I_25073 (I429315,I3042);
DFFARX1 I_25074 (I338302,I3035,I429315,I429341,);
not I_25075 (I429349,I429341);
nand I_25076 (I429366,I338305,I338302);
and I_25077 (I429383,I429366,I338314);
DFFARX1 I_25078 (I429383,I3035,I429315,I429409,);
DFFARX1 I_25079 (I429409,I3035,I429315,I429304,);
DFFARX1 I_25080 (I338311,I3035,I429315,I429440,);
nand I_25081 (I429448,I429440,I338317);
not I_25082 (I429465,I429448);
DFFARX1 I_25083 (I429465,I3035,I429315,I429491,);
not I_25084 (I429499,I429491);
nor I_25085 (I429307,I429349,I429499);
DFFARX1 I_25086 (I338326,I3035,I429315,I429539,);
nor I_25087 (I429298,I429539,I429409);
nor I_25088 (I429289,I429539,I429465);
nand I_25089 (I429575,I338320,I338308);
and I_25090 (I429592,I429575,I338305);
DFFARX1 I_25091 (I429592,I3035,I429315,I429618,);
not I_25092 (I429626,I429618);
nand I_25093 (I429643,I429626,I429539);
nand I_25094 (I429292,I429626,I429448);
nor I_25095 (I429674,I338323,I338308);
and I_25096 (I429691,I429539,I429674);
nor I_25097 (I429708,I429626,I429691);
DFFARX1 I_25098 (I429708,I3035,I429315,I429301,);
nor I_25099 (I429739,I429341,I429674);
DFFARX1 I_25100 (I429739,I3035,I429315,I429286,);
nor I_25101 (I429770,I429618,I429674);
not I_25102 (I429787,I429770);
nand I_25103 (I429295,I429787,I429643);
not I_25104 (I429842,I3042);
DFFARX1 I_25105 (I590804,I3035,I429842,I429868,);
not I_25106 (I429876,I429868);
nand I_25107 (I429893,I590786,I590786);
and I_25108 (I429910,I429893,I590792);
DFFARX1 I_25109 (I429910,I3035,I429842,I429936,);
DFFARX1 I_25110 (I429936,I3035,I429842,I429831,);
DFFARX1 I_25111 (I590789,I3035,I429842,I429967,);
nand I_25112 (I429975,I429967,I590798);
not I_25113 (I429992,I429975);
DFFARX1 I_25114 (I429992,I3035,I429842,I430018,);
not I_25115 (I430026,I430018);
nor I_25116 (I429834,I429876,I430026);
DFFARX1 I_25117 (I590810,I3035,I429842,I430066,);
nor I_25118 (I429825,I430066,I429936);
nor I_25119 (I429816,I430066,I429992);
nand I_25120 (I430102,I590801,I590795);
and I_25121 (I430119,I430102,I590789);
DFFARX1 I_25122 (I430119,I3035,I429842,I430145,);
not I_25123 (I430153,I430145);
nand I_25124 (I430170,I430153,I430066);
nand I_25125 (I429819,I430153,I429975);
nor I_25126 (I430201,I590807,I590795);
and I_25127 (I430218,I430066,I430201);
nor I_25128 (I430235,I430153,I430218);
DFFARX1 I_25129 (I430235,I3035,I429842,I429828,);
nor I_25130 (I430266,I429868,I430201);
DFFARX1 I_25131 (I430266,I3035,I429842,I429813,);
nor I_25132 (I430297,I430145,I430201);
not I_25133 (I430314,I430297);
nand I_25134 (I429822,I430314,I430170);
not I_25135 (I430369,I3042);
DFFARX1 I_25136 (I140190,I3035,I430369,I430395,);
not I_25137 (I430403,I430395);
nand I_25138 (I430420,I140187,I140205);
and I_25139 (I430437,I430420,I140196);
DFFARX1 I_25140 (I430437,I3035,I430369,I430463,);
DFFARX1 I_25141 (I430463,I3035,I430369,I430358,);
DFFARX1 I_25142 (I140202,I3035,I430369,I430494,);
nand I_25143 (I430502,I430494,I140199);
not I_25144 (I430519,I430502);
DFFARX1 I_25145 (I430519,I3035,I430369,I430545,);
not I_25146 (I430553,I430545);
nor I_25147 (I430361,I430403,I430553);
DFFARX1 I_25148 (I140193,I3035,I430369,I430593,);
nor I_25149 (I430352,I430593,I430463);
nor I_25150 (I430343,I430593,I430519);
nand I_25151 (I430629,I140184,I140208);
and I_25152 (I430646,I430629,I140187);
DFFARX1 I_25153 (I430646,I3035,I430369,I430672,);
not I_25154 (I430680,I430672);
nand I_25155 (I430697,I430680,I430593);
nand I_25156 (I430346,I430680,I430502);
nor I_25157 (I430728,I140184,I140208);
and I_25158 (I430745,I430593,I430728);
nor I_25159 (I430762,I430680,I430745);
DFFARX1 I_25160 (I430762,I3035,I430369,I430355,);
nor I_25161 (I430793,I430395,I430728);
DFFARX1 I_25162 (I430793,I3035,I430369,I430340,);
nor I_25163 (I430824,I430672,I430728);
not I_25164 (I430841,I430824);
nand I_25165 (I430349,I430841,I430697);
not I_25166 (I430896,I3042);
DFFARX1 I_25167 (I556030,I3035,I430896,I430922,);
not I_25168 (I430930,I430922);
nand I_25169 (I430947,I556039,I556027);
and I_25170 (I430964,I430947,I556024);
DFFARX1 I_25171 (I430964,I3035,I430896,I430990,);
DFFARX1 I_25172 (I430990,I3035,I430896,I430885,);
DFFARX1 I_25173 (I556024,I3035,I430896,I431021,);
nand I_25174 (I431029,I431021,I556021);
not I_25175 (I431046,I431029);
DFFARX1 I_25176 (I431046,I3035,I430896,I431072,);
not I_25177 (I431080,I431072);
nor I_25178 (I430888,I430930,I431080);
DFFARX1 I_25179 (I556027,I3035,I430896,I431120,);
nor I_25180 (I430879,I431120,I430990);
nor I_25181 (I430870,I431120,I431046);
nand I_25182 (I431156,I556042,I556033);
and I_25183 (I431173,I431156,I556036);
DFFARX1 I_25184 (I431173,I3035,I430896,I431199,);
not I_25185 (I431207,I431199);
nand I_25186 (I431224,I431207,I431120);
nand I_25187 (I430873,I431207,I431029);
nor I_25188 (I431255,I556021,I556033);
and I_25189 (I431272,I431120,I431255);
nor I_25190 (I431289,I431207,I431272);
DFFARX1 I_25191 (I431289,I3035,I430896,I430882,);
nor I_25192 (I431320,I430922,I431255);
DFFARX1 I_25193 (I431320,I3035,I430896,I430867,);
nor I_25194 (I431351,I431199,I431255);
not I_25195 (I431368,I431351);
nand I_25196 (I430876,I431368,I431224);
not I_25197 (I431423,I3042);
DFFARX1 I_25198 (I33652,I3035,I431423,I431449,);
not I_25199 (I431457,I431449);
nand I_25200 (I431474,I33628,I33637);
and I_25201 (I431491,I431474,I33631);
DFFARX1 I_25202 (I431491,I3035,I431423,I431517,);
DFFARX1 I_25203 (I431517,I3035,I431423,I431412,);
DFFARX1 I_25204 (I33649,I3035,I431423,I431548,);
nand I_25205 (I431556,I431548,I33640);
not I_25206 (I431573,I431556);
DFFARX1 I_25207 (I431573,I3035,I431423,I431599,);
not I_25208 (I431607,I431599);
nor I_25209 (I431415,I431457,I431607);
DFFARX1 I_25210 (I33634,I3035,I431423,I431647,);
nor I_25211 (I431406,I431647,I431517);
nor I_25212 (I431397,I431647,I431573);
nand I_25213 (I431683,I33646,I33643);
and I_25214 (I431700,I431683,I33631);
DFFARX1 I_25215 (I431700,I3035,I431423,I431726,);
not I_25216 (I431734,I431726);
nand I_25217 (I431751,I431734,I431647);
nand I_25218 (I431400,I431734,I431556);
nor I_25219 (I431782,I33628,I33643);
and I_25220 (I431799,I431647,I431782);
nor I_25221 (I431816,I431734,I431799);
DFFARX1 I_25222 (I431816,I3035,I431423,I431409,);
nor I_25223 (I431847,I431449,I431782);
DFFARX1 I_25224 (I431847,I3035,I431423,I431394,);
nor I_25225 (I431878,I431726,I431782);
not I_25226 (I431895,I431878);
nand I_25227 (I431403,I431895,I431751);
not I_25228 (I431950,I3042);
DFFARX1 I_25229 (I182982,I3035,I431950,I431976,);
not I_25230 (I431984,I431976);
nand I_25231 (I432001,I182973,I182973);
and I_25232 (I432018,I432001,I182991);
DFFARX1 I_25233 (I432018,I3035,I431950,I432044,);
DFFARX1 I_25234 (I432044,I3035,I431950,I431939,);
DFFARX1 I_25235 (I182994,I3035,I431950,I432075,);
nand I_25236 (I432083,I432075,I182976);
not I_25237 (I432100,I432083);
DFFARX1 I_25238 (I432100,I3035,I431950,I432126,);
not I_25239 (I432134,I432126);
nor I_25240 (I431942,I431984,I432134);
DFFARX1 I_25241 (I182988,I3035,I431950,I432174,);
nor I_25242 (I431933,I432174,I432044);
nor I_25243 (I431924,I432174,I432100);
nand I_25244 (I432210,I183000,I182979);
and I_25245 (I432227,I432210,I182985);
DFFARX1 I_25246 (I432227,I3035,I431950,I432253,);
not I_25247 (I432261,I432253);
nand I_25248 (I432278,I432261,I432174);
nand I_25249 (I431927,I432261,I432083);
nor I_25250 (I432309,I182997,I182979);
and I_25251 (I432326,I432174,I432309);
nor I_25252 (I432343,I432261,I432326);
DFFARX1 I_25253 (I432343,I3035,I431950,I431936,);
nor I_25254 (I432374,I431976,I432309);
DFFARX1 I_25255 (I432374,I3035,I431950,I431921,);
nor I_25256 (I432405,I432253,I432309);
not I_25257 (I432422,I432405);
nand I_25258 (I431930,I432422,I432278);
not I_25259 (I432477,I3042);
DFFARX1 I_25260 (I727583,I3035,I432477,I432503,);
not I_25261 (I432511,I432503);
nand I_25262 (I432528,I727580,I727589);
and I_25263 (I432545,I432528,I727568);
DFFARX1 I_25264 (I432545,I3035,I432477,I432571,);
DFFARX1 I_25265 (I432571,I3035,I432477,I432466,);
DFFARX1 I_25266 (I727571,I3035,I432477,I432602,);
nand I_25267 (I432610,I432602,I727586);
not I_25268 (I432627,I432610);
DFFARX1 I_25269 (I432627,I3035,I432477,I432653,);
not I_25270 (I432661,I432653);
nor I_25271 (I432469,I432511,I432661);
DFFARX1 I_25272 (I727592,I3035,I432477,I432701,);
nor I_25273 (I432460,I432701,I432571);
nor I_25274 (I432451,I432701,I432627);
nand I_25275 (I432737,I727574,I727595);
and I_25276 (I432754,I432737,I727577);
DFFARX1 I_25277 (I432754,I3035,I432477,I432780,);
not I_25278 (I432788,I432780);
nand I_25279 (I432805,I432788,I432701);
nand I_25280 (I432454,I432788,I432610);
nor I_25281 (I432836,I727568,I727595);
and I_25282 (I432853,I432701,I432836);
nor I_25283 (I432870,I432788,I432853);
DFFARX1 I_25284 (I432870,I3035,I432477,I432463,);
nor I_25285 (I432901,I432503,I432836);
DFFARX1 I_25286 (I432901,I3035,I432477,I432448,);
nor I_25287 (I432932,I432780,I432836);
not I_25288 (I432949,I432932);
nand I_25289 (I432457,I432949,I432805);
not I_25290 (I433004,I3042);
DFFARX1 I_25291 (I696668,I3035,I433004,I433030,);
not I_25292 (I433038,I433030);
nand I_25293 (I433055,I696662,I696680);
and I_25294 (I433072,I433055,I696665);
DFFARX1 I_25295 (I433072,I3035,I433004,I433098,);
DFFARX1 I_25296 (I433098,I3035,I433004,I432993,);
DFFARX1 I_25297 (I696686,I3035,I433004,I433129,);
nand I_25298 (I433137,I433129,I696671);
not I_25299 (I433154,I433137);
DFFARX1 I_25300 (I433154,I3035,I433004,I433180,);
not I_25301 (I433188,I433180);
nor I_25302 (I432996,I433038,I433188);
DFFARX1 I_25303 (I696683,I3035,I433004,I433228,);
nor I_25304 (I432987,I433228,I433098);
nor I_25305 (I432978,I433228,I433154);
nand I_25306 (I433264,I696674,I696689);
and I_25307 (I433281,I433264,I696677);
DFFARX1 I_25308 (I433281,I3035,I433004,I433307,);
not I_25309 (I433315,I433307);
nand I_25310 (I433332,I433315,I433228);
nand I_25311 (I432981,I433315,I433137);
nor I_25312 (I433363,I696662,I696689);
and I_25313 (I433380,I433228,I433363);
nor I_25314 (I433397,I433315,I433380);
DFFARX1 I_25315 (I433397,I3035,I433004,I432990,);
nor I_25316 (I433428,I433030,I433363);
DFFARX1 I_25317 (I433428,I3035,I433004,I432975,);
nor I_25318 (I433459,I433307,I433363);
not I_25319 (I433476,I433459);
nand I_25320 (I432984,I433476,I433332);
not I_25321 (I433531,I3042);
DFFARX1 I_25322 (I340036,I3035,I433531,I433557,);
not I_25323 (I433565,I433557);
nand I_25324 (I433582,I340039,I340036);
and I_25325 (I433599,I433582,I340048);
DFFARX1 I_25326 (I433599,I3035,I433531,I433625,);
DFFARX1 I_25327 (I433625,I3035,I433531,I433520,);
DFFARX1 I_25328 (I340045,I3035,I433531,I433656,);
nand I_25329 (I433664,I433656,I340051);
not I_25330 (I433681,I433664);
DFFARX1 I_25331 (I433681,I3035,I433531,I433707,);
not I_25332 (I433715,I433707);
nor I_25333 (I433523,I433565,I433715);
DFFARX1 I_25334 (I340060,I3035,I433531,I433755,);
nor I_25335 (I433514,I433755,I433625);
nor I_25336 (I433505,I433755,I433681);
nand I_25337 (I433791,I340054,I340042);
and I_25338 (I433808,I433791,I340039);
DFFARX1 I_25339 (I433808,I3035,I433531,I433834,);
not I_25340 (I433842,I433834);
nand I_25341 (I433859,I433842,I433755);
nand I_25342 (I433508,I433842,I433664);
nor I_25343 (I433890,I340057,I340042);
and I_25344 (I433907,I433755,I433890);
nor I_25345 (I433924,I433842,I433907);
DFFARX1 I_25346 (I433924,I3035,I433531,I433517,);
nor I_25347 (I433955,I433557,I433890);
DFFARX1 I_25348 (I433955,I3035,I433531,I433502,);
nor I_25349 (I433986,I433834,I433890);
not I_25350 (I434003,I433986);
nand I_25351 (I433511,I434003,I433859);
not I_25352 (I434058,I3042);
DFFARX1 I_25353 (I586758,I3035,I434058,I434084,);
not I_25354 (I434092,I434084);
nand I_25355 (I434109,I586740,I586740);
and I_25356 (I434126,I434109,I586746);
DFFARX1 I_25357 (I434126,I3035,I434058,I434152,);
DFFARX1 I_25358 (I434152,I3035,I434058,I434047,);
DFFARX1 I_25359 (I586743,I3035,I434058,I434183,);
nand I_25360 (I434191,I434183,I586752);
not I_25361 (I434208,I434191);
DFFARX1 I_25362 (I434208,I3035,I434058,I434234,);
not I_25363 (I434242,I434234);
nor I_25364 (I434050,I434092,I434242);
DFFARX1 I_25365 (I586764,I3035,I434058,I434282,);
nor I_25366 (I434041,I434282,I434152);
nor I_25367 (I434032,I434282,I434208);
nand I_25368 (I434318,I586755,I586749);
and I_25369 (I434335,I434318,I586743);
DFFARX1 I_25370 (I434335,I3035,I434058,I434361,);
not I_25371 (I434369,I434361);
nand I_25372 (I434386,I434369,I434282);
nand I_25373 (I434035,I434369,I434191);
nor I_25374 (I434417,I586761,I586749);
and I_25375 (I434434,I434282,I434417);
nor I_25376 (I434451,I434369,I434434);
DFFARX1 I_25377 (I434451,I3035,I434058,I434044,);
nor I_25378 (I434482,I434084,I434417);
DFFARX1 I_25379 (I434482,I3035,I434058,I434029,);
nor I_25380 (I434513,I434361,I434417);
not I_25381 (I434530,I434513);
nand I_25382 (I434038,I434530,I434386);
not I_25383 (I434585,I3042);
DFFARX1 I_25384 (I736508,I3035,I434585,I434611,);
not I_25385 (I434619,I434611);
nand I_25386 (I434636,I736505,I736514);
and I_25387 (I434653,I434636,I736493);
DFFARX1 I_25388 (I434653,I3035,I434585,I434679,);
DFFARX1 I_25389 (I434679,I3035,I434585,I434574,);
DFFARX1 I_25390 (I736496,I3035,I434585,I434710,);
nand I_25391 (I434718,I434710,I736511);
not I_25392 (I434735,I434718);
DFFARX1 I_25393 (I434735,I3035,I434585,I434761,);
not I_25394 (I434769,I434761);
nor I_25395 (I434577,I434619,I434769);
DFFARX1 I_25396 (I736517,I3035,I434585,I434809,);
nor I_25397 (I434568,I434809,I434679);
nor I_25398 (I434559,I434809,I434735);
nand I_25399 (I434845,I736499,I736520);
and I_25400 (I434862,I434845,I736502);
DFFARX1 I_25401 (I434862,I3035,I434585,I434888,);
not I_25402 (I434896,I434888);
nand I_25403 (I434913,I434896,I434809);
nand I_25404 (I434562,I434896,I434718);
nor I_25405 (I434944,I736493,I736520);
and I_25406 (I434961,I434809,I434944);
nor I_25407 (I434978,I434896,I434961);
DFFARX1 I_25408 (I434978,I3035,I434585,I434571,);
nor I_25409 (I435009,I434611,I434944);
DFFARX1 I_25410 (I435009,I3035,I434585,I434556,);
nor I_25411 (I435040,I434888,I434944);
not I_25412 (I435057,I435040);
nand I_25413 (I434565,I435057,I434913);
not I_25414 (I435112,I3042);
DFFARX1 I_25415 (I514187,I3035,I435112,I435138,);
not I_25416 (I435146,I435138);
nand I_25417 (I435163,I514202,I514184);
and I_25418 (I435180,I435163,I514184);
DFFARX1 I_25419 (I435180,I3035,I435112,I435206,);
DFFARX1 I_25420 (I435206,I3035,I435112,I435101,);
DFFARX1 I_25421 (I514193,I3035,I435112,I435237,);
nand I_25422 (I435245,I435237,I514211);
not I_25423 (I435262,I435245);
DFFARX1 I_25424 (I435262,I3035,I435112,I435288,);
not I_25425 (I435296,I435288);
nor I_25426 (I435104,I435146,I435296);
DFFARX1 I_25427 (I514208,I3035,I435112,I435336,);
nor I_25428 (I435095,I435336,I435206);
nor I_25429 (I435086,I435336,I435262);
nand I_25430 (I435372,I514205,I514196);
and I_25431 (I435389,I435372,I514190);
DFFARX1 I_25432 (I435389,I3035,I435112,I435415,);
not I_25433 (I435423,I435415);
nand I_25434 (I435440,I435423,I435336);
nand I_25435 (I435089,I435423,I435245);
nor I_25436 (I435471,I514199,I514196);
and I_25437 (I435488,I435336,I435471);
nor I_25438 (I435505,I435423,I435488);
DFFARX1 I_25439 (I435505,I3035,I435112,I435098,);
nor I_25440 (I435536,I435138,I435471);
DFFARX1 I_25441 (I435536,I3035,I435112,I435083,);
nor I_25442 (I435567,I435415,I435471);
not I_25443 (I435584,I435567);
nand I_25444 (I435092,I435584,I435440);
not I_25445 (I435639,I3042);
DFFARX1 I_25446 (I256011,I3035,I435639,I435665,);
not I_25447 (I435673,I435665);
nand I_25448 (I435690,I256008,I256017);
and I_25449 (I435707,I435690,I256026);
DFFARX1 I_25450 (I435707,I3035,I435639,I435733,);
DFFARX1 I_25451 (I435733,I3035,I435639,I435628,);
DFFARX1 I_25452 (I256029,I3035,I435639,I435764,);
nand I_25453 (I435772,I435764,I256032);
not I_25454 (I435789,I435772);
DFFARX1 I_25455 (I435789,I3035,I435639,I435815,);
not I_25456 (I435823,I435815);
nor I_25457 (I435631,I435673,I435823);
DFFARX1 I_25458 (I256005,I3035,I435639,I435863,);
nor I_25459 (I435622,I435863,I435733);
nor I_25460 (I435613,I435863,I435789);
nand I_25461 (I435899,I256020,I256023);
and I_25462 (I435916,I435899,I256014);
DFFARX1 I_25463 (I435916,I3035,I435639,I435942,);
not I_25464 (I435950,I435942);
nand I_25465 (I435967,I435950,I435863);
nand I_25466 (I435616,I435950,I435772);
nor I_25467 (I435998,I256005,I256023);
and I_25468 (I436015,I435863,I435998);
nor I_25469 (I436032,I435950,I436015);
DFFARX1 I_25470 (I436032,I3035,I435639,I435625,);
nor I_25471 (I436063,I435665,I435998);
DFFARX1 I_25472 (I436063,I3035,I435639,I435610,);
nor I_25473 (I436094,I435942,I435998);
not I_25474 (I436111,I436094);
nand I_25475 (I435619,I436111,I435967);
not I_25476 (I436166,I3042);
DFFARX1 I_25477 (I125315,I3035,I436166,I436192,);
not I_25478 (I436200,I436192);
nand I_25479 (I436217,I125312,I125330);
and I_25480 (I436234,I436217,I125321);
DFFARX1 I_25481 (I436234,I3035,I436166,I436260,);
DFFARX1 I_25482 (I436260,I3035,I436166,I436155,);
DFFARX1 I_25483 (I125327,I3035,I436166,I436291,);
nand I_25484 (I436299,I436291,I125324);
not I_25485 (I436316,I436299);
DFFARX1 I_25486 (I436316,I3035,I436166,I436342,);
not I_25487 (I436350,I436342);
nor I_25488 (I436158,I436200,I436350);
DFFARX1 I_25489 (I125318,I3035,I436166,I436390,);
nor I_25490 (I436149,I436390,I436260);
nor I_25491 (I436140,I436390,I436316);
nand I_25492 (I436426,I125309,I125333);
and I_25493 (I436443,I436426,I125312);
DFFARX1 I_25494 (I436443,I3035,I436166,I436469,);
not I_25495 (I436477,I436469);
nand I_25496 (I436494,I436477,I436390);
nand I_25497 (I436143,I436477,I436299);
nor I_25498 (I436525,I125309,I125333);
and I_25499 (I436542,I436390,I436525);
nor I_25500 (I436559,I436477,I436542);
DFFARX1 I_25501 (I436559,I3035,I436166,I436152,);
nor I_25502 (I436590,I436192,I436525);
DFFARX1 I_25503 (I436590,I3035,I436166,I436137,);
nor I_25504 (I436621,I436469,I436525);
not I_25505 (I436638,I436621);
nand I_25506 (I436146,I436638,I436494);
not I_25507 (I436693,I3042);
DFFARX1 I_25508 (I81880,I3035,I436693,I436719,);
not I_25509 (I436727,I436719);
nand I_25510 (I436744,I81877,I81895);
and I_25511 (I436761,I436744,I81886);
DFFARX1 I_25512 (I436761,I3035,I436693,I436787,);
DFFARX1 I_25513 (I436787,I3035,I436693,I436682,);
DFFARX1 I_25514 (I81892,I3035,I436693,I436818,);
nand I_25515 (I436826,I436818,I81889);
not I_25516 (I436843,I436826);
DFFARX1 I_25517 (I436843,I3035,I436693,I436869,);
not I_25518 (I436877,I436869);
nor I_25519 (I436685,I436727,I436877);
DFFARX1 I_25520 (I81883,I3035,I436693,I436917,);
nor I_25521 (I436676,I436917,I436787);
nor I_25522 (I436667,I436917,I436843);
nand I_25523 (I436953,I81874,I81898);
and I_25524 (I436970,I436953,I81877);
DFFARX1 I_25525 (I436970,I3035,I436693,I436996,);
not I_25526 (I437004,I436996);
nand I_25527 (I437021,I437004,I436917);
nand I_25528 (I436670,I437004,I436826);
nor I_25529 (I437052,I81874,I81898);
and I_25530 (I437069,I436917,I437052);
nor I_25531 (I437086,I437004,I437069);
DFFARX1 I_25532 (I437086,I3035,I436693,I436679,);
nor I_25533 (I437117,I436719,I437052);
DFFARX1 I_25534 (I437117,I3035,I436693,I436664,);
nor I_25535 (I437148,I436996,I437052);
not I_25536 (I437165,I437148);
nand I_25537 (I436673,I437165,I437021);
not I_25538 (I437220,I3042);
DFFARX1 I_25539 (I476719,I3035,I437220,I437246,);
not I_25540 (I437254,I437246);
nand I_25541 (I437271,I476734,I476716);
and I_25542 (I437288,I437271,I476716);
DFFARX1 I_25543 (I437288,I3035,I437220,I437314,);
DFFARX1 I_25544 (I437314,I3035,I437220,I437209,);
DFFARX1 I_25545 (I476725,I3035,I437220,I437345,);
nand I_25546 (I437353,I437345,I476743);
not I_25547 (I437370,I437353);
DFFARX1 I_25548 (I437370,I3035,I437220,I437396,);
not I_25549 (I437404,I437396);
nor I_25550 (I437212,I437254,I437404);
DFFARX1 I_25551 (I476740,I3035,I437220,I437444,);
nor I_25552 (I437203,I437444,I437314);
nor I_25553 (I437194,I437444,I437370);
nand I_25554 (I437480,I476737,I476728);
and I_25555 (I437497,I437480,I476722);
DFFARX1 I_25556 (I437497,I3035,I437220,I437523,);
not I_25557 (I437531,I437523);
nand I_25558 (I437548,I437531,I437444);
nand I_25559 (I437197,I437531,I437353);
nor I_25560 (I437579,I476731,I476728);
and I_25561 (I437596,I437444,I437579);
nor I_25562 (I437613,I437531,I437596);
DFFARX1 I_25563 (I437613,I3035,I437220,I437206,);
nor I_25564 (I437644,I437246,I437579);
DFFARX1 I_25565 (I437644,I3035,I437220,I437191,);
nor I_25566 (I437675,I437523,I437579);
not I_25567 (I437692,I437675);
nand I_25568 (I437200,I437692,I437548);
not I_25569 (I437747,I3042);
DFFARX1 I_25570 (I551542,I3035,I437747,I437773,);
not I_25571 (I437781,I437773);
nand I_25572 (I437798,I551551,I551539);
and I_25573 (I437815,I437798,I551536);
DFFARX1 I_25574 (I437815,I3035,I437747,I437841,);
DFFARX1 I_25575 (I437841,I3035,I437747,I437736,);
DFFARX1 I_25576 (I551536,I3035,I437747,I437872,);
nand I_25577 (I437880,I437872,I551533);
not I_25578 (I437897,I437880);
DFFARX1 I_25579 (I437897,I3035,I437747,I437923,);
not I_25580 (I437931,I437923);
nor I_25581 (I437739,I437781,I437931);
DFFARX1 I_25582 (I551539,I3035,I437747,I437971,);
nor I_25583 (I437730,I437971,I437841);
nor I_25584 (I437721,I437971,I437897);
nand I_25585 (I438007,I551554,I551545);
and I_25586 (I438024,I438007,I551548);
DFFARX1 I_25587 (I438024,I3035,I437747,I438050,);
not I_25588 (I438058,I438050);
nand I_25589 (I438075,I438058,I437971);
nand I_25590 (I437724,I438058,I437880);
nor I_25591 (I438106,I551533,I551545);
and I_25592 (I438123,I437971,I438106);
nor I_25593 (I438140,I438058,I438123);
DFFARX1 I_25594 (I438140,I3035,I437747,I437733,);
nor I_25595 (I438171,I437773,I438106);
DFFARX1 I_25596 (I438171,I3035,I437747,I437718,);
nor I_25597 (I438202,I438050,I438106);
not I_25598 (I438219,I438202);
nand I_25599 (I437727,I438219,I438075);
not I_25600 (I438274,I3042);
DFFARX1 I_25601 (I324445,I3035,I438274,I438300,);
not I_25602 (I438308,I438300);
nand I_25603 (I438325,I324430,I324451);
and I_25604 (I438342,I438325,I324439);
DFFARX1 I_25605 (I438342,I3035,I438274,I438368,);
DFFARX1 I_25606 (I438368,I3035,I438274,I438263,);
DFFARX1 I_25607 (I324433,I3035,I438274,I438399,);
nand I_25608 (I438407,I438399,I324442);
not I_25609 (I438424,I438407);
DFFARX1 I_25610 (I438424,I3035,I438274,I438450,);
not I_25611 (I438458,I438450);
nor I_25612 (I438266,I438308,I438458);
DFFARX1 I_25613 (I324448,I3035,I438274,I438498,);
nor I_25614 (I438257,I438498,I438368);
nor I_25615 (I438248,I438498,I438424);
nand I_25616 (I438534,I324430,I324433);
and I_25617 (I438551,I438534,I324454);
DFFARX1 I_25618 (I438551,I3035,I438274,I438577,);
not I_25619 (I438585,I438577);
nand I_25620 (I438602,I438585,I438498);
nand I_25621 (I438251,I438585,I438407);
nor I_25622 (I438633,I324436,I324433);
and I_25623 (I438650,I438498,I438633);
nor I_25624 (I438667,I438585,I438650);
DFFARX1 I_25625 (I438667,I3035,I438274,I438260,);
nor I_25626 (I438698,I438300,I438633);
DFFARX1 I_25627 (I438698,I3035,I438274,I438245,);
nor I_25628 (I438729,I438577,I438633);
not I_25629 (I438746,I438729);
nand I_25630 (I438254,I438746,I438602);
not I_25631 (I438801,I3042);
DFFARX1 I_25632 (I282922,I3035,I438801,I438827,);
not I_25633 (I438835,I438827);
nand I_25634 (I438852,I282940,I282931);
and I_25635 (I438869,I438852,I282934);
DFFARX1 I_25636 (I438869,I3035,I438801,I438895,);
DFFARX1 I_25637 (I438895,I3035,I438801,I438790,);
DFFARX1 I_25638 (I282928,I3035,I438801,I438926,);
nand I_25639 (I438934,I438926,I282919);
not I_25640 (I438951,I438934);
DFFARX1 I_25641 (I438951,I3035,I438801,I438977,);
not I_25642 (I438985,I438977);
nor I_25643 (I438793,I438835,I438985);
DFFARX1 I_25644 (I282925,I3035,I438801,I439025,);
nor I_25645 (I438784,I439025,I438895);
nor I_25646 (I438775,I439025,I438951);
nand I_25647 (I439061,I282919,I282916);
and I_25648 (I439078,I439061,I282937);
DFFARX1 I_25649 (I439078,I3035,I438801,I439104,);
not I_25650 (I439112,I439104);
nand I_25651 (I439129,I439112,I439025);
nand I_25652 (I438778,I439112,I438934);
nor I_25653 (I439160,I282916,I282916);
and I_25654 (I439177,I439025,I439160);
nor I_25655 (I439194,I439112,I439177);
DFFARX1 I_25656 (I439194,I3035,I438801,I438787,);
nor I_25657 (I439225,I438827,I439160);
DFFARX1 I_25658 (I439225,I3035,I438801,I438772,);
nor I_25659 (I439256,I439104,I439160);
not I_25660 (I439273,I439256);
nand I_25661 (I438781,I439273,I439129);
not I_25662 (I439328,I3042);
DFFARX1 I_25663 (I81285,I3035,I439328,I439354,);
not I_25664 (I439362,I439354);
nand I_25665 (I439379,I81282,I81300);
and I_25666 (I439396,I439379,I81291);
DFFARX1 I_25667 (I439396,I3035,I439328,I439422,);
DFFARX1 I_25668 (I439422,I3035,I439328,I439317,);
DFFARX1 I_25669 (I81297,I3035,I439328,I439453,);
nand I_25670 (I439461,I439453,I81294);
not I_25671 (I439478,I439461);
DFFARX1 I_25672 (I439478,I3035,I439328,I439504,);
not I_25673 (I439512,I439504);
nor I_25674 (I439320,I439362,I439512);
DFFARX1 I_25675 (I81288,I3035,I439328,I439552,);
nor I_25676 (I439311,I439552,I439422);
nor I_25677 (I439302,I439552,I439478);
nand I_25678 (I439588,I81279,I81303);
and I_25679 (I439605,I439588,I81282);
DFFARX1 I_25680 (I439605,I3035,I439328,I439631,);
not I_25681 (I439639,I439631);
nand I_25682 (I439656,I439639,I439552);
nand I_25683 (I439305,I439639,I439461);
nor I_25684 (I439687,I81279,I81303);
and I_25685 (I439704,I439552,I439687);
nor I_25686 (I439721,I439639,I439704);
DFFARX1 I_25687 (I439721,I3035,I439328,I439314,);
nor I_25688 (I439752,I439354,I439687);
DFFARX1 I_25689 (I439752,I3035,I439328,I439299,);
nor I_25690 (I439783,I439631,I439687);
not I_25691 (I439800,I439783);
nand I_25692 (I439308,I439800,I439656);
not I_25693 (I439855,I3042);
DFFARX1 I_25694 (I321555,I3035,I439855,I439881,);
not I_25695 (I439889,I439881);
nand I_25696 (I439906,I321540,I321561);
and I_25697 (I439923,I439906,I321549);
DFFARX1 I_25698 (I439923,I3035,I439855,I439949,);
DFFARX1 I_25699 (I439949,I3035,I439855,I439844,);
DFFARX1 I_25700 (I321543,I3035,I439855,I439980,);
nand I_25701 (I439988,I439980,I321552);
not I_25702 (I440005,I439988);
DFFARX1 I_25703 (I440005,I3035,I439855,I440031,);
not I_25704 (I440039,I440031);
nor I_25705 (I439847,I439889,I440039);
DFFARX1 I_25706 (I321558,I3035,I439855,I440079,);
nor I_25707 (I439838,I440079,I439949);
nor I_25708 (I439829,I440079,I440005);
nand I_25709 (I440115,I321540,I321543);
and I_25710 (I440132,I440115,I321564);
DFFARX1 I_25711 (I440132,I3035,I439855,I440158,);
not I_25712 (I440166,I440158);
nand I_25713 (I440183,I440166,I440079);
nand I_25714 (I439832,I440166,I439988);
nor I_25715 (I440214,I321546,I321543);
and I_25716 (I440231,I440079,I440214);
nor I_25717 (I440248,I440166,I440231);
DFFARX1 I_25718 (I440248,I3035,I439855,I439841,);
nor I_25719 (I440279,I439881,I440214);
DFFARX1 I_25720 (I440279,I3035,I439855,I439826,);
nor I_25721 (I440310,I440158,I440214);
not I_25722 (I440327,I440310);
nand I_25723 (I439835,I440327,I440183);
not I_25724 (I440382,I3042);
DFFARX1 I_25725 (I583868,I3035,I440382,I440408,);
not I_25726 (I440416,I440408);
nand I_25727 (I440433,I583850,I583850);
and I_25728 (I440450,I440433,I583856);
DFFARX1 I_25729 (I440450,I3035,I440382,I440476,);
DFFARX1 I_25730 (I440476,I3035,I440382,I440371,);
DFFARX1 I_25731 (I583853,I3035,I440382,I440507,);
nand I_25732 (I440515,I440507,I583862);
not I_25733 (I440532,I440515);
DFFARX1 I_25734 (I440532,I3035,I440382,I440558,);
not I_25735 (I440566,I440558);
nor I_25736 (I440374,I440416,I440566);
DFFARX1 I_25737 (I583874,I3035,I440382,I440606,);
nor I_25738 (I440365,I440606,I440476);
nor I_25739 (I440356,I440606,I440532);
nand I_25740 (I440642,I583865,I583859);
and I_25741 (I440659,I440642,I583853);
DFFARX1 I_25742 (I440659,I3035,I440382,I440685,);
not I_25743 (I440693,I440685);
nand I_25744 (I440710,I440693,I440606);
nand I_25745 (I440359,I440693,I440515);
nor I_25746 (I440741,I583871,I583859);
and I_25747 (I440758,I440606,I440741);
nor I_25748 (I440775,I440693,I440758);
DFFARX1 I_25749 (I440775,I3035,I440382,I440368,);
nor I_25750 (I440806,I440408,I440741);
DFFARX1 I_25751 (I440806,I3035,I440382,I440353,);
nor I_25752 (I440837,I440685,I440741);
not I_25753 (I440854,I440837);
nand I_25754 (I440362,I440854,I440710);
not I_25755 (I440909,I3042);
DFFARX1 I_25756 (I80095,I3035,I440909,I440935,);
not I_25757 (I440943,I440935);
nand I_25758 (I440960,I80092,I80110);
and I_25759 (I440977,I440960,I80101);
DFFARX1 I_25760 (I440977,I3035,I440909,I441003,);
DFFARX1 I_25761 (I441003,I3035,I440909,I440898,);
DFFARX1 I_25762 (I80107,I3035,I440909,I441034,);
nand I_25763 (I441042,I441034,I80104);
not I_25764 (I441059,I441042);
DFFARX1 I_25765 (I441059,I3035,I440909,I441085,);
not I_25766 (I441093,I441085);
nor I_25767 (I440901,I440943,I441093);
DFFARX1 I_25768 (I80098,I3035,I440909,I441133,);
nor I_25769 (I440892,I441133,I441003);
nor I_25770 (I440883,I441133,I441059);
nand I_25771 (I441169,I80089,I80113);
and I_25772 (I441186,I441169,I80092);
DFFARX1 I_25773 (I441186,I3035,I440909,I441212,);
not I_25774 (I441220,I441212);
nand I_25775 (I441237,I441220,I441133);
nand I_25776 (I440886,I441220,I441042);
nor I_25777 (I441268,I80089,I80113);
and I_25778 (I441285,I441133,I441268);
nor I_25779 (I441302,I441220,I441285);
DFFARX1 I_25780 (I441302,I3035,I440909,I440895,);
nor I_25781 (I441333,I440935,I441268);
DFFARX1 I_25782 (I441333,I3035,I440909,I440880,);
nor I_25783 (I441364,I441212,I441268);
not I_25784 (I441381,I441364);
nand I_25785 (I440889,I441381,I441237);
not I_25786 (I441436,I3042);
DFFARX1 I_25787 (I653426,I3035,I441436,I441462,);
not I_25788 (I441470,I441462);
nand I_25789 (I441487,I653432,I653414);
and I_25790 (I441504,I441487,I653423);
DFFARX1 I_25791 (I441504,I3035,I441436,I441530,);
DFFARX1 I_25792 (I441530,I3035,I441436,I441425,);
DFFARX1 I_25793 (I653429,I3035,I441436,I441561,);
nand I_25794 (I441569,I441561,I653417);
not I_25795 (I441586,I441569);
DFFARX1 I_25796 (I441586,I3035,I441436,I441612,);
not I_25797 (I441620,I441612);
nor I_25798 (I441428,I441470,I441620);
DFFARX1 I_25799 (I653435,I3035,I441436,I441660,);
nor I_25800 (I441419,I441660,I441530);
nor I_25801 (I441410,I441660,I441586);
nand I_25802 (I441696,I653414,I653420);
and I_25803 (I441713,I441696,I653438);
DFFARX1 I_25804 (I441713,I3035,I441436,I441739,);
not I_25805 (I441747,I441739);
nand I_25806 (I441764,I441747,I441660);
nand I_25807 (I441413,I441747,I441569);
nor I_25808 (I441795,I653417,I653420);
and I_25809 (I441812,I441660,I441795);
nor I_25810 (I441829,I441747,I441812);
DFFARX1 I_25811 (I441829,I3035,I441436,I441422,);
nor I_25812 (I441860,I441462,I441795);
DFFARX1 I_25813 (I441860,I3035,I441436,I441407,);
nor I_25814 (I441891,I441739,I441795);
not I_25815 (I441908,I441891);
nand I_25816 (I441416,I441908,I441764);
not I_25817 (I441963,I3042);
DFFARX1 I_25818 (I741863,I3035,I441963,I441989,);
not I_25819 (I441997,I441989);
nand I_25820 (I442014,I741860,I741869);
and I_25821 (I442031,I442014,I741848);
DFFARX1 I_25822 (I442031,I3035,I441963,I442057,);
DFFARX1 I_25823 (I442057,I3035,I441963,I441952,);
DFFARX1 I_25824 (I741851,I3035,I441963,I442088,);
nand I_25825 (I442096,I442088,I741866);
not I_25826 (I442113,I442096);
DFFARX1 I_25827 (I442113,I3035,I441963,I442139,);
not I_25828 (I442147,I442139);
nor I_25829 (I441955,I441997,I442147);
DFFARX1 I_25830 (I741872,I3035,I441963,I442187,);
nor I_25831 (I441946,I442187,I442057);
nor I_25832 (I441937,I442187,I442113);
nand I_25833 (I442223,I741854,I741875);
and I_25834 (I442240,I442223,I741857);
DFFARX1 I_25835 (I442240,I3035,I441963,I442266,);
not I_25836 (I442274,I442266);
nand I_25837 (I442291,I442274,I442187);
nand I_25838 (I441940,I442274,I442096);
nor I_25839 (I442322,I741848,I741875);
and I_25840 (I442339,I442187,I442322);
nor I_25841 (I442356,I442274,I442339);
DFFARX1 I_25842 (I442356,I3035,I441963,I441949,);
nor I_25843 (I442387,I441989,I442322);
DFFARX1 I_25844 (I442387,I3035,I441963,I441934,);
nor I_25845 (I442418,I442266,I442322);
not I_25846 (I442435,I442418);
nand I_25847 (I441943,I442435,I442291);
not I_25848 (I442490,I3042);
DFFARX1 I_25849 (I649618,I3035,I442490,I442516,);
not I_25850 (I442524,I442516);
nand I_25851 (I442541,I649624,I649606);
and I_25852 (I442558,I442541,I649615);
DFFARX1 I_25853 (I442558,I3035,I442490,I442584,);
DFFARX1 I_25854 (I442584,I3035,I442490,I442479,);
DFFARX1 I_25855 (I649621,I3035,I442490,I442615,);
nand I_25856 (I442623,I442615,I649609);
not I_25857 (I442640,I442623);
DFFARX1 I_25858 (I442640,I3035,I442490,I442666,);
not I_25859 (I442674,I442666);
nor I_25860 (I442482,I442524,I442674);
DFFARX1 I_25861 (I649627,I3035,I442490,I442714,);
nor I_25862 (I442473,I442714,I442584);
nor I_25863 (I442464,I442714,I442640);
nand I_25864 (I442750,I649606,I649612);
and I_25865 (I442767,I442750,I649630);
DFFARX1 I_25866 (I442767,I3035,I442490,I442793,);
not I_25867 (I442801,I442793);
nand I_25868 (I442818,I442801,I442714);
nand I_25869 (I442467,I442801,I442623);
nor I_25870 (I442849,I649609,I649612);
and I_25871 (I442866,I442714,I442849);
nor I_25872 (I442883,I442801,I442866);
DFFARX1 I_25873 (I442883,I3035,I442490,I442476,);
nor I_25874 (I442914,I442516,I442849);
DFFARX1 I_25875 (I442914,I3035,I442490,I442461,);
nor I_25876 (I442945,I442793,I442849);
not I_25877 (I442962,I442945);
nand I_25878 (I442470,I442962,I442818);
not I_25879 (I443017,I3042);
DFFARX1 I_25880 (I375872,I3035,I443017,I443043,);
not I_25881 (I443051,I443043);
nand I_25882 (I443068,I375875,I375872);
and I_25883 (I443085,I443068,I375884);
DFFARX1 I_25884 (I443085,I3035,I443017,I443111,);
DFFARX1 I_25885 (I443111,I3035,I443017,I443006,);
DFFARX1 I_25886 (I375881,I3035,I443017,I443142,);
nand I_25887 (I443150,I443142,I375887);
not I_25888 (I443167,I443150);
DFFARX1 I_25889 (I443167,I3035,I443017,I443193,);
not I_25890 (I443201,I443193);
nor I_25891 (I443009,I443051,I443201);
DFFARX1 I_25892 (I375896,I3035,I443017,I443241,);
nor I_25893 (I443000,I443241,I443111);
nor I_25894 (I442991,I443241,I443167);
nand I_25895 (I443277,I375890,I375878);
and I_25896 (I443294,I443277,I375875);
DFFARX1 I_25897 (I443294,I3035,I443017,I443320,);
not I_25898 (I443328,I443320);
nand I_25899 (I443345,I443328,I443241);
nand I_25900 (I442994,I443328,I443150);
nor I_25901 (I443376,I375893,I375878);
and I_25902 (I443393,I443241,I443376);
nor I_25903 (I443410,I443328,I443393);
DFFARX1 I_25904 (I443410,I3035,I443017,I443003,);
nor I_25905 (I443441,I443043,I443376);
DFFARX1 I_25906 (I443441,I3035,I443017,I442988,);
nor I_25907 (I443472,I443320,I443376);
not I_25908 (I443489,I443472);
nand I_25909 (I442997,I443489,I443345);
not I_25910 (I443544,I3042);
DFFARX1 I_25911 (I646870,I3035,I443544,I443570,);
not I_25912 (I443578,I443570);
nand I_25913 (I443595,I646852,I646852);
and I_25914 (I443612,I443595,I646858);
DFFARX1 I_25915 (I443612,I3035,I443544,I443638,);
DFFARX1 I_25916 (I443638,I3035,I443544,I443533,);
DFFARX1 I_25917 (I646855,I3035,I443544,I443669,);
nand I_25918 (I443677,I443669,I646864);
not I_25919 (I443694,I443677);
DFFARX1 I_25920 (I443694,I3035,I443544,I443720,);
not I_25921 (I443728,I443720);
nor I_25922 (I443536,I443578,I443728);
DFFARX1 I_25923 (I646876,I3035,I443544,I443768,);
nor I_25924 (I443527,I443768,I443638);
nor I_25925 (I443518,I443768,I443694);
nand I_25926 (I443804,I646867,I646861);
and I_25927 (I443821,I443804,I646855);
DFFARX1 I_25928 (I443821,I3035,I443544,I443847,);
not I_25929 (I443855,I443847);
nand I_25930 (I443872,I443855,I443768);
nand I_25931 (I443521,I443855,I443677);
nor I_25932 (I443903,I646873,I646861);
and I_25933 (I443920,I443768,I443903);
nor I_25934 (I443937,I443855,I443920);
DFFARX1 I_25935 (I443937,I3035,I443544,I443530,);
nor I_25936 (I443968,I443570,I443903);
DFFARX1 I_25937 (I443968,I3035,I443544,I443515,);
nor I_25938 (I443999,I443847,I443903);
not I_25939 (I444016,I443999);
nand I_25940 (I443524,I444016,I443872);
not I_25941 (I444071,I3042);
DFFARX1 I_25942 (I265259,I3035,I444071,I444097,);
not I_25943 (I444105,I444097);
nand I_25944 (I444122,I265256,I265265);
and I_25945 (I444139,I444122,I265274);
DFFARX1 I_25946 (I444139,I3035,I444071,I444165,);
DFFARX1 I_25947 (I444165,I3035,I444071,I444060,);
DFFARX1 I_25948 (I265277,I3035,I444071,I444196,);
nand I_25949 (I444204,I444196,I265280);
not I_25950 (I444221,I444204);
DFFARX1 I_25951 (I444221,I3035,I444071,I444247,);
not I_25952 (I444255,I444247);
nor I_25953 (I444063,I444105,I444255);
DFFARX1 I_25954 (I265253,I3035,I444071,I444295,);
nor I_25955 (I444054,I444295,I444165);
nor I_25956 (I444045,I444295,I444221);
nand I_25957 (I444331,I265268,I265271);
and I_25958 (I444348,I444331,I265262);
DFFARX1 I_25959 (I444348,I3035,I444071,I444374,);
not I_25960 (I444382,I444374);
nand I_25961 (I444399,I444382,I444295);
nand I_25962 (I444048,I444382,I444204);
nor I_25963 (I444430,I265253,I265271);
and I_25964 (I444447,I444295,I444430);
nor I_25965 (I444464,I444382,I444447);
DFFARX1 I_25966 (I444464,I3035,I444071,I444057,);
nor I_25967 (I444495,I444097,I444430);
DFFARX1 I_25968 (I444495,I3035,I444071,I444042,);
nor I_25969 (I444526,I444374,I444430);
not I_25970 (I444543,I444526);
nand I_25971 (I444051,I444543,I444399);
not I_25972 (I444598,I3042);
DFFARX1 I_25973 (I596584,I3035,I444598,I444624,);
not I_25974 (I444632,I444624);
nand I_25975 (I444649,I596566,I596566);
and I_25976 (I444666,I444649,I596572);
DFFARX1 I_25977 (I444666,I3035,I444598,I444692,);
DFFARX1 I_25978 (I444692,I3035,I444598,I444587,);
DFFARX1 I_25979 (I596569,I3035,I444598,I444723,);
nand I_25980 (I444731,I444723,I596578);
not I_25981 (I444748,I444731);
DFFARX1 I_25982 (I444748,I3035,I444598,I444774,);
not I_25983 (I444782,I444774);
nor I_25984 (I444590,I444632,I444782);
DFFARX1 I_25985 (I596590,I3035,I444598,I444822,);
nor I_25986 (I444581,I444822,I444692);
nor I_25987 (I444572,I444822,I444748);
nand I_25988 (I444858,I596581,I596575);
and I_25989 (I444875,I444858,I596569);
DFFARX1 I_25990 (I444875,I3035,I444598,I444901,);
not I_25991 (I444909,I444901);
nand I_25992 (I444926,I444909,I444822);
nand I_25993 (I444575,I444909,I444731);
nor I_25994 (I444957,I596587,I596575);
and I_25995 (I444974,I444822,I444957);
nor I_25996 (I444991,I444909,I444974);
DFFARX1 I_25997 (I444991,I3035,I444598,I444584,);
nor I_25998 (I445022,I444624,I444957);
DFFARX1 I_25999 (I445022,I3035,I444598,I444569,);
nor I_26000 (I445053,I444901,I444957);
not I_26001 (I445070,I445053);
nand I_26002 (I444578,I445070,I444926);
not I_26003 (I445125,I3042);
DFFARX1 I_26004 (I514833,I3035,I445125,I445151,);
not I_26005 (I445159,I445151);
nand I_26006 (I445176,I514848,I514830);
and I_26007 (I445193,I445176,I514830);
DFFARX1 I_26008 (I445193,I3035,I445125,I445219,);
DFFARX1 I_26009 (I445219,I3035,I445125,I445114,);
DFFARX1 I_26010 (I514839,I3035,I445125,I445250,);
nand I_26011 (I445258,I445250,I514857);
not I_26012 (I445275,I445258);
DFFARX1 I_26013 (I445275,I3035,I445125,I445301,);
not I_26014 (I445309,I445301);
nor I_26015 (I445117,I445159,I445309);
DFFARX1 I_26016 (I514854,I3035,I445125,I445349,);
nor I_26017 (I445108,I445349,I445219);
nor I_26018 (I445099,I445349,I445275);
nand I_26019 (I445385,I514851,I514842);
and I_26020 (I445402,I445385,I514836);
DFFARX1 I_26021 (I445402,I3035,I445125,I445428,);
not I_26022 (I445436,I445428);
nand I_26023 (I445453,I445436,I445349);
nand I_26024 (I445102,I445436,I445258);
nor I_26025 (I445484,I514845,I514842);
and I_26026 (I445501,I445349,I445484);
nor I_26027 (I445518,I445436,I445501);
DFFARX1 I_26028 (I445518,I3035,I445125,I445111,);
nor I_26029 (I445549,I445151,I445484);
DFFARX1 I_26030 (I445549,I3035,I445125,I445096,);
nor I_26031 (I445580,I445428,I445484);
not I_26032 (I445597,I445580);
nand I_26033 (I445105,I445597,I445453);
not I_26034 (I445652,I3042);
DFFARX1 I_26035 (I615658,I3035,I445652,I445678,);
not I_26036 (I445686,I445678);
nand I_26037 (I445703,I615640,I615640);
and I_26038 (I445720,I445703,I615646);
DFFARX1 I_26039 (I445720,I3035,I445652,I445746,);
DFFARX1 I_26040 (I445746,I3035,I445652,I445641,);
DFFARX1 I_26041 (I615643,I3035,I445652,I445777,);
nand I_26042 (I445785,I445777,I615652);
not I_26043 (I445802,I445785);
DFFARX1 I_26044 (I445802,I3035,I445652,I445828,);
not I_26045 (I445836,I445828);
nor I_26046 (I445644,I445686,I445836);
DFFARX1 I_26047 (I615664,I3035,I445652,I445876,);
nor I_26048 (I445635,I445876,I445746);
nor I_26049 (I445626,I445876,I445802);
nand I_26050 (I445912,I615655,I615649);
and I_26051 (I445929,I445912,I615643);
DFFARX1 I_26052 (I445929,I3035,I445652,I445955,);
not I_26053 (I445963,I445955);
nand I_26054 (I445980,I445963,I445876);
nand I_26055 (I445629,I445963,I445785);
nor I_26056 (I446011,I615661,I615649);
and I_26057 (I446028,I445876,I446011);
nor I_26058 (I446045,I445963,I446028);
DFFARX1 I_26059 (I446045,I3035,I445652,I445638,);
nor I_26060 (I446076,I445678,I446011);
DFFARX1 I_26061 (I446076,I3035,I445652,I445623,);
nor I_26062 (I446107,I445955,I446011);
not I_26063 (I446124,I446107);
nand I_26064 (I445632,I446124,I445980);
not I_26065 (I446179,I3042);
DFFARX1 I_26066 (I277771,I3035,I446179,I446205,);
not I_26067 (I446213,I446205);
nand I_26068 (I446230,I277768,I277777);
and I_26069 (I446247,I446230,I277786);
DFFARX1 I_26070 (I446247,I3035,I446179,I446273,);
DFFARX1 I_26071 (I446273,I3035,I446179,I446168,);
DFFARX1 I_26072 (I277789,I3035,I446179,I446304,);
nand I_26073 (I446312,I446304,I277792);
not I_26074 (I446329,I446312);
DFFARX1 I_26075 (I446329,I3035,I446179,I446355,);
not I_26076 (I446363,I446355);
nor I_26077 (I446171,I446213,I446363);
DFFARX1 I_26078 (I277765,I3035,I446179,I446403,);
nor I_26079 (I446162,I446403,I446273);
nor I_26080 (I446153,I446403,I446329);
nand I_26081 (I446439,I277780,I277783);
and I_26082 (I446456,I446439,I277774);
DFFARX1 I_26083 (I446456,I3035,I446179,I446482,);
not I_26084 (I446490,I446482);
nand I_26085 (I446507,I446490,I446403);
nand I_26086 (I446156,I446490,I446312);
nor I_26087 (I446538,I277765,I277783);
and I_26088 (I446555,I446403,I446538);
nor I_26089 (I446572,I446490,I446555);
DFFARX1 I_26090 (I446572,I3035,I446179,I446165,);
nor I_26091 (I446603,I446205,I446538);
DFFARX1 I_26092 (I446603,I3035,I446179,I446150,);
nor I_26093 (I446634,I446482,I446538);
not I_26094 (I446651,I446634);
nand I_26095 (I446159,I446651,I446507);
not I_26096 (I446706,I3042);
DFFARX1 I_26097 (I388010,I3035,I446706,I446732,);
not I_26098 (I446740,I446732);
nand I_26099 (I446757,I388013,I388010);
and I_26100 (I446774,I446757,I388022);
DFFARX1 I_26101 (I446774,I3035,I446706,I446800,);
DFFARX1 I_26102 (I446800,I3035,I446706,I446695,);
DFFARX1 I_26103 (I388019,I3035,I446706,I446831,);
nand I_26104 (I446839,I446831,I388025);
not I_26105 (I446856,I446839);
DFFARX1 I_26106 (I446856,I3035,I446706,I446882,);
not I_26107 (I446890,I446882);
nor I_26108 (I446698,I446740,I446890);
DFFARX1 I_26109 (I388034,I3035,I446706,I446930,);
nor I_26110 (I446689,I446930,I446800);
nor I_26111 (I446680,I446930,I446856);
nand I_26112 (I446966,I388028,I388016);
and I_26113 (I446983,I446966,I388013);
DFFARX1 I_26114 (I446983,I3035,I446706,I447009,);
not I_26115 (I447017,I447009);
nand I_26116 (I447034,I447017,I446930);
nand I_26117 (I446683,I447017,I446839);
nor I_26118 (I447065,I388031,I388016);
and I_26119 (I447082,I446930,I447065);
nor I_26120 (I447099,I447017,I447082);
DFFARX1 I_26121 (I447099,I3035,I446706,I446692,);
nor I_26122 (I447130,I446732,I447065);
DFFARX1 I_26123 (I447130,I3035,I446706,I446677,);
nor I_26124 (I447161,I447009,I447065);
not I_26125 (I447178,I447161);
nand I_26126 (I446686,I447178,I447034);
not I_26127 (I447233,I3042);
DFFARX1 I_26128 (I84855,I3035,I447233,I447259,);
not I_26129 (I447267,I447259);
nand I_26130 (I447284,I84852,I84870);
and I_26131 (I447301,I447284,I84861);
DFFARX1 I_26132 (I447301,I3035,I447233,I447327,);
DFFARX1 I_26133 (I447327,I3035,I447233,I447222,);
DFFARX1 I_26134 (I84867,I3035,I447233,I447358,);
nand I_26135 (I447366,I447358,I84864);
not I_26136 (I447383,I447366);
DFFARX1 I_26137 (I447383,I3035,I447233,I447409,);
not I_26138 (I447417,I447409);
nor I_26139 (I447225,I447267,I447417);
DFFARX1 I_26140 (I84858,I3035,I447233,I447457,);
nor I_26141 (I447216,I447457,I447327);
nor I_26142 (I447207,I447457,I447383);
nand I_26143 (I447493,I84849,I84873);
and I_26144 (I447510,I447493,I84852);
DFFARX1 I_26145 (I447510,I3035,I447233,I447536,);
not I_26146 (I447544,I447536);
nand I_26147 (I447561,I447544,I447457);
nand I_26148 (I447210,I447544,I447366);
nor I_26149 (I447592,I84849,I84873);
and I_26150 (I447609,I447457,I447592);
nor I_26151 (I447626,I447544,I447609);
DFFARX1 I_26152 (I447626,I3035,I447233,I447219,);
nor I_26153 (I447657,I447259,I447592);
DFFARX1 I_26154 (I447657,I3035,I447233,I447204,);
nor I_26155 (I447688,I447536,I447592);
not I_26156 (I447705,I447688);
nand I_26157 (I447213,I447705,I447561);
not I_26158 (I447760,I3042);
DFFARX1 I_26159 (I504497,I3035,I447760,I447786,);
not I_26160 (I447794,I447786);
nand I_26161 (I447811,I504512,I504494);
and I_26162 (I447828,I447811,I504494);
DFFARX1 I_26163 (I447828,I3035,I447760,I447854,);
DFFARX1 I_26164 (I447854,I3035,I447760,I447749,);
DFFARX1 I_26165 (I504503,I3035,I447760,I447885,);
nand I_26166 (I447893,I447885,I504521);
not I_26167 (I447910,I447893);
DFFARX1 I_26168 (I447910,I3035,I447760,I447936,);
not I_26169 (I447944,I447936);
nor I_26170 (I447752,I447794,I447944);
DFFARX1 I_26171 (I504518,I3035,I447760,I447984,);
nor I_26172 (I447743,I447984,I447854);
nor I_26173 (I447734,I447984,I447910);
nand I_26174 (I448020,I504515,I504506);
and I_26175 (I448037,I448020,I504500);
DFFARX1 I_26176 (I448037,I3035,I447760,I448063,);
not I_26177 (I448071,I448063);
nand I_26178 (I448088,I448071,I447984);
nand I_26179 (I447737,I448071,I447893);
nor I_26180 (I448119,I504509,I504506);
and I_26181 (I448136,I447984,I448119);
nor I_26182 (I448153,I448071,I448136);
DFFARX1 I_26183 (I448153,I3035,I447760,I447746,);
nor I_26184 (I448184,I447786,I448119);
DFFARX1 I_26185 (I448184,I3035,I447760,I447731,);
nor I_26186 (I448215,I448063,I448119);
not I_26187 (I448232,I448215);
nand I_26188 (I447740,I448232,I448088);
not I_26189 (I448287,I3042);
DFFARX1 I_26190 (I686956,I3035,I448287,I448313,);
not I_26191 (I448321,I448313);
nand I_26192 (I448338,I686938,I686941);
and I_26193 (I448355,I448338,I686953);
DFFARX1 I_26194 (I448355,I3035,I448287,I448381,);
DFFARX1 I_26195 (I448381,I3035,I448287,I448276,);
DFFARX1 I_26196 (I686962,I3035,I448287,I448412,);
nand I_26197 (I448420,I448412,I686947);
not I_26198 (I448437,I448420);
DFFARX1 I_26199 (I448437,I3035,I448287,I448463,);
not I_26200 (I448471,I448463);
nor I_26201 (I448279,I448321,I448471);
DFFARX1 I_26202 (I686959,I3035,I448287,I448511,);
nor I_26203 (I448270,I448511,I448381);
nor I_26204 (I448261,I448511,I448437);
nand I_26205 (I448547,I686950,I686944);
and I_26206 (I448564,I448547,I686938);
DFFARX1 I_26207 (I448564,I3035,I448287,I448590,);
not I_26208 (I448598,I448590);
nand I_26209 (I448615,I448598,I448511);
nand I_26210 (I448264,I448598,I448420);
nor I_26211 (I448646,I686941,I686944);
and I_26212 (I448663,I448511,I448646);
nor I_26213 (I448680,I448598,I448663);
DFFARX1 I_26214 (I448680,I3035,I448287,I448273,);
nor I_26215 (I448711,I448313,I448646);
DFFARX1 I_26216 (I448711,I3035,I448287,I448258,);
nor I_26217 (I448742,I448590,I448646);
not I_26218 (I448759,I448742);
nand I_26219 (I448267,I448759,I448615);
not I_26220 (I448814,I3042);
DFFARX1 I_26221 (I284707,I3035,I448814,I448840,);
not I_26222 (I448848,I448840);
nand I_26223 (I448865,I284725,I284716);
and I_26224 (I448882,I448865,I284719);
DFFARX1 I_26225 (I448882,I3035,I448814,I448908,);
DFFARX1 I_26226 (I448908,I3035,I448814,I448803,);
DFFARX1 I_26227 (I284713,I3035,I448814,I448939,);
nand I_26228 (I448947,I448939,I284704);
not I_26229 (I448964,I448947);
DFFARX1 I_26230 (I448964,I3035,I448814,I448990,);
not I_26231 (I448998,I448990);
nor I_26232 (I448806,I448848,I448998);
DFFARX1 I_26233 (I284710,I3035,I448814,I449038,);
nor I_26234 (I448797,I449038,I448908);
nor I_26235 (I448788,I449038,I448964);
nand I_26236 (I449074,I284704,I284701);
and I_26237 (I449091,I449074,I284722);
DFFARX1 I_26238 (I449091,I3035,I448814,I449117,);
not I_26239 (I449125,I449117);
nand I_26240 (I449142,I449125,I449038);
nand I_26241 (I448791,I449125,I448947);
nor I_26242 (I449173,I284701,I284701);
and I_26243 (I449190,I449038,I449173);
nor I_26244 (I449207,I449125,I449190);
DFFARX1 I_26245 (I449207,I3035,I448814,I448800,);
nor I_26246 (I449238,I448840,I449173);
DFFARX1 I_26247 (I449238,I3035,I448814,I448785,);
nor I_26248 (I449269,I449117,I449173);
not I_26249 (I449286,I449269);
nand I_26250 (I448794,I449286,I449142);
not I_26251 (I449341,I3042);
DFFARX1 I_26252 (I619126,I3035,I449341,I449367,);
not I_26253 (I449375,I449367);
nand I_26254 (I449392,I619108,I619108);
and I_26255 (I449409,I449392,I619114);
DFFARX1 I_26256 (I449409,I3035,I449341,I449435,);
DFFARX1 I_26257 (I449435,I3035,I449341,I449330,);
DFFARX1 I_26258 (I619111,I3035,I449341,I449466,);
nand I_26259 (I449474,I449466,I619120);
not I_26260 (I449491,I449474);
DFFARX1 I_26261 (I449491,I3035,I449341,I449517,);
not I_26262 (I449525,I449517);
nor I_26263 (I449333,I449375,I449525);
DFFARX1 I_26264 (I619132,I3035,I449341,I449565,);
nor I_26265 (I449324,I449565,I449435);
nor I_26266 (I449315,I449565,I449491);
nand I_26267 (I449601,I619123,I619117);
and I_26268 (I449618,I449601,I619111);
DFFARX1 I_26269 (I449618,I3035,I449341,I449644,);
not I_26270 (I449652,I449644);
nand I_26271 (I449669,I449652,I449565);
nand I_26272 (I449318,I449652,I449474);
nor I_26273 (I449700,I619129,I619117);
and I_26274 (I449717,I449565,I449700);
nor I_26275 (I449734,I449652,I449717);
DFFARX1 I_26276 (I449734,I3035,I449341,I449327,);
nor I_26277 (I449765,I449367,I449700);
DFFARX1 I_26278 (I449765,I3035,I449341,I449312,);
nor I_26279 (I449796,I449644,I449700);
not I_26280 (I449813,I449796);
nand I_26281 (I449321,I449813,I449669);
not I_26282 (I449868,I3042);
DFFARX1 I_26283 (I298392,I3035,I449868,I449894,);
not I_26284 (I449902,I449894);
nand I_26285 (I449919,I298410,I298401);
and I_26286 (I449936,I449919,I298404);
DFFARX1 I_26287 (I449936,I3035,I449868,I449962,);
DFFARX1 I_26288 (I449962,I3035,I449868,I449857,);
DFFARX1 I_26289 (I298398,I3035,I449868,I449993,);
nand I_26290 (I450001,I449993,I298389);
not I_26291 (I450018,I450001);
DFFARX1 I_26292 (I450018,I3035,I449868,I450044,);
not I_26293 (I450052,I450044);
nor I_26294 (I449860,I449902,I450052);
DFFARX1 I_26295 (I298395,I3035,I449868,I450092,);
nor I_26296 (I449851,I450092,I449962);
nor I_26297 (I449842,I450092,I450018);
nand I_26298 (I450128,I298389,I298386);
and I_26299 (I450145,I450128,I298407);
DFFARX1 I_26300 (I450145,I3035,I449868,I450171,);
not I_26301 (I450179,I450171);
nand I_26302 (I450196,I450179,I450092);
nand I_26303 (I449845,I450179,I450001);
nor I_26304 (I450227,I298386,I298386);
and I_26305 (I450244,I450092,I450227);
nor I_26306 (I450261,I450179,I450244);
DFFARX1 I_26307 (I450261,I3035,I449868,I449854,);
nor I_26308 (I450292,I449894,I450227);
DFFARX1 I_26309 (I450292,I3035,I449868,I449839,);
nor I_26310 (I450323,I450171,I450227);
not I_26311 (I450340,I450323);
nand I_26312 (I449848,I450340,I450196);
not I_26313 (I450395,I3042);
DFFARX1 I_26314 (I631264,I3035,I450395,I450421,);
not I_26315 (I450429,I450421);
nand I_26316 (I450446,I631246,I631246);
and I_26317 (I450463,I450446,I631252);
DFFARX1 I_26318 (I450463,I3035,I450395,I450489,);
DFFARX1 I_26319 (I450489,I3035,I450395,I450384,);
DFFARX1 I_26320 (I631249,I3035,I450395,I450520,);
nand I_26321 (I450528,I450520,I631258);
not I_26322 (I450545,I450528);
DFFARX1 I_26323 (I450545,I3035,I450395,I450571,);
not I_26324 (I450579,I450571);
nor I_26325 (I450387,I450429,I450579);
DFFARX1 I_26326 (I631270,I3035,I450395,I450619,);
nor I_26327 (I450378,I450619,I450489);
nor I_26328 (I450369,I450619,I450545);
nand I_26329 (I450655,I631261,I631255);
and I_26330 (I450672,I450655,I631249);
DFFARX1 I_26331 (I450672,I3035,I450395,I450698,);
not I_26332 (I450706,I450698);
nand I_26333 (I450723,I450706,I450619);
nand I_26334 (I450372,I450706,I450528);
nor I_26335 (I450754,I631267,I631255);
and I_26336 (I450771,I450619,I450754);
nor I_26337 (I450788,I450706,I450771);
DFFARX1 I_26338 (I450788,I3035,I450395,I450381,);
nor I_26339 (I450819,I450421,I450754);
DFFARX1 I_26340 (I450819,I3035,I450395,I450366,);
nor I_26341 (I450850,I450698,I450754);
not I_26342 (I450867,I450850);
nand I_26343 (I450375,I450867,I450723);
not I_26344 (I450922,I3042);
DFFARX1 I_26345 (I407662,I3035,I450922,I450948,);
not I_26346 (I450956,I450948);
nand I_26347 (I450973,I407665,I407662);
and I_26348 (I450990,I450973,I407674);
DFFARX1 I_26349 (I450990,I3035,I450922,I451016,);
DFFARX1 I_26350 (I451016,I3035,I450922,I450911,);
DFFARX1 I_26351 (I407671,I3035,I450922,I451047,);
nand I_26352 (I451055,I451047,I407677);
not I_26353 (I451072,I451055);
DFFARX1 I_26354 (I451072,I3035,I450922,I451098,);
not I_26355 (I451106,I451098);
nor I_26356 (I450914,I450956,I451106);
DFFARX1 I_26357 (I407686,I3035,I450922,I451146,);
nor I_26358 (I450905,I451146,I451016);
nor I_26359 (I450896,I451146,I451072);
nand I_26360 (I451182,I407680,I407668);
and I_26361 (I451199,I451182,I407665);
DFFARX1 I_26362 (I451199,I3035,I450922,I451225,);
not I_26363 (I451233,I451225);
nand I_26364 (I451250,I451233,I451146);
nand I_26365 (I450899,I451233,I451055);
nor I_26366 (I451281,I407683,I407668);
and I_26367 (I451298,I451146,I451281);
nor I_26368 (I451315,I451233,I451298);
DFFARX1 I_26369 (I451315,I3035,I450922,I450908,);
nor I_26370 (I451346,I450948,I451281);
DFFARX1 I_26371 (I451346,I3035,I450922,I450893,);
nor I_26372 (I451377,I451225,I451281);
not I_26373 (I451394,I451377);
nand I_26374 (I450902,I451394,I451250);
not I_26375 (I451449,I3042);
DFFARX1 I_26376 (I487701,I3035,I451449,I451475,);
not I_26377 (I451483,I451475);
nand I_26378 (I451500,I487716,I487698);
and I_26379 (I451517,I451500,I487698);
DFFARX1 I_26380 (I451517,I3035,I451449,I451543,);
DFFARX1 I_26381 (I451543,I3035,I451449,I451438,);
DFFARX1 I_26382 (I487707,I3035,I451449,I451574,);
nand I_26383 (I451582,I451574,I487725);
not I_26384 (I451599,I451582);
DFFARX1 I_26385 (I451599,I3035,I451449,I451625,);
not I_26386 (I451633,I451625);
nor I_26387 (I451441,I451483,I451633);
DFFARX1 I_26388 (I487722,I3035,I451449,I451673,);
nor I_26389 (I451432,I451673,I451543);
nor I_26390 (I451423,I451673,I451599);
nand I_26391 (I451709,I487719,I487710);
and I_26392 (I451726,I451709,I487704);
DFFARX1 I_26393 (I451726,I3035,I451449,I451752,);
not I_26394 (I451760,I451752);
nand I_26395 (I451777,I451760,I451673);
nand I_26396 (I451426,I451760,I451582);
nor I_26397 (I451808,I487713,I487710);
and I_26398 (I451825,I451673,I451808);
nor I_26399 (I451842,I451760,I451825);
DFFARX1 I_26400 (I451842,I3035,I451449,I451435,);
nor I_26401 (I451873,I451475,I451808);
DFFARX1 I_26402 (I451873,I3035,I451449,I451420,);
nor I_26403 (I451904,I451752,I451808);
not I_26404 (I451921,I451904);
nand I_26405 (I451429,I451921,I451777);
not I_26406 (I451976,I3042);
DFFARX1 I_26407 (I488993,I3035,I451976,I452002,);
not I_26408 (I452010,I452002);
nand I_26409 (I452027,I489008,I488990);
and I_26410 (I452044,I452027,I488990);
DFFARX1 I_26411 (I452044,I3035,I451976,I452070,);
DFFARX1 I_26412 (I452070,I3035,I451976,I451965,);
DFFARX1 I_26413 (I488999,I3035,I451976,I452101,);
nand I_26414 (I452109,I452101,I489017);
not I_26415 (I452126,I452109);
DFFARX1 I_26416 (I452126,I3035,I451976,I452152,);
not I_26417 (I452160,I452152);
nor I_26418 (I451968,I452010,I452160);
DFFARX1 I_26419 (I489014,I3035,I451976,I452200,);
nor I_26420 (I451959,I452200,I452070);
nor I_26421 (I451950,I452200,I452126);
nand I_26422 (I452236,I489011,I489002);
and I_26423 (I452253,I452236,I488996);
DFFARX1 I_26424 (I452253,I3035,I451976,I452279,);
not I_26425 (I452287,I452279);
nand I_26426 (I452304,I452287,I452200);
nand I_26427 (I451953,I452287,I452109);
nor I_26428 (I452335,I489005,I489002);
and I_26429 (I452352,I452200,I452335);
nor I_26430 (I452369,I452287,I452352);
DFFARX1 I_26431 (I452369,I3035,I451976,I451962,);
nor I_26432 (I452400,I452002,I452335);
DFFARX1 I_26433 (I452400,I3035,I451976,I451947,);
nor I_26434 (I452431,I452279,I452335);
not I_26435 (I452448,I452431);
nand I_26436 (I451956,I452448,I452304);
not I_26437 (I452503,I3042);
DFFARX1 I_26438 (I611612,I3035,I452503,I452529,);
not I_26439 (I452537,I452529);
nand I_26440 (I452554,I611594,I611594);
and I_26441 (I452571,I452554,I611600);
DFFARX1 I_26442 (I452571,I3035,I452503,I452597,);
DFFARX1 I_26443 (I452597,I3035,I452503,I452492,);
DFFARX1 I_26444 (I611597,I3035,I452503,I452628,);
nand I_26445 (I452636,I452628,I611606);
not I_26446 (I452653,I452636);
DFFARX1 I_26447 (I452653,I3035,I452503,I452679,);
not I_26448 (I452687,I452679);
nor I_26449 (I452495,I452537,I452687);
DFFARX1 I_26450 (I611618,I3035,I452503,I452727,);
nor I_26451 (I452486,I452727,I452597);
nor I_26452 (I452477,I452727,I452653);
nand I_26453 (I452763,I611609,I611603);
and I_26454 (I452780,I452763,I611597);
DFFARX1 I_26455 (I452780,I3035,I452503,I452806,);
not I_26456 (I452814,I452806);
nand I_26457 (I452831,I452814,I452727);
nand I_26458 (I452480,I452814,I452636);
nor I_26459 (I452862,I611615,I611603);
and I_26460 (I452879,I452727,I452862);
nor I_26461 (I452896,I452814,I452879);
DFFARX1 I_26462 (I452896,I3035,I452503,I452489,);
nor I_26463 (I452927,I452529,I452862);
DFFARX1 I_26464 (I452927,I3035,I452503,I452474,);
nor I_26465 (I452958,I452806,I452862);
not I_26466 (I452975,I452958);
nand I_26467 (I452483,I452975,I452831);
not I_26468 (I453030,I3042);
DFFARX1 I_26469 (I360844,I3035,I453030,I453056,);
not I_26470 (I453064,I453056);
nand I_26471 (I453081,I360847,I360844);
and I_26472 (I453098,I453081,I360856);
DFFARX1 I_26473 (I453098,I3035,I453030,I453124,);
DFFARX1 I_26474 (I453124,I3035,I453030,I453019,);
DFFARX1 I_26475 (I360853,I3035,I453030,I453155,);
nand I_26476 (I453163,I453155,I360859);
not I_26477 (I453180,I453163);
DFFARX1 I_26478 (I453180,I3035,I453030,I453206,);
not I_26479 (I453214,I453206);
nor I_26480 (I453022,I453064,I453214);
DFFARX1 I_26481 (I360868,I3035,I453030,I453254,);
nor I_26482 (I453013,I453254,I453124);
nor I_26483 (I453004,I453254,I453180);
nand I_26484 (I453290,I360862,I360850);
and I_26485 (I453307,I453290,I360847);
DFFARX1 I_26486 (I453307,I3035,I453030,I453333,);
not I_26487 (I453341,I453333);
nand I_26488 (I453358,I453341,I453254);
nand I_26489 (I453007,I453341,I453163);
nor I_26490 (I453389,I360865,I360850);
and I_26491 (I453406,I453254,I453389);
nor I_26492 (I453423,I453341,I453406);
DFFARX1 I_26493 (I453423,I3035,I453030,I453016,);
nor I_26494 (I453454,I453056,I453389);
DFFARX1 I_26495 (I453454,I3035,I453030,I453001,);
nor I_26496 (I453485,I453333,I453389);
not I_26497 (I453502,I453485);
nand I_26498 (I453010,I453502,I453358);
not I_26499 (I453557,I3042);
DFFARX1 I_26500 (I638200,I3035,I453557,I453583,);
not I_26501 (I453591,I453583);
nand I_26502 (I453608,I638182,I638182);
and I_26503 (I453625,I453608,I638188);
DFFARX1 I_26504 (I453625,I3035,I453557,I453651,);
DFFARX1 I_26505 (I453651,I3035,I453557,I453546,);
DFFARX1 I_26506 (I638185,I3035,I453557,I453682,);
nand I_26507 (I453690,I453682,I638194);
not I_26508 (I453707,I453690);
DFFARX1 I_26509 (I453707,I3035,I453557,I453733,);
not I_26510 (I453741,I453733);
nor I_26511 (I453549,I453591,I453741);
DFFARX1 I_26512 (I638206,I3035,I453557,I453781,);
nor I_26513 (I453540,I453781,I453651);
nor I_26514 (I453531,I453781,I453707);
nand I_26515 (I453817,I638197,I638191);
and I_26516 (I453834,I453817,I638185);
DFFARX1 I_26517 (I453834,I3035,I453557,I453860,);
not I_26518 (I453868,I453860);
nand I_26519 (I453885,I453868,I453781);
nand I_26520 (I453534,I453868,I453690);
nor I_26521 (I453916,I638203,I638191);
and I_26522 (I453933,I453781,I453916);
nor I_26523 (I453950,I453868,I453933);
DFFARX1 I_26524 (I453950,I3035,I453557,I453543,);
nor I_26525 (I453981,I453583,I453916);
DFFARX1 I_26526 (I453981,I3035,I453557,I453528,);
nor I_26527 (I454012,I453860,I453916);
not I_26528 (I454029,I454012);
nand I_26529 (I453537,I454029,I453885);
not I_26530 (I454084,I3042);
DFFARX1 I_26531 (I414598,I3035,I454084,I454110,);
not I_26532 (I454118,I454110);
nand I_26533 (I454135,I414601,I414598);
and I_26534 (I454152,I454135,I414610);
DFFARX1 I_26535 (I454152,I3035,I454084,I454178,);
DFFARX1 I_26536 (I454178,I3035,I454084,I454073,);
DFFARX1 I_26537 (I414607,I3035,I454084,I454209,);
nand I_26538 (I454217,I454209,I414613);
not I_26539 (I454234,I454217);
DFFARX1 I_26540 (I454234,I3035,I454084,I454260,);
not I_26541 (I454268,I454260);
nor I_26542 (I454076,I454118,I454268);
DFFARX1 I_26543 (I414622,I3035,I454084,I454308,);
nor I_26544 (I454067,I454308,I454178);
nor I_26545 (I454058,I454308,I454234);
nand I_26546 (I454344,I414616,I414604);
and I_26547 (I454361,I454344,I414601);
DFFARX1 I_26548 (I454361,I3035,I454084,I454387,);
not I_26549 (I454395,I454387);
nand I_26550 (I454412,I454395,I454308);
nand I_26551 (I454061,I454395,I454217);
nor I_26552 (I454443,I414619,I414604);
and I_26553 (I454460,I454308,I454443);
nor I_26554 (I454477,I454395,I454460);
DFFARX1 I_26555 (I454477,I3035,I454084,I454070,);
nor I_26556 (I454508,I454110,I454443);
DFFARX1 I_26557 (I454508,I3035,I454084,I454055,);
nor I_26558 (I454539,I454387,I454443);
not I_26559 (I454556,I454539);
nand I_26560 (I454064,I454556,I454412);
not I_26561 (I454611,I3042);
DFFARX1 I_26562 (I112820,I3035,I454611,I454637,);
not I_26563 (I454645,I454637);
nand I_26564 (I454662,I112817,I112835);
and I_26565 (I454679,I454662,I112826);
DFFARX1 I_26566 (I454679,I3035,I454611,I454705,);
DFFARX1 I_26567 (I454705,I3035,I454611,I454600,);
DFFARX1 I_26568 (I112832,I3035,I454611,I454736,);
nand I_26569 (I454744,I454736,I112829);
not I_26570 (I454761,I454744);
DFFARX1 I_26571 (I454761,I3035,I454611,I454787,);
not I_26572 (I454795,I454787);
nor I_26573 (I454603,I454645,I454795);
DFFARX1 I_26574 (I112823,I3035,I454611,I454835,);
nor I_26575 (I454594,I454835,I454705);
nor I_26576 (I454585,I454835,I454761);
nand I_26577 (I454871,I112814,I112838);
and I_26578 (I454888,I454871,I112817);
DFFARX1 I_26579 (I454888,I3035,I454611,I454914,);
not I_26580 (I454922,I454914);
nand I_26581 (I454939,I454922,I454835);
nand I_26582 (I454588,I454922,I454744);
nor I_26583 (I454970,I112814,I112838);
and I_26584 (I454987,I454835,I454970);
nor I_26585 (I455004,I454922,I454987);
DFFARX1 I_26586 (I455004,I3035,I454611,I454597,);
nor I_26587 (I455035,I454637,I454970);
DFFARX1 I_26588 (I455035,I3035,I454611,I454582,);
nor I_26589 (I455066,I454914,I454970);
not I_26590 (I455083,I455066);
nand I_26591 (I454591,I455083,I454939);
not I_26592 (I455138,I3042);
DFFARX1 I_26593 (I418644,I3035,I455138,I455164,);
not I_26594 (I455172,I455164);
nand I_26595 (I455189,I418647,I418644);
and I_26596 (I455206,I455189,I418656);
DFFARX1 I_26597 (I455206,I3035,I455138,I455232,);
DFFARX1 I_26598 (I455232,I3035,I455138,I455127,);
DFFARX1 I_26599 (I418653,I3035,I455138,I455263,);
nand I_26600 (I455271,I455263,I418659);
not I_26601 (I455288,I455271);
DFFARX1 I_26602 (I455288,I3035,I455138,I455314,);
not I_26603 (I455322,I455314);
nor I_26604 (I455130,I455172,I455322);
DFFARX1 I_26605 (I418668,I3035,I455138,I455362,);
nor I_26606 (I455121,I455362,I455232);
nor I_26607 (I455112,I455362,I455288);
nand I_26608 (I455398,I418662,I418650);
and I_26609 (I455415,I455398,I418647);
DFFARX1 I_26610 (I455415,I3035,I455138,I455441,);
not I_26611 (I455449,I455441);
nand I_26612 (I455466,I455449,I455362);
nand I_26613 (I455115,I455449,I455271);
nor I_26614 (I455497,I418665,I418650);
and I_26615 (I455514,I455362,I455497);
nor I_26616 (I455531,I455449,I455514);
DFFARX1 I_26617 (I455531,I3035,I455138,I455124,);
nor I_26618 (I455562,I455164,I455497);
DFFARX1 I_26619 (I455562,I3035,I455138,I455109,);
nor I_26620 (I455593,I455441,I455497);
not I_26621 (I455610,I455593);
nand I_26622 (I455118,I455610,I455466);
not I_26623 (I455665,I3042);
DFFARX1 I_26624 (I128290,I3035,I455665,I455691,);
not I_26625 (I455699,I455691);
nand I_26626 (I455716,I128287,I128305);
and I_26627 (I455733,I455716,I128296);
DFFARX1 I_26628 (I455733,I3035,I455665,I455759,);
DFFARX1 I_26629 (I455759,I3035,I455665,I455654,);
DFFARX1 I_26630 (I128302,I3035,I455665,I455790,);
nand I_26631 (I455798,I455790,I128299);
not I_26632 (I455815,I455798);
DFFARX1 I_26633 (I455815,I3035,I455665,I455841,);
not I_26634 (I455849,I455841);
nor I_26635 (I455657,I455699,I455849);
DFFARX1 I_26636 (I128293,I3035,I455665,I455889,);
nor I_26637 (I455648,I455889,I455759);
nor I_26638 (I455639,I455889,I455815);
nand I_26639 (I455925,I128284,I128308);
and I_26640 (I455942,I455925,I128287);
DFFARX1 I_26641 (I455942,I3035,I455665,I455968,);
not I_26642 (I455976,I455968);
nand I_26643 (I455993,I455976,I455889);
nand I_26644 (I455642,I455976,I455798);
nor I_26645 (I456024,I128284,I128308);
and I_26646 (I456041,I455889,I456024);
nor I_26647 (I456058,I455976,I456041);
DFFARX1 I_26648 (I456058,I3035,I455665,I455651,);
nor I_26649 (I456089,I455691,I456024);
DFFARX1 I_26650 (I456089,I3035,I455665,I455636,);
nor I_26651 (I456120,I455968,I456024);
not I_26652 (I456137,I456120);
nand I_26653 (I455645,I456137,I455993);
not I_26654 (I456192,I3042);
DFFARX1 I_26655 (I122935,I3035,I456192,I456218,);
not I_26656 (I456226,I456218);
nand I_26657 (I456243,I122932,I122950);
and I_26658 (I456260,I456243,I122941);
DFFARX1 I_26659 (I456260,I3035,I456192,I456286,);
DFFARX1 I_26660 (I456286,I3035,I456192,I456181,);
DFFARX1 I_26661 (I122947,I3035,I456192,I456317,);
nand I_26662 (I456325,I456317,I122944);
not I_26663 (I456342,I456325);
DFFARX1 I_26664 (I456342,I3035,I456192,I456368,);
not I_26665 (I456376,I456368);
nor I_26666 (I456184,I456226,I456376);
DFFARX1 I_26667 (I122938,I3035,I456192,I456416,);
nor I_26668 (I456175,I456416,I456286);
nor I_26669 (I456166,I456416,I456342);
nand I_26670 (I456452,I122929,I122953);
and I_26671 (I456469,I456452,I122932);
DFFARX1 I_26672 (I456469,I3035,I456192,I456495,);
not I_26673 (I456503,I456495);
nand I_26674 (I456520,I456503,I456416);
nand I_26675 (I456169,I456503,I456325);
nor I_26676 (I456551,I122929,I122953);
and I_26677 (I456568,I456416,I456551);
nor I_26678 (I456585,I456503,I456568);
DFFARX1 I_26679 (I456585,I3035,I456192,I456178,);
nor I_26680 (I456616,I456218,I456551);
DFFARX1 I_26681 (I456616,I3035,I456192,I456163,);
nor I_26682 (I456647,I456495,I456551);
not I_26683 (I456664,I456647);
nand I_26684 (I456172,I456664,I456520);
not I_26685 (I456719,I3042);
DFFARX1 I_26686 (I276139,I3035,I456719,I456745,);
not I_26687 (I456753,I456745);
nand I_26688 (I456770,I276136,I276145);
and I_26689 (I456787,I456770,I276154);
DFFARX1 I_26690 (I456787,I3035,I456719,I456813,);
DFFARX1 I_26691 (I456813,I3035,I456719,I456708,);
DFFARX1 I_26692 (I276157,I3035,I456719,I456844,);
nand I_26693 (I456852,I456844,I276160);
not I_26694 (I456869,I456852);
DFFARX1 I_26695 (I456869,I3035,I456719,I456895,);
not I_26696 (I456903,I456895);
nor I_26697 (I456711,I456753,I456903);
DFFARX1 I_26698 (I276133,I3035,I456719,I456943,);
nor I_26699 (I456702,I456943,I456813);
nor I_26700 (I456693,I456943,I456869);
nand I_26701 (I456979,I276148,I276151);
and I_26702 (I456996,I456979,I276142);
DFFARX1 I_26703 (I456996,I3035,I456719,I457022,);
not I_26704 (I457030,I457022);
nand I_26705 (I457047,I457030,I456943);
nand I_26706 (I456696,I457030,I456852);
nor I_26707 (I457078,I276133,I276151);
and I_26708 (I457095,I456943,I457078);
nor I_26709 (I457112,I457030,I457095);
DFFARX1 I_26710 (I457112,I3035,I456719,I456705,);
nor I_26711 (I457143,I456745,I457078);
DFFARX1 I_26712 (I457143,I3035,I456719,I456690,);
nor I_26713 (I457174,I457022,I457078);
not I_26714 (I457191,I457174);
nand I_26715 (I456699,I457191,I457047);
not I_26716 (I457246,I3042);
DFFARX1 I_26717 (I585024,I3035,I457246,I457272,);
not I_26718 (I457280,I457272);
nand I_26719 (I457297,I585006,I585006);
and I_26720 (I457314,I457297,I585012);
DFFARX1 I_26721 (I457314,I3035,I457246,I457340,);
DFFARX1 I_26722 (I457340,I3035,I457246,I457235,);
DFFARX1 I_26723 (I585009,I3035,I457246,I457371,);
nand I_26724 (I457379,I457371,I585018);
not I_26725 (I457396,I457379);
DFFARX1 I_26726 (I457396,I3035,I457246,I457422,);
not I_26727 (I457430,I457422);
nor I_26728 (I457238,I457280,I457430);
DFFARX1 I_26729 (I585030,I3035,I457246,I457470,);
nor I_26730 (I457229,I457470,I457340);
nor I_26731 (I457220,I457470,I457396);
nand I_26732 (I457506,I585021,I585015);
and I_26733 (I457523,I457506,I585009);
DFFARX1 I_26734 (I457523,I3035,I457246,I457549,);
not I_26735 (I457557,I457549);
nand I_26736 (I457574,I457557,I457470);
nand I_26737 (I457223,I457557,I457379);
nor I_26738 (I457605,I585027,I585015);
and I_26739 (I457622,I457470,I457605);
nor I_26740 (I457639,I457557,I457622);
DFFARX1 I_26741 (I457639,I3035,I457246,I457232,);
nor I_26742 (I457670,I457272,I457605);
DFFARX1 I_26743 (I457670,I3035,I457246,I457217,);
nor I_26744 (I457701,I457549,I457605);
not I_26745 (I457718,I457701);
nand I_26746 (I457226,I457718,I457574);
not I_26747 (I457773,I3042);
DFFARX1 I_26748 (I250027,I3035,I457773,I457799,);
not I_26749 (I457807,I457799);
nand I_26750 (I457824,I250024,I250033);
and I_26751 (I457841,I457824,I250042);
DFFARX1 I_26752 (I457841,I3035,I457773,I457867,);
DFFARX1 I_26753 (I457867,I3035,I457773,I457762,);
DFFARX1 I_26754 (I250045,I3035,I457773,I457898,);
nand I_26755 (I457906,I457898,I250048);
not I_26756 (I457923,I457906);
DFFARX1 I_26757 (I457923,I3035,I457773,I457949,);
not I_26758 (I457957,I457949);
nor I_26759 (I457765,I457807,I457957);
DFFARX1 I_26760 (I250021,I3035,I457773,I457997,);
nor I_26761 (I457756,I457997,I457867);
nor I_26762 (I457747,I457997,I457923);
nand I_26763 (I458033,I250036,I250039);
and I_26764 (I458050,I458033,I250030);
DFFARX1 I_26765 (I458050,I3035,I457773,I458076,);
not I_26766 (I458084,I458076);
nand I_26767 (I458101,I458084,I457997);
nand I_26768 (I457750,I458084,I457906);
nor I_26769 (I458132,I250021,I250039);
and I_26770 (I458149,I457997,I458132);
nor I_26771 (I458166,I458084,I458149);
DFFARX1 I_26772 (I458166,I3035,I457773,I457759,);
nor I_26773 (I458197,I457799,I458132);
DFFARX1 I_26774 (I458197,I3035,I457773,I457744,);
nor I_26775 (I458228,I458076,I458132);
not I_26776 (I458245,I458228);
nand I_26777 (I457753,I458245,I458101);
not I_26778 (I458300,I3042);
DFFARX1 I_26779 (I644558,I3035,I458300,I458326,);
not I_26780 (I458334,I458326);
nand I_26781 (I458351,I644540,I644540);
and I_26782 (I458368,I458351,I644546);
DFFARX1 I_26783 (I458368,I3035,I458300,I458394,);
DFFARX1 I_26784 (I458394,I3035,I458300,I458289,);
DFFARX1 I_26785 (I644543,I3035,I458300,I458425,);
nand I_26786 (I458433,I458425,I644552);
not I_26787 (I458450,I458433);
DFFARX1 I_26788 (I458450,I3035,I458300,I458476,);
not I_26789 (I458484,I458476);
nor I_26790 (I458292,I458334,I458484);
DFFARX1 I_26791 (I644564,I3035,I458300,I458524,);
nor I_26792 (I458283,I458524,I458394);
nor I_26793 (I458274,I458524,I458450);
nand I_26794 (I458560,I644555,I644549);
and I_26795 (I458577,I458560,I644543);
DFFARX1 I_26796 (I458577,I3035,I458300,I458603,);
not I_26797 (I458611,I458603);
nand I_26798 (I458628,I458611,I458524);
nand I_26799 (I458277,I458611,I458433);
nor I_26800 (I458659,I644561,I644549);
and I_26801 (I458676,I458524,I458659);
nor I_26802 (I458693,I458611,I458676);
DFFARX1 I_26803 (I458693,I3035,I458300,I458286,);
nor I_26804 (I458724,I458326,I458659);
DFFARX1 I_26805 (I458724,I3035,I458300,I458271,);
nor I_26806 (I458755,I458603,I458659);
not I_26807 (I458772,I458755);
nand I_26808 (I458280,I458772,I458628);
not I_26809 (I458827,I3042);
DFFARX1 I_26810 (I496745,I3035,I458827,I458853,);
not I_26811 (I458861,I458853);
nand I_26812 (I458878,I496760,I496742);
and I_26813 (I458895,I458878,I496742);
DFFARX1 I_26814 (I458895,I3035,I458827,I458921,);
DFFARX1 I_26815 (I458921,I3035,I458827,I458816,);
DFFARX1 I_26816 (I496751,I3035,I458827,I458952,);
nand I_26817 (I458960,I458952,I496769);
not I_26818 (I458977,I458960);
DFFARX1 I_26819 (I458977,I3035,I458827,I459003,);
not I_26820 (I459011,I459003);
nor I_26821 (I458819,I458861,I459011);
DFFARX1 I_26822 (I496766,I3035,I458827,I459051,);
nor I_26823 (I458810,I459051,I458921);
nor I_26824 (I458801,I459051,I458977);
nand I_26825 (I459087,I496763,I496754);
and I_26826 (I459104,I459087,I496748);
DFFARX1 I_26827 (I459104,I3035,I458827,I459130,);
not I_26828 (I459138,I459130);
nand I_26829 (I459155,I459138,I459051);
nand I_26830 (I458804,I459138,I458960);
nor I_26831 (I459186,I496757,I496754);
and I_26832 (I459203,I459051,I459186);
nor I_26833 (I459220,I459138,I459203);
DFFARX1 I_26834 (I459220,I3035,I458827,I458813,);
nor I_26835 (I459251,I458853,I459186);
DFFARX1 I_26836 (I459251,I3035,I458827,I458798,);
nor I_26837 (I459282,I459130,I459186);
not I_26838 (I459299,I459282);
nand I_26839 (I458807,I459299,I459155);
not I_26840 (I459354,I3042);
DFFARX1 I_26841 (I646292,I3035,I459354,I459380,);
not I_26842 (I459388,I459380);
nand I_26843 (I459405,I646274,I646274);
and I_26844 (I459422,I459405,I646280);
DFFARX1 I_26845 (I459422,I3035,I459354,I459448,);
DFFARX1 I_26846 (I459448,I3035,I459354,I459343,);
DFFARX1 I_26847 (I646277,I3035,I459354,I459479,);
nand I_26848 (I459487,I459479,I646286);
not I_26849 (I459504,I459487);
DFFARX1 I_26850 (I459504,I3035,I459354,I459530,);
not I_26851 (I459538,I459530);
nor I_26852 (I459346,I459388,I459538);
DFFARX1 I_26853 (I646298,I3035,I459354,I459578,);
nor I_26854 (I459337,I459578,I459448);
nor I_26855 (I459328,I459578,I459504);
nand I_26856 (I459614,I646289,I646283);
and I_26857 (I459631,I459614,I646277);
DFFARX1 I_26858 (I459631,I3035,I459354,I459657,);
not I_26859 (I459665,I459657);
nand I_26860 (I459682,I459665,I459578);
nand I_26861 (I459331,I459665,I459487);
nor I_26862 (I459713,I646295,I646283);
and I_26863 (I459730,I459578,I459713);
nor I_26864 (I459747,I459665,I459730);
DFFARX1 I_26865 (I459747,I3035,I459354,I459340,);
nor I_26866 (I459778,I459380,I459713);
DFFARX1 I_26867 (I459778,I3035,I459354,I459325,);
nor I_26868 (I459809,I459657,I459713);
not I_26869 (I459826,I459809);
nand I_26870 (I459334,I459826,I459682);
not I_26871 (I459881,I3042);
DFFARX1 I_26872 (I139000,I3035,I459881,I459907,);
not I_26873 (I459915,I459907);
nand I_26874 (I459932,I138997,I139015);
and I_26875 (I459949,I459932,I139006);
DFFARX1 I_26876 (I459949,I3035,I459881,I459975,);
DFFARX1 I_26877 (I459975,I3035,I459881,I459870,);
DFFARX1 I_26878 (I139012,I3035,I459881,I460006,);
nand I_26879 (I460014,I460006,I139009);
not I_26880 (I460031,I460014);
DFFARX1 I_26881 (I460031,I3035,I459881,I460057,);
not I_26882 (I460065,I460057);
nor I_26883 (I459873,I459915,I460065);
DFFARX1 I_26884 (I139003,I3035,I459881,I460105,);
nor I_26885 (I459864,I460105,I459975);
nor I_26886 (I459855,I460105,I460031);
nand I_26887 (I460141,I138994,I139018);
and I_26888 (I460158,I460141,I138997);
DFFARX1 I_26889 (I460158,I3035,I459881,I460184,);
not I_26890 (I460192,I460184);
nand I_26891 (I460209,I460192,I460105);
nand I_26892 (I459858,I460192,I460014);
nor I_26893 (I460240,I138994,I139018);
and I_26894 (I460257,I460105,I460240);
nor I_26895 (I460274,I460192,I460257);
DFFARX1 I_26896 (I460274,I3035,I459881,I459867,);
nor I_26897 (I460305,I459907,I460240);
DFFARX1 I_26898 (I460305,I3035,I459881,I459852,);
nor I_26899 (I460336,I460184,I460240);
not I_26900 (I460353,I460336);
nand I_26901 (I459861,I460353,I460209);
not I_26902 (I460408,I3042);
DFFARX1 I_26903 (I525815,I3035,I460408,I460434,);
not I_26904 (I460442,I460434);
nand I_26905 (I460459,I525830,I525812);
and I_26906 (I460476,I460459,I525812);
DFFARX1 I_26907 (I460476,I3035,I460408,I460502,);
DFFARX1 I_26908 (I460502,I3035,I460408,I460397,);
DFFARX1 I_26909 (I525821,I3035,I460408,I460533,);
nand I_26910 (I460541,I460533,I525839);
not I_26911 (I460558,I460541);
DFFARX1 I_26912 (I460558,I3035,I460408,I460584,);
not I_26913 (I460592,I460584);
nor I_26914 (I460400,I460442,I460592);
DFFARX1 I_26915 (I525836,I3035,I460408,I460632,);
nor I_26916 (I460391,I460632,I460502);
nor I_26917 (I460382,I460632,I460558);
nand I_26918 (I460668,I525833,I525824);
and I_26919 (I460685,I460668,I525818);
DFFARX1 I_26920 (I460685,I3035,I460408,I460711,);
not I_26921 (I460719,I460711);
nand I_26922 (I460736,I460719,I460632);
nand I_26923 (I460385,I460719,I460541);
nor I_26924 (I460767,I525827,I525824);
and I_26925 (I460784,I460632,I460767);
nor I_26926 (I460801,I460719,I460784);
DFFARX1 I_26927 (I460801,I3035,I460408,I460394,);
nor I_26928 (I460832,I460434,I460767);
DFFARX1 I_26929 (I460832,I3035,I460408,I460379,);
nor I_26930 (I460863,I460711,I460767);
not I_26931 (I460880,I460863);
nand I_26932 (I460388,I460880,I460736);
not I_26933 (I460935,I3042);
DFFARX1 I_26934 (I617970,I3035,I460935,I460961,);
not I_26935 (I460969,I460961);
nand I_26936 (I460986,I617952,I617952);
and I_26937 (I461003,I460986,I617958);
DFFARX1 I_26938 (I461003,I3035,I460935,I461029,);
DFFARX1 I_26939 (I461029,I3035,I460935,I460924,);
DFFARX1 I_26940 (I617955,I3035,I460935,I461060,);
nand I_26941 (I461068,I461060,I617964);
not I_26942 (I461085,I461068);
DFFARX1 I_26943 (I461085,I3035,I460935,I461111,);
not I_26944 (I461119,I461111);
nor I_26945 (I460927,I460969,I461119);
DFFARX1 I_26946 (I617976,I3035,I460935,I461159,);
nor I_26947 (I460918,I461159,I461029);
nor I_26948 (I460909,I461159,I461085);
nand I_26949 (I461195,I617967,I617961);
and I_26950 (I461212,I461195,I617955);
DFFARX1 I_26951 (I461212,I3035,I460935,I461238,);
not I_26952 (I461246,I461238);
nand I_26953 (I461263,I461246,I461159);
nand I_26954 (I460912,I461246,I461068);
nor I_26955 (I461294,I617973,I617961);
and I_26956 (I461311,I461159,I461294);
nor I_26957 (I461328,I461246,I461311);
DFFARX1 I_26958 (I461328,I3035,I460935,I460921,);
nor I_26959 (I461359,I460961,I461294);
DFFARX1 I_26960 (I461359,I3035,I460935,I460906,);
nor I_26961 (I461390,I461238,I461294);
not I_26962 (I461407,I461390);
nand I_26963 (I460915,I461407,I461263);
not I_26964 (I461462,I3042);
DFFARX1 I_26965 (I176131,I3035,I461462,I461488,);
not I_26966 (I461496,I461488);
nand I_26967 (I461513,I176122,I176122);
and I_26968 (I461530,I461513,I176140);
DFFARX1 I_26969 (I461530,I3035,I461462,I461556,);
DFFARX1 I_26970 (I461556,I3035,I461462,I461451,);
DFFARX1 I_26971 (I176143,I3035,I461462,I461587,);
nand I_26972 (I461595,I461587,I176125);
not I_26973 (I461612,I461595);
DFFARX1 I_26974 (I461612,I3035,I461462,I461638,);
not I_26975 (I461646,I461638);
nor I_26976 (I461454,I461496,I461646);
DFFARX1 I_26977 (I176137,I3035,I461462,I461686,);
nor I_26978 (I461445,I461686,I461556);
nor I_26979 (I461436,I461686,I461612);
nand I_26980 (I461722,I176149,I176128);
and I_26981 (I461739,I461722,I176134);
DFFARX1 I_26982 (I461739,I3035,I461462,I461765,);
not I_26983 (I461773,I461765);
nand I_26984 (I461790,I461773,I461686);
nand I_26985 (I461439,I461773,I461595);
nor I_26986 (I461821,I176146,I176128);
and I_26987 (I461838,I461686,I461821);
nor I_26988 (I461855,I461773,I461838);
DFFARX1 I_26989 (I461855,I3035,I461462,I461448,);
nor I_26990 (I461886,I461488,I461821);
DFFARX1 I_26991 (I461886,I3035,I461462,I461433,);
nor I_26992 (I461917,I461765,I461821);
not I_26993 (I461934,I461917);
nand I_26994 (I461442,I461934,I461790);
not I_26995 (I461989,I3042);
DFFARX1 I_26996 (I12557,I3035,I461989,I462015,);
not I_26997 (I462023,I462015);
nand I_26998 (I462040,I12569,I12572);
and I_26999 (I462057,I462040,I12548);
DFFARX1 I_27000 (I462057,I3035,I461989,I462083,);
DFFARX1 I_27001 (I462083,I3035,I461989,I461978,);
DFFARX1 I_27002 (I12566,I3035,I461989,I462114,);
nand I_27003 (I462122,I462114,I12554);
not I_27004 (I462139,I462122);
DFFARX1 I_27005 (I462139,I3035,I461989,I462165,);
not I_27006 (I462173,I462165);
nor I_27007 (I461981,I462023,I462173);
DFFARX1 I_27008 (I12551,I3035,I461989,I462213,);
nor I_27009 (I461972,I462213,I462083);
nor I_27010 (I461963,I462213,I462139);
nand I_27011 (I462249,I12560,I12551);
and I_27012 (I462266,I462249,I12548);
DFFARX1 I_27013 (I462266,I3035,I461989,I462292,);
not I_27014 (I462300,I462292);
nand I_27015 (I462317,I462300,I462213);
nand I_27016 (I461966,I462300,I462122);
nor I_27017 (I462348,I12563,I12551);
and I_27018 (I462365,I462213,I462348);
nor I_27019 (I462382,I462300,I462365);
DFFARX1 I_27020 (I462382,I3035,I461989,I461975,);
nor I_27021 (I462413,I462015,I462348);
DFFARX1 I_27022 (I462413,I3035,I461989,I461960,);
nor I_27023 (I462444,I462292,I462348);
not I_27024 (I462461,I462444);
nand I_27025 (I461969,I462461,I462317);
not I_27026 (I462516,I3042);
DFFARX1 I_27027 (I142570,I3035,I462516,I462542,);
not I_27028 (I462550,I462542);
nand I_27029 (I462567,I142567,I142585);
and I_27030 (I462584,I462567,I142576);
DFFARX1 I_27031 (I462584,I3035,I462516,I462610,);
DFFARX1 I_27032 (I462610,I3035,I462516,I462505,);
DFFARX1 I_27033 (I142582,I3035,I462516,I462641,);
nand I_27034 (I462649,I462641,I142579);
not I_27035 (I462666,I462649);
DFFARX1 I_27036 (I462666,I3035,I462516,I462692,);
not I_27037 (I462700,I462692);
nor I_27038 (I462508,I462550,I462700);
DFFARX1 I_27039 (I142573,I3035,I462516,I462740,);
nor I_27040 (I462499,I462740,I462610);
nor I_27041 (I462490,I462740,I462666);
nand I_27042 (I462776,I142564,I142588);
and I_27043 (I462793,I462776,I142567);
DFFARX1 I_27044 (I462793,I3035,I462516,I462819,);
not I_27045 (I462827,I462819);
nand I_27046 (I462844,I462827,I462740);
nand I_27047 (I462493,I462827,I462649);
nor I_27048 (I462875,I142564,I142588);
and I_27049 (I462892,I462740,I462875);
nor I_27050 (I462909,I462827,I462892);
DFFARX1 I_27051 (I462909,I3035,I462516,I462502,);
nor I_27052 (I462940,I462542,I462875);
DFFARX1 I_27053 (I462940,I3035,I462516,I462487,);
nor I_27054 (I462971,I462819,I462875);
not I_27055 (I462988,I462971);
nand I_27056 (I462496,I462988,I462844);
not I_27057 (I463043,I3042);
DFFARX1 I_27058 (I151362,I3035,I463043,I463069,);
not I_27059 (I463077,I463069);
nand I_27060 (I463094,I151353,I151353);
and I_27061 (I463111,I463094,I151371);
DFFARX1 I_27062 (I463111,I3035,I463043,I463137,);
DFFARX1 I_27063 (I463137,I3035,I463043,I463032,);
DFFARX1 I_27064 (I151374,I3035,I463043,I463168,);
nand I_27065 (I463176,I463168,I151356);
not I_27066 (I463193,I463176);
DFFARX1 I_27067 (I463193,I3035,I463043,I463219,);
not I_27068 (I463227,I463219);
nor I_27069 (I463035,I463077,I463227);
DFFARX1 I_27070 (I151368,I3035,I463043,I463267,);
nor I_27071 (I463026,I463267,I463137);
nor I_27072 (I463017,I463267,I463193);
nand I_27073 (I463303,I151380,I151359);
and I_27074 (I463320,I463303,I151365);
DFFARX1 I_27075 (I463320,I3035,I463043,I463346,);
not I_27076 (I463354,I463346);
nand I_27077 (I463371,I463354,I463267);
nand I_27078 (I463020,I463354,I463176);
nor I_27079 (I463402,I151377,I151359);
and I_27080 (I463419,I463267,I463402);
nor I_27081 (I463436,I463354,I463419);
DFFARX1 I_27082 (I463436,I3035,I463043,I463029,);
nor I_27083 (I463467,I463069,I463402);
DFFARX1 I_27084 (I463467,I3035,I463043,I463014,);
nor I_27085 (I463498,I463346,I463402);
not I_27086 (I463515,I463498);
nand I_27087 (I463023,I463515,I463371);
not I_27088 (I463570,I3042);
DFFARX1 I_27089 (I1724,I3035,I463570,I463596,);
not I_27090 (I463604,I463596);
nand I_27091 (I463621,I2932,I2028);
and I_27092 (I463638,I463621,I2668);
DFFARX1 I_27093 (I463638,I3035,I463570,I463664,);
DFFARX1 I_27094 (I463664,I3035,I463570,I463559,);
DFFARX1 I_27095 (I1580,I3035,I463570,I463695,);
nand I_27096 (I463703,I463695,I1940);
not I_27097 (I463720,I463703);
DFFARX1 I_27098 (I463720,I3035,I463570,I463746,);
not I_27099 (I463754,I463746);
nor I_27100 (I463562,I463604,I463754);
DFFARX1 I_27101 (I2884,I3035,I463570,I463794,);
nor I_27102 (I463553,I463794,I463664);
nor I_27103 (I463544,I463794,I463720);
nand I_27104 (I463830,I1532,I2660);
and I_27105 (I463847,I463830,I1780);
DFFARX1 I_27106 (I463847,I3035,I463570,I463873,);
not I_27107 (I463881,I463873);
nand I_27108 (I463898,I463881,I463794);
nand I_27109 (I463547,I463881,I463703);
nor I_27110 (I463929,I1404,I2660);
and I_27111 (I463946,I463794,I463929);
nor I_27112 (I463963,I463881,I463946);
DFFARX1 I_27113 (I463963,I3035,I463570,I463556,);
nor I_27114 (I463994,I463596,I463929);
DFFARX1 I_27115 (I463994,I3035,I463570,I463541,);
nor I_27116 (I464025,I463873,I463929);
not I_27117 (I464042,I464025);
nand I_27118 (I463550,I464042,I463898);
not I_27119 (I464097,I3042);
DFFARX1 I_27120 (I563323,I3035,I464097,I464123,);
not I_27121 (I464131,I464123);
nand I_27122 (I464148,I563332,I563320);
and I_27123 (I464165,I464148,I563317);
DFFARX1 I_27124 (I464165,I3035,I464097,I464191,);
DFFARX1 I_27125 (I464191,I3035,I464097,I464086,);
DFFARX1 I_27126 (I563317,I3035,I464097,I464222,);
nand I_27127 (I464230,I464222,I563314);
not I_27128 (I464247,I464230);
DFFARX1 I_27129 (I464247,I3035,I464097,I464273,);
not I_27130 (I464281,I464273);
nor I_27131 (I464089,I464131,I464281);
DFFARX1 I_27132 (I563320,I3035,I464097,I464321,);
nor I_27133 (I464080,I464321,I464191);
nor I_27134 (I464071,I464321,I464247);
nand I_27135 (I464357,I563335,I563326);
and I_27136 (I464374,I464357,I563329);
DFFARX1 I_27137 (I464374,I3035,I464097,I464400,);
not I_27138 (I464408,I464400);
nand I_27139 (I464425,I464408,I464321);
nand I_27140 (I464074,I464408,I464230);
nor I_27141 (I464456,I563314,I563326);
and I_27142 (I464473,I464321,I464456);
nor I_27143 (I464490,I464408,I464473);
DFFARX1 I_27144 (I464490,I3035,I464097,I464083,);
nor I_27145 (I464521,I464123,I464456);
DFFARX1 I_27146 (I464521,I3035,I464097,I464068,);
nor I_27147 (I464552,I464400,I464456);
not I_27148 (I464569,I464552);
nand I_27149 (I464077,I464569,I464425);
not I_27150 (I464624,I3042);
DFFARX1 I_27151 (I59475,I3035,I464624,I464650,);
not I_27152 (I464658,I464650);
nand I_27153 (I464675,I59451,I59460);
and I_27154 (I464692,I464675,I59454);
DFFARX1 I_27155 (I464692,I3035,I464624,I464718,);
DFFARX1 I_27156 (I464718,I3035,I464624,I464613,);
DFFARX1 I_27157 (I59472,I3035,I464624,I464749,);
nand I_27158 (I464757,I464749,I59463);
not I_27159 (I464774,I464757);
DFFARX1 I_27160 (I464774,I3035,I464624,I464800,);
not I_27161 (I464808,I464800);
nor I_27162 (I464616,I464658,I464808);
DFFARX1 I_27163 (I59457,I3035,I464624,I464848,);
nor I_27164 (I464607,I464848,I464718);
nor I_27165 (I464598,I464848,I464774);
nand I_27166 (I464884,I59469,I59466);
and I_27167 (I464901,I464884,I59454);
DFFARX1 I_27168 (I464901,I3035,I464624,I464927,);
not I_27169 (I464935,I464927);
nand I_27170 (I464952,I464935,I464848);
nand I_27171 (I464601,I464935,I464757);
nor I_27172 (I464983,I59451,I59466);
and I_27173 (I465000,I464848,I464983);
nor I_27174 (I465017,I464935,I465000);
DFFARX1 I_27175 (I465017,I3035,I464624,I464610,);
nor I_27176 (I465048,I464650,I464983);
DFFARX1 I_27177 (I465048,I3035,I464624,I464595,);
nor I_27178 (I465079,I464927,I464983);
not I_27179 (I465096,I465079);
nand I_27180 (I464604,I465096,I464952);
not I_27181 (I465151,I3042);
DFFARX1 I_27182 (I66326,I3035,I465151,I465177,);
not I_27183 (I465185,I465177);
nand I_27184 (I465202,I66302,I66311);
and I_27185 (I465219,I465202,I66305);
DFFARX1 I_27186 (I465219,I3035,I465151,I465245,);
DFFARX1 I_27187 (I465245,I3035,I465151,I465140,);
DFFARX1 I_27188 (I66323,I3035,I465151,I465276,);
nand I_27189 (I465284,I465276,I66314);
not I_27190 (I465301,I465284);
DFFARX1 I_27191 (I465301,I3035,I465151,I465327,);
not I_27192 (I465335,I465327);
nor I_27193 (I465143,I465185,I465335);
DFFARX1 I_27194 (I66308,I3035,I465151,I465375,);
nor I_27195 (I465134,I465375,I465245);
nor I_27196 (I465125,I465375,I465301);
nand I_27197 (I465411,I66320,I66317);
and I_27198 (I465428,I465411,I66305);
DFFARX1 I_27199 (I465428,I3035,I465151,I465454,);
not I_27200 (I465462,I465454);
nand I_27201 (I465479,I465462,I465375);
nand I_27202 (I465128,I465462,I465284);
nor I_27203 (I465510,I66302,I66317);
and I_27204 (I465527,I465375,I465510);
nor I_27205 (I465544,I465462,I465527);
DFFARX1 I_27206 (I465544,I3035,I465151,I465137,);
nor I_27207 (I465575,I465177,I465510);
DFFARX1 I_27208 (I465575,I3035,I465151,I465122,);
nor I_27209 (I465606,I465454,I465510);
not I_27210 (I465623,I465606);
nand I_27211 (I465131,I465623,I465479);
not I_27212 (I465678,I3042);
DFFARX1 I_27213 (I52097,I3035,I465678,I465704,);
not I_27214 (I465712,I465704);
nand I_27215 (I465729,I52073,I52082);
and I_27216 (I465746,I465729,I52076);
DFFARX1 I_27217 (I465746,I3035,I465678,I465772,);
DFFARX1 I_27218 (I465772,I3035,I465678,I465667,);
DFFARX1 I_27219 (I52094,I3035,I465678,I465803,);
nand I_27220 (I465811,I465803,I52085);
not I_27221 (I465828,I465811);
DFFARX1 I_27222 (I465828,I3035,I465678,I465854,);
not I_27223 (I465862,I465854);
nor I_27224 (I465670,I465712,I465862);
DFFARX1 I_27225 (I52079,I3035,I465678,I465902,);
nor I_27226 (I465661,I465902,I465772);
nor I_27227 (I465652,I465902,I465828);
nand I_27228 (I465938,I52091,I52088);
and I_27229 (I465955,I465938,I52076);
DFFARX1 I_27230 (I465955,I3035,I465678,I465981,);
not I_27231 (I465989,I465981);
nand I_27232 (I466006,I465989,I465902);
nand I_27233 (I465655,I465989,I465811);
nor I_27234 (I466037,I52073,I52088);
and I_27235 (I466054,I465902,I466037);
nor I_27236 (I466071,I465989,I466054);
DFFARX1 I_27237 (I466071,I3035,I465678,I465664,);
nor I_27238 (I466102,I465704,I466037);
DFFARX1 I_27239 (I466102,I3035,I465678,I465649,);
nor I_27240 (I466133,I465981,I466037);
not I_27241 (I466150,I466133);
nand I_27242 (I465658,I466150,I466006);
not I_27243 (I466205,I3042);
DFFARX1 I_27244 (I712113,I3035,I466205,I466231,);
not I_27245 (I466239,I466231);
nand I_27246 (I466256,I712110,I712119);
and I_27247 (I466273,I466256,I712098);
DFFARX1 I_27248 (I466273,I3035,I466205,I466299,);
DFFARX1 I_27249 (I466299,I3035,I466205,I466194,);
DFFARX1 I_27250 (I712101,I3035,I466205,I466330,);
nand I_27251 (I466338,I466330,I712116);
not I_27252 (I466355,I466338);
DFFARX1 I_27253 (I466355,I3035,I466205,I466381,);
not I_27254 (I466389,I466381);
nor I_27255 (I466197,I466239,I466389);
DFFARX1 I_27256 (I712122,I3035,I466205,I466429,);
nor I_27257 (I466188,I466429,I466299);
nor I_27258 (I466179,I466429,I466355);
nand I_27259 (I466465,I712104,I712125);
and I_27260 (I466482,I466465,I712107);
DFFARX1 I_27261 (I466482,I3035,I466205,I466508,);
not I_27262 (I466516,I466508);
nand I_27263 (I466533,I466516,I466429);
nand I_27264 (I466182,I466516,I466338);
nor I_27265 (I466564,I712098,I712125);
and I_27266 (I466581,I466429,I466564);
nor I_27267 (I466598,I466516,I466581);
DFFARX1 I_27268 (I466598,I3035,I466205,I466191,);
nor I_27269 (I466629,I466231,I466564);
DFFARX1 I_27270 (I466629,I3035,I466205,I466176,);
nor I_27271 (I466660,I466508,I466564);
not I_27272 (I466677,I466660);
nand I_27273 (I466185,I466677,I466533);
not I_27274 (I466732,I3042);
DFFARX1 I_27275 (I2212,I3035,I466732,I466758,);
not I_27276 (I466766,I466758);
nand I_27277 (I466783,I1868,I2940);
and I_27278 (I466800,I466783,I2532);
DFFARX1 I_27279 (I466800,I3035,I466732,I466826,);
DFFARX1 I_27280 (I466826,I3035,I466732,I466721,);
DFFARX1 I_27281 (I1452,I3035,I466732,I466857,);
nand I_27282 (I466865,I466857,I2708);
not I_27283 (I466882,I466865);
DFFARX1 I_27284 (I466882,I3035,I466732,I466908,);
not I_27285 (I466916,I466908);
nor I_27286 (I466724,I466766,I466916);
DFFARX1 I_27287 (I2740,I3035,I466732,I466956,);
nor I_27288 (I466715,I466956,I466826);
nor I_27289 (I466706,I466956,I466882);
nand I_27290 (I466992,I2428,I1420);
and I_27291 (I467009,I466992,I2252);
DFFARX1 I_27292 (I467009,I3035,I466732,I467035,);
not I_27293 (I467043,I467035);
nand I_27294 (I467060,I467043,I466956);
nand I_27295 (I466709,I467043,I466865);
nor I_27296 (I467091,I1964,I1420);
and I_27297 (I467108,I466956,I467091);
nor I_27298 (I467125,I467043,I467108);
DFFARX1 I_27299 (I467125,I3035,I466732,I466718,);
nor I_27300 (I467156,I466758,I467091);
DFFARX1 I_27301 (I467156,I3035,I466732,I466703,);
nor I_27302 (I467187,I467035,I467091);
not I_27303 (I467204,I467187);
nand I_27304 (I466712,I467204,I467060);
not I_27305 (I467259,I3042);
DFFARX1 I_27306 (I111630,I3035,I467259,I467285,);
not I_27307 (I467293,I467285);
nand I_27308 (I467310,I111627,I111645);
and I_27309 (I467327,I467310,I111636);
DFFARX1 I_27310 (I467327,I3035,I467259,I467353,);
DFFARX1 I_27311 (I467353,I3035,I467259,I467248,);
DFFARX1 I_27312 (I111642,I3035,I467259,I467384,);
nand I_27313 (I467392,I467384,I111639);
not I_27314 (I467409,I467392);
DFFARX1 I_27315 (I467409,I3035,I467259,I467435,);
not I_27316 (I467443,I467435);
nor I_27317 (I467251,I467293,I467443);
DFFARX1 I_27318 (I111633,I3035,I467259,I467483,);
nor I_27319 (I467242,I467483,I467353);
nor I_27320 (I467233,I467483,I467409);
nand I_27321 (I467519,I111624,I111648);
and I_27322 (I467536,I467519,I111627);
DFFARX1 I_27323 (I467536,I3035,I467259,I467562,);
not I_27324 (I467570,I467562);
nand I_27325 (I467587,I467570,I467483);
nand I_27326 (I467236,I467570,I467392);
nor I_27327 (I467618,I111624,I111648);
and I_27328 (I467635,I467483,I467618);
nor I_27329 (I467652,I467570,I467635);
DFFARX1 I_27330 (I467652,I3035,I467259,I467245,);
nor I_27331 (I467683,I467285,I467618);
DFFARX1 I_27332 (I467683,I3035,I467259,I467230,);
nor I_27333 (I467714,I467562,I467618);
not I_27334 (I467731,I467714);
nand I_27335 (I467239,I467731,I467587);
not I_27336 (I467786,I3042);
DFFARX1 I_27337 (I500621,I3035,I467786,I467812,);
not I_27338 (I467820,I467812);
nand I_27339 (I467837,I500636,I500618);
and I_27340 (I467854,I467837,I500618);
DFFARX1 I_27341 (I467854,I3035,I467786,I467880,);
DFFARX1 I_27342 (I467880,I3035,I467786,I467775,);
DFFARX1 I_27343 (I500627,I3035,I467786,I467911,);
nand I_27344 (I467919,I467911,I500645);
not I_27345 (I467936,I467919);
DFFARX1 I_27346 (I467936,I3035,I467786,I467962,);
not I_27347 (I467970,I467962);
nor I_27348 (I467778,I467820,I467970);
DFFARX1 I_27349 (I500642,I3035,I467786,I468010,);
nor I_27350 (I467769,I468010,I467880);
nor I_27351 (I467760,I468010,I467936);
nand I_27352 (I468046,I500639,I500630);
and I_27353 (I468063,I468046,I500624);
DFFARX1 I_27354 (I468063,I3035,I467786,I468089,);
not I_27355 (I468097,I468089);
nand I_27356 (I468114,I468097,I468010);
nand I_27357 (I467763,I468097,I467919);
nor I_27358 (I468145,I500633,I500630);
and I_27359 (I468162,I468010,I468145);
nor I_27360 (I468179,I468097,I468162);
DFFARX1 I_27361 (I468179,I3035,I467786,I467772,);
nor I_27362 (I468210,I467812,I468145);
DFFARX1 I_27363 (I468210,I3035,I467786,I467757,);
nor I_27364 (I468241,I468089,I468145);
not I_27365 (I468258,I468241);
nand I_27366 (I467766,I468258,I468114);
not I_27367 (I468313,I3042);
DFFARX1 I_27368 (I294227,I3035,I468313,I468339,);
not I_27369 (I468347,I468339);
nand I_27370 (I468364,I294245,I294236);
and I_27371 (I468381,I468364,I294239);
DFFARX1 I_27372 (I468381,I3035,I468313,I468407,);
DFFARX1 I_27373 (I468407,I3035,I468313,I468302,);
DFFARX1 I_27374 (I294233,I3035,I468313,I468438,);
nand I_27375 (I468446,I468438,I294224);
not I_27376 (I468463,I468446);
DFFARX1 I_27377 (I468463,I3035,I468313,I468489,);
not I_27378 (I468497,I468489);
nor I_27379 (I468305,I468347,I468497);
DFFARX1 I_27380 (I294230,I3035,I468313,I468537,);
nor I_27381 (I468296,I468537,I468407);
nor I_27382 (I468287,I468537,I468463);
nand I_27383 (I468573,I294224,I294221);
and I_27384 (I468590,I468573,I294242);
DFFARX1 I_27385 (I468590,I3035,I468313,I468616,);
not I_27386 (I468624,I468616);
nand I_27387 (I468641,I468624,I468537);
nand I_27388 (I468290,I468624,I468446);
nor I_27389 (I468672,I294221,I294221);
and I_27390 (I468689,I468537,I468672);
nor I_27391 (I468706,I468624,I468689);
DFFARX1 I_27392 (I468706,I3035,I468313,I468299,);
nor I_27393 (I468737,I468339,I468672);
DFFARX1 I_27394 (I468737,I3035,I468313,I468284,);
nor I_27395 (I468768,I468616,I468672);
not I_27396 (I468785,I468768);
nand I_27397 (I468293,I468785,I468641);
not I_27398 (I468840,I3042);
DFFARX1 I_27399 (I344082,I3035,I468840,I468866,);
not I_27400 (I468874,I468866);
nand I_27401 (I468891,I344085,I344082);
and I_27402 (I468908,I468891,I344094);
DFFARX1 I_27403 (I468908,I3035,I468840,I468934,);
DFFARX1 I_27404 (I468934,I3035,I468840,I468829,);
DFFARX1 I_27405 (I344091,I3035,I468840,I468965,);
nand I_27406 (I468973,I468965,I344097);
not I_27407 (I468990,I468973);
DFFARX1 I_27408 (I468990,I3035,I468840,I469016,);
not I_27409 (I469024,I469016);
nor I_27410 (I468832,I468874,I469024);
DFFARX1 I_27411 (I344106,I3035,I468840,I469064,);
nor I_27412 (I468823,I469064,I468934);
nor I_27413 (I468814,I469064,I468990);
nand I_27414 (I469100,I344100,I344088);
and I_27415 (I469117,I469100,I344085);
DFFARX1 I_27416 (I469117,I3035,I468840,I469143,);
not I_27417 (I469151,I469143);
nand I_27418 (I469168,I469151,I469064);
nand I_27419 (I468817,I469151,I468973);
nor I_27420 (I469199,I344103,I344088);
and I_27421 (I469216,I469064,I469199);
nor I_27422 (I469233,I469151,I469216);
DFFARX1 I_27423 (I469233,I3035,I468840,I468826,);
nor I_27424 (I469264,I468866,I469199);
DFFARX1 I_27425 (I469264,I3035,I468840,I468811,);
nor I_27426 (I469295,I469143,I469199);
not I_27427 (I469312,I469295);
nand I_27428 (I468820,I469312,I469168);
not I_27429 (I469367,I3042);
DFFARX1 I_27430 (I710923,I3035,I469367,I469393,);
not I_27431 (I469401,I469393);
nand I_27432 (I469418,I710920,I710929);
and I_27433 (I469435,I469418,I710908);
DFFARX1 I_27434 (I469435,I3035,I469367,I469461,);
DFFARX1 I_27435 (I469461,I3035,I469367,I469356,);
DFFARX1 I_27436 (I710911,I3035,I469367,I469492,);
nand I_27437 (I469500,I469492,I710926);
not I_27438 (I469517,I469500);
DFFARX1 I_27439 (I469517,I3035,I469367,I469543,);
not I_27440 (I469551,I469543);
nor I_27441 (I469359,I469401,I469551);
DFFARX1 I_27442 (I710932,I3035,I469367,I469591,);
nor I_27443 (I469350,I469591,I469461);
nor I_27444 (I469341,I469591,I469517);
nand I_27445 (I469627,I710914,I710935);
and I_27446 (I469644,I469627,I710917);
DFFARX1 I_27447 (I469644,I3035,I469367,I469670,);
not I_27448 (I469678,I469670);
nand I_27449 (I469695,I469678,I469591);
nand I_27450 (I469344,I469678,I469500);
nor I_27451 (I469726,I710908,I710935);
and I_27452 (I469743,I469591,I469726);
nor I_27453 (I469760,I469678,I469743);
DFFARX1 I_27454 (I469760,I3035,I469367,I469353,);
nor I_27455 (I469791,I469393,I469726);
DFFARX1 I_27456 (I469791,I3035,I469367,I469338,);
nor I_27457 (I469822,I469670,I469726);
not I_27458 (I469839,I469822);
nand I_27459 (I469347,I469839,I469695);
not I_27460 (I469894,I3042);
DFFARX1 I_27461 (I334271,I3035,I469894,I469920,);
not I_27462 (I469928,I469920);
nand I_27463 (I469945,I334256,I334277);
and I_27464 (I469962,I469945,I334265);
DFFARX1 I_27465 (I469962,I3035,I469894,I469988,);
DFFARX1 I_27466 (I469988,I3035,I469894,I469883,);
DFFARX1 I_27467 (I334259,I3035,I469894,I470019,);
nand I_27468 (I470027,I470019,I334268);
not I_27469 (I470044,I470027);
DFFARX1 I_27470 (I470044,I3035,I469894,I470070,);
not I_27471 (I470078,I470070);
nor I_27472 (I469886,I469928,I470078);
DFFARX1 I_27473 (I334274,I3035,I469894,I470118,);
nor I_27474 (I469877,I470118,I469988);
nor I_27475 (I469868,I470118,I470044);
nand I_27476 (I470154,I334256,I334259);
and I_27477 (I470171,I470154,I334280);
DFFARX1 I_27478 (I470171,I3035,I469894,I470197,);
not I_27479 (I470205,I470197);
nand I_27480 (I470222,I470205,I470118);
nand I_27481 (I469871,I470205,I470027);
nor I_27482 (I470253,I334262,I334259);
and I_27483 (I470270,I470118,I470253);
nor I_27484 (I470287,I470205,I470270);
DFFARX1 I_27485 (I470287,I3035,I469894,I469880,);
nor I_27486 (I470318,I469920,I470253);
DFFARX1 I_27487 (I470318,I3035,I469894,I469865,);
nor I_27488 (I470349,I470197,I470253);
not I_27489 (I470366,I470349);
nand I_27490 (I469874,I470366,I470222);
not I_27491 (I470421,I3042);
DFFARX1 I_27492 (I322133,I3035,I470421,I470447,);
not I_27493 (I470455,I470447);
nand I_27494 (I470472,I322118,I322139);
and I_27495 (I470489,I470472,I322127);
DFFARX1 I_27496 (I470489,I3035,I470421,I470515,);
DFFARX1 I_27497 (I470515,I3035,I470421,I470410,);
DFFARX1 I_27498 (I322121,I3035,I470421,I470546,);
nand I_27499 (I470554,I470546,I322130);
not I_27500 (I470571,I470554);
DFFARX1 I_27501 (I470571,I3035,I470421,I470597,);
not I_27502 (I470605,I470597);
nor I_27503 (I470413,I470455,I470605);
DFFARX1 I_27504 (I322136,I3035,I470421,I470645,);
nor I_27505 (I470404,I470645,I470515);
nor I_27506 (I470395,I470645,I470571);
nand I_27507 (I470681,I322118,I322121);
and I_27508 (I470698,I470681,I322142);
DFFARX1 I_27509 (I470698,I3035,I470421,I470724,);
not I_27510 (I470732,I470724);
nand I_27511 (I470749,I470732,I470645);
nand I_27512 (I470398,I470732,I470554);
nor I_27513 (I470780,I322124,I322121);
and I_27514 (I470797,I470645,I470780);
nor I_27515 (I470814,I470732,I470797);
DFFARX1 I_27516 (I470814,I3035,I470421,I470407,);
nor I_27517 (I470845,I470447,I470780);
DFFARX1 I_27518 (I470845,I3035,I470421,I470392,);
nor I_27519 (I470876,I470724,I470780);
not I_27520 (I470893,I470876);
nand I_27521 (I470401,I470893,I470749);
not I_27522 (I470948,I3042);
DFFARX1 I_27523 (I700808,I3035,I470948,I470974,);
not I_27524 (I470982,I470974);
nand I_27525 (I470999,I700805,I700814);
and I_27526 (I471016,I470999,I700793);
DFFARX1 I_27527 (I471016,I3035,I470948,I471042,);
DFFARX1 I_27528 (I471042,I3035,I470948,I470937,);
DFFARX1 I_27529 (I700796,I3035,I470948,I471073,);
nand I_27530 (I471081,I471073,I700811);
not I_27531 (I471098,I471081);
DFFARX1 I_27532 (I471098,I3035,I470948,I471124,);
not I_27533 (I471132,I471124);
nor I_27534 (I470940,I470982,I471132);
DFFARX1 I_27535 (I700817,I3035,I470948,I471172,);
nor I_27536 (I470931,I471172,I471042);
nor I_27537 (I470922,I471172,I471098);
nand I_27538 (I471208,I700799,I700820);
and I_27539 (I471225,I471208,I700802);
DFFARX1 I_27540 (I471225,I3035,I470948,I471251,);
not I_27541 (I471259,I471251);
nand I_27542 (I471276,I471259,I471172);
nand I_27543 (I470925,I471259,I471081);
nor I_27544 (I471307,I700793,I700820);
and I_27545 (I471324,I471172,I471307);
nor I_27546 (I471341,I471259,I471324);
DFFARX1 I_27547 (I471341,I3035,I470948,I470934,);
nor I_27548 (I471372,I470974,I471307);
DFFARX1 I_27549 (I471372,I3035,I470948,I470919,);
nor I_27550 (I471403,I471251,I471307);
not I_27551 (I471420,I471403);
nand I_27552 (I470928,I471420,I471276);
not I_27553 (I471475,I3042);
DFFARX1 I_27554 (I532275,I3035,I471475,I471501,);
not I_27555 (I471509,I471501);
nand I_27556 (I471526,I532290,I532272);
and I_27557 (I471543,I471526,I532272);
DFFARX1 I_27558 (I471543,I3035,I471475,I471569,);
DFFARX1 I_27559 (I471569,I3035,I471475,I471464,);
DFFARX1 I_27560 (I532281,I3035,I471475,I471600,);
nand I_27561 (I471608,I471600,I532299);
not I_27562 (I471625,I471608);
DFFARX1 I_27563 (I471625,I3035,I471475,I471651,);
not I_27564 (I471659,I471651);
nor I_27565 (I471467,I471509,I471659);
DFFARX1 I_27566 (I532296,I3035,I471475,I471699,);
nor I_27567 (I471458,I471699,I471569);
nor I_27568 (I471449,I471699,I471625);
nand I_27569 (I471735,I532293,I532284);
and I_27570 (I471752,I471735,I532278);
DFFARX1 I_27571 (I471752,I3035,I471475,I471778,);
not I_27572 (I471786,I471778);
nand I_27573 (I471803,I471786,I471699);
nand I_27574 (I471452,I471786,I471608);
nor I_27575 (I471834,I532287,I532284);
and I_27576 (I471851,I471699,I471834);
nor I_27577 (I471868,I471786,I471851);
DFFARX1 I_27578 (I471868,I3035,I471475,I471461,);
nor I_27579 (I471899,I471501,I471834);
DFFARX1 I_27580 (I471899,I3035,I471475,I471446,);
nor I_27581 (I471930,I471778,I471834);
not I_27582 (I471947,I471930);
nand I_27583 (I471455,I471947,I471803);
not I_27584 (I472002,I3042);
DFFARX1 I_27585 (I615080,I3035,I472002,I472028,);
not I_27586 (I472036,I472028);
nand I_27587 (I472053,I615062,I615062);
and I_27588 (I472070,I472053,I615068);
DFFARX1 I_27589 (I472070,I3035,I472002,I472096,);
DFFARX1 I_27590 (I472096,I3035,I472002,I471991,);
DFFARX1 I_27591 (I615065,I3035,I472002,I472127,);
nand I_27592 (I472135,I472127,I615074);
not I_27593 (I472152,I472135);
DFFARX1 I_27594 (I472152,I3035,I472002,I472178,);
not I_27595 (I472186,I472178);
nor I_27596 (I471994,I472036,I472186);
DFFARX1 I_27597 (I615086,I3035,I472002,I472226,);
nor I_27598 (I471985,I472226,I472096);
nor I_27599 (I471976,I472226,I472152);
nand I_27600 (I472262,I615077,I615071);
and I_27601 (I472279,I472262,I615065);
DFFARX1 I_27602 (I472279,I3035,I472002,I472305,);
not I_27603 (I472313,I472305);
nand I_27604 (I472330,I472313,I472226);
nand I_27605 (I471979,I472313,I472135);
nor I_27606 (I472361,I615083,I615071);
and I_27607 (I472378,I472226,I472361);
nor I_27608 (I472395,I472313,I472378);
DFFARX1 I_27609 (I472395,I3035,I472002,I471988,);
nor I_27610 (I472426,I472028,I472361);
DFFARX1 I_27611 (I472426,I3035,I472002,I471973,);
nor I_27612 (I472457,I472305,I472361);
not I_27613 (I472474,I472457);
nand I_27614 (I471982,I472474,I472330);
not I_27615 (I472529,I3042);
DFFARX1 I_27616 (I22570,I3035,I472529,I472555,);
not I_27617 (I472563,I472555);
nand I_27618 (I472580,I22582,I22585);
and I_27619 (I472597,I472580,I22561);
DFFARX1 I_27620 (I472597,I3035,I472529,I472623,);
DFFARX1 I_27621 (I472623,I3035,I472529,I472518,);
DFFARX1 I_27622 (I22579,I3035,I472529,I472654,);
nand I_27623 (I472662,I472654,I22567);
not I_27624 (I472679,I472662);
DFFARX1 I_27625 (I472679,I3035,I472529,I472705,);
not I_27626 (I472713,I472705);
nor I_27627 (I472521,I472563,I472713);
DFFARX1 I_27628 (I22564,I3035,I472529,I472753,);
nor I_27629 (I472512,I472753,I472623);
nor I_27630 (I472503,I472753,I472679);
nand I_27631 (I472789,I22573,I22564);
and I_27632 (I472806,I472789,I22561);
DFFARX1 I_27633 (I472806,I3035,I472529,I472832,);
not I_27634 (I472840,I472832);
nand I_27635 (I472857,I472840,I472753);
nand I_27636 (I472506,I472840,I472662);
nor I_27637 (I472888,I22576,I22564);
and I_27638 (I472905,I472753,I472888);
nor I_27639 (I472922,I472840,I472905);
DFFARX1 I_27640 (I472922,I3035,I472529,I472515,);
nor I_27641 (I472953,I472555,I472888);
DFFARX1 I_27642 (I472953,I3035,I472529,I472500,);
nor I_27643 (I472984,I472832,I472888);
not I_27644 (I473001,I472984);
nand I_27645 (I472509,I473001,I472857);
not I_27646 (I473056,I3042);
DFFARX1 I_27647 (I336583,I3035,I473056,I473082,);
not I_27648 (I473090,I473082);
nand I_27649 (I473107,I336568,I336589);
and I_27650 (I473124,I473107,I336577);
DFFARX1 I_27651 (I473124,I3035,I473056,I473150,);
DFFARX1 I_27652 (I473150,I3035,I473056,I473045,);
DFFARX1 I_27653 (I336571,I3035,I473056,I473181,);
nand I_27654 (I473189,I473181,I336580);
not I_27655 (I473206,I473189);
DFFARX1 I_27656 (I473206,I3035,I473056,I473232,);
not I_27657 (I473240,I473232);
nor I_27658 (I473048,I473090,I473240);
DFFARX1 I_27659 (I336586,I3035,I473056,I473280,);
nor I_27660 (I473039,I473280,I473150);
nor I_27661 (I473030,I473280,I473206);
nand I_27662 (I473316,I336568,I336571);
and I_27663 (I473333,I473316,I336592);
DFFARX1 I_27664 (I473333,I3035,I473056,I473359,);
not I_27665 (I473367,I473359);
nand I_27666 (I473384,I473367,I473280);
nand I_27667 (I473033,I473367,I473189);
nor I_27668 (I473415,I336574,I336571);
and I_27669 (I473432,I473280,I473415);
nor I_27670 (I473449,I473367,I473432);
DFFARX1 I_27671 (I473449,I3035,I473056,I473042,);
nor I_27672 (I473480,I473082,I473415);
DFFARX1 I_27673 (I473480,I3035,I473056,I473027,);
nor I_27674 (I473511,I473359,I473415);
not I_27675 (I473528,I473511);
nand I_27676 (I473036,I473528,I473384);
not I_27677 (I473583,I3042);
DFFARX1 I_27678 (I14138,I3035,I473583,I473609,);
not I_27679 (I473617,I473609);
nand I_27680 (I473634,I14150,I14153);
and I_27681 (I473651,I473634,I14129);
DFFARX1 I_27682 (I473651,I3035,I473583,I473677,);
DFFARX1 I_27683 (I473677,I3035,I473583,I473572,);
DFFARX1 I_27684 (I14147,I3035,I473583,I473708,);
nand I_27685 (I473716,I473708,I14135);
not I_27686 (I473733,I473716);
DFFARX1 I_27687 (I473733,I3035,I473583,I473759,);
not I_27688 (I473767,I473759);
nor I_27689 (I473575,I473617,I473767);
DFFARX1 I_27690 (I14132,I3035,I473583,I473807,);
nor I_27691 (I473566,I473807,I473677);
nor I_27692 (I473557,I473807,I473733);
nand I_27693 (I473843,I14141,I14132);
and I_27694 (I473860,I473843,I14129);
DFFARX1 I_27695 (I473860,I3035,I473583,I473886,);
not I_27696 (I473894,I473886);
nand I_27697 (I473911,I473894,I473807);
nand I_27698 (I473560,I473894,I473716);
nor I_27699 (I473942,I14144,I14132);
and I_27700 (I473959,I473807,I473942);
nor I_27701 (I473976,I473894,I473959);
DFFARX1 I_27702 (I473976,I3035,I473583,I473569,);
nor I_27703 (I474007,I473609,I473942);
DFFARX1 I_27704 (I474007,I3035,I473583,I473554,);
nor I_27705 (I474038,I473886,I473942);
not I_27706 (I474055,I474038);
nand I_27707 (I473563,I474055,I473911);
not I_27708 (I474110,I3042);
DFFARX1 I_27709 (I638778,I3035,I474110,I474136,);
not I_27710 (I474144,I474136);
nand I_27711 (I474161,I638760,I638760);
and I_27712 (I474178,I474161,I638766);
DFFARX1 I_27713 (I474178,I3035,I474110,I474204,);
DFFARX1 I_27714 (I474204,I3035,I474110,I474099,);
DFFARX1 I_27715 (I638763,I3035,I474110,I474235,);
nand I_27716 (I474243,I474235,I638772);
not I_27717 (I474260,I474243);
DFFARX1 I_27718 (I474260,I3035,I474110,I474286,);
not I_27719 (I474294,I474286);
nor I_27720 (I474102,I474144,I474294);
DFFARX1 I_27721 (I638784,I3035,I474110,I474334,);
nor I_27722 (I474093,I474334,I474204);
nor I_27723 (I474084,I474334,I474260);
nand I_27724 (I474370,I638775,I638769);
and I_27725 (I474387,I474370,I638763);
DFFARX1 I_27726 (I474387,I3035,I474110,I474413,);
not I_27727 (I474421,I474413);
nand I_27728 (I474438,I474421,I474334);
nand I_27729 (I474087,I474421,I474243);
nor I_27730 (I474469,I638781,I638769);
and I_27731 (I474486,I474334,I474469);
nor I_27732 (I474503,I474421,I474486);
DFFARX1 I_27733 (I474503,I3035,I474110,I474096,);
nor I_27734 (I474534,I474136,I474469);
DFFARX1 I_27735 (I474534,I3035,I474110,I474081,);
nor I_27736 (I474565,I474413,I474469);
not I_27737 (I474582,I474565);
nand I_27738 (I474090,I474582,I474438);
not I_27739 (I474637,I3042);
DFFARX1 I_27740 (I346394,I3035,I474637,I474663,);
not I_27741 (I474671,I474663);
nand I_27742 (I474688,I346397,I346394);
and I_27743 (I474705,I474688,I346406);
DFFARX1 I_27744 (I474705,I3035,I474637,I474731,);
DFFARX1 I_27745 (I474731,I3035,I474637,I474626,);
DFFARX1 I_27746 (I346403,I3035,I474637,I474762,);
nand I_27747 (I474770,I474762,I346409);
not I_27748 (I474787,I474770);
DFFARX1 I_27749 (I474787,I3035,I474637,I474813,);
not I_27750 (I474821,I474813);
nor I_27751 (I474629,I474671,I474821);
DFFARX1 I_27752 (I346418,I3035,I474637,I474861,);
nor I_27753 (I474620,I474861,I474731);
nor I_27754 (I474611,I474861,I474787);
nand I_27755 (I474897,I346412,I346400);
and I_27756 (I474914,I474897,I346397);
DFFARX1 I_27757 (I474914,I3035,I474637,I474940,);
not I_27758 (I474948,I474940);
nand I_27759 (I474965,I474948,I474861);
nand I_27760 (I474614,I474948,I474770);
nor I_27761 (I474996,I346415,I346400);
and I_27762 (I475013,I474861,I474996);
nor I_27763 (I475030,I474948,I475013);
DFFARX1 I_27764 (I475030,I3035,I474637,I474623,);
nor I_27765 (I475061,I474663,I474996);
DFFARX1 I_27766 (I475061,I3035,I474637,I474608,);
nor I_27767 (I475092,I474940,I474996);
not I_27768 (I475109,I475092);
nand I_27769 (I474617,I475109,I474965);
not I_27770 (I475164,I3042);
DFFARX1 I_27771 (I498037,I3035,I475164,I475190,);
not I_27772 (I475198,I475190);
nand I_27773 (I475215,I498052,I498034);
and I_27774 (I475232,I475215,I498034);
DFFARX1 I_27775 (I475232,I3035,I475164,I475258,);
DFFARX1 I_27776 (I475258,I3035,I475164,I475153,);
DFFARX1 I_27777 (I498043,I3035,I475164,I475289,);
nand I_27778 (I475297,I475289,I498061);
not I_27779 (I475314,I475297);
DFFARX1 I_27780 (I475314,I3035,I475164,I475340,);
not I_27781 (I475348,I475340);
nor I_27782 (I475156,I475198,I475348);
DFFARX1 I_27783 (I498058,I3035,I475164,I475388,);
nor I_27784 (I475147,I475388,I475258);
nor I_27785 (I475138,I475388,I475314);
nand I_27786 (I475424,I498055,I498046);
and I_27787 (I475441,I475424,I498040);
DFFARX1 I_27788 (I475441,I3035,I475164,I475467,);
not I_27789 (I475475,I475467);
nand I_27790 (I475492,I475475,I475388);
nand I_27791 (I475141,I475475,I475297);
nor I_27792 (I475523,I498049,I498046);
and I_27793 (I475540,I475388,I475523);
nor I_27794 (I475557,I475475,I475540);
DFFARX1 I_27795 (I475557,I3035,I475164,I475150,);
nor I_27796 (I475588,I475190,I475523);
DFFARX1 I_27797 (I475588,I3035,I475164,I475135,);
nor I_27798 (I475619,I475467,I475523);
not I_27799 (I475636,I475619);
nand I_27800 (I475144,I475636,I475492);
not I_27801 (I475691,I3042);
DFFARX1 I_27802 (I200373,I3035,I475691,I475717,);
not I_27803 (I475725,I475717);
nand I_27804 (I475742,I200364,I200364);
and I_27805 (I475759,I475742,I200382);
DFFARX1 I_27806 (I475759,I3035,I475691,I475785,);
DFFARX1 I_27807 (I475785,I3035,I475691,I475680,);
DFFARX1 I_27808 (I200385,I3035,I475691,I475816,);
nand I_27809 (I475824,I475816,I200367);
not I_27810 (I475841,I475824);
DFFARX1 I_27811 (I475841,I3035,I475691,I475867,);
not I_27812 (I475875,I475867);
nor I_27813 (I475683,I475725,I475875);
DFFARX1 I_27814 (I200379,I3035,I475691,I475915,);
nor I_27815 (I475674,I475915,I475785);
nor I_27816 (I475665,I475915,I475841);
nand I_27817 (I475951,I200391,I200370);
and I_27818 (I475968,I475951,I200376);
DFFARX1 I_27819 (I475968,I3035,I475691,I475994,);
not I_27820 (I476002,I475994);
nand I_27821 (I476019,I476002,I475915);
nand I_27822 (I475668,I476002,I475824);
nor I_27823 (I476050,I200388,I200370);
and I_27824 (I476067,I475915,I476050);
nor I_27825 (I476084,I476002,I476067);
DFFARX1 I_27826 (I476084,I3035,I475691,I475677,);
nor I_27827 (I476115,I475717,I476050);
DFFARX1 I_27828 (I476115,I3035,I475691,I475662,);
nor I_27829 (I476146,I475994,I476050);
not I_27830 (I476163,I476146);
nand I_27831 (I475671,I476163,I476019);
not I_27832 (I476218,I3042);
DFFARX1 I_27833 (I622594,I3035,I476218,I476244,);
not I_27834 (I476252,I476244);
nand I_27835 (I476269,I622576,I622576);
and I_27836 (I476286,I476269,I622582);
DFFARX1 I_27837 (I476286,I3035,I476218,I476312,);
DFFARX1 I_27838 (I476312,I3035,I476218,I476207,);
DFFARX1 I_27839 (I622579,I3035,I476218,I476343,);
nand I_27840 (I476351,I476343,I622588);
not I_27841 (I476368,I476351);
DFFARX1 I_27842 (I476368,I3035,I476218,I476394,);
not I_27843 (I476402,I476394);
nor I_27844 (I476210,I476252,I476402);
DFFARX1 I_27845 (I622600,I3035,I476218,I476442,);
nor I_27846 (I476201,I476442,I476312);
nor I_27847 (I476192,I476442,I476368);
nand I_27848 (I476478,I622591,I622585);
and I_27849 (I476495,I476478,I622579);
DFFARX1 I_27850 (I476495,I3035,I476218,I476521,);
not I_27851 (I476529,I476521);
nand I_27852 (I476546,I476529,I476442);
nand I_27853 (I476195,I476529,I476351);
nor I_27854 (I476577,I622597,I622585);
and I_27855 (I476594,I476442,I476577);
nor I_27856 (I476611,I476529,I476594);
DFFARX1 I_27857 (I476611,I3035,I476218,I476204,);
nor I_27858 (I476642,I476244,I476577);
DFFARX1 I_27859 (I476642,I3035,I476218,I476189,);
nor I_27860 (I476673,I476521,I476577);
not I_27861 (I476690,I476673);
nand I_27862 (I476198,I476690,I476546);
not I_27863 (I476751,I3042);
DFFARX1 I_27864 (I34155,I3035,I476751,I476777,);
DFFARX1 I_27865 (I34161,I3035,I476751,I476794,);
not I_27866 (I476802,I476794);
not I_27867 (I476819,I34179);
nor I_27868 (I476836,I476819,I34158);
not I_27869 (I476853,I34164);
nor I_27870 (I476870,I476836,I34170);
nor I_27871 (I476887,I476794,I476870);
DFFARX1 I_27872 (I476887,I3035,I476751,I476737,);
nor I_27873 (I476918,I34170,I34158);
nand I_27874 (I476935,I476918,I34179);
DFFARX1 I_27875 (I476935,I3035,I476751,I476740,);
nor I_27876 (I476966,I476853,I34170);
nand I_27877 (I476983,I476966,I34176);
nor I_27878 (I477000,I476777,I476983);
DFFARX1 I_27879 (I477000,I3035,I476751,I476716,);
not I_27880 (I477031,I476983);
nand I_27881 (I476728,I476794,I477031);
DFFARX1 I_27882 (I476983,I3035,I476751,I477071,);
not I_27883 (I477079,I477071);
not I_27884 (I477096,I34170);
not I_27885 (I477113,I34158);
nor I_27886 (I477130,I477113,I34164);
nor I_27887 (I476743,I477079,I477130);
nor I_27888 (I477161,I477113,I34167);
and I_27889 (I477178,I477161,I34155);
or I_27890 (I477195,I477178,I34173);
DFFARX1 I_27891 (I477195,I3035,I476751,I477221,);
nor I_27892 (I476731,I477221,I476777);
not I_27893 (I477243,I477221);
and I_27894 (I477260,I477243,I476777);
nor I_27895 (I476725,I476802,I477260);
nand I_27896 (I477291,I477243,I476853);
nor I_27897 (I476719,I477113,I477291);
nand I_27898 (I476722,I477243,I477031);
nand I_27899 (I477336,I476853,I34158);
nor I_27900 (I476734,I477096,I477336);
not I_27901 (I477397,I3042);
DFFARX1 I_27902 (I168744,I3035,I477397,I477423,);
DFFARX1 I_27903 (I168750,I3035,I477397,I477440,);
not I_27904 (I477448,I477440);
not I_27905 (I477465,I168771);
nor I_27906 (I477482,I477465,I168759);
not I_27907 (I477499,I168768);
nor I_27908 (I477516,I477482,I168753);
nor I_27909 (I477533,I477440,I477516);
DFFARX1 I_27910 (I477533,I3035,I477397,I477383,);
nor I_27911 (I477564,I168753,I168759);
nand I_27912 (I477581,I477564,I168771);
DFFARX1 I_27913 (I477581,I3035,I477397,I477386,);
nor I_27914 (I477612,I477499,I168753);
nand I_27915 (I477629,I477612,I168744);
nor I_27916 (I477646,I477423,I477629);
DFFARX1 I_27917 (I477646,I3035,I477397,I477362,);
not I_27918 (I477677,I477629);
nand I_27919 (I477374,I477440,I477677);
DFFARX1 I_27920 (I477629,I3035,I477397,I477717,);
not I_27921 (I477725,I477717);
not I_27922 (I477742,I168753);
not I_27923 (I477759,I168756);
nor I_27924 (I477776,I477759,I168768);
nor I_27925 (I477389,I477725,I477776);
nor I_27926 (I477807,I477759,I168765);
and I_27927 (I477824,I477807,I168747);
or I_27928 (I477841,I477824,I168762);
DFFARX1 I_27929 (I477841,I3035,I477397,I477867,);
nor I_27930 (I477377,I477867,I477423);
not I_27931 (I477889,I477867);
and I_27932 (I477906,I477889,I477423);
nor I_27933 (I477371,I477448,I477906);
nand I_27934 (I477937,I477889,I477499);
nor I_27935 (I477365,I477759,I477937);
nand I_27936 (I477368,I477889,I477677);
nand I_27937 (I477982,I477499,I168756);
nor I_27938 (I477380,I477742,I477982);
not I_27939 (I478043,I3042);
DFFARX1 I_27940 (I10967,I3035,I478043,I478069,);
DFFARX1 I_27941 (I10973,I3035,I478043,I478086,);
not I_27942 (I478094,I478086);
not I_27943 (I478111,I10967);
nor I_27944 (I478128,I478111,I10979);
not I_27945 (I478145,I10991);
nor I_27946 (I478162,I478128,I10985);
nor I_27947 (I478179,I478086,I478162);
DFFARX1 I_27948 (I478179,I3035,I478043,I478029,);
nor I_27949 (I478210,I10985,I10979);
nand I_27950 (I478227,I478210,I10967);
DFFARX1 I_27951 (I478227,I3035,I478043,I478032,);
nor I_27952 (I478258,I478145,I10985);
nand I_27953 (I478275,I478258,I10970);
nor I_27954 (I478292,I478069,I478275);
DFFARX1 I_27955 (I478292,I3035,I478043,I478008,);
not I_27956 (I478323,I478275);
nand I_27957 (I478020,I478086,I478323);
DFFARX1 I_27958 (I478275,I3035,I478043,I478363,);
not I_27959 (I478371,I478363);
not I_27960 (I478388,I10985);
not I_27961 (I478405,I10970);
nor I_27962 (I478422,I478405,I10991);
nor I_27963 (I478035,I478371,I478422);
nor I_27964 (I478453,I478405,I10988);
and I_27965 (I478470,I478453,I10982);
or I_27966 (I478487,I478470,I10976);
DFFARX1 I_27967 (I478487,I3035,I478043,I478513,);
nor I_27968 (I478023,I478513,I478069);
not I_27969 (I478535,I478513);
and I_27970 (I478552,I478535,I478069);
nor I_27971 (I478017,I478094,I478552);
nand I_27972 (I478583,I478535,I478145);
nor I_27973 (I478011,I478405,I478583);
nand I_27974 (I478014,I478535,I478323);
nand I_27975 (I478628,I478145,I10970);
nor I_27976 (I478026,I478388,I478628);
not I_27977 (I478689,I3042);
DFFARX1 I_27978 (I32047,I3035,I478689,I478715,);
DFFARX1 I_27979 (I32053,I3035,I478689,I478732,);
not I_27980 (I478740,I478732);
not I_27981 (I478757,I32071);
nor I_27982 (I478774,I478757,I32050);
not I_27983 (I478791,I32056);
nor I_27984 (I478808,I478774,I32062);
nor I_27985 (I478825,I478732,I478808);
DFFARX1 I_27986 (I478825,I3035,I478689,I478675,);
nor I_27987 (I478856,I32062,I32050);
nand I_27988 (I478873,I478856,I32071);
DFFARX1 I_27989 (I478873,I3035,I478689,I478678,);
nor I_27990 (I478904,I478791,I32062);
nand I_27991 (I478921,I478904,I32068);
nor I_27992 (I478938,I478715,I478921);
DFFARX1 I_27993 (I478938,I3035,I478689,I478654,);
not I_27994 (I478969,I478921);
nand I_27995 (I478666,I478732,I478969);
DFFARX1 I_27996 (I478921,I3035,I478689,I479009,);
not I_27997 (I479017,I479009);
not I_27998 (I479034,I32062);
not I_27999 (I479051,I32050);
nor I_28000 (I479068,I479051,I32056);
nor I_28001 (I478681,I479017,I479068);
nor I_28002 (I479099,I479051,I32059);
and I_28003 (I479116,I479099,I32047);
or I_28004 (I479133,I479116,I32065);
DFFARX1 I_28005 (I479133,I3035,I478689,I479159,);
nor I_28006 (I478669,I479159,I478715);
not I_28007 (I479181,I479159);
and I_28008 (I479198,I479181,I478715);
nor I_28009 (I478663,I478740,I479198);
nand I_28010 (I479229,I479181,I478791);
nor I_28011 (I478657,I479051,I479229);
nand I_28012 (I478660,I479181,I478969);
nand I_28013 (I479274,I478791,I32050);
nor I_28014 (I478672,I479034,I479274);
not I_28015 (I479335,I3042);
DFFARX1 I_28016 (I186135,I3035,I479335,I479361,);
DFFARX1 I_28017 (I186141,I3035,I479335,I479378,);
not I_28018 (I479386,I479378);
not I_28019 (I479403,I186162);
nor I_28020 (I479420,I479403,I186150);
not I_28021 (I479437,I186159);
nor I_28022 (I479454,I479420,I186144);
nor I_28023 (I479471,I479378,I479454);
DFFARX1 I_28024 (I479471,I3035,I479335,I479321,);
nor I_28025 (I479502,I186144,I186150);
nand I_28026 (I479519,I479502,I186162);
DFFARX1 I_28027 (I479519,I3035,I479335,I479324,);
nor I_28028 (I479550,I479437,I186144);
nand I_28029 (I479567,I479550,I186135);
nor I_28030 (I479584,I479361,I479567);
DFFARX1 I_28031 (I479584,I3035,I479335,I479300,);
not I_28032 (I479615,I479567);
nand I_28033 (I479312,I479378,I479615);
DFFARX1 I_28034 (I479567,I3035,I479335,I479655,);
not I_28035 (I479663,I479655);
not I_28036 (I479680,I186144);
not I_28037 (I479697,I186147);
nor I_28038 (I479714,I479697,I186159);
nor I_28039 (I479327,I479663,I479714);
nor I_28040 (I479745,I479697,I186156);
and I_28041 (I479762,I479745,I186138);
or I_28042 (I479779,I479762,I186153);
DFFARX1 I_28043 (I479779,I3035,I479335,I479805,);
nor I_28044 (I479315,I479805,I479361);
not I_28045 (I479827,I479805);
and I_28046 (I479844,I479827,I479361);
nor I_28047 (I479309,I479386,I479844);
nand I_28048 (I479875,I479827,I479437);
nor I_28049 (I479303,I479697,I479875);
nand I_28050 (I479306,I479827,I479615);
nand I_28051 (I479920,I479437,I186147);
nor I_28052 (I479318,I479680,I479920);
not I_28053 (I479981,I3042);
DFFARX1 I_28054 (I77727,I3035,I479981,I480007,);
DFFARX1 I_28055 (I77730,I3035,I479981,I480024,);
not I_28056 (I480032,I480024);
not I_28057 (I480049,I77715);
nor I_28058 (I480066,I480049,I77709);
not I_28059 (I480083,I77718);
nor I_28060 (I480100,I480066,I77733);
nor I_28061 (I480117,I480024,I480100);
DFFARX1 I_28062 (I480117,I3035,I479981,I479967,);
nor I_28063 (I480148,I77733,I77709);
nand I_28064 (I480165,I480148,I77715);
DFFARX1 I_28065 (I480165,I3035,I479981,I479970,);
nor I_28066 (I480196,I480083,I77733);
nand I_28067 (I480213,I480196,I77736);
nor I_28068 (I480230,I480007,I480213);
DFFARX1 I_28069 (I480230,I3035,I479981,I479946,);
not I_28070 (I480261,I480213);
nand I_28071 (I479958,I480024,I480261);
DFFARX1 I_28072 (I480213,I3035,I479981,I480301,);
not I_28073 (I480309,I480301);
not I_28074 (I480326,I77733);
not I_28075 (I480343,I77712);
nor I_28076 (I480360,I480343,I77718);
nor I_28077 (I479973,I480309,I480360);
nor I_28078 (I480391,I480343,I77721);
and I_28079 (I480408,I480391,I77709);
or I_28080 (I480425,I480408,I77724);
DFFARX1 I_28081 (I480425,I3035,I479981,I480451,);
nor I_28082 (I479961,I480451,I480007);
not I_28083 (I480473,I480451);
and I_28084 (I480490,I480473,I480007);
nor I_28085 (I479955,I480032,I480490);
nand I_28086 (I480521,I480473,I480083);
nor I_28087 (I479949,I480343,I480521);
nand I_28088 (I479952,I480473,I480261);
nand I_28089 (I480566,I480083,I77712);
nor I_28090 (I479964,I480326,I480566);
not I_28091 (I480627,I3042);
DFFARX1 I_28092 (I214066,I3035,I480627,I480653,);
DFFARX1 I_28093 (I214072,I3035,I480627,I480670,);
not I_28094 (I480678,I480670);
not I_28095 (I480695,I214093);
nor I_28096 (I480712,I480695,I214081);
not I_28097 (I480729,I214090);
nor I_28098 (I480746,I480712,I214075);
nor I_28099 (I480763,I480670,I480746);
DFFARX1 I_28100 (I480763,I3035,I480627,I480613,);
nor I_28101 (I480794,I214075,I214081);
nand I_28102 (I480811,I480794,I214093);
DFFARX1 I_28103 (I480811,I3035,I480627,I480616,);
nor I_28104 (I480842,I480729,I214075);
nand I_28105 (I480859,I480842,I214066);
nor I_28106 (I480876,I480653,I480859);
DFFARX1 I_28107 (I480876,I3035,I480627,I480592,);
not I_28108 (I480907,I480859);
nand I_28109 (I480604,I480670,I480907);
DFFARX1 I_28110 (I480859,I3035,I480627,I480947,);
not I_28111 (I480955,I480947);
not I_28112 (I480972,I214075);
not I_28113 (I480989,I214078);
nor I_28114 (I481006,I480989,I214090);
nor I_28115 (I480619,I480955,I481006);
nor I_28116 (I481037,I480989,I214087);
and I_28117 (I481054,I481037,I214069);
or I_28118 (I481071,I481054,I214084);
DFFARX1 I_28119 (I481071,I3035,I480627,I481097,);
nor I_28120 (I480607,I481097,I480653);
not I_28121 (I481119,I481097);
and I_28122 (I481136,I481119,I480653);
nor I_28123 (I480601,I480678,I481136);
nand I_28124 (I481167,I481119,I480729);
nor I_28125 (I480595,I480989,I481167);
nand I_28126 (I480598,I481119,I480907);
nand I_28127 (I481212,I480729,I214078);
nor I_28128 (I480610,I480972,I481212);
not I_28129 (I481273,I3042);
DFFARX1 I_28130 (I285894,I3035,I481273,I481299,);
DFFARX1 I_28131 (I285906,I3035,I481273,I481316,);
not I_28132 (I481324,I481316);
not I_28133 (I481341,I285891);
nor I_28134 (I481358,I481341,I285909);
not I_28135 (I481375,I285915);
nor I_28136 (I481392,I481358,I285897);
nor I_28137 (I481409,I481316,I481392);
DFFARX1 I_28138 (I481409,I3035,I481273,I481259,);
nor I_28139 (I481440,I285897,I285909);
nand I_28140 (I481457,I481440,I285891);
DFFARX1 I_28141 (I481457,I3035,I481273,I481262,);
nor I_28142 (I481488,I481375,I285897);
nand I_28143 (I481505,I481488,I285900);
nor I_28144 (I481522,I481299,I481505);
DFFARX1 I_28145 (I481522,I3035,I481273,I481238,);
not I_28146 (I481553,I481505);
nand I_28147 (I481250,I481316,I481553);
DFFARX1 I_28148 (I481505,I3035,I481273,I481593,);
not I_28149 (I481601,I481593);
not I_28150 (I481618,I285897);
not I_28151 (I481635,I285903);
nor I_28152 (I481652,I481635,I285915);
nor I_28153 (I481265,I481601,I481652);
nor I_28154 (I481683,I481635,I285912);
and I_28155 (I481700,I481683,I285891);
or I_28156 (I481717,I481700,I285894);
DFFARX1 I_28157 (I481717,I3035,I481273,I481743,);
nor I_28158 (I481253,I481743,I481299);
not I_28159 (I481765,I481743);
and I_28160 (I481782,I481765,I481299);
nor I_28161 (I481247,I481324,I481782);
nand I_28162 (I481813,I481765,I481375);
nor I_28163 (I481241,I481635,I481813);
nand I_28164 (I481244,I481765,I481553);
nand I_28165 (I481858,I481375,I285903);
nor I_28166 (I481256,I481618,I481858);
not I_28167 (I481919,I3042);
DFFARX1 I_28168 (I246219,I3035,I481919,I481945,);
DFFARX1 I_28169 (I246216,I3035,I481919,I481962,);
not I_28170 (I481970,I481962);
not I_28171 (I481987,I246231);
nor I_28172 (I482004,I481987,I246234);
not I_28173 (I482021,I246222);
nor I_28174 (I482038,I482004,I246228);
nor I_28175 (I482055,I481962,I482038);
DFFARX1 I_28176 (I482055,I3035,I481919,I481905,);
nor I_28177 (I482086,I246228,I246234);
nand I_28178 (I482103,I482086,I246231);
DFFARX1 I_28179 (I482103,I3035,I481919,I481908,);
nor I_28180 (I482134,I482021,I246228);
nand I_28181 (I482151,I482134,I246240);
nor I_28182 (I482168,I481945,I482151);
DFFARX1 I_28183 (I482168,I3035,I481919,I481884,);
not I_28184 (I482199,I482151);
nand I_28185 (I481896,I481962,I482199);
DFFARX1 I_28186 (I482151,I3035,I481919,I482239,);
not I_28187 (I482247,I482239);
not I_28188 (I482264,I246228);
not I_28189 (I482281,I246213);
nor I_28190 (I482298,I482281,I246222);
nor I_28191 (I481911,I482247,I482298);
nor I_28192 (I482329,I482281,I246225);
and I_28193 (I482346,I482329,I246213);
or I_28194 (I482363,I482346,I246237);
DFFARX1 I_28195 (I482363,I3035,I481919,I482389,);
nor I_28196 (I481899,I482389,I481945);
not I_28197 (I482411,I482389);
and I_28198 (I482428,I482411,I481945);
nor I_28199 (I481893,I481970,I482428);
nand I_28200 (I482459,I482411,I482021);
nor I_28201 (I481887,I482281,I482459);
nand I_28202 (I481890,I482411,I482199);
nand I_28203 (I482504,I482021,I246213);
nor I_28204 (I481902,I482264,I482504);
not I_28205 (I482565,I3042);
DFFARX1 I_28206 (I554338,I3035,I482565,I482591,);
DFFARX1 I_28207 (I554341,I3035,I482565,I482608,);
not I_28208 (I482616,I482608);
not I_28209 (I482633,I554338);
nor I_28210 (I482650,I482633,I554350);
not I_28211 (I482667,I554359);
nor I_28212 (I482684,I482650,I554347);
nor I_28213 (I482701,I482608,I482684);
DFFARX1 I_28214 (I482701,I3035,I482565,I482551,);
nor I_28215 (I482732,I554347,I554350);
nand I_28216 (I482749,I482732,I554338);
DFFARX1 I_28217 (I482749,I3035,I482565,I482554,);
nor I_28218 (I482780,I482667,I554347);
nand I_28219 (I482797,I482780,I554353);
nor I_28220 (I482814,I482591,I482797);
DFFARX1 I_28221 (I482814,I3035,I482565,I482530,);
not I_28222 (I482845,I482797);
nand I_28223 (I482542,I482608,I482845);
DFFARX1 I_28224 (I482797,I3035,I482565,I482885,);
not I_28225 (I482893,I482885);
not I_28226 (I482910,I554347);
not I_28227 (I482927,I554344);
nor I_28228 (I482944,I482927,I554359);
nor I_28229 (I482557,I482893,I482944);
nor I_28230 (I482975,I482927,I554356);
and I_28231 (I482992,I482975,I554344);
or I_28232 (I483009,I482992,I554341);
DFFARX1 I_28233 (I483009,I3035,I482565,I483035,);
nor I_28234 (I482545,I483035,I482591);
not I_28235 (I483057,I483035);
and I_28236 (I483074,I483057,I482591);
nor I_28237 (I482539,I482616,I483074);
nand I_28238 (I483105,I483057,I482667);
nor I_28239 (I482533,I482927,I483105);
nand I_28240 (I482536,I483057,I482845);
nand I_28241 (I483150,I482667,I554344);
nor I_28242 (I482548,I482910,I483150);
not I_28243 (I483211,I3042);
DFFARX1 I_28244 (I309405,I3035,I483211,I483237,);
DFFARX1 I_28245 (I309417,I3035,I483211,I483254,);
not I_28246 (I483262,I483254);
not I_28247 (I483279,I309426);
nor I_28248 (I483296,I483279,I309402);
not I_28249 (I483313,I309420);
nor I_28250 (I483330,I483296,I309414);
nor I_28251 (I483347,I483254,I483330);
DFFARX1 I_28252 (I483347,I3035,I483211,I483197,);
nor I_28253 (I483378,I309414,I309402);
nand I_28254 (I483395,I483378,I309426);
DFFARX1 I_28255 (I483395,I3035,I483211,I483200,);
nor I_28256 (I483426,I483313,I309414);
nand I_28257 (I483443,I483426,I309408);
nor I_28258 (I483460,I483237,I483443);
DFFARX1 I_28259 (I483460,I3035,I483211,I483176,);
not I_28260 (I483491,I483443);
nand I_28261 (I483188,I483254,I483491);
DFFARX1 I_28262 (I483443,I3035,I483211,I483531,);
not I_28263 (I483539,I483531);
not I_28264 (I483556,I309414);
not I_28265 (I483573,I309423);
nor I_28266 (I483590,I483573,I309420);
nor I_28267 (I483203,I483539,I483590);
nor I_28268 (I483621,I483573,I309405);
and I_28269 (I483638,I483621,I309402);
or I_28270 (I483655,I483638,I309411);
DFFARX1 I_28271 (I483655,I3035,I483211,I483681,);
nor I_28272 (I483191,I483681,I483237);
not I_28273 (I483703,I483681);
and I_28274 (I483720,I483703,I483237);
nor I_28275 (I483185,I483262,I483720);
nand I_28276 (I483751,I483703,I483313);
nor I_28277 (I483179,I483573,I483751);
nand I_28278 (I483182,I483703,I483491);
nand I_28279 (I483796,I483313,I309423);
nor I_28280 (I483194,I483556,I483796);
not I_28281 (I483857,I3042);
DFFARX1 I_28282 (I159785,I3035,I483857,I483883,);
DFFARX1 I_28283 (I159791,I3035,I483857,I483900,);
not I_28284 (I483908,I483900);
not I_28285 (I483925,I159812);
nor I_28286 (I483942,I483925,I159800);
not I_28287 (I483959,I159809);
nor I_28288 (I483976,I483942,I159794);
nor I_28289 (I483993,I483900,I483976);
DFFARX1 I_28290 (I483993,I3035,I483857,I483843,);
nor I_28291 (I484024,I159794,I159800);
nand I_28292 (I484041,I484024,I159812);
DFFARX1 I_28293 (I484041,I3035,I483857,I483846,);
nor I_28294 (I484072,I483959,I159794);
nand I_28295 (I484089,I484072,I159785);
nor I_28296 (I484106,I483883,I484089);
DFFARX1 I_28297 (I484106,I3035,I483857,I483822,);
not I_28298 (I484137,I484089);
nand I_28299 (I483834,I483900,I484137);
DFFARX1 I_28300 (I484089,I3035,I483857,I484177,);
not I_28301 (I484185,I484177);
not I_28302 (I484202,I159794);
not I_28303 (I484219,I159797);
nor I_28304 (I484236,I484219,I159809);
nor I_28305 (I483849,I484185,I484236);
nor I_28306 (I484267,I484219,I159806);
and I_28307 (I484284,I484267,I159788);
or I_28308 (I484301,I484284,I159803);
DFFARX1 I_28309 (I484301,I3035,I483857,I484327,);
nor I_28310 (I483837,I484327,I483883);
not I_28311 (I484349,I484327);
and I_28312 (I484366,I484349,I483883);
nor I_28313 (I483831,I483908,I484366);
nand I_28314 (I484397,I484349,I483959);
nor I_28315 (I483825,I484219,I484397);
nand I_28316 (I483828,I484349,I484137);
nand I_28317 (I484442,I483959,I159797);
nor I_28318 (I483840,I484202,I484442);
not I_28319 (I484503,I3042);
DFFARX1 I_28320 (I51019,I3035,I484503,I484529,);
DFFARX1 I_28321 (I51025,I3035,I484503,I484546,);
not I_28322 (I484554,I484546);
not I_28323 (I484571,I51043);
nor I_28324 (I484588,I484571,I51022);
not I_28325 (I484605,I51028);
nor I_28326 (I484622,I484588,I51034);
nor I_28327 (I484639,I484546,I484622);
DFFARX1 I_28328 (I484639,I3035,I484503,I484489,);
nor I_28329 (I484670,I51034,I51022);
nand I_28330 (I484687,I484670,I51043);
DFFARX1 I_28331 (I484687,I3035,I484503,I484492,);
nor I_28332 (I484718,I484605,I51034);
nand I_28333 (I484735,I484718,I51040);
nor I_28334 (I484752,I484529,I484735);
DFFARX1 I_28335 (I484752,I3035,I484503,I484468,);
not I_28336 (I484783,I484735);
nand I_28337 (I484480,I484546,I484783);
DFFARX1 I_28338 (I484735,I3035,I484503,I484823,);
not I_28339 (I484831,I484823);
not I_28340 (I484848,I51034);
not I_28341 (I484865,I51022);
nor I_28342 (I484882,I484865,I51028);
nor I_28343 (I484495,I484831,I484882);
nor I_28344 (I484913,I484865,I51031);
and I_28345 (I484930,I484913,I51019);
or I_28346 (I484947,I484930,I51037);
DFFARX1 I_28347 (I484947,I3035,I484503,I484973,);
nor I_28348 (I484483,I484973,I484529);
not I_28349 (I484995,I484973);
and I_28350 (I485012,I484995,I484529);
nor I_28351 (I484477,I484554,I485012);
nand I_28352 (I485043,I484995,I484605);
nor I_28353 (I484471,I484865,I485043);
nand I_28354 (I484474,I484995,I484783);
nand I_28355 (I485088,I484605,I51022);
nor I_28356 (I484486,I484848,I485088);
not I_28357 (I485149,I3042);
DFFARX1 I_28358 (I206688,I3035,I485149,I485175,);
DFFARX1 I_28359 (I206694,I3035,I485149,I485192,);
not I_28360 (I485200,I485192);
not I_28361 (I485217,I206715);
nor I_28362 (I485234,I485217,I206703);
not I_28363 (I485251,I206712);
nor I_28364 (I485268,I485234,I206697);
nor I_28365 (I485285,I485192,I485268);
DFFARX1 I_28366 (I485285,I3035,I485149,I485135,);
nor I_28367 (I485316,I206697,I206703);
nand I_28368 (I485333,I485316,I206715);
DFFARX1 I_28369 (I485333,I3035,I485149,I485138,);
nor I_28370 (I485364,I485251,I206697);
nand I_28371 (I485381,I485364,I206688);
nor I_28372 (I485398,I485175,I485381);
DFFARX1 I_28373 (I485398,I3035,I485149,I485114,);
not I_28374 (I485429,I485381);
nand I_28375 (I485126,I485192,I485429);
DFFARX1 I_28376 (I485381,I3035,I485149,I485469,);
not I_28377 (I485477,I485469);
not I_28378 (I485494,I206697);
not I_28379 (I485511,I206700);
nor I_28380 (I485528,I485511,I206712);
nor I_28381 (I485141,I485477,I485528);
nor I_28382 (I485559,I485511,I206709);
and I_28383 (I485576,I485559,I206691);
or I_28384 (I485593,I485576,I206706);
DFFARX1 I_28385 (I485593,I3035,I485149,I485619,);
nor I_28386 (I485129,I485619,I485175);
not I_28387 (I485641,I485619);
and I_28388 (I485658,I485641,I485175);
nor I_28389 (I485123,I485200,I485658);
nand I_28390 (I485689,I485641,I485251);
nor I_28391 (I485117,I485511,I485689);
nand I_28392 (I485120,I485641,I485429);
nand I_28393 (I485734,I485251,I206700);
nor I_28394 (I485132,I485494,I485734);
not I_28395 (I485795,I3042);
DFFARX1 I_28396 (I549850,I3035,I485795,I485821,);
DFFARX1 I_28397 (I549853,I3035,I485795,I485838,);
not I_28398 (I485846,I485838);
not I_28399 (I485863,I549850);
nor I_28400 (I485880,I485863,I549862);
not I_28401 (I485897,I549871);
nor I_28402 (I485914,I485880,I549859);
nor I_28403 (I485931,I485838,I485914);
DFFARX1 I_28404 (I485931,I3035,I485795,I485781,);
nor I_28405 (I485962,I549859,I549862);
nand I_28406 (I485979,I485962,I549850);
DFFARX1 I_28407 (I485979,I3035,I485795,I485784,);
nor I_28408 (I486010,I485897,I549859);
nand I_28409 (I486027,I486010,I549865);
nor I_28410 (I486044,I485821,I486027);
DFFARX1 I_28411 (I486044,I3035,I485795,I485760,);
not I_28412 (I486075,I486027);
nand I_28413 (I485772,I485838,I486075);
DFFARX1 I_28414 (I486027,I3035,I485795,I486115,);
not I_28415 (I486123,I486115);
not I_28416 (I486140,I549859);
not I_28417 (I486157,I549856);
nor I_28418 (I486174,I486157,I549871);
nor I_28419 (I485787,I486123,I486174);
nor I_28420 (I486205,I486157,I549868);
and I_28421 (I486222,I486205,I549856);
or I_28422 (I486239,I486222,I549853);
DFFARX1 I_28423 (I486239,I3035,I485795,I486265,);
nor I_28424 (I485775,I486265,I485821);
not I_28425 (I486287,I486265);
and I_28426 (I486304,I486287,I485821);
nor I_28427 (I485769,I485846,I486304);
nand I_28428 (I486335,I486287,I485897);
nor I_28429 (I485763,I486157,I486335);
nand I_28430 (I485766,I486287,I486075);
nand I_28431 (I486380,I485897,I549856);
nor I_28432 (I485778,I486140,I486380);
not I_28433 (I486441,I3042);
DFFARX1 I_28434 (I548728,I3035,I486441,I486467,);
DFFARX1 I_28435 (I548731,I3035,I486441,I486484,);
not I_28436 (I486492,I486484);
not I_28437 (I486509,I548728);
nor I_28438 (I486526,I486509,I548740);
not I_28439 (I486543,I548749);
nor I_28440 (I486560,I486526,I548737);
nor I_28441 (I486577,I486484,I486560);
DFFARX1 I_28442 (I486577,I3035,I486441,I486427,);
nor I_28443 (I486608,I548737,I548740);
nand I_28444 (I486625,I486608,I548728);
DFFARX1 I_28445 (I486625,I3035,I486441,I486430,);
nor I_28446 (I486656,I486543,I548737);
nand I_28447 (I486673,I486656,I548743);
nor I_28448 (I486690,I486467,I486673);
DFFARX1 I_28449 (I486690,I3035,I486441,I486406,);
not I_28450 (I486721,I486673);
nand I_28451 (I486418,I486484,I486721);
DFFARX1 I_28452 (I486673,I3035,I486441,I486761,);
not I_28453 (I486769,I486761);
not I_28454 (I486786,I548737);
not I_28455 (I486803,I548734);
nor I_28456 (I486820,I486803,I548749);
nor I_28457 (I486433,I486769,I486820);
nor I_28458 (I486851,I486803,I548746);
and I_28459 (I486868,I486851,I548734);
or I_28460 (I486885,I486868,I548731);
DFFARX1 I_28461 (I486885,I3035,I486441,I486911,);
nor I_28462 (I486421,I486911,I486467);
not I_28463 (I486933,I486911);
and I_28464 (I486950,I486933,I486467);
nor I_28465 (I486415,I486492,I486950);
nand I_28466 (I486981,I486933,I486543);
nor I_28467 (I486409,I486803,I486981);
nand I_28468 (I486412,I486933,I486721);
nand I_28469 (I487026,I486543,I548734);
nor I_28470 (I486424,I486786,I487026);
not I_28471 (I487087,I3042);
DFFARX1 I_28472 (I412292,I3035,I487087,I487113,);
DFFARX1 I_28473 (I412286,I3035,I487087,I487130,);
not I_28474 (I487138,I487130);
not I_28475 (I487155,I412301);
nor I_28476 (I487172,I487155,I412286);
not I_28477 (I487189,I412295);
nor I_28478 (I487206,I487172,I412304);
nor I_28479 (I487223,I487130,I487206);
DFFARX1 I_28480 (I487223,I3035,I487087,I487073,);
nor I_28481 (I487254,I412304,I412286);
nand I_28482 (I487271,I487254,I412301);
DFFARX1 I_28483 (I487271,I3035,I487087,I487076,);
nor I_28484 (I487302,I487189,I412304);
nand I_28485 (I487319,I487302,I412289);
nor I_28486 (I487336,I487113,I487319);
DFFARX1 I_28487 (I487336,I3035,I487087,I487052,);
not I_28488 (I487367,I487319);
nand I_28489 (I487064,I487130,I487367);
DFFARX1 I_28490 (I487319,I3035,I487087,I487407,);
not I_28491 (I487415,I487407);
not I_28492 (I487432,I412304);
not I_28493 (I487449,I412298);
nor I_28494 (I487466,I487449,I412295);
nor I_28495 (I487079,I487415,I487466);
nor I_28496 (I487497,I487449,I412307);
and I_28497 (I487514,I487497,I412310);
or I_28498 (I487531,I487514,I412289);
DFFARX1 I_28499 (I487531,I3035,I487087,I487557,);
nor I_28500 (I487067,I487557,I487113);
not I_28501 (I487579,I487557);
and I_28502 (I487596,I487579,I487113);
nor I_28503 (I487061,I487138,I487596);
nand I_28504 (I487627,I487579,I487189);
nor I_28505 (I487055,I487449,I487627);
nand I_28506 (I487058,I487579,I487367);
nand I_28507 (I487672,I487189,I412298);
nor I_28508 (I487070,I487432,I487672);
not I_28509 (I487733,I3042);
DFFARX1 I_28510 (I220390,I3035,I487733,I487759,);
DFFARX1 I_28511 (I220396,I3035,I487733,I487776,);
not I_28512 (I487784,I487776);
not I_28513 (I487801,I220417);
nor I_28514 (I487818,I487801,I220405);
not I_28515 (I487835,I220414);
nor I_28516 (I487852,I487818,I220399);
nor I_28517 (I487869,I487776,I487852);
DFFARX1 I_28518 (I487869,I3035,I487733,I487719,);
nor I_28519 (I487900,I220399,I220405);
nand I_28520 (I487917,I487900,I220417);
DFFARX1 I_28521 (I487917,I3035,I487733,I487722,);
nor I_28522 (I487948,I487835,I220399);
nand I_28523 (I487965,I487948,I220390);
nor I_28524 (I487982,I487759,I487965);
DFFARX1 I_28525 (I487982,I3035,I487733,I487698,);
not I_28526 (I488013,I487965);
nand I_28527 (I487710,I487776,I488013);
DFFARX1 I_28528 (I487965,I3035,I487733,I488053,);
not I_28529 (I488061,I488053);
not I_28530 (I488078,I220399);
not I_28531 (I488095,I220402);
nor I_28532 (I488112,I488095,I220414);
nor I_28533 (I487725,I488061,I488112);
nor I_28534 (I488143,I488095,I220411);
and I_28535 (I488160,I488143,I220393);
or I_28536 (I488177,I488160,I220408);
DFFARX1 I_28537 (I488177,I3035,I487733,I488203,);
nor I_28538 (I487713,I488203,I487759);
not I_28539 (I488225,I488203);
and I_28540 (I488242,I488225,I487759);
nor I_28541 (I487707,I487784,I488242);
nand I_28542 (I488273,I488225,I487835);
nor I_28543 (I487701,I488095,I488273);
nand I_28544 (I487704,I488225,I488013);
nand I_28545 (I488318,I487835,I220402);
nor I_28546 (I487716,I488078,I488318);
not I_28547 (I488379,I3042);
DFFARX1 I_28548 (I309983,I3035,I488379,I488405,);
DFFARX1 I_28549 (I309995,I3035,I488379,I488422,);
not I_28550 (I488430,I488422);
not I_28551 (I488447,I310004);
nor I_28552 (I488464,I488447,I309980);
not I_28553 (I488481,I309998);
nor I_28554 (I488498,I488464,I309992);
nor I_28555 (I488515,I488422,I488498);
DFFARX1 I_28556 (I488515,I3035,I488379,I488365,);
nor I_28557 (I488546,I309992,I309980);
nand I_28558 (I488563,I488546,I310004);
DFFARX1 I_28559 (I488563,I3035,I488379,I488368,);
nor I_28560 (I488594,I488481,I309992);
nand I_28561 (I488611,I488594,I309986);
nor I_28562 (I488628,I488405,I488611);
DFFARX1 I_28563 (I488628,I3035,I488379,I488344,);
not I_28564 (I488659,I488611);
nand I_28565 (I488356,I488422,I488659);
DFFARX1 I_28566 (I488611,I3035,I488379,I488699,);
not I_28567 (I488707,I488699);
not I_28568 (I488724,I309992);
not I_28569 (I488741,I310001);
nor I_28570 (I488758,I488741,I309998);
nor I_28571 (I488371,I488707,I488758);
nor I_28572 (I488789,I488741,I309983);
and I_28573 (I488806,I488789,I309980);
or I_28574 (I488823,I488806,I309989);
DFFARX1 I_28575 (I488823,I3035,I488379,I488849,);
nor I_28576 (I488359,I488849,I488405);
not I_28577 (I488871,I488849);
and I_28578 (I488888,I488871,I488405);
nor I_28579 (I488353,I488430,I488888);
nand I_28580 (I488919,I488871,I488481);
nor I_28581 (I488347,I488741,I488919);
nand I_28582 (I488350,I488871,I488659);
nand I_28583 (I488964,I488481,I310001);
nor I_28584 (I488362,I488724,I488964);
not I_28585 (I489025,I3042);
DFFARX1 I_28586 (I601786,I3035,I489025,I489051,);
DFFARX1 I_28587 (I601768,I3035,I489025,I489068,);
not I_28588 (I489076,I489068);
not I_28589 (I489093,I601777);
nor I_28590 (I489110,I489093,I601789);
not I_28591 (I489127,I601771);
nor I_28592 (I489144,I489110,I601780);
nor I_28593 (I489161,I489068,I489144);
DFFARX1 I_28594 (I489161,I3035,I489025,I489011,);
nor I_28595 (I489192,I601780,I601789);
nand I_28596 (I489209,I489192,I601777);
DFFARX1 I_28597 (I489209,I3035,I489025,I489014,);
nor I_28598 (I489240,I489127,I601780);
nand I_28599 (I489257,I489240,I601792);
nor I_28600 (I489274,I489051,I489257);
DFFARX1 I_28601 (I489274,I3035,I489025,I488990,);
not I_28602 (I489305,I489257);
nand I_28603 (I489002,I489068,I489305);
DFFARX1 I_28604 (I489257,I3035,I489025,I489345,);
not I_28605 (I489353,I489345);
not I_28606 (I489370,I601780);
not I_28607 (I489387,I601768);
nor I_28608 (I489404,I489387,I601771);
nor I_28609 (I489017,I489353,I489404);
nor I_28610 (I489435,I489387,I601774);
and I_28611 (I489452,I489435,I601783);
or I_28612 (I489469,I489452,I601771);
DFFARX1 I_28613 (I489469,I3035,I489025,I489495,);
nor I_28614 (I489005,I489495,I489051);
not I_28615 (I489517,I489495);
and I_28616 (I489534,I489517,I489051);
nor I_28617 (I488999,I489076,I489534);
nand I_28618 (I489565,I489517,I489127);
nor I_28619 (I488993,I489387,I489565);
nand I_28620 (I488996,I489517,I489305);
nand I_28621 (I489610,I489127,I601768);
nor I_28622 (I489008,I489370,I489610);
not I_28623 (I489671,I3042);
DFFARX1 I_28624 (I601208,I3035,I489671,I489697,);
DFFARX1 I_28625 (I601190,I3035,I489671,I489714,);
not I_28626 (I489722,I489714);
not I_28627 (I489739,I601199);
nor I_28628 (I489756,I489739,I601211);
not I_28629 (I489773,I601193);
nor I_28630 (I489790,I489756,I601202);
nor I_28631 (I489807,I489714,I489790);
DFFARX1 I_28632 (I489807,I3035,I489671,I489657,);
nor I_28633 (I489838,I601202,I601211);
nand I_28634 (I489855,I489838,I601199);
DFFARX1 I_28635 (I489855,I3035,I489671,I489660,);
nor I_28636 (I489886,I489773,I601202);
nand I_28637 (I489903,I489886,I601214);
nor I_28638 (I489920,I489697,I489903);
DFFARX1 I_28639 (I489920,I3035,I489671,I489636,);
not I_28640 (I489951,I489903);
nand I_28641 (I489648,I489714,I489951);
DFFARX1 I_28642 (I489903,I3035,I489671,I489991,);
not I_28643 (I489999,I489991);
not I_28644 (I490016,I601202);
not I_28645 (I490033,I601190);
nor I_28646 (I490050,I490033,I601193);
nor I_28647 (I489663,I489999,I490050);
nor I_28648 (I490081,I490033,I601196);
and I_28649 (I490098,I490081,I601205);
or I_28650 (I490115,I490098,I601193);
DFFARX1 I_28651 (I490115,I3035,I489671,I490141,);
nor I_28652 (I489651,I490141,I489697);
not I_28653 (I490163,I490141);
and I_28654 (I490180,I490163,I489697);
nor I_28655 (I489645,I489722,I490180);
nand I_28656 (I490211,I490163,I489773);
nor I_28657 (I489639,I490033,I490211);
nand I_28658 (I489642,I490163,I489951);
nand I_28659 (I490256,I489773,I601190);
nor I_28660 (I489654,I490016,I490256);
not I_28661 (I490317,I3042);
DFFARX1 I_28662 (I102110,I3035,I490317,I490343,);
DFFARX1 I_28663 (I102122,I3035,I490317,I490360,);
not I_28664 (I490368,I490360);
not I_28665 (I490385,I102128);
nor I_28666 (I490402,I490385,I102113);
not I_28667 (I490419,I102104);
nor I_28668 (I490436,I490402,I102125);
nor I_28669 (I490453,I490360,I490436);
DFFARX1 I_28670 (I490453,I3035,I490317,I490303,);
nor I_28671 (I490484,I102125,I102113);
nand I_28672 (I490501,I490484,I102128);
DFFARX1 I_28673 (I490501,I3035,I490317,I490306,);
nor I_28674 (I490532,I490419,I102125);
nand I_28675 (I490549,I490532,I102107);
nor I_28676 (I490566,I490343,I490549);
DFFARX1 I_28677 (I490566,I3035,I490317,I490282,);
not I_28678 (I490597,I490549);
nand I_28679 (I490294,I490360,I490597);
DFFARX1 I_28680 (I490549,I3035,I490317,I490637,);
not I_28681 (I490645,I490637);
not I_28682 (I490662,I102125);
not I_28683 (I490679,I102116);
nor I_28684 (I490696,I490679,I102104);
nor I_28685 (I490309,I490645,I490696);
nor I_28686 (I490727,I490679,I102119);
and I_28687 (I490744,I490727,I102107);
or I_28688 (I490761,I490744,I102104);
DFFARX1 I_28689 (I490761,I3035,I490317,I490787,);
nor I_28690 (I490297,I490787,I490343);
not I_28691 (I490809,I490787);
and I_28692 (I490826,I490809,I490343);
nor I_28693 (I490291,I490368,I490826);
nand I_28694 (I490857,I490809,I490419);
nor I_28695 (I490285,I490679,I490857);
nand I_28696 (I490288,I490809,I490597);
nand I_28697 (I490902,I490419,I102116);
nor I_28698 (I490300,I490662,I490902);
not I_28699 (I490963,I3042);
DFFARX1 I_28700 (I568924,I3035,I490963,I490989,);
DFFARX1 I_28701 (I568927,I3035,I490963,I491006,);
not I_28702 (I491014,I491006);
not I_28703 (I491031,I568924);
nor I_28704 (I491048,I491031,I568936);
not I_28705 (I491065,I568945);
nor I_28706 (I491082,I491048,I568933);
nor I_28707 (I491099,I491006,I491082);
DFFARX1 I_28708 (I491099,I3035,I490963,I490949,);
nor I_28709 (I491130,I568933,I568936);
nand I_28710 (I491147,I491130,I568924);
DFFARX1 I_28711 (I491147,I3035,I490963,I490952,);
nor I_28712 (I491178,I491065,I568933);
nand I_28713 (I491195,I491178,I568939);
nor I_28714 (I491212,I490989,I491195);
DFFARX1 I_28715 (I491212,I3035,I490963,I490928,);
not I_28716 (I491243,I491195);
nand I_28717 (I490940,I491006,I491243);
DFFARX1 I_28718 (I491195,I3035,I490963,I491283,);
not I_28719 (I491291,I491283);
not I_28720 (I491308,I568933);
not I_28721 (I491325,I568930);
nor I_28722 (I491342,I491325,I568945);
nor I_28723 (I490955,I491291,I491342);
nor I_28724 (I491373,I491325,I568942);
and I_28725 (I491390,I491373,I568930);
or I_28726 (I491407,I491390,I568927);
DFFARX1 I_28727 (I491407,I3035,I490963,I491433,);
nor I_28728 (I490943,I491433,I490989);
not I_28729 (I491455,I491433);
and I_28730 (I491472,I491455,I490989);
nor I_28731 (I490937,I491014,I491472);
nand I_28732 (I491503,I491455,I491065);
nor I_28733 (I490931,I491325,I491503);
nand I_28734 (I490934,I491455,I491243);
nand I_28735 (I491548,I491065,I568930);
nor I_28736 (I490946,I491308,I491548);
not I_28737 (I491609,I3042);
DFFARX1 I_28738 (I240235,I3035,I491609,I491635,);
DFFARX1 I_28739 (I240232,I3035,I491609,I491652,);
not I_28740 (I491660,I491652);
not I_28741 (I491677,I240247);
nor I_28742 (I491694,I491677,I240250);
not I_28743 (I491711,I240238);
nor I_28744 (I491728,I491694,I240244);
nor I_28745 (I491745,I491652,I491728);
DFFARX1 I_28746 (I491745,I3035,I491609,I491595,);
nor I_28747 (I491776,I240244,I240250);
nand I_28748 (I491793,I491776,I240247);
DFFARX1 I_28749 (I491793,I3035,I491609,I491598,);
nor I_28750 (I491824,I491711,I240244);
nand I_28751 (I491841,I491824,I240256);
nor I_28752 (I491858,I491635,I491841);
DFFARX1 I_28753 (I491858,I3035,I491609,I491574,);
not I_28754 (I491889,I491841);
nand I_28755 (I491586,I491652,I491889);
DFFARX1 I_28756 (I491841,I3035,I491609,I491929,);
not I_28757 (I491937,I491929);
not I_28758 (I491954,I240244);
not I_28759 (I491971,I240229);
nor I_28760 (I491988,I491971,I240238);
nor I_28761 (I491601,I491937,I491988);
nor I_28762 (I492019,I491971,I240241);
and I_28763 (I492036,I492019,I240229);
or I_28764 (I492053,I492036,I240253);
DFFARX1 I_28765 (I492053,I3035,I491609,I492079,);
nor I_28766 (I491589,I492079,I491635);
not I_28767 (I492101,I492079);
and I_28768 (I492118,I492101,I491635);
nor I_28769 (I491583,I491660,I492118);
nand I_28770 (I492149,I492101,I491711);
nor I_28771 (I491577,I491971,I492149);
nand I_28772 (I491580,I492101,I491889);
nand I_28773 (I492194,I491711,I240229);
nor I_28774 (I491592,I491954,I492194);
not I_28775 (I492255,I3042);
DFFARX1 I_28776 (I9913,I3035,I492255,I492281,);
DFFARX1 I_28777 (I9919,I3035,I492255,I492298,);
not I_28778 (I492306,I492298);
not I_28779 (I492323,I9913);
nor I_28780 (I492340,I492323,I9925);
not I_28781 (I492357,I9937);
nor I_28782 (I492374,I492340,I9931);
nor I_28783 (I492391,I492298,I492374);
DFFARX1 I_28784 (I492391,I3035,I492255,I492241,);
nor I_28785 (I492422,I9931,I9925);
nand I_28786 (I492439,I492422,I9913);
DFFARX1 I_28787 (I492439,I3035,I492255,I492244,);
nor I_28788 (I492470,I492357,I9931);
nand I_28789 (I492487,I492470,I9916);
nor I_28790 (I492504,I492281,I492487);
DFFARX1 I_28791 (I492504,I3035,I492255,I492220,);
not I_28792 (I492535,I492487);
nand I_28793 (I492232,I492298,I492535);
DFFARX1 I_28794 (I492487,I3035,I492255,I492575,);
not I_28795 (I492583,I492575);
not I_28796 (I492600,I9931);
not I_28797 (I492617,I9916);
nor I_28798 (I492634,I492617,I9937);
nor I_28799 (I492247,I492583,I492634);
nor I_28800 (I492665,I492617,I9934);
and I_28801 (I492682,I492665,I9928);
or I_28802 (I492699,I492682,I9922);
DFFARX1 I_28803 (I492699,I3035,I492255,I492725,);
nor I_28804 (I492235,I492725,I492281);
not I_28805 (I492747,I492725);
and I_28806 (I492764,I492747,I492281);
nor I_28807 (I492229,I492306,I492764);
nand I_28808 (I492795,I492747,I492357);
nor I_28809 (I492223,I492617,I492795);
nand I_28810 (I492226,I492747,I492535);
nand I_28811 (I492840,I492357,I9916);
nor I_28812 (I492238,I492600,I492840);
not I_28813 (I492901,I3042);
DFFARX1 I_28814 (I682901,I3035,I492901,I492927,);
DFFARX1 I_28815 (I682895,I3035,I492901,I492944,);
not I_28816 (I492952,I492944);
not I_28817 (I492969,I682904);
nor I_28818 (I492986,I492969,I682916);
not I_28819 (I493003,I682898);
nor I_28820 (I493020,I492986,I682895);
nor I_28821 (I493037,I492944,I493020);
DFFARX1 I_28822 (I493037,I3035,I492901,I492887,);
nor I_28823 (I493068,I682895,I682916);
nand I_28824 (I493085,I493068,I682904);
DFFARX1 I_28825 (I493085,I3035,I492901,I492890,);
nor I_28826 (I493116,I493003,I682895);
nand I_28827 (I493133,I493116,I682892);
nor I_28828 (I493150,I492927,I493133);
DFFARX1 I_28829 (I493150,I3035,I492901,I492866,);
not I_28830 (I493181,I493133);
nand I_28831 (I492878,I492944,I493181);
DFFARX1 I_28832 (I493133,I3035,I492901,I493221,);
not I_28833 (I493229,I493221);
not I_28834 (I493246,I682895);
not I_28835 (I493263,I682913);
nor I_28836 (I493280,I493263,I682898);
nor I_28837 (I492893,I493229,I493280);
nor I_28838 (I493311,I493263,I682907);
and I_28839 (I493328,I493311,I682892);
or I_28840 (I493345,I493328,I682910);
DFFARX1 I_28841 (I493345,I3035,I492901,I493371,);
nor I_28842 (I492881,I493371,I492927);
not I_28843 (I493393,I493371);
and I_28844 (I493410,I493393,I492927);
nor I_28845 (I492875,I492952,I493410);
nand I_28846 (I493441,I493393,I493003);
nor I_28847 (I492869,I493263,I493441);
nand I_28848 (I492872,I493393,I493181);
nand I_28849 (I493486,I493003,I682913);
nor I_28850 (I492884,I493246,I493486);
not I_28851 (I493547,I3042);
DFFARX1 I_28852 (I430873,I3035,I493547,I493573,);
DFFARX1 I_28853 (I430870,I3035,I493547,I493590,);
not I_28854 (I493598,I493590);
not I_28855 (I493615,I430870);
nor I_28856 (I493632,I493615,I430873);
not I_28857 (I493649,I430885);
nor I_28858 (I493666,I493632,I430879);
nor I_28859 (I493683,I493590,I493666);
DFFARX1 I_28860 (I493683,I3035,I493547,I493533,);
nor I_28861 (I493714,I430879,I430873);
nand I_28862 (I493731,I493714,I430870);
DFFARX1 I_28863 (I493731,I3035,I493547,I493536,);
nor I_28864 (I493762,I493649,I430879);
nand I_28865 (I493779,I493762,I430867);
nor I_28866 (I493796,I493573,I493779);
DFFARX1 I_28867 (I493796,I3035,I493547,I493512,);
not I_28868 (I493827,I493779);
nand I_28869 (I493524,I493590,I493827);
DFFARX1 I_28870 (I493779,I3035,I493547,I493867,);
not I_28871 (I493875,I493867);
not I_28872 (I493892,I430879);
not I_28873 (I493909,I430876);
nor I_28874 (I493926,I493909,I430885);
nor I_28875 (I493539,I493875,I493926);
nor I_28876 (I493957,I493909,I430882);
and I_28877 (I493974,I493957,I430888);
or I_28878 (I493991,I493974,I430867);
DFFARX1 I_28879 (I493991,I3035,I493547,I494017,);
nor I_28880 (I493527,I494017,I493573);
not I_28881 (I494039,I494017);
and I_28882 (I494056,I494039,I493573);
nor I_28883 (I493521,I493598,I494056);
nand I_28884 (I494087,I494039,I493649);
nor I_28885 (I493515,I493909,I494087);
nand I_28886 (I493518,I494039,I493827);
nand I_28887 (I494132,I493649,I430876);
nor I_28888 (I493530,I493892,I494132);
not I_28889 (I494193,I3042);
DFFARX1 I_28890 (I647448,I3035,I494193,I494219,);
DFFARX1 I_28891 (I647454,I3035,I494193,I494236,);
not I_28892 (I494244,I494236);
not I_28893 (I494261,I647451);
nor I_28894 (I494278,I494261,I647430);
not I_28895 (I494295,I647433);
nor I_28896 (I494312,I494278,I647439);
nor I_28897 (I494329,I494236,I494312);
DFFARX1 I_28898 (I494329,I3035,I494193,I494179,);
nor I_28899 (I494360,I647439,I647430);
nand I_28900 (I494377,I494360,I647451);
DFFARX1 I_28901 (I494377,I3035,I494193,I494182,);
nor I_28902 (I494408,I494295,I647439);
nand I_28903 (I494425,I494408,I647433);
nor I_28904 (I494442,I494219,I494425);
DFFARX1 I_28905 (I494442,I3035,I494193,I494158,);
not I_28906 (I494473,I494425);
nand I_28907 (I494170,I494236,I494473);
DFFARX1 I_28908 (I494425,I3035,I494193,I494513,);
not I_28909 (I494521,I494513);
not I_28910 (I494538,I647439);
not I_28911 (I494555,I647442);
nor I_28912 (I494572,I494555,I647433);
nor I_28913 (I494185,I494521,I494572);
nor I_28914 (I494603,I494555,I647430);
and I_28915 (I494620,I494603,I647436);
or I_28916 (I494637,I494620,I647445);
DFFARX1 I_28917 (I494637,I3035,I494193,I494663,);
nor I_28918 (I494173,I494663,I494219);
not I_28919 (I494685,I494663);
and I_28920 (I494702,I494685,I494219);
nor I_28921 (I494167,I494244,I494702);
nand I_28922 (I494733,I494685,I494295);
nor I_28923 (I494161,I494555,I494733);
nand I_28924 (I494164,I494685,I494473);
nand I_28925 (I494778,I494295,I647442);
nor I_28926 (I494176,I494538,I494778);
not I_28927 (I494839,I3042);
DFFARX1 I_28928 (I408824,I3035,I494839,I494865,);
DFFARX1 I_28929 (I408818,I3035,I494839,I494882,);
not I_28930 (I494890,I494882);
not I_28931 (I494907,I408833);
nor I_28932 (I494924,I494907,I408818);
not I_28933 (I494941,I408827);
nor I_28934 (I494958,I494924,I408836);
nor I_28935 (I494975,I494882,I494958);
DFFARX1 I_28936 (I494975,I3035,I494839,I494825,);
nor I_28937 (I495006,I408836,I408818);
nand I_28938 (I495023,I495006,I408833);
DFFARX1 I_28939 (I495023,I3035,I494839,I494828,);
nor I_28940 (I495054,I494941,I408836);
nand I_28941 (I495071,I495054,I408821);
nor I_28942 (I495088,I494865,I495071);
DFFARX1 I_28943 (I495088,I3035,I494839,I494804,);
not I_28944 (I495119,I495071);
nand I_28945 (I494816,I494882,I495119);
DFFARX1 I_28946 (I495071,I3035,I494839,I495159,);
not I_28947 (I495167,I495159);
not I_28948 (I495184,I408836);
not I_28949 (I495201,I408830);
nor I_28950 (I495218,I495201,I408827);
nor I_28951 (I494831,I495167,I495218);
nor I_28952 (I495249,I495201,I408839);
and I_28953 (I495266,I495249,I408842);
or I_28954 (I495283,I495266,I408821);
DFFARX1 I_28955 (I495283,I3035,I494839,I495309,);
nor I_28956 (I494819,I495309,I494865);
not I_28957 (I495331,I495309);
and I_28958 (I495348,I495331,I494865);
nor I_28959 (I494813,I494890,I495348);
nand I_28960 (I495379,I495331,I494941);
nor I_28961 (I494807,I495201,I495379);
nand I_28962 (I494810,I495331,I495119);
nand I_28963 (I495424,I494941,I408830);
nor I_28964 (I494822,I495184,I495424);
not I_28965 (I495485,I3042);
DFFARX1 I_28966 (I250571,I3035,I495485,I495511,);
DFFARX1 I_28967 (I250568,I3035,I495485,I495528,);
not I_28968 (I495536,I495528);
not I_28969 (I495553,I250583);
nor I_28970 (I495570,I495553,I250586);
not I_28971 (I495587,I250574);
nor I_28972 (I495604,I495570,I250580);
nor I_28973 (I495621,I495528,I495604);
DFFARX1 I_28974 (I495621,I3035,I495485,I495471,);
nor I_28975 (I495652,I250580,I250586);
nand I_28976 (I495669,I495652,I250583);
DFFARX1 I_28977 (I495669,I3035,I495485,I495474,);
nor I_28978 (I495700,I495587,I250580);
nand I_28979 (I495717,I495700,I250592);
nor I_28980 (I495734,I495511,I495717);
DFFARX1 I_28981 (I495734,I3035,I495485,I495450,);
not I_28982 (I495765,I495717);
nand I_28983 (I495462,I495528,I495765);
DFFARX1 I_28984 (I495717,I3035,I495485,I495805,);
not I_28985 (I495813,I495805);
not I_28986 (I495830,I250580);
not I_28987 (I495847,I250565);
nor I_28988 (I495864,I495847,I250574);
nor I_28989 (I495477,I495813,I495864);
nor I_28990 (I495895,I495847,I250577);
and I_28991 (I495912,I495895,I250565);
or I_28992 (I495929,I495912,I250589);
DFFARX1 I_28993 (I495929,I3035,I495485,I495955,);
nor I_28994 (I495465,I495955,I495511);
not I_28995 (I495977,I495955);
and I_28996 (I495994,I495977,I495511);
nor I_28997 (I495459,I495536,I495994);
nand I_28998 (I496025,I495977,I495587);
nor I_28999 (I495453,I495847,I496025);
nand I_29000 (I495456,I495977,I495765);
nand I_29001 (I496070,I495587,I250565);
nor I_29002 (I495468,I495830,I496070);
not I_29003 (I496131,I3042);
DFFARX1 I_29004 (I726973,I3035,I496131,I496157,);
DFFARX1 I_29005 (I726997,I3035,I496131,I496174,);
not I_29006 (I496182,I496174);
not I_29007 (I496199,I726979);
nor I_29008 (I496216,I496199,I726988);
not I_29009 (I496233,I726973);
nor I_29010 (I496250,I496216,I726994);
nor I_29011 (I496267,I496174,I496250);
DFFARX1 I_29012 (I496267,I3035,I496131,I496117,);
nor I_29013 (I496298,I726994,I726988);
nand I_29014 (I496315,I496298,I726979);
DFFARX1 I_29015 (I496315,I3035,I496131,I496120,);
nor I_29016 (I496346,I496233,I726994);
nand I_29017 (I496363,I496346,I726991);
nor I_29018 (I496380,I496157,I496363);
DFFARX1 I_29019 (I496380,I3035,I496131,I496096,);
not I_29020 (I496411,I496363);
nand I_29021 (I496108,I496174,I496411);
DFFARX1 I_29022 (I496363,I3035,I496131,I496451,);
not I_29023 (I496459,I496451);
not I_29024 (I496476,I726994);
not I_29025 (I496493,I726985);
nor I_29026 (I496510,I496493,I726973);
nor I_29027 (I496123,I496459,I496510);
nor I_29028 (I496541,I496493,I726976);
and I_29029 (I496558,I496541,I727000);
or I_29030 (I496575,I496558,I726982);
DFFARX1 I_29031 (I496575,I3035,I496131,I496601,);
nor I_29032 (I496111,I496601,I496157);
not I_29033 (I496623,I496601);
and I_29034 (I496640,I496623,I496157);
nor I_29035 (I496105,I496182,I496640);
nand I_29036 (I496671,I496623,I496233);
nor I_29037 (I496099,I496493,I496671);
nand I_29038 (I496102,I496623,I496411);
nand I_29039 (I496716,I496233,I726985);
nor I_29040 (I496114,I496476,I496716);
not I_29041 (I496777,I3042);
DFFARX1 I_29042 (I16237,I3035,I496777,I496803,);
DFFARX1 I_29043 (I16243,I3035,I496777,I496820,);
not I_29044 (I496828,I496820);
not I_29045 (I496845,I16237);
nor I_29046 (I496862,I496845,I16249);
not I_29047 (I496879,I16261);
nor I_29048 (I496896,I496862,I16255);
nor I_29049 (I496913,I496820,I496896);
DFFARX1 I_29050 (I496913,I3035,I496777,I496763,);
nor I_29051 (I496944,I16255,I16249);
nand I_29052 (I496961,I496944,I16237);
DFFARX1 I_29053 (I496961,I3035,I496777,I496766,);
nor I_29054 (I496992,I496879,I16255);
nand I_29055 (I497009,I496992,I16240);
nor I_29056 (I497026,I496803,I497009);
DFFARX1 I_29057 (I497026,I3035,I496777,I496742,);
not I_29058 (I497057,I497009);
nand I_29059 (I496754,I496820,I497057);
DFFARX1 I_29060 (I497009,I3035,I496777,I497097,);
not I_29061 (I497105,I497097);
not I_29062 (I497122,I16255);
not I_29063 (I497139,I16240);
nor I_29064 (I497156,I497139,I16261);
nor I_29065 (I496769,I497105,I497156);
nor I_29066 (I497187,I497139,I16258);
and I_29067 (I497204,I497187,I16252);
or I_29068 (I497221,I497204,I16246);
DFFARX1 I_29069 (I497221,I3035,I496777,I497247,);
nor I_29070 (I496757,I497247,I496803);
not I_29071 (I497269,I497247);
and I_29072 (I497286,I497269,I496803);
nor I_29073 (I496751,I496828,I497286);
nand I_29074 (I497317,I497269,I496879);
nor I_29075 (I496745,I497139,I497317);
nand I_29076 (I496748,I497269,I497057);
nand I_29077 (I497362,I496879,I16240);
nor I_29078 (I496760,I497122,I497362);
not I_29079 (I497423,I3042);
DFFARX1 I_29080 (I251115,I3035,I497423,I497449,);
DFFARX1 I_29081 (I251112,I3035,I497423,I497466,);
not I_29082 (I497474,I497466);
not I_29083 (I497491,I251127);
nor I_29084 (I497508,I497491,I251130);
not I_29085 (I497525,I251118);
nor I_29086 (I497542,I497508,I251124);
nor I_29087 (I497559,I497466,I497542);
DFFARX1 I_29088 (I497559,I3035,I497423,I497409,);
nor I_29089 (I497590,I251124,I251130);
nand I_29090 (I497607,I497590,I251127);
DFFARX1 I_29091 (I497607,I3035,I497423,I497412,);
nor I_29092 (I497638,I497525,I251124);
nand I_29093 (I497655,I497638,I251136);
nor I_29094 (I497672,I497449,I497655);
DFFARX1 I_29095 (I497672,I3035,I497423,I497388,);
not I_29096 (I497703,I497655);
nand I_29097 (I497400,I497466,I497703);
DFFARX1 I_29098 (I497655,I3035,I497423,I497743,);
not I_29099 (I497751,I497743);
not I_29100 (I497768,I251124);
not I_29101 (I497785,I251109);
nor I_29102 (I497802,I497785,I251118);
nor I_29103 (I497415,I497751,I497802);
nor I_29104 (I497833,I497785,I251121);
and I_29105 (I497850,I497833,I251109);
or I_29106 (I497867,I497850,I251133);
DFFARX1 I_29107 (I497867,I3035,I497423,I497893,);
nor I_29108 (I497403,I497893,I497449);
not I_29109 (I497915,I497893);
and I_29110 (I497932,I497915,I497449);
nor I_29111 (I497397,I497474,I497932);
nand I_29112 (I497963,I497915,I497525);
nor I_29113 (I497391,I497785,I497963);
nand I_29114 (I497394,I497915,I497703);
nand I_29115 (I498008,I497525,I251109);
nor I_29116 (I497406,I497768,I498008);
not I_29117 (I498069,I3042);
DFFARX1 I_29118 (I208796,I3035,I498069,I498095,);
DFFARX1 I_29119 (I208802,I3035,I498069,I498112,);
not I_29120 (I498120,I498112);
not I_29121 (I498137,I208823);
nor I_29122 (I498154,I498137,I208811);
not I_29123 (I498171,I208820);
nor I_29124 (I498188,I498154,I208805);
nor I_29125 (I498205,I498112,I498188);
DFFARX1 I_29126 (I498205,I3035,I498069,I498055,);
nor I_29127 (I498236,I208805,I208811);
nand I_29128 (I498253,I498236,I208823);
DFFARX1 I_29129 (I498253,I3035,I498069,I498058,);
nor I_29130 (I498284,I498171,I208805);
nand I_29131 (I498301,I498284,I208796);
nor I_29132 (I498318,I498095,I498301);
DFFARX1 I_29133 (I498318,I3035,I498069,I498034,);
not I_29134 (I498349,I498301);
nand I_29135 (I498046,I498112,I498349);
DFFARX1 I_29136 (I498301,I3035,I498069,I498389,);
not I_29137 (I498397,I498389);
not I_29138 (I498414,I208805);
not I_29139 (I498431,I208808);
nor I_29140 (I498448,I498431,I208820);
nor I_29141 (I498061,I498397,I498448);
nor I_29142 (I498479,I498431,I208817);
and I_29143 (I498496,I498479,I208799);
or I_29144 (I498513,I498496,I208814);
DFFARX1 I_29145 (I498513,I3035,I498069,I498539,);
nor I_29146 (I498049,I498539,I498095);
not I_29147 (I498561,I498539);
and I_29148 (I498578,I498561,I498095);
nor I_29149 (I498043,I498120,I498578);
nand I_29150 (I498609,I498561,I498171);
nor I_29151 (I498037,I498431,I498609);
nand I_29152 (I498040,I498561,I498349);
nand I_29153 (I498654,I498171,I208808);
nor I_29154 (I498052,I498414,I498654);
not I_29155 (I498715,I3042);
DFFARX1 I_29156 (I280539,I3035,I498715,I498741,);
DFFARX1 I_29157 (I280551,I3035,I498715,I498758,);
not I_29158 (I498766,I498758);
not I_29159 (I498783,I280536);
nor I_29160 (I498800,I498783,I280554);
not I_29161 (I498817,I280560);
nor I_29162 (I498834,I498800,I280542);
nor I_29163 (I498851,I498758,I498834);
DFFARX1 I_29164 (I498851,I3035,I498715,I498701,);
nor I_29165 (I498882,I280542,I280554);
nand I_29166 (I498899,I498882,I280536);
DFFARX1 I_29167 (I498899,I3035,I498715,I498704,);
nor I_29168 (I498930,I498817,I280542);
nand I_29169 (I498947,I498930,I280545);
nor I_29170 (I498964,I498741,I498947);
DFFARX1 I_29171 (I498964,I3035,I498715,I498680,);
not I_29172 (I498995,I498947);
nand I_29173 (I498692,I498758,I498995);
DFFARX1 I_29174 (I498947,I3035,I498715,I499035,);
not I_29175 (I499043,I499035);
not I_29176 (I499060,I280542);
not I_29177 (I499077,I280548);
nor I_29178 (I499094,I499077,I280560);
nor I_29179 (I498707,I499043,I499094);
nor I_29180 (I499125,I499077,I280557);
and I_29181 (I499142,I499125,I280536);
or I_29182 (I499159,I499142,I280539);
DFFARX1 I_29183 (I499159,I3035,I498715,I499185,);
nor I_29184 (I498695,I499185,I498741);
not I_29185 (I499207,I499185);
and I_29186 (I499224,I499207,I498741);
nor I_29187 (I498689,I498766,I499224);
nand I_29188 (I499255,I499207,I498817);
nor I_29189 (I498683,I499077,I499255);
nand I_29190 (I498686,I499207,I498995);
nand I_29191 (I499300,I498817,I280548);
nor I_29192 (I498698,I499060,I499300);
not I_29193 (I499361,I3042);
DFFARX1 I_29194 (I141380,I3035,I499361,I499387,);
DFFARX1 I_29195 (I141392,I3035,I499361,I499404,);
not I_29196 (I499412,I499404);
not I_29197 (I499429,I141398);
nor I_29198 (I499446,I499429,I141383);
not I_29199 (I499463,I141374);
nor I_29200 (I499480,I499446,I141395);
nor I_29201 (I499497,I499404,I499480);
DFFARX1 I_29202 (I499497,I3035,I499361,I499347,);
nor I_29203 (I499528,I141395,I141383);
nand I_29204 (I499545,I499528,I141398);
DFFARX1 I_29205 (I499545,I3035,I499361,I499350,);
nor I_29206 (I499576,I499463,I141395);
nand I_29207 (I499593,I499576,I141377);
nor I_29208 (I499610,I499387,I499593);
DFFARX1 I_29209 (I499610,I3035,I499361,I499326,);
not I_29210 (I499641,I499593);
nand I_29211 (I499338,I499404,I499641);
DFFARX1 I_29212 (I499593,I3035,I499361,I499681,);
not I_29213 (I499689,I499681);
not I_29214 (I499706,I141395);
not I_29215 (I499723,I141386);
nor I_29216 (I499740,I499723,I141374);
nor I_29217 (I499353,I499689,I499740);
nor I_29218 (I499771,I499723,I141389);
and I_29219 (I499788,I499771,I141377);
or I_29220 (I499805,I499788,I141374);
DFFARX1 I_29221 (I499805,I3035,I499361,I499831,);
nor I_29222 (I499341,I499831,I499387);
not I_29223 (I499853,I499831);
and I_29224 (I499870,I499853,I499387);
nor I_29225 (I499335,I499412,I499870);
nand I_29226 (I499901,I499853,I499463);
nor I_29227 (I499329,I499723,I499901);
nand I_29228 (I499332,I499853,I499641);
nand I_29229 (I499946,I499463,I141386);
nor I_29230 (I499344,I499706,I499946);
not I_29231 (I500007,I3042);
DFFARX1 I_29232 (I153461,I3035,I500007,I500033,);
DFFARX1 I_29233 (I153467,I3035,I500007,I500050,);
not I_29234 (I500058,I500050);
not I_29235 (I500075,I153488);
nor I_29236 (I500092,I500075,I153476);
not I_29237 (I500109,I153485);
nor I_29238 (I500126,I500092,I153470);
nor I_29239 (I500143,I500050,I500126);
DFFARX1 I_29240 (I500143,I3035,I500007,I499993,);
nor I_29241 (I500174,I153470,I153476);
nand I_29242 (I500191,I500174,I153488);
DFFARX1 I_29243 (I500191,I3035,I500007,I499996,);
nor I_29244 (I500222,I500109,I153470);
nand I_29245 (I500239,I500222,I153461);
nor I_29246 (I500256,I500033,I500239);
DFFARX1 I_29247 (I500256,I3035,I500007,I499972,);
not I_29248 (I500287,I500239);
nand I_29249 (I499984,I500050,I500287);
DFFARX1 I_29250 (I500239,I3035,I500007,I500327,);
not I_29251 (I500335,I500327);
not I_29252 (I500352,I153470);
not I_29253 (I500369,I153473);
nor I_29254 (I500386,I500369,I153485);
nor I_29255 (I499999,I500335,I500386);
nor I_29256 (I500417,I500369,I153482);
and I_29257 (I500434,I500417,I153464);
or I_29258 (I500451,I500434,I153479);
DFFARX1 I_29259 (I500451,I3035,I500007,I500477,);
nor I_29260 (I499987,I500477,I500033);
not I_29261 (I500499,I500477);
and I_29262 (I500516,I500499,I500033);
nor I_29263 (I499981,I500058,I500516);
nand I_29264 (I500547,I500499,I500109);
nor I_29265 (I499975,I500369,I500547);
nand I_29266 (I499978,I500499,I500287);
nand I_29267 (I500592,I500109,I153473);
nor I_29268 (I499990,I500352,I500592);
not I_29269 (I500653,I3042);
DFFARX1 I_29270 (I381658,I3035,I500653,I500679,);
DFFARX1 I_29271 (I381652,I3035,I500653,I500696,);
not I_29272 (I500704,I500696);
not I_29273 (I500721,I381667);
nor I_29274 (I500738,I500721,I381652);
not I_29275 (I500755,I381661);
nor I_29276 (I500772,I500738,I381670);
nor I_29277 (I500789,I500696,I500772);
DFFARX1 I_29278 (I500789,I3035,I500653,I500639,);
nor I_29279 (I500820,I381670,I381652);
nand I_29280 (I500837,I500820,I381667);
DFFARX1 I_29281 (I500837,I3035,I500653,I500642,);
nor I_29282 (I500868,I500755,I381670);
nand I_29283 (I500885,I500868,I381655);
nor I_29284 (I500902,I500679,I500885);
DFFARX1 I_29285 (I500902,I3035,I500653,I500618,);
not I_29286 (I500933,I500885);
nand I_29287 (I500630,I500696,I500933);
DFFARX1 I_29288 (I500885,I3035,I500653,I500973,);
not I_29289 (I500981,I500973);
not I_29290 (I500998,I381670);
not I_29291 (I501015,I381664);
nor I_29292 (I501032,I501015,I381661);
nor I_29293 (I500645,I500981,I501032);
nor I_29294 (I501063,I501015,I381673);
and I_29295 (I501080,I501063,I381676);
or I_29296 (I501097,I501080,I381655);
DFFARX1 I_29297 (I501097,I3035,I500653,I501123,);
nor I_29298 (I500633,I501123,I500679);
not I_29299 (I501145,I501123);
and I_29300 (I501162,I501145,I500679);
nor I_29301 (I500627,I500704,I501162);
nand I_29302 (I501193,I501145,I500755);
nor I_29303 (I500621,I501015,I501193);
nand I_29304 (I500624,I501145,I500933);
nand I_29305 (I501238,I500755,I381664);
nor I_29306 (I500636,I500998,I501238);
not I_29307 (I501299,I3042);
DFFARX1 I_29308 (I120555,I3035,I501299,I501325,);
DFFARX1 I_29309 (I120567,I3035,I501299,I501342,);
not I_29310 (I501350,I501342);
not I_29311 (I501367,I120573);
nor I_29312 (I501384,I501367,I120558);
not I_29313 (I501401,I120549);
nor I_29314 (I501418,I501384,I120570);
nor I_29315 (I501435,I501342,I501418);
DFFARX1 I_29316 (I501435,I3035,I501299,I501285,);
nor I_29317 (I501466,I120570,I120558);
nand I_29318 (I501483,I501466,I120573);
DFFARX1 I_29319 (I501483,I3035,I501299,I501288,);
nor I_29320 (I501514,I501401,I120570);
nand I_29321 (I501531,I501514,I120552);
nor I_29322 (I501548,I501325,I501531);
DFFARX1 I_29323 (I501548,I3035,I501299,I501264,);
not I_29324 (I501579,I501531);
nand I_29325 (I501276,I501342,I501579);
DFFARX1 I_29326 (I501531,I3035,I501299,I501619,);
not I_29327 (I501627,I501619);
not I_29328 (I501644,I120570);
not I_29329 (I501661,I120561);
nor I_29330 (I501678,I501661,I120549);
nor I_29331 (I501291,I501627,I501678);
nor I_29332 (I501709,I501661,I120564);
and I_29333 (I501726,I501709,I120552);
or I_29334 (I501743,I501726,I120549);
DFFARX1 I_29335 (I501743,I3035,I501299,I501769,);
nor I_29336 (I501279,I501769,I501325);
not I_29337 (I501791,I501769);
and I_29338 (I501808,I501791,I501325);
nor I_29339 (I501273,I501350,I501808);
nand I_29340 (I501839,I501791,I501401);
nor I_29341 (I501267,I501661,I501839);
nand I_29342 (I501270,I501791,I501579);
nand I_29343 (I501884,I501401,I120561);
nor I_29344 (I501282,I501644,I501884);
not I_29345 (I501945,I3042);
DFFARX1 I_29346 (I228295,I3035,I501945,I501971,);
DFFARX1 I_29347 (I228301,I3035,I501945,I501988,);
not I_29348 (I501996,I501988);
not I_29349 (I502013,I228322);
nor I_29350 (I502030,I502013,I228310);
not I_29351 (I502047,I228319);
nor I_29352 (I502064,I502030,I228304);
nor I_29353 (I502081,I501988,I502064);
DFFARX1 I_29354 (I502081,I3035,I501945,I501931,);
nor I_29355 (I502112,I228304,I228310);
nand I_29356 (I502129,I502112,I228322);
DFFARX1 I_29357 (I502129,I3035,I501945,I501934,);
nor I_29358 (I502160,I502047,I228304);
nand I_29359 (I502177,I502160,I228295);
nor I_29360 (I502194,I501971,I502177);
DFFARX1 I_29361 (I502194,I3035,I501945,I501910,);
not I_29362 (I502225,I502177);
nand I_29363 (I501922,I501988,I502225);
DFFARX1 I_29364 (I502177,I3035,I501945,I502265,);
not I_29365 (I502273,I502265);
not I_29366 (I502290,I228304);
not I_29367 (I502307,I228307);
nor I_29368 (I502324,I502307,I228319);
nor I_29369 (I501937,I502273,I502324);
nor I_29370 (I502355,I502307,I228316);
and I_29371 (I502372,I502355,I228298);
or I_29372 (I502389,I502372,I228313);
DFFARX1 I_29373 (I502389,I3035,I501945,I502415,);
nor I_29374 (I501925,I502415,I501971);
not I_29375 (I502437,I502415);
and I_29376 (I502454,I502437,I501971);
nor I_29377 (I501919,I501996,I502454);
nand I_29378 (I502485,I502437,I502047);
nor I_29379 (I501913,I502307,I502485);
nand I_29380 (I501916,I502437,I502225);
nand I_29381 (I502530,I502047,I228307);
nor I_29382 (I501928,I502290,I502530);
not I_29383 (I502591,I3042);
DFFARX1 I_29384 (I345244,I3035,I502591,I502617,);
DFFARX1 I_29385 (I345238,I3035,I502591,I502634,);
not I_29386 (I502642,I502634);
not I_29387 (I502659,I345253);
nor I_29388 (I502676,I502659,I345238);
not I_29389 (I502693,I345247);
nor I_29390 (I502710,I502676,I345256);
nor I_29391 (I502727,I502634,I502710);
DFFARX1 I_29392 (I502727,I3035,I502591,I502577,);
nor I_29393 (I502758,I345256,I345238);
nand I_29394 (I502775,I502758,I345253);
DFFARX1 I_29395 (I502775,I3035,I502591,I502580,);
nor I_29396 (I502806,I502693,I345256);
nand I_29397 (I502823,I502806,I345241);
nor I_29398 (I502840,I502617,I502823);
DFFARX1 I_29399 (I502840,I3035,I502591,I502556,);
not I_29400 (I502871,I502823);
nand I_29401 (I502568,I502634,I502871);
DFFARX1 I_29402 (I502823,I3035,I502591,I502911,);
not I_29403 (I502919,I502911);
not I_29404 (I502936,I345256);
not I_29405 (I502953,I345250);
nor I_29406 (I502970,I502953,I345247);
nor I_29407 (I502583,I502919,I502970);
nor I_29408 (I503001,I502953,I345259);
and I_29409 (I503018,I503001,I345262);
or I_29410 (I503035,I503018,I345241);
DFFARX1 I_29411 (I503035,I3035,I502591,I503061,);
nor I_29412 (I502571,I503061,I502617);
not I_29413 (I503083,I503061);
and I_29414 (I503100,I503083,I502617);
nor I_29415 (I502565,I502642,I503100);
nand I_29416 (I503131,I503083,I502693);
nor I_29417 (I502559,I502953,I503131);
nand I_29418 (I502562,I503083,I502871);
nand I_29419 (I503176,I502693,I345250);
nor I_29420 (I502574,I502936,I503176);
not I_29421 (I503237,I3042);
DFFARX1 I_29422 (I6023,I3035,I503237,I503263,);
DFFARX1 I_29423 (I6020,I3035,I503237,I503280,);
not I_29424 (I503288,I503280);
not I_29425 (I503305,I6032);
nor I_29426 (I503322,I503305,I6029);
not I_29427 (I503339,I6038);
nor I_29428 (I503356,I503322,I6035);
nor I_29429 (I503373,I503280,I503356);
DFFARX1 I_29430 (I503373,I3035,I503237,I503223,);
nor I_29431 (I503404,I6035,I6029);
nand I_29432 (I503421,I503404,I6032);
DFFARX1 I_29433 (I503421,I3035,I503237,I503226,);
nor I_29434 (I503452,I503339,I6035);
nand I_29435 (I503469,I503452,I6026);
nor I_29436 (I503486,I503263,I503469);
DFFARX1 I_29437 (I503486,I3035,I503237,I503202,);
not I_29438 (I503517,I503469);
nand I_29439 (I503214,I503280,I503517);
DFFARX1 I_29440 (I503469,I3035,I503237,I503557,);
not I_29441 (I503565,I503557);
not I_29442 (I503582,I6035);
not I_29443 (I503599,I6026);
nor I_29444 (I503616,I503599,I6038);
nor I_29445 (I503229,I503565,I503616);
nor I_29446 (I503647,I503599,I6020);
and I_29447 (I503664,I503647,I6041);
or I_29448 (I503681,I503664,I6023);
DFFARX1 I_29449 (I503681,I3035,I503237,I503707,);
nor I_29450 (I503217,I503707,I503263);
not I_29451 (I503729,I503707);
and I_29452 (I503746,I503729,I503263);
nor I_29453 (I503211,I503288,I503746);
nand I_29454 (I503777,I503729,I503339);
nor I_29455 (I503205,I503599,I503777);
nand I_29456 (I503208,I503729,I503517);
nand I_29457 (I503822,I503339,I6026);
nor I_29458 (I503220,I503582,I503822);
not I_29459 (I503883,I3042);
DFFARX1 I_29460 (I331369,I3035,I503883,I503909,);
DFFARX1 I_29461 (I331381,I3035,I503883,I503926,);
not I_29462 (I503934,I503926);
not I_29463 (I503951,I331390);
nor I_29464 (I503968,I503951,I331366);
not I_29465 (I503985,I331384);
nor I_29466 (I504002,I503968,I331378);
nor I_29467 (I504019,I503926,I504002);
DFFARX1 I_29468 (I504019,I3035,I503883,I503869,);
nor I_29469 (I504050,I331378,I331366);
nand I_29470 (I504067,I504050,I331390);
DFFARX1 I_29471 (I504067,I3035,I503883,I503872,);
nor I_29472 (I504098,I503985,I331378);
nand I_29473 (I504115,I504098,I331372);
nor I_29474 (I504132,I503909,I504115);
DFFARX1 I_29475 (I504132,I3035,I503883,I503848,);
not I_29476 (I504163,I504115);
nand I_29477 (I503860,I503926,I504163);
DFFARX1 I_29478 (I504115,I3035,I503883,I504203,);
not I_29479 (I504211,I504203);
not I_29480 (I504228,I331378);
not I_29481 (I504245,I331387);
nor I_29482 (I504262,I504245,I331384);
nor I_29483 (I503875,I504211,I504262);
nor I_29484 (I504293,I504245,I331369);
and I_29485 (I504310,I504293,I331366);
or I_29486 (I504327,I504310,I331375);
DFFARX1 I_29487 (I504327,I3035,I503883,I504353,);
nor I_29488 (I503863,I504353,I503909);
not I_29489 (I504375,I504353);
and I_29490 (I504392,I504375,I503909);
nor I_29491 (I503857,I503934,I504392);
nand I_29492 (I504423,I504375,I503985);
nor I_29493 (I503851,I504245,I504423);
nand I_29494 (I503854,I504375,I504163);
nand I_29495 (I504468,I503985,I331387);
nor I_29496 (I503866,I504228,I504468);
not I_29497 (I504529,I3042);
DFFARX1 I_29498 (I241323,I3035,I504529,I504555,);
DFFARX1 I_29499 (I241320,I3035,I504529,I504572,);
not I_29500 (I504580,I504572);
not I_29501 (I504597,I241335);
nor I_29502 (I504614,I504597,I241338);
not I_29503 (I504631,I241326);
nor I_29504 (I504648,I504614,I241332);
nor I_29505 (I504665,I504572,I504648);
DFFARX1 I_29506 (I504665,I3035,I504529,I504515,);
nor I_29507 (I504696,I241332,I241338);
nand I_29508 (I504713,I504696,I241335);
DFFARX1 I_29509 (I504713,I3035,I504529,I504518,);
nor I_29510 (I504744,I504631,I241332);
nand I_29511 (I504761,I504744,I241344);
nor I_29512 (I504778,I504555,I504761);
DFFARX1 I_29513 (I504778,I3035,I504529,I504494,);
not I_29514 (I504809,I504761);
nand I_29515 (I504506,I504572,I504809);
DFFARX1 I_29516 (I504761,I3035,I504529,I504849,);
not I_29517 (I504857,I504849);
not I_29518 (I504874,I241332);
not I_29519 (I504891,I241317);
nor I_29520 (I504908,I504891,I241326);
nor I_29521 (I504521,I504857,I504908);
nor I_29522 (I504939,I504891,I241329);
and I_29523 (I504956,I504939,I241317);
or I_29524 (I504973,I504956,I241341);
DFFARX1 I_29525 (I504973,I3035,I504529,I504999,);
nor I_29526 (I504509,I504999,I504555);
not I_29527 (I505021,I504999);
and I_29528 (I505038,I505021,I504555);
nor I_29529 (I504503,I504580,I505038);
nand I_29530 (I505069,I505021,I504631);
nor I_29531 (I504497,I504891,I505069);
nand I_29532 (I504500,I505021,I504809);
nand I_29533 (I505114,I504631,I241317);
nor I_29534 (I504512,I504874,I505114);
not I_29535 (I505175,I3042);
DFFARX1 I_29536 (I335415,I3035,I505175,I505201,);
DFFARX1 I_29537 (I335427,I3035,I505175,I505218,);
not I_29538 (I505226,I505218);
not I_29539 (I505243,I335436);
nor I_29540 (I505260,I505243,I335412);
not I_29541 (I505277,I335430);
nor I_29542 (I505294,I505260,I335424);
nor I_29543 (I505311,I505218,I505294);
DFFARX1 I_29544 (I505311,I3035,I505175,I505161,);
nor I_29545 (I505342,I335424,I335412);
nand I_29546 (I505359,I505342,I335436);
DFFARX1 I_29547 (I505359,I3035,I505175,I505164,);
nor I_29548 (I505390,I505277,I335424);
nand I_29549 (I505407,I505390,I335418);
nor I_29550 (I505424,I505201,I505407);
DFFARX1 I_29551 (I505424,I3035,I505175,I505140,);
not I_29552 (I505455,I505407);
nand I_29553 (I505152,I505218,I505455);
DFFARX1 I_29554 (I505407,I3035,I505175,I505495,);
not I_29555 (I505503,I505495);
not I_29556 (I505520,I335424);
not I_29557 (I505537,I335433);
nor I_29558 (I505554,I505537,I335430);
nor I_29559 (I505167,I505503,I505554);
nor I_29560 (I505585,I505537,I335415);
and I_29561 (I505602,I505585,I335412);
or I_29562 (I505619,I505602,I335421);
DFFARX1 I_29563 (I505619,I3035,I505175,I505645,);
nor I_29564 (I505155,I505645,I505201);
not I_29565 (I505667,I505645);
and I_29566 (I505684,I505667,I505201);
nor I_29567 (I505149,I505226,I505684);
nand I_29568 (I505715,I505667,I505277);
nor I_29569 (I505143,I505537,I505715);
nand I_29570 (I505146,I505667,I505455);
nand I_29571 (I505760,I505277,I335433);
nor I_29572 (I505158,I505520,I505760);
not I_29573 (I505821,I3042);
DFFARX1 I_29574 (I156623,I3035,I505821,I505847,);
DFFARX1 I_29575 (I156629,I3035,I505821,I505864,);
not I_29576 (I505872,I505864);
not I_29577 (I505889,I156650);
nor I_29578 (I505906,I505889,I156638);
not I_29579 (I505923,I156647);
nor I_29580 (I505940,I505906,I156632);
nor I_29581 (I505957,I505864,I505940);
DFFARX1 I_29582 (I505957,I3035,I505821,I505807,);
nor I_29583 (I505988,I156632,I156638);
nand I_29584 (I506005,I505988,I156650);
DFFARX1 I_29585 (I506005,I3035,I505821,I505810,);
nor I_29586 (I506036,I505923,I156632);
nand I_29587 (I506053,I506036,I156623);
nor I_29588 (I506070,I505847,I506053);
DFFARX1 I_29589 (I506070,I3035,I505821,I505786,);
not I_29590 (I506101,I506053);
nand I_29591 (I505798,I505864,I506101);
DFFARX1 I_29592 (I506053,I3035,I505821,I506141,);
not I_29593 (I506149,I506141);
not I_29594 (I506166,I156632);
not I_29595 (I506183,I156635);
nor I_29596 (I506200,I506183,I156647);
nor I_29597 (I505813,I506149,I506200);
nor I_29598 (I506231,I506183,I156644);
and I_29599 (I506248,I506231,I156626);
or I_29600 (I506265,I506248,I156641);
DFFARX1 I_29601 (I506265,I3035,I505821,I506291,);
nor I_29602 (I505801,I506291,I505847);
not I_29603 (I506313,I506291);
and I_29604 (I506330,I506313,I505847);
nor I_29605 (I505795,I505872,I506330);
nand I_29606 (I506361,I506313,I505923);
nor I_29607 (I505789,I506183,I506361);
nand I_29608 (I505792,I506313,I506101);
nand I_29609 (I506406,I505923,I156635);
nor I_29610 (I505804,I506166,I506406);
not I_29611 (I506467,I3042);
DFFARX1 I_29612 (I383970,I3035,I506467,I506493,);
DFFARX1 I_29613 (I383964,I3035,I506467,I506510,);
not I_29614 (I506518,I506510);
not I_29615 (I506535,I383979);
nor I_29616 (I506552,I506535,I383964);
not I_29617 (I506569,I383973);
nor I_29618 (I506586,I506552,I383982);
nor I_29619 (I506603,I506510,I506586);
DFFARX1 I_29620 (I506603,I3035,I506467,I506453,);
nor I_29621 (I506634,I383982,I383964);
nand I_29622 (I506651,I506634,I383979);
DFFARX1 I_29623 (I506651,I3035,I506467,I506456,);
nor I_29624 (I506682,I506569,I383982);
nand I_29625 (I506699,I506682,I383967);
nor I_29626 (I506716,I506493,I506699);
DFFARX1 I_29627 (I506716,I3035,I506467,I506432,);
not I_29628 (I506747,I506699);
nand I_29629 (I506444,I506510,I506747);
DFFARX1 I_29630 (I506699,I3035,I506467,I506787,);
not I_29631 (I506795,I506787);
not I_29632 (I506812,I383982);
not I_29633 (I506829,I383976);
nor I_29634 (I506846,I506829,I383973);
nor I_29635 (I506459,I506795,I506846);
nor I_29636 (I506877,I506829,I383985);
and I_29637 (I506894,I506877,I383988);
or I_29638 (I506911,I506894,I383967);
DFFARX1 I_29639 (I506911,I3035,I506467,I506937,);
nor I_29640 (I506447,I506937,I506493);
not I_29641 (I506959,I506937);
and I_29642 (I506976,I506959,I506493);
nor I_29643 (I506441,I506518,I506976);
nand I_29644 (I507007,I506959,I506569);
nor I_29645 (I506435,I506829,I507007);
nand I_29646 (I506438,I506959,I506747);
nand I_29647 (I507052,I506569,I383976);
nor I_29648 (I506450,I506812,I507052);
not I_29649 (I507113,I3042);
DFFARX1 I_29650 (I174541,I3035,I507113,I507139,);
DFFARX1 I_29651 (I174547,I3035,I507113,I507156,);
not I_29652 (I507164,I507156);
not I_29653 (I507181,I174568);
nor I_29654 (I507198,I507181,I174556);
not I_29655 (I507215,I174565);
nor I_29656 (I507232,I507198,I174550);
nor I_29657 (I507249,I507156,I507232);
DFFARX1 I_29658 (I507249,I3035,I507113,I507099,);
nor I_29659 (I507280,I174550,I174556);
nand I_29660 (I507297,I507280,I174568);
DFFARX1 I_29661 (I507297,I3035,I507113,I507102,);
nor I_29662 (I507328,I507215,I174550);
nand I_29663 (I507345,I507328,I174541);
nor I_29664 (I507362,I507139,I507345);
DFFARX1 I_29665 (I507362,I3035,I507113,I507078,);
not I_29666 (I507393,I507345);
nand I_29667 (I507090,I507156,I507393);
DFFARX1 I_29668 (I507345,I3035,I507113,I507433,);
not I_29669 (I507441,I507433);
not I_29670 (I507458,I174550);
not I_29671 (I507475,I174553);
nor I_29672 (I507492,I507475,I174565);
nor I_29673 (I507105,I507441,I507492);
nor I_29674 (I507523,I507475,I174562);
and I_29675 (I507540,I507523,I174544);
or I_29676 (I507557,I507540,I174559);
DFFARX1 I_29677 (I507557,I3035,I507113,I507583,);
nor I_29678 (I507093,I507583,I507139);
not I_29679 (I507605,I507583);
and I_29680 (I507622,I507605,I507139);
nor I_29681 (I507087,I507164,I507622);
nand I_29682 (I507653,I507605,I507215);
nor I_29683 (I507081,I507475,I507653);
nand I_29684 (I507084,I507605,I507393);
nand I_29685 (I507698,I507215,I174553);
nor I_29686 (I507096,I507458,I507698);
not I_29687 (I507759,I3042);
DFFARX1 I_29688 (I202999,I3035,I507759,I507785,);
DFFARX1 I_29689 (I203005,I3035,I507759,I507802,);
not I_29690 (I507810,I507802);
not I_29691 (I507827,I203026);
nor I_29692 (I507844,I507827,I203014);
not I_29693 (I507861,I203023);
nor I_29694 (I507878,I507844,I203008);
nor I_29695 (I507895,I507802,I507878);
DFFARX1 I_29696 (I507895,I3035,I507759,I507745,);
nor I_29697 (I507926,I203008,I203014);
nand I_29698 (I507943,I507926,I203026);
DFFARX1 I_29699 (I507943,I3035,I507759,I507748,);
nor I_29700 (I507974,I507861,I203008);
nand I_29701 (I507991,I507974,I202999);
nor I_29702 (I508008,I507785,I507991);
DFFARX1 I_29703 (I508008,I3035,I507759,I507724,);
not I_29704 (I508039,I507991);
nand I_29705 (I507736,I507802,I508039);
DFFARX1 I_29706 (I507991,I3035,I507759,I508079,);
not I_29707 (I508087,I508079);
not I_29708 (I508104,I203008);
not I_29709 (I508121,I203011);
nor I_29710 (I508138,I508121,I203023);
nor I_29711 (I507751,I508087,I508138);
nor I_29712 (I508169,I508121,I203020);
and I_29713 (I508186,I508169,I203002);
or I_29714 (I508203,I508186,I203017);
DFFARX1 I_29715 (I508203,I3035,I507759,I508229,);
nor I_29716 (I507739,I508229,I507785);
not I_29717 (I508251,I508229);
and I_29718 (I508268,I508251,I507785);
nor I_29719 (I507733,I507810,I508268);
nand I_29720 (I508299,I508251,I507861);
nor I_29721 (I507727,I508121,I508299);
nand I_29722 (I507730,I508251,I508039);
nand I_29723 (I508344,I507861,I203011);
nor I_29724 (I507742,I508104,I508344);
not I_29725 (I508405,I3042);
DFFARX1 I_29726 (I743038,I3035,I508405,I508431,);
DFFARX1 I_29727 (I743062,I3035,I508405,I508448,);
not I_29728 (I508456,I508448);
not I_29729 (I508473,I743044);
nor I_29730 (I508490,I508473,I743053);
not I_29731 (I508507,I743038);
nor I_29732 (I508524,I508490,I743059);
nor I_29733 (I508541,I508448,I508524);
DFFARX1 I_29734 (I508541,I3035,I508405,I508391,);
nor I_29735 (I508572,I743059,I743053);
nand I_29736 (I508589,I508572,I743044);
DFFARX1 I_29737 (I508589,I3035,I508405,I508394,);
nor I_29738 (I508620,I508507,I743059);
nand I_29739 (I508637,I508620,I743056);
nor I_29740 (I508654,I508431,I508637);
DFFARX1 I_29741 (I508654,I3035,I508405,I508370,);
not I_29742 (I508685,I508637);
nand I_29743 (I508382,I508448,I508685);
DFFARX1 I_29744 (I508637,I3035,I508405,I508725,);
not I_29745 (I508733,I508725);
not I_29746 (I508750,I743059);
not I_29747 (I508767,I743050);
nor I_29748 (I508784,I508767,I743038);
nor I_29749 (I508397,I508733,I508784);
nor I_29750 (I508815,I508767,I743041);
and I_29751 (I508832,I508815,I743065);
or I_29752 (I508849,I508832,I743047);
DFFARX1 I_29753 (I508849,I3035,I508405,I508875,);
nor I_29754 (I508385,I508875,I508431);
not I_29755 (I508897,I508875);
and I_29756 (I508914,I508897,I508431);
nor I_29757 (I508379,I508456,I508914);
nand I_29758 (I508945,I508897,I508507);
nor I_29759 (I508373,I508767,I508945);
nand I_29760 (I508376,I508897,I508685);
nand I_29761 (I508990,I508507,I743050);
nor I_29762 (I508388,I508750,I508990);
not I_29763 (I509051,I3042);
DFFARX1 I_29764 (I190878,I3035,I509051,I509077,);
DFFARX1 I_29765 (I190884,I3035,I509051,I509094,);
not I_29766 (I509102,I509094);
not I_29767 (I509119,I190905);
nor I_29768 (I509136,I509119,I190893);
not I_29769 (I509153,I190902);
nor I_29770 (I509170,I509136,I190887);
nor I_29771 (I509187,I509094,I509170);
DFFARX1 I_29772 (I509187,I3035,I509051,I509037,);
nor I_29773 (I509218,I190887,I190893);
nand I_29774 (I509235,I509218,I190905);
DFFARX1 I_29775 (I509235,I3035,I509051,I509040,);
nor I_29776 (I509266,I509153,I190887);
nand I_29777 (I509283,I509266,I190878);
nor I_29778 (I509300,I509077,I509283);
DFFARX1 I_29779 (I509300,I3035,I509051,I509016,);
not I_29780 (I509331,I509283);
nand I_29781 (I509028,I509094,I509331);
DFFARX1 I_29782 (I509283,I3035,I509051,I509371,);
not I_29783 (I509379,I509371);
not I_29784 (I509396,I190887);
not I_29785 (I509413,I190890);
nor I_29786 (I509430,I509413,I190902);
nor I_29787 (I509043,I509379,I509430);
nor I_29788 (I509461,I509413,I190899);
and I_29789 (I509478,I509461,I190881);
or I_29790 (I509495,I509478,I190896);
DFFARX1 I_29791 (I509495,I3035,I509051,I509521,);
nor I_29792 (I509031,I509521,I509077);
not I_29793 (I509543,I509521);
and I_29794 (I509560,I509543,I509077);
nor I_29795 (I509025,I509102,I509560);
nand I_29796 (I509591,I509543,I509153);
nor I_29797 (I509019,I509413,I509591);
nand I_29798 (I509022,I509543,I509331);
nand I_29799 (I509636,I509153,I190890);
nor I_29800 (I509034,I509396,I509636);
not I_29801 (I509697,I3042);
DFFARX1 I_29802 (I364896,I3035,I509697,I509723,);
DFFARX1 I_29803 (I364890,I3035,I509697,I509740,);
not I_29804 (I509748,I509740);
not I_29805 (I509765,I364905);
nor I_29806 (I509782,I509765,I364890);
not I_29807 (I509799,I364899);
nor I_29808 (I509816,I509782,I364908);
nor I_29809 (I509833,I509740,I509816);
DFFARX1 I_29810 (I509833,I3035,I509697,I509683,);
nor I_29811 (I509864,I364908,I364890);
nand I_29812 (I509881,I509864,I364905);
DFFARX1 I_29813 (I509881,I3035,I509697,I509686,);
nor I_29814 (I509912,I509799,I364908);
nand I_29815 (I509929,I509912,I364893);
nor I_29816 (I509946,I509723,I509929);
DFFARX1 I_29817 (I509946,I3035,I509697,I509662,);
not I_29818 (I509977,I509929);
nand I_29819 (I509674,I509740,I509977);
DFFARX1 I_29820 (I509929,I3035,I509697,I510017,);
not I_29821 (I510025,I510017);
not I_29822 (I510042,I364908);
not I_29823 (I510059,I364902);
nor I_29824 (I510076,I510059,I364899);
nor I_29825 (I509689,I510025,I510076);
nor I_29826 (I510107,I510059,I364911);
and I_29827 (I510124,I510107,I364914);
or I_29828 (I510141,I510124,I364893);
DFFARX1 I_29829 (I510141,I3035,I509697,I510167,);
nor I_29830 (I509677,I510167,I509723);
not I_29831 (I510189,I510167);
and I_29832 (I510206,I510189,I509723);
nor I_29833 (I509671,I509748,I510206);
nand I_29834 (I510237,I510189,I509799);
nor I_29835 (I509665,I510059,I510237);
nand I_29836 (I509668,I510189,I509977);
nand I_29837 (I510282,I509799,I364902);
nor I_29838 (I509680,I510042,I510282);
not I_29839 (I510343,I3042);
DFFARX1 I_29840 (I100325,I3035,I510343,I510369,);
DFFARX1 I_29841 (I100337,I3035,I510343,I510386,);
not I_29842 (I510394,I510386);
not I_29843 (I510411,I100343);
nor I_29844 (I510428,I510411,I100328);
not I_29845 (I510445,I100319);
nor I_29846 (I510462,I510428,I100340);
nor I_29847 (I510479,I510386,I510462);
DFFARX1 I_29848 (I510479,I3035,I510343,I510329,);
nor I_29849 (I510510,I100340,I100328);
nand I_29850 (I510527,I510510,I100343);
DFFARX1 I_29851 (I510527,I3035,I510343,I510332,);
nor I_29852 (I510558,I510445,I100340);
nand I_29853 (I510575,I510558,I100322);
nor I_29854 (I510592,I510369,I510575);
DFFARX1 I_29855 (I510592,I3035,I510343,I510308,);
not I_29856 (I510623,I510575);
nand I_29857 (I510320,I510386,I510623);
DFFARX1 I_29858 (I510575,I3035,I510343,I510663,);
not I_29859 (I510671,I510663);
not I_29860 (I510688,I100340);
not I_29861 (I510705,I100331);
nor I_29862 (I510722,I510705,I100319);
nor I_29863 (I510335,I510671,I510722);
nor I_29864 (I510753,I510705,I100334);
and I_29865 (I510770,I510753,I100322);
or I_29866 (I510787,I510770,I100319);
DFFARX1 I_29867 (I510787,I3035,I510343,I510813,);
nor I_29868 (I510323,I510813,I510369);
not I_29869 (I510835,I510813);
and I_29870 (I510852,I510835,I510369);
nor I_29871 (I510317,I510394,I510852);
nand I_29872 (I510883,I510835,I510445);
nor I_29873 (I510311,I510705,I510883);
nand I_29874 (I510314,I510835,I510623);
nand I_29875 (I510928,I510445,I100331);
nor I_29876 (I510326,I510688,I510928);
not I_29877 (I510989,I3042);
DFFARX1 I_29878 (I566680,I3035,I510989,I511015,);
DFFARX1 I_29879 (I566683,I3035,I510989,I511032,);
not I_29880 (I511040,I511032);
not I_29881 (I511057,I566680);
nor I_29882 (I511074,I511057,I566692);
not I_29883 (I511091,I566701);
nor I_29884 (I511108,I511074,I566689);
nor I_29885 (I511125,I511032,I511108);
DFFARX1 I_29886 (I511125,I3035,I510989,I510975,);
nor I_29887 (I511156,I566689,I566692);
nand I_29888 (I511173,I511156,I566680);
DFFARX1 I_29889 (I511173,I3035,I510989,I510978,);
nor I_29890 (I511204,I511091,I566689);
nand I_29891 (I511221,I511204,I566695);
nor I_29892 (I511238,I511015,I511221);
DFFARX1 I_29893 (I511238,I3035,I510989,I510954,);
not I_29894 (I511269,I511221);
nand I_29895 (I510966,I511032,I511269);
DFFARX1 I_29896 (I511221,I3035,I510989,I511309,);
not I_29897 (I511317,I511309);
not I_29898 (I511334,I566689);
not I_29899 (I511351,I566686);
nor I_29900 (I511368,I511351,I566701);
nor I_29901 (I510981,I511317,I511368);
nor I_29902 (I511399,I511351,I566698);
and I_29903 (I511416,I511399,I566686);
or I_29904 (I511433,I511416,I566683);
DFFARX1 I_29905 (I511433,I3035,I510989,I511459,);
nor I_29906 (I510969,I511459,I511015);
not I_29907 (I511481,I511459);
and I_29908 (I511498,I511481,I511015);
nor I_29909 (I510963,I511040,I511498);
nand I_29910 (I511529,I511481,I511091);
nor I_29911 (I510957,I511351,I511529);
nand I_29912 (I510960,I511481,I511269);
nand I_29913 (I511574,I511091,I566686);
nor I_29914 (I510972,I511334,I511574);
not I_29915 (I511635,I3042);
DFFARX1 I_29916 (I199837,I3035,I511635,I511661,);
DFFARX1 I_29917 (I199843,I3035,I511635,I511678,);
not I_29918 (I511686,I511678);
not I_29919 (I511703,I199864);
nor I_29920 (I511720,I511703,I199852);
not I_29921 (I511737,I199861);
nor I_29922 (I511754,I511720,I199846);
nor I_29923 (I511771,I511678,I511754);
DFFARX1 I_29924 (I511771,I3035,I511635,I511621,);
nor I_29925 (I511802,I199846,I199852);
nand I_29926 (I511819,I511802,I199864);
DFFARX1 I_29927 (I511819,I3035,I511635,I511624,);
nor I_29928 (I511850,I511737,I199846);
nand I_29929 (I511867,I511850,I199837);
nor I_29930 (I511884,I511661,I511867);
DFFARX1 I_29931 (I511884,I3035,I511635,I511600,);
not I_29932 (I511915,I511867);
nand I_29933 (I511612,I511678,I511915);
DFFARX1 I_29934 (I511867,I3035,I511635,I511955,);
not I_29935 (I511963,I511955);
not I_29936 (I511980,I199846);
not I_29937 (I511997,I199849);
nor I_29938 (I512014,I511997,I199861);
nor I_29939 (I511627,I511963,I512014);
nor I_29940 (I512045,I511997,I199858);
and I_29941 (I512062,I512045,I199840);
or I_29942 (I512079,I512062,I199855);
DFFARX1 I_29943 (I512079,I3035,I511635,I512105,);
nor I_29944 (I511615,I512105,I511661);
not I_29945 (I512127,I512105);
and I_29946 (I512144,I512127,I511661);
nor I_29947 (I511609,I511686,I512144);
nand I_29948 (I512175,I512127,I511737);
nor I_29949 (I511603,I511997,I512175);
nand I_29950 (I511606,I512127,I511915);
nand I_29951 (I512220,I511737,I199849);
nor I_29952 (I511618,I511980,I512220);
not I_29953 (I512281,I3042);
DFFARX1 I_29954 (I724593,I3035,I512281,I512307,);
DFFARX1 I_29955 (I724617,I3035,I512281,I512324,);
not I_29956 (I512332,I512324);
not I_29957 (I512349,I724599);
nor I_29958 (I512366,I512349,I724608);
not I_29959 (I512383,I724593);
nor I_29960 (I512400,I512366,I724614);
nor I_29961 (I512417,I512324,I512400);
DFFARX1 I_29962 (I512417,I3035,I512281,I512267,);
nor I_29963 (I512448,I724614,I724608);
nand I_29964 (I512465,I512448,I724599);
DFFARX1 I_29965 (I512465,I3035,I512281,I512270,);
nor I_29966 (I512496,I512383,I724614);
nand I_29967 (I512513,I512496,I724611);
nor I_29968 (I512530,I512307,I512513);
DFFARX1 I_29969 (I512530,I3035,I512281,I512246,);
not I_29970 (I512561,I512513);
nand I_29971 (I512258,I512324,I512561);
DFFARX1 I_29972 (I512513,I3035,I512281,I512601,);
not I_29973 (I512609,I512601);
not I_29974 (I512626,I724614);
not I_29975 (I512643,I724605);
nor I_29976 (I512660,I512643,I724593);
nor I_29977 (I512273,I512609,I512660);
nor I_29978 (I512691,I512643,I724596);
and I_29979 (I512708,I512691,I724620);
or I_29980 (I512725,I512708,I724602);
DFFARX1 I_29981 (I512725,I3035,I512281,I512751,);
nor I_29982 (I512261,I512751,I512307);
not I_29983 (I512773,I512751);
and I_29984 (I512790,I512773,I512307);
nor I_29985 (I512255,I512332,I512790);
nand I_29986 (I512821,I512773,I512383);
nor I_29987 (I512249,I512643,I512821);
nand I_29988 (I512252,I512773,I512561);
nand I_29989 (I512866,I512383,I724605);
nor I_29990 (I512264,I512626,I512866);
not I_29991 (I512927,I3042);
DFFARX1 I_29992 (I444575,I3035,I512927,I512953,);
DFFARX1 I_29993 (I444572,I3035,I512927,I512970,);
not I_29994 (I512978,I512970);
not I_29995 (I512995,I444572);
nor I_29996 (I513012,I512995,I444575);
not I_29997 (I513029,I444587);
nor I_29998 (I513046,I513012,I444581);
nor I_29999 (I513063,I512970,I513046);
DFFARX1 I_30000 (I513063,I3035,I512927,I512913,);
nor I_30001 (I513094,I444581,I444575);
nand I_30002 (I513111,I513094,I444572);
DFFARX1 I_30003 (I513111,I3035,I512927,I512916,);
nor I_30004 (I513142,I513029,I444581);
nand I_30005 (I513159,I513142,I444569);
nor I_30006 (I513176,I512953,I513159);
DFFARX1 I_30007 (I513176,I3035,I512927,I512892,);
not I_30008 (I513207,I513159);
nand I_30009 (I512904,I512970,I513207);
DFFARX1 I_30010 (I513159,I3035,I512927,I513247,);
not I_30011 (I513255,I513247);
not I_30012 (I513272,I444581);
not I_30013 (I513289,I444578);
nor I_30014 (I513306,I513289,I444587);
nor I_30015 (I512919,I513255,I513306);
nor I_30016 (I513337,I513289,I444584);
and I_30017 (I513354,I513337,I444590);
or I_30018 (I513371,I513354,I444569);
DFFARX1 I_30019 (I513371,I3035,I512927,I513397,);
nor I_30020 (I512907,I513397,I512953);
not I_30021 (I513419,I513397);
and I_30022 (I513436,I513419,I512953);
nor I_30023 (I512901,I512978,I513436);
nand I_30024 (I513467,I513419,I513029);
nor I_30025 (I512895,I513289,I513467);
nand I_30026 (I512898,I513419,I513207);
nand I_30027 (I513512,I513029,I444578);
nor I_30028 (I512910,I513272,I513512);
not I_30029 (I513573,I3042);
DFFARX1 I_30030 (I327323,I3035,I513573,I513599,);
DFFARX1 I_30031 (I327335,I3035,I513573,I513616,);
not I_30032 (I513624,I513616);
not I_30033 (I513641,I327344);
nor I_30034 (I513658,I513641,I327320);
not I_30035 (I513675,I327338);
nor I_30036 (I513692,I513658,I327332);
nor I_30037 (I513709,I513616,I513692);
DFFARX1 I_30038 (I513709,I3035,I513573,I513559,);
nor I_30039 (I513740,I327332,I327320);
nand I_30040 (I513757,I513740,I327344);
DFFARX1 I_30041 (I513757,I3035,I513573,I513562,);
nor I_30042 (I513788,I513675,I327332);
nand I_30043 (I513805,I513788,I327326);
nor I_30044 (I513822,I513599,I513805);
DFFARX1 I_30045 (I513822,I3035,I513573,I513538,);
not I_30046 (I513853,I513805);
nand I_30047 (I513550,I513616,I513853);
DFFARX1 I_30048 (I513805,I3035,I513573,I513893,);
not I_30049 (I513901,I513893);
not I_30050 (I513918,I327332);
not I_30051 (I513935,I327341);
nor I_30052 (I513952,I513935,I327338);
nor I_30053 (I513565,I513901,I513952);
nor I_30054 (I513983,I513935,I327323);
and I_30055 (I514000,I513983,I327320);
or I_30056 (I514017,I514000,I327329);
DFFARX1 I_30057 (I514017,I3035,I513573,I514043,);
nor I_30058 (I513553,I514043,I513599);
not I_30059 (I514065,I514043);
and I_30060 (I514082,I514065,I513599);
nor I_30061 (I513547,I513624,I514082);
nand I_30062 (I514113,I514065,I513675);
nor I_30063 (I513541,I513935,I514113);
nand I_30064 (I513544,I514065,I513853);
nand I_30065 (I514158,I513675,I327341);
nor I_30066 (I513556,I513918,I514158);
not I_30067 (I514219,I3042);
DFFARX1 I_30068 (I67883,I3035,I514219,I514245,);
DFFARX1 I_30069 (I67889,I3035,I514219,I514262,);
not I_30070 (I514270,I514262);
not I_30071 (I514287,I67907);
nor I_30072 (I514304,I514287,I67886);
not I_30073 (I514321,I67892);
nor I_30074 (I514338,I514304,I67898);
nor I_30075 (I514355,I514262,I514338);
DFFARX1 I_30076 (I514355,I3035,I514219,I514205,);
nor I_30077 (I514386,I67898,I67886);
nand I_30078 (I514403,I514386,I67907);
DFFARX1 I_30079 (I514403,I3035,I514219,I514208,);
nor I_30080 (I514434,I514321,I67898);
nand I_30081 (I514451,I514434,I67904);
nor I_30082 (I514468,I514245,I514451);
DFFARX1 I_30083 (I514468,I3035,I514219,I514184,);
not I_30084 (I514499,I514451);
nand I_30085 (I514196,I514262,I514499);
DFFARX1 I_30086 (I514451,I3035,I514219,I514539,);
not I_30087 (I514547,I514539);
not I_30088 (I514564,I67898);
not I_30089 (I514581,I67886);
nor I_30090 (I514598,I514581,I67892);
nor I_30091 (I514211,I514547,I514598);
nor I_30092 (I514629,I514581,I67895);
and I_30093 (I514646,I514629,I67883);
or I_30094 (I514663,I514646,I67901);
DFFARX1 I_30095 (I514663,I3035,I514219,I514689,);
nor I_30096 (I514199,I514689,I514245);
not I_30097 (I514711,I514689);
and I_30098 (I514728,I514711,I514245);
nor I_30099 (I514193,I514270,I514728);
nand I_30100 (I514759,I514711,I514321);
nor I_30101 (I514187,I514581,I514759);
nand I_30102 (I514190,I514711,I514499);
nand I_30103 (I514804,I514321,I67886);
nor I_30104 (I514202,I514564,I514804);
not I_30105 (I514865,I3042);
DFFARX1 I_30106 (I626640,I3035,I514865,I514891,);
DFFARX1 I_30107 (I626622,I3035,I514865,I514908,);
not I_30108 (I514916,I514908);
not I_30109 (I514933,I626631);
nor I_30110 (I514950,I514933,I626643);
not I_30111 (I514967,I626625);
nor I_30112 (I514984,I514950,I626634);
nor I_30113 (I515001,I514908,I514984);
DFFARX1 I_30114 (I515001,I3035,I514865,I514851,);
nor I_30115 (I515032,I626634,I626643);
nand I_30116 (I515049,I515032,I626631);
DFFARX1 I_30117 (I515049,I3035,I514865,I514854,);
nor I_30118 (I515080,I514967,I626634);
nand I_30119 (I515097,I515080,I626646);
nor I_30120 (I515114,I514891,I515097);
DFFARX1 I_30121 (I515114,I3035,I514865,I514830,);
not I_30122 (I515145,I515097);
nand I_30123 (I514842,I514908,I515145);
DFFARX1 I_30124 (I515097,I3035,I514865,I515185,);
not I_30125 (I515193,I515185);
not I_30126 (I515210,I626634);
not I_30127 (I515227,I626622);
nor I_30128 (I515244,I515227,I626625);
nor I_30129 (I514857,I515193,I515244);
nor I_30130 (I515275,I515227,I626628);
and I_30131 (I515292,I515275,I626637);
or I_30132 (I515309,I515292,I626625);
DFFARX1 I_30133 (I515309,I3035,I514865,I515335,);
nor I_30134 (I514845,I515335,I514891);
not I_30135 (I515357,I515335);
and I_30136 (I515374,I515357,I514891);
nor I_30137 (I514839,I514916,I515374);
nand I_30138 (I515405,I515357,I514967);
nor I_30139 (I514833,I515227,I515405);
nand I_30140 (I514836,I515357,I515145);
nand I_30141 (I515450,I514967,I626622);
nor I_30142 (I514848,I515210,I515450);
not I_30143 (I515511,I3042);
DFFARX1 I_30144 (I668664,I3035,I515511,I515537,);
DFFARX1 I_30145 (I668670,I3035,I515511,I515554,);
not I_30146 (I515562,I515554);
not I_30147 (I515579,I668667);
nor I_30148 (I515596,I515579,I668646);
not I_30149 (I515613,I668649);
nor I_30150 (I515630,I515596,I668655);
nor I_30151 (I515647,I515554,I515630);
DFFARX1 I_30152 (I515647,I3035,I515511,I515497,);
nor I_30153 (I515678,I668655,I668646);
nand I_30154 (I515695,I515678,I668667);
DFFARX1 I_30155 (I515695,I3035,I515511,I515500,);
nor I_30156 (I515726,I515613,I668655);
nand I_30157 (I515743,I515726,I668649);
nor I_30158 (I515760,I515537,I515743);
DFFARX1 I_30159 (I515760,I3035,I515511,I515476,);
not I_30160 (I515791,I515743);
nand I_30161 (I515488,I515554,I515791);
DFFARX1 I_30162 (I515743,I3035,I515511,I515831,);
not I_30163 (I515839,I515831);
not I_30164 (I515856,I668655);
not I_30165 (I515873,I668658);
nor I_30166 (I515890,I515873,I668649);
nor I_30167 (I515503,I515839,I515890);
nor I_30168 (I515921,I515873,I668646);
and I_30169 (I515938,I515921,I668652);
or I_30170 (I515955,I515938,I668661);
DFFARX1 I_30171 (I515955,I3035,I515511,I515981,);
nor I_30172 (I515491,I515981,I515537);
not I_30173 (I516003,I515981);
and I_30174 (I516020,I516003,I515537);
nor I_30175 (I515485,I515562,I516020);
nand I_30176 (I516051,I516003,I515613);
nor I_30177 (I515479,I515873,I516051);
nand I_30178 (I515482,I516003,I515791);
nand I_30179 (I516096,I515613,I668658);
nor I_30180 (I515494,I515856,I516096);
not I_30181 (I516157,I3042);
DFFARX1 I_30182 (I455642,I3035,I516157,I516183,);
DFFARX1 I_30183 (I455639,I3035,I516157,I516200,);
not I_30184 (I516208,I516200);
not I_30185 (I516225,I455639);
nor I_30186 (I516242,I516225,I455642);
not I_30187 (I516259,I455654);
nor I_30188 (I516276,I516242,I455648);
nor I_30189 (I516293,I516200,I516276);
DFFARX1 I_30190 (I516293,I3035,I516157,I516143,);
nor I_30191 (I516324,I455648,I455642);
nand I_30192 (I516341,I516324,I455639);
DFFARX1 I_30193 (I516341,I3035,I516157,I516146,);
nor I_30194 (I516372,I516259,I455648);
nand I_30195 (I516389,I516372,I455636);
nor I_30196 (I516406,I516183,I516389);
DFFARX1 I_30197 (I516406,I3035,I516157,I516122,);
not I_30198 (I516437,I516389);
nand I_30199 (I516134,I516200,I516437);
DFFARX1 I_30200 (I516389,I3035,I516157,I516477,);
not I_30201 (I516485,I516477);
not I_30202 (I516502,I455648);
not I_30203 (I516519,I455645);
nor I_30204 (I516536,I516519,I455654);
nor I_30205 (I516149,I516485,I516536);
nor I_30206 (I516567,I516519,I455651);
and I_30207 (I516584,I516567,I455657);
or I_30208 (I516601,I516584,I455636);
DFFARX1 I_30209 (I516601,I3035,I516157,I516627,);
nor I_30210 (I516137,I516627,I516183);
not I_30211 (I516649,I516627);
and I_30212 (I516666,I516649,I516183);
nor I_30213 (I516131,I516208,I516666);
nand I_30214 (I516697,I516649,I516259);
nor I_30215 (I516125,I516519,I516697);
nand I_30216 (I516128,I516649,I516437);
nand I_30217 (I516742,I516259,I455645);
nor I_30218 (I516140,I516502,I516742);
not I_30219 (I516803,I3042);
DFFARX1 I_30220 (I93780,I3035,I516803,I516829,);
DFFARX1 I_30221 (I93792,I3035,I516803,I516846,);
not I_30222 (I516854,I516846);
not I_30223 (I516871,I93798);
nor I_30224 (I516888,I516871,I93783);
not I_30225 (I516905,I93774);
nor I_30226 (I516922,I516888,I93795);
nor I_30227 (I516939,I516846,I516922);
DFFARX1 I_30228 (I516939,I3035,I516803,I516789,);
nor I_30229 (I516970,I93795,I93783);
nand I_30230 (I516987,I516970,I93798);
DFFARX1 I_30231 (I516987,I3035,I516803,I516792,);
nor I_30232 (I517018,I516905,I93795);
nand I_30233 (I517035,I517018,I93777);
nor I_30234 (I517052,I516829,I517035);
DFFARX1 I_30235 (I517052,I3035,I516803,I516768,);
not I_30236 (I517083,I517035);
nand I_30237 (I516780,I516846,I517083);
DFFARX1 I_30238 (I517035,I3035,I516803,I517123,);
not I_30239 (I517131,I517123);
not I_30240 (I517148,I93795);
not I_30241 (I517165,I93786);
nor I_30242 (I517182,I517165,I93774);
nor I_30243 (I516795,I517131,I517182);
nor I_30244 (I517213,I517165,I93789);
and I_30245 (I517230,I517213,I93777);
or I_30246 (I517247,I517230,I93774);
DFFARX1 I_30247 (I517247,I3035,I516803,I517273,);
nor I_30248 (I516783,I517273,I516829);
not I_30249 (I517295,I517273);
and I_30250 (I517312,I517295,I516829);
nor I_30251 (I516777,I516854,I517312);
nand I_30252 (I517343,I517295,I516905);
nor I_30253 (I516771,I517165,I517343);
nand I_30254 (I516774,I517295,I517083);
nand I_30255 (I517388,I516905,I93786);
nor I_30256 (I516786,I517148,I517388);
not I_30257 (I517449,I3042);
DFFARX1 I_30258 (I716263,I3035,I517449,I517475,);
DFFARX1 I_30259 (I716287,I3035,I517449,I517492,);
not I_30260 (I517500,I517492);
not I_30261 (I517517,I716269);
nor I_30262 (I517534,I517517,I716278);
not I_30263 (I517551,I716263);
nor I_30264 (I517568,I517534,I716284);
nor I_30265 (I517585,I517492,I517568);
DFFARX1 I_30266 (I517585,I3035,I517449,I517435,);
nor I_30267 (I517616,I716284,I716278);
nand I_30268 (I517633,I517616,I716269);
DFFARX1 I_30269 (I517633,I3035,I517449,I517438,);
nor I_30270 (I517664,I517551,I716284);
nand I_30271 (I517681,I517664,I716281);
nor I_30272 (I517698,I517475,I517681);
DFFARX1 I_30273 (I517698,I3035,I517449,I517414,);
not I_30274 (I517729,I517681);
nand I_30275 (I517426,I517492,I517729);
DFFARX1 I_30276 (I517681,I3035,I517449,I517769,);
not I_30277 (I517777,I517769);
not I_30278 (I517794,I716284);
not I_30279 (I517811,I716275);
nor I_30280 (I517828,I517811,I716263);
nor I_30281 (I517441,I517777,I517828);
nor I_30282 (I517859,I517811,I716266);
and I_30283 (I517876,I517859,I716290);
or I_30284 (I517893,I517876,I716272);
DFFARX1 I_30285 (I517893,I3035,I517449,I517919,);
nor I_30286 (I517429,I517919,I517475);
not I_30287 (I517941,I517919);
and I_30288 (I517958,I517941,I517475);
nor I_30289 (I517423,I517500,I517958);
nand I_30290 (I517989,I517941,I517551);
nor I_30291 (I517417,I517811,I517989);
nand I_30292 (I517420,I517941,I517729);
nand I_30293 (I518034,I517551,I716275);
nor I_30294 (I517432,I517794,I518034);
not I_30295 (I518095,I3042);
DFFARX1 I_30296 (I342354,I3035,I518095,I518121,);
DFFARX1 I_30297 (I342348,I3035,I518095,I518138,);
not I_30298 (I518146,I518138);
not I_30299 (I518163,I342363);
nor I_30300 (I518180,I518163,I342348);
not I_30301 (I518197,I342357);
nor I_30302 (I518214,I518180,I342366);
nor I_30303 (I518231,I518138,I518214);
DFFARX1 I_30304 (I518231,I3035,I518095,I518081,);
nor I_30305 (I518262,I342366,I342348);
nand I_30306 (I518279,I518262,I342363);
DFFARX1 I_30307 (I518279,I3035,I518095,I518084,);
nor I_30308 (I518310,I518197,I342366);
nand I_30309 (I518327,I518310,I342351);
nor I_30310 (I518344,I518121,I518327);
DFFARX1 I_30311 (I518344,I3035,I518095,I518060,);
not I_30312 (I518375,I518327);
nand I_30313 (I518072,I518138,I518375);
DFFARX1 I_30314 (I518327,I3035,I518095,I518415,);
not I_30315 (I518423,I518415);
not I_30316 (I518440,I342366);
not I_30317 (I518457,I342360);
nor I_30318 (I518474,I518457,I342357);
nor I_30319 (I518087,I518423,I518474);
nor I_30320 (I518505,I518457,I342369);
and I_30321 (I518522,I518505,I342372);
or I_30322 (I518539,I518522,I342351);
DFFARX1 I_30323 (I518539,I3035,I518095,I518565,);
nor I_30324 (I518075,I518565,I518121);
not I_30325 (I518587,I518565);
and I_30326 (I518604,I518587,I518121);
nor I_30327 (I518069,I518146,I518604);
nand I_30328 (I518635,I518587,I518197);
nor I_30329 (I518063,I518457,I518635);
nand I_30330 (I518066,I518587,I518375);
nand I_30331 (I518680,I518197,I342360);
nor I_30332 (I518078,I518440,I518680);
not I_30333 (I518741,I3042);
DFFARX1 I_30334 (I197729,I3035,I518741,I518767,);
DFFARX1 I_30335 (I197735,I3035,I518741,I518784,);
not I_30336 (I518792,I518784);
not I_30337 (I518809,I197756);
nor I_30338 (I518826,I518809,I197744);
not I_30339 (I518843,I197753);
nor I_30340 (I518860,I518826,I197738);
nor I_30341 (I518877,I518784,I518860);
DFFARX1 I_30342 (I518877,I3035,I518741,I518727,);
nor I_30343 (I518908,I197738,I197744);
nand I_30344 (I518925,I518908,I197756);
DFFARX1 I_30345 (I518925,I3035,I518741,I518730,);
nor I_30346 (I518956,I518843,I197738);
nand I_30347 (I518973,I518956,I197729);
nor I_30348 (I518990,I518767,I518973);
DFFARX1 I_30349 (I518990,I3035,I518741,I518706,);
not I_30350 (I519021,I518973);
nand I_30351 (I518718,I518784,I519021);
DFFARX1 I_30352 (I518973,I3035,I518741,I519061,);
not I_30353 (I519069,I519061);
not I_30354 (I519086,I197738);
not I_30355 (I519103,I197741);
nor I_30356 (I519120,I519103,I197753);
nor I_30357 (I518733,I519069,I519120);
nor I_30358 (I519151,I519103,I197750);
and I_30359 (I519168,I519151,I197732);
or I_30360 (I519185,I519168,I197747);
DFFARX1 I_30361 (I519185,I3035,I518741,I519211,);
nor I_30362 (I518721,I519211,I518767);
not I_30363 (I519233,I519211);
and I_30364 (I519250,I519233,I518767);
nor I_30365 (I518715,I518792,I519250);
nand I_30366 (I519281,I519233,I518843);
nor I_30367 (I518709,I519103,I519281);
nand I_30368 (I518712,I519233,I519021);
nand I_30369 (I519326,I518843,I197741);
nor I_30370 (I518724,I519086,I519326);
not I_30371 (I519387,I3042);
DFFARX1 I_30372 (I269611,I3035,I519387,I519413,);
DFFARX1 I_30373 (I269608,I3035,I519387,I519430,);
not I_30374 (I519438,I519430);
not I_30375 (I519455,I269623);
nor I_30376 (I519472,I519455,I269626);
not I_30377 (I519489,I269614);
nor I_30378 (I519506,I519472,I269620);
nor I_30379 (I519523,I519430,I519506);
DFFARX1 I_30380 (I519523,I3035,I519387,I519373,);
nor I_30381 (I519554,I269620,I269626);
nand I_30382 (I519571,I519554,I269623);
DFFARX1 I_30383 (I519571,I3035,I519387,I519376,);
nor I_30384 (I519602,I519489,I269620);
nand I_30385 (I519619,I519602,I269632);
nor I_30386 (I519636,I519413,I519619);
DFFARX1 I_30387 (I519636,I3035,I519387,I519352,);
not I_30388 (I519667,I519619);
nand I_30389 (I519364,I519430,I519667);
DFFARX1 I_30390 (I519619,I3035,I519387,I519707,);
not I_30391 (I519715,I519707);
not I_30392 (I519732,I269620);
not I_30393 (I519749,I269605);
nor I_30394 (I519766,I519749,I269614);
nor I_30395 (I519379,I519715,I519766);
nor I_30396 (I519797,I519749,I269617);
and I_30397 (I519814,I519797,I269605);
or I_30398 (I519831,I519814,I269629);
DFFARX1 I_30399 (I519831,I3035,I519387,I519857,);
nor I_30400 (I519367,I519857,I519413);
not I_30401 (I519879,I519857);
and I_30402 (I519896,I519879,I519413);
nor I_30403 (I519361,I519438,I519896);
nand I_30404 (I519927,I519879,I519489);
nor I_30405 (I519355,I519749,I519927);
nand I_30406 (I519358,I519879,I519667);
nand I_30407 (I519972,I519489,I269605);
nor I_30408 (I519370,I519732,I519972);
not I_30409 (I520033,I3042);
DFFARX1 I_30410 (I28885,I3035,I520033,I520059,);
DFFARX1 I_30411 (I28891,I3035,I520033,I520076,);
not I_30412 (I520084,I520076);
not I_30413 (I520101,I28909);
nor I_30414 (I520118,I520101,I28888);
not I_30415 (I520135,I28894);
nor I_30416 (I520152,I520118,I28900);
nor I_30417 (I520169,I520076,I520152);
DFFARX1 I_30418 (I520169,I3035,I520033,I520019,);
nor I_30419 (I520200,I28900,I28888);
nand I_30420 (I520217,I520200,I28909);
DFFARX1 I_30421 (I520217,I3035,I520033,I520022,);
nor I_30422 (I520248,I520135,I28900);
nand I_30423 (I520265,I520248,I28906);
nor I_30424 (I520282,I520059,I520265);
DFFARX1 I_30425 (I520282,I3035,I520033,I519998,);
not I_30426 (I520313,I520265);
nand I_30427 (I520010,I520076,I520313);
DFFARX1 I_30428 (I520265,I3035,I520033,I520353,);
not I_30429 (I520361,I520353);
not I_30430 (I520378,I28900);
not I_30431 (I520395,I28888);
nor I_30432 (I520412,I520395,I28894);
nor I_30433 (I520025,I520361,I520412);
nor I_30434 (I520443,I520395,I28897);
and I_30435 (I520460,I520443,I28885);
or I_30436 (I520477,I520460,I28903);
DFFARX1 I_30437 (I520477,I3035,I520033,I520503,);
nor I_30438 (I520013,I520503,I520059);
not I_30439 (I520525,I520503);
and I_30440 (I520542,I520525,I520059);
nor I_30441 (I520007,I520084,I520542);
nand I_30442 (I520573,I520525,I520135);
nor I_30443 (I520001,I520395,I520573);
nand I_30444 (I520004,I520525,I520313);
nand I_30445 (I520618,I520135,I28888);
nor I_30446 (I520016,I520378,I520618);
not I_30447 (I520679,I3042);
DFFARX1 I_30448 (I8332,I3035,I520679,I520705,);
DFFARX1 I_30449 (I8338,I3035,I520679,I520722,);
not I_30450 (I520730,I520722);
not I_30451 (I520747,I8332);
nor I_30452 (I520764,I520747,I8344);
not I_30453 (I520781,I8356);
nor I_30454 (I520798,I520764,I8350);
nor I_30455 (I520815,I520722,I520798);
DFFARX1 I_30456 (I520815,I3035,I520679,I520665,);
nor I_30457 (I520846,I8350,I8344);
nand I_30458 (I520863,I520846,I8332);
DFFARX1 I_30459 (I520863,I3035,I520679,I520668,);
nor I_30460 (I520894,I520781,I8350);
nand I_30461 (I520911,I520894,I8335);
nor I_30462 (I520928,I520705,I520911);
DFFARX1 I_30463 (I520928,I3035,I520679,I520644,);
not I_30464 (I520959,I520911);
nand I_30465 (I520656,I520722,I520959);
DFFARX1 I_30466 (I520911,I3035,I520679,I520999,);
not I_30467 (I521007,I520999);
not I_30468 (I521024,I8350);
not I_30469 (I521041,I8335);
nor I_30470 (I521058,I521041,I8356);
nor I_30471 (I520671,I521007,I521058);
nor I_30472 (I521089,I521041,I8353);
and I_30473 (I521106,I521089,I8347);
or I_30474 (I521123,I521106,I8341);
DFFARX1 I_30475 (I521123,I3035,I520679,I521149,);
nor I_30476 (I520659,I521149,I520705);
not I_30477 (I521171,I521149);
and I_30478 (I521188,I521171,I520705);
nor I_30479 (I520653,I520730,I521188);
nand I_30480 (I521219,I521171,I520781);
nor I_30481 (I520647,I521041,I521219);
nand I_30482 (I520650,I521171,I520959);
nand I_30483 (I521264,I520781,I8335);
nor I_30484 (I520662,I521024,I521264);
not I_30485 (I521325,I3042);
DFFARX1 I_30486 (I611034,I3035,I521325,I521351,);
DFFARX1 I_30487 (I611016,I3035,I521325,I521368,);
not I_30488 (I521376,I521368);
not I_30489 (I521393,I611025);
nor I_30490 (I521410,I521393,I611037);
not I_30491 (I521427,I611019);
nor I_30492 (I521444,I521410,I611028);
nor I_30493 (I521461,I521368,I521444);
DFFARX1 I_30494 (I521461,I3035,I521325,I521311,);
nor I_30495 (I521492,I611028,I611037);
nand I_30496 (I521509,I521492,I611025);
DFFARX1 I_30497 (I521509,I3035,I521325,I521314,);
nor I_30498 (I521540,I521427,I611028);
nand I_30499 (I521557,I521540,I611040);
nor I_30500 (I521574,I521351,I521557);
DFFARX1 I_30501 (I521574,I3035,I521325,I521290,);
not I_30502 (I521605,I521557);
nand I_30503 (I521302,I521368,I521605);
DFFARX1 I_30504 (I521557,I3035,I521325,I521645,);
not I_30505 (I521653,I521645);
not I_30506 (I521670,I611028);
not I_30507 (I521687,I611016);
nor I_30508 (I521704,I521687,I611019);
nor I_30509 (I521317,I521653,I521704);
nor I_30510 (I521735,I521687,I611022);
and I_30511 (I521752,I521735,I611031);
or I_30512 (I521769,I521752,I611019);
DFFARX1 I_30513 (I521769,I3035,I521325,I521795,);
nor I_30514 (I521305,I521795,I521351);
not I_30515 (I521817,I521795);
and I_30516 (I521834,I521817,I521351);
nor I_30517 (I521299,I521376,I521834);
nand I_30518 (I521865,I521817,I521427);
nor I_30519 (I521293,I521687,I521865);
nand I_30520 (I521296,I521817,I521605);
nand I_30521 (I521910,I521427,I611016);
nor I_30522 (I521308,I521670,I521910);
not I_30523 (I521971,I3042);
DFFARX1 I_30524 (I131860,I3035,I521971,I521997,);
DFFARX1 I_30525 (I131872,I3035,I521971,I522014,);
not I_30526 (I522022,I522014);
not I_30527 (I522039,I131878);
nor I_30528 (I522056,I522039,I131863);
not I_30529 (I522073,I131854);
nor I_30530 (I522090,I522056,I131875);
nor I_30531 (I522107,I522014,I522090);
DFFARX1 I_30532 (I522107,I3035,I521971,I521957,);
nor I_30533 (I522138,I131875,I131863);
nand I_30534 (I522155,I522138,I131878);
DFFARX1 I_30535 (I522155,I3035,I521971,I521960,);
nor I_30536 (I522186,I522073,I131875);
nand I_30537 (I522203,I522186,I131857);
nor I_30538 (I522220,I521997,I522203);
DFFARX1 I_30539 (I522220,I3035,I521971,I521936,);
not I_30540 (I522251,I522203);
nand I_30541 (I521948,I522014,I522251);
DFFARX1 I_30542 (I522203,I3035,I521971,I522291,);
not I_30543 (I522299,I522291);
not I_30544 (I522316,I131875);
not I_30545 (I522333,I131866);
nor I_30546 (I522350,I522333,I131854);
nor I_30547 (I521963,I522299,I522350);
nor I_30548 (I522381,I522333,I131869);
and I_30549 (I522398,I522381,I131857);
or I_30550 (I522415,I522398,I131854);
DFFARX1 I_30551 (I522415,I3035,I521971,I522441,);
nor I_30552 (I521951,I522441,I521997);
not I_30553 (I522463,I522441);
and I_30554 (I522480,I522463,I521997);
nor I_30555 (I521945,I522022,I522480);
nand I_30556 (I522511,I522463,I522073);
nor I_30557 (I521939,I522333,I522511);
nand I_30558 (I521942,I522463,I522251);
nand I_30559 (I522556,I522073,I131866);
nor I_30560 (I521954,I522316,I522556);
not I_30561 (I522617,I3042);
DFFARX1 I_30562 (I577510,I3035,I522617,I522643,);
DFFARX1 I_30563 (I577492,I3035,I522617,I522660,);
not I_30564 (I522668,I522660);
not I_30565 (I522685,I577501);
nor I_30566 (I522702,I522685,I577513);
not I_30567 (I522719,I577495);
nor I_30568 (I522736,I522702,I577504);
nor I_30569 (I522753,I522660,I522736);
DFFARX1 I_30570 (I522753,I3035,I522617,I522603,);
nor I_30571 (I522784,I577504,I577513);
nand I_30572 (I522801,I522784,I577501);
DFFARX1 I_30573 (I522801,I3035,I522617,I522606,);
nor I_30574 (I522832,I522719,I577504);
nand I_30575 (I522849,I522832,I577516);
nor I_30576 (I522866,I522643,I522849);
DFFARX1 I_30577 (I522866,I3035,I522617,I522582,);
not I_30578 (I522897,I522849);
nand I_30579 (I522594,I522660,I522897);
DFFARX1 I_30580 (I522849,I3035,I522617,I522937,);
not I_30581 (I522945,I522937);
not I_30582 (I522962,I577504);
not I_30583 (I522979,I577492);
nor I_30584 (I522996,I522979,I577495);
nor I_30585 (I522609,I522945,I522996);
nor I_30586 (I523027,I522979,I577498);
and I_30587 (I523044,I523027,I577507);
or I_30588 (I523061,I523044,I577495);
DFFARX1 I_30589 (I523061,I3035,I522617,I523087,);
nor I_30590 (I522597,I523087,I522643);
not I_30591 (I523109,I523087);
and I_30592 (I523126,I523109,I522643);
nor I_30593 (I522591,I522668,I523126);
nand I_30594 (I523157,I523109,I522719);
nor I_30595 (I522585,I522979,I523157);
nand I_30596 (I522588,I523109,I522897);
nand I_30597 (I523202,I522719,I577492);
nor I_30598 (I522600,I522962,I523202);
not I_30599 (I523263,I3042);
DFFARX1 I_30600 (I439305,I3035,I523263,I523289,);
DFFARX1 I_30601 (I439302,I3035,I523263,I523306,);
not I_30602 (I523314,I523306);
not I_30603 (I523331,I439302);
nor I_30604 (I523348,I523331,I439305);
not I_30605 (I523365,I439317);
nor I_30606 (I523382,I523348,I439311);
nor I_30607 (I523399,I523306,I523382);
DFFARX1 I_30608 (I523399,I3035,I523263,I523249,);
nor I_30609 (I523430,I439311,I439305);
nand I_30610 (I523447,I523430,I439302);
DFFARX1 I_30611 (I523447,I3035,I523263,I523252,);
nor I_30612 (I523478,I523365,I439311);
nand I_30613 (I523495,I523478,I439299);
nor I_30614 (I523512,I523289,I523495);
DFFARX1 I_30615 (I523512,I3035,I523263,I523228,);
not I_30616 (I523543,I523495);
nand I_30617 (I523240,I523306,I523543);
DFFARX1 I_30618 (I523495,I3035,I523263,I523583,);
not I_30619 (I523591,I523583);
not I_30620 (I523608,I439311);
not I_30621 (I523625,I439308);
nor I_30622 (I523642,I523625,I439317);
nor I_30623 (I523255,I523591,I523642);
nor I_30624 (I523673,I523625,I439314);
and I_30625 (I523690,I523673,I439320);
or I_30626 (I523707,I523690,I439299);
DFFARX1 I_30627 (I523707,I3035,I523263,I523733,);
nor I_30628 (I523243,I523733,I523289);
not I_30629 (I523755,I523733);
and I_30630 (I523772,I523755,I523289);
nor I_30631 (I523237,I523314,I523772);
nand I_30632 (I523803,I523755,I523365);
nor I_30633 (I523231,I523625,I523803);
nand I_30634 (I523234,I523755,I523543);
nand I_30635 (I523848,I523365,I439308);
nor I_30636 (I523246,I523608,I523848);
not I_30637 (I523909,I3042);
DFFARX1 I_30638 (I110440,I3035,I523909,I523935,);
DFFARX1 I_30639 (I110452,I3035,I523909,I523952,);
not I_30640 (I523960,I523952);
not I_30641 (I523977,I110458);
nor I_30642 (I523994,I523977,I110443);
not I_30643 (I524011,I110434);
nor I_30644 (I524028,I523994,I110455);
nor I_30645 (I524045,I523952,I524028);
DFFARX1 I_30646 (I524045,I3035,I523909,I523895,);
nor I_30647 (I524076,I110455,I110443);
nand I_30648 (I524093,I524076,I110458);
DFFARX1 I_30649 (I524093,I3035,I523909,I523898,);
nor I_30650 (I524124,I524011,I110455);
nand I_30651 (I524141,I524124,I110437);
nor I_30652 (I524158,I523935,I524141);
DFFARX1 I_30653 (I524158,I3035,I523909,I523874,);
not I_30654 (I524189,I524141);
nand I_30655 (I523886,I523952,I524189);
DFFARX1 I_30656 (I524141,I3035,I523909,I524229,);
not I_30657 (I524237,I524229);
not I_30658 (I524254,I110455);
not I_30659 (I524271,I110446);
nor I_30660 (I524288,I524271,I110434);
nor I_30661 (I523901,I524237,I524288);
nor I_30662 (I524319,I524271,I110449);
and I_30663 (I524336,I524319,I110437);
or I_30664 (I524353,I524336,I110434);
DFFARX1 I_30665 (I524353,I3035,I523909,I524379,);
nor I_30666 (I523889,I524379,I523935);
not I_30667 (I524401,I524379);
and I_30668 (I524418,I524401,I523935);
nor I_30669 (I523883,I523960,I524418);
nand I_30670 (I524449,I524401,I524011);
nor I_30671 (I523877,I524271,I524449);
nand I_30672 (I523880,I524401,I524189);
nand I_30673 (I524494,I524011,I110446);
nor I_30674 (I523892,I524254,I524494);
not I_30675 (I524555,I3042);
DFFARX1 I_30676 (I391484,I3035,I524555,I524581,);
DFFARX1 I_30677 (I391478,I3035,I524555,I524598,);
not I_30678 (I524606,I524598);
not I_30679 (I524623,I391493);
nor I_30680 (I524640,I524623,I391478);
not I_30681 (I524657,I391487);
nor I_30682 (I524674,I524640,I391496);
nor I_30683 (I524691,I524598,I524674);
DFFARX1 I_30684 (I524691,I3035,I524555,I524541,);
nor I_30685 (I524722,I391496,I391478);
nand I_30686 (I524739,I524722,I391493);
DFFARX1 I_30687 (I524739,I3035,I524555,I524544,);
nor I_30688 (I524770,I524657,I391496);
nand I_30689 (I524787,I524770,I391481);
nor I_30690 (I524804,I524581,I524787);
DFFARX1 I_30691 (I524804,I3035,I524555,I524520,);
not I_30692 (I524835,I524787);
nand I_30693 (I524532,I524598,I524835);
DFFARX1 I_30694 (I524787,I3035,I524555,I524875,);
not I_30695 (I524883,I524875);
not I_30696 (I524900,I391496);
not I_30697 (I524917,I391490);
nor I_30698 (I524934,I524917,I391487);
nor I_30699 (I524547,I524883,I524934);
nor I_30700 (I524965,I524917,I391499);
and I_30701 (I524982,I524965,I391502);
or I_30702 (I524999,I524982,I391481);
DFFARX1 I_30703 (I524999,I3035,I524555,I525025,);
nor I_30704 (I524535,I525025,I524581);
not I_30705 (I525047,I525025);
and I_30706 (I525064,I525047,I524581);
nor I_30707 (I524529,I524606,I525064);
nand I_30708 (I525095,I525047,I524657);
nor I_30709 (I524523,I524917,I525095);
nand I_30710 (I524526,I525047,I524835);
nand I_30711 (I525140,I524657,I391490);
nor I_30712 (I524538,I524900,I525140);
not I_30713 (I525201,I3042);
DFFARX1 I_30714 (I614502,I3035,I525201,I525227,);
DFFARX1 I_30715 (I614484,I3035,I525201,I525244,);
not I_30716 (I525252,I525244);
not I_30717 (I525269,I614493);
nor I_30718 (I525286,I525269,I614505);
not I_30719 (I525303,I614487);
nor I_30720 (I525320,I525286,I614496);
nor I_30721 (I525337,I525244,I525320);
DFFARX1 I_30722 (I525337,I3035,I525201,I525187,);
nor I_30723 (I525368,I614496,I614505);
nand I_30724 (I525385,I525368,I614493);
DFFARX1 I_30725 (I525385,I3035,I525201,I525190,);
nor I_30726 (I525416,I525303,I614496);
nand I_30727 (I525433,I525416,I614508);
nor I_30728 (I525450,I525227,I525433);
DFFARX1 I_30729 (I525450,I3035,I525201,I525166,);
not I_30730 (I525481,I525433);
nand I_30731 (I525178,I525244,I525481);
DFFARX1 I_30732 (I525433,I3035,I525201,I525521,);
not I_30733 (I525529,I525521);
not I_30734 (I525546,I614496);
not I_30735 (I525563,I614484);
nor I_30736 (I525580,I525563,I614487);
nor I_30737 (I525193,I525529,I525580);
nor I_30738 (I525611,I525563,I614490);
and I_30739 (I525628,I525611,I614499);
or I_30740 (I525645,I525628,I614487);
DFFARX1 I_30741 (I525645,I3035,I525201,I525671,);
nor I_30742 (I525181,I525671,I525227);
not I_30743 (I525693,I525671);
and I_30744 (I525710,I525693,I525227);
nor I_30745 (I525175,I525252,I525710);
nand I_30746 (I525741,I525693,I525303);
nor I_30747 (I525169,I525563,I525741);
nand I_30748 (I525172,I525693,I525481);
nand I_30749 (I525786,I525303,I614484);
nor I_30750 (I525184,I525546,I525786);
not I_30751 (I525847,I3042);
DFFARX1 I_30752 (I94970,I3035,I525847,I525873,);
DFFARX1 I_30753 (I94982,I3035,I525847,I525890,);
not I_30754 (I525898,I525890);
not I_30755 (I525915,I94988);
nor I_30756 (I525932,I525915,I94973);
not I_30757 (I525949,I94964);
nor I_30758 (I525966,I525932,I94985);
nor I_30759 (I525983,I525890,I525966);
DFFARX1 I_30760 (I525983,I3035,I525847,I525833,);
nor I_30761 (I526014,I94985,I94973);
nand I_30762 (I526031,I526014,I94988);
DFFARX1 I_30763 (I526031,I3035,I525847,I525836,);
nor I_30764 (I526062,I525949,I94985);
nand I_30765 (I526079,I526062,I94967);
nor I_30766 (I526096,I525873,I526079);
DFFARX1 I_30767 (I526096,I3035,I525847,I525812,);
not I_30768 (I526127,I526079);
nand I_30769 (I525824,I525890,I526127);
DFFARX1 I_30770 (I526079,I3035,I525847,I526167,);
not I_30771 (I526175,I526167);
not I_30772 (I526192,I94985);
not I_30773 (I526209,I94976);
nor I_30774 (I526226,I526209,I94964);
nor I_30775 (I525839,I526175,I526226);
nor I_30776 (I526257,I526209,I94979);
and I_30777 (I526274,I526257,I94967);
or I_30778 (I526291,I526274,I94964);
DFFARX1 I_30779 (I526291,I3035,I525847,I526317,);
nor I_30780 (I525827,I526317,I525873);
not I_30781 (I526339,I526317);
and I_30782 (I526356,I526339,I525873);
nor I_30783 (I525821,I525898,I526356);
nand I_30784 (I526387,I526339,I525949);
nor I_30785 (I525815,I526209,I526387);
nand I_30786 (I525818,I526339,I526127);
nand I_30787 (I526432,I525949,I94976);
nor I_30788 (I525830,I526192,I526432);
not I_30789 (I526493,I3042);
DFFARX1 I_30790 (I694433,I3035,I526493,I526519,);
DFFARX1 I_30791 (I694430,I3035,I526493,I526536,);
not I_30792 (I526544,I526536);
not I_30793 (I526561,I694427);
nor I_30794 (I526578,I526561,I694418);
not I_30795 (I526595,I694439);
nor I_30796 (I526612,I526578,I694418);
nor I_30797 (I526629,I526536,I526612);
DFFARX1 I_30798 (I526629,I3035,I526493,I526479,);
nor I_30799 (I526660,I694418,I694418);
nand I_30800 (I526677,I526660,I694427);
DFFARX1 I_30801 (I526677,I3035,I526493,I526482,);
nor I_30802 (I526708,I526595,I694418);
nand I_30803 (I526725,I526708,I694442);
nor I_30804 (I526742,I526519,I526725);
DFFARX1 I_30805 (I526742,I3035,I526493,I526458,);
not I_30806 (I526773,I526725);
nand I_30807 (I526470,I526536,I526773);
DFFARX1 I_30808 (I526725,I3035,I526493,I526813,);
not I_30809 (I526821,I526813);
not I_30810 (I526838,I694418);
not I_30811 (I526855,I694421);
nor I_30812 (I526872,I526855,I694439);
nor I_30813 (I526485,I526821,I526872);
nor I_30814 (I526903,I526855,I694424);
and I_30815 (I526920,I526903,I694445);
or I_30816 (I526937,I526920,I694436);
DFFARX1 I_30817 (I526937,I3035,I526493,I526963,);
nor I_30818 (I526473,I526963,I526519);
not I_30819 (I526985,I526963);
and I_30820 (I527002,I526985,I526519);
nor I_30821 (I526467,I526544,I527002);
nand I_30822 (I527033,I526985,I526595);
nor I_30823 (I526461,I526855,I527033);
nand I_30824 (I526464,I526985,I526773);
nand I_30825 (I527078,I526595,I694421);
nor I_30826 (I526476,I526838,I527078);
not I_30827 (I527139,I3042);
DFFARX1 I_30828 (I1788,I3035,I527139,I527165,);
DFFARX1 I_30829 (I2180,I3035,I527139,I527182,);
not I_30830 (I527190,I527182);
not I_30831 (I527207,I2308);
nor I_30832 (I527224,I527207,I2244);
not I_30833 (I527241,I2004);
nor I_30834 (I527258,I527224,I2348);
nor I_30835 (I527275,I527182,I527258);
DFFARX1 I_30836 (I527275,I3035,I527139,I527125,);
nor I_30837 (I527306,I2348,I2244);
nand I_30838 (I527323,I527306,I2308);
DFFARX1 I_30839 (I527323,I3035,I527139,I527128,);
nor I_30840 (I527354,I527241,I2348);
nand I_30841 (I527371,I527354,I1692);
nor I_30842 (I527388,I527165,I527371);
DFFARX1 I_30843 (I527388,I3035,I527139,I527104,);
not I_30844 (I527419,I527371);
nand I_30845 (I527116,I527182,I527419);
DFFARX1 I_30846 (I527371,I3035,I527139,I527459,);
not I_30847 (I527467,I527459);
not I_30848 (I527484,I2348);
not I_30849 (I527501,I1796);
nor I_30850 (I527518,I527501,I2004);
nor I_30851 (I527131,I527467,I527518);
nor I_30852 (I527549,I527501,I2852);
and I_30853 (I527566,I527549,I2372);
or I_30854 (I527583,I527566,I1812);
DFFARX1 I_30855 (I527583,I3035,I527139,I527609,);
nor I_30856 (I527119,I527609,I527165);
not I_30857 (I527631,I527609);
and I_30858 (I527648,I527631,I527165);
nor I_30859 (I527113,I527190,I527648);
nand I_30860 (I527679,I527631,I527241);
nor I_30861 (I527107,I527501,I527679);
nand I_30862 (I527110,I527631,I527419);
nand I_30863 (I527724,I527241,I1796);
nor I_30864 (I527122,I527484,I527724);
not I_30865 (I527785,I3042);
DFFARX1 I_30866 (I58397,I3035,I527785,I527811,);
DFFARX1 I_30867 (I58403,I3035,I527785,I527828,);
not I_30868 (I527836,I527828);
not I_30869 (I527853,I58421);
nor I_30870 (I527870,I527853,I58400);
not I_30871 (I527887,I58406);
nor I_30872 (I527904,I527870,I58412);
nor I_30873 (I527921,I527828,I527904);
DFFARX1 I_30874 (I527921,I3035,I527785,I527771,);
nor I_30875 (I527952,I58412,I58400);
nand I_30876 (I527969,I527952,I58421);
DFFARX1 I_30877 (I527969,I3035,I527785,I527774,);
nor I_30878 (I528000,I527887,I58412);
nand I_30879 (I528017,I528000,I58418);
nor I_30880 (I528034,I527811,I528017);
DFFARX1 I_30881 (I528034,I3035,I527785,I527750,);
not I_30882 (I528065,I528017);
nand I_30883 (I527762,I527828,I528065);
DFFARX1 I_30884 (I528017,I3035,I527785,I528105,);
not I_30885 (I528113,I528105);
not I_30886 (I528130,I58412);
not I_30887 (I528147,I58400);
nor I_30888 (I528164,I528147,I58406);
nor I_30889 (I527777,I528113,I528164);
nor I_30890 (I528195,I528147,I58409);
and I_30891 (I528212,I528195,I58397);
or I_30892 (I528229,I528212,I58415);
DFFARX1 I_30893 (I528229,I3035,I527785,I528255,);
nor I_30894 (I527765,I528255,I527811);
not I_30895 (I528277,I528255);
and I_30896 (I528294,I528277,I527811);
nor I_30897 (I527759,I527836,I528294);
nand I_30898 (I528325,I528277,I527887);
nor I_30899 (I527753,I528147,I528325);
nand I_30900 (I527756,I528277,I528065);
nand I_30901 (I528370,I527887,I58400);
nor I_30902 (I527768,I528130,I528370);
not I_30903 (I528431,I3042);
DFFARX1 I_30904 (I186662,I3035,I528431,I528457,);
DFFARX1 I_30905 (I186668,I3035,I528431,I528474,);
not I_30906 (I528482,I528474);
not I_30907 (I528499,I186689);
nor I_30908 (I528516,I528499,I186677);
not I_30909 (I528533,I186686);
nor I_30910 (I528550,I528516,I186671);
nor I_30911 (I528567,I528474,I528550);
DFFARX1 I_30912 (I528567,I3035,I528431,I528417,);
nor I_30913 (I528598,I186671,I186677);
nand I_30914 (I528615,I528598,I186689);
DFFARX1 I_30915 (I528615,I3035,I528431,I528420,);
nor I_30916 (I528646,I528533,I186671);
nand I_30917 (I528663,I528646,I186662);
nor I_30918 (I528680,I528457,I528663);
DFFARX1 I_30919 (I528680,I3035,I528431,I528396,);
not I_30920 (I528711,I528663);
nand I_30921 (I528408,I528474,I528711);
DFFARX1 I_30922 (I528663,I3035,I528431,I528751,);
not I_30923 (I528759,I528751);
not I_30924 (I528776,I186671);
not I_30925 (I528793,I186674);
nor I_30926 (I528810,I528793,I186686);
nor I_30927 (I528423,I528759,I528810);
nor I_30928 (I528841,I528793,I186683);
and I_30929 (I528858,I528841,I186665);
or I_30930 (I528875,I528858,I186680);
DFFARX1 I_30931 (I528875,I3035,I528431,I528901,);
nor I_30932 (I528411,I528901,I528457);
not I_30933 (I528923,I528901);
and I_30934 (I528940,I528923,I528457);
nor I_30935 (I528405,I528482,I528940);
nand I_30936 (I528971,I528923,I528533);
nor I_30937 (I528399,I528793,I528971);
nand I_30938 (I528402,I528923,I528711);
nand I_30939 (I529016,I528533,I186674);
nor I_30940 (I528414,I528776,I529016);
not I_30941 (I529077,I3042);
DFFARX1 I_30942 (I427184,I3035,I529077,I529103,);
DFFARX1 I_30943 (I427181,I3035,I529077,I529120,);
not I_30944 (I529128,I529120);
not I_30945 (I529145,I427181);
nor I_30946 (I529162,I529145,I427184);
not I_30947 (I529179,I427196);
nor I_30948 (I529196,I529162,I427190);
nor I_30949 (I529213,I529120,I529196);
DFFARX1 I_30950 (I529213,I3035,I529077,I529063,);
nor I_30951 (I529244,I427190,I427184);
nand I_30952 (I529261,I529244,I427181);
DFFARX1 I_30953 (I529261,I3035,I529077,I529066,);
nor I_30954 (I529292,I529179,I427190);
nand I_30955 (I529309,I529292,I427178);
nor I_30956 (I529326,I529103,I529309);
DFFARX1 I_30957 (I529326,I3035,I529077,I529042,);
not I_30958 (I529357,I529309);
nand I_30959 (I529054,I529120,I529357);
DFFARX1 I_30960 (I529309,I3035,I529077,I529397,);
not I_30961 (I529405,I529397);
not I_30962 (I529422,I427190);
not I_30963 (I529439,I427187);
nor I_30964 (I529456,I529439,I427196);
nor I_30965 (I529069,I529405,I529456);
nor I_30966 (I529487,I529439,I427193);
and I_30967 (I529504,I529487,I427199);
or I_30968 (I529521,I529504,I427178);
DFFARX1 I_30969 (I529521,I3035,I529077,I529547,);
nor I_30970 (I529057,I529547,I529103);
not I_30971 (I529569,I529547);
and I_30972 (I529586,I529569,I529103);
nor I_30973 (I529051,I529128,I529586);
nand I_30974 (I529617,I529569,I529179);
nor I_30975 (I529045,I529439,I529617);
nand I_30976 (I529048,I529569,I529357);
nand I_30977 (I529662,I529179,I427187);
nor I_30978 (I529060,I529422,I529662);
not I_30979 (I529723,I3042);
DFFARX1 I_30980 (I278859,I3035,I529723,I529749,);
DFFARX1 I_30981 (I278856,I3035,I529723,I529766,);
not I_30982 (I529774,I529766);
not I_30983 (I529791,I278871);
nor I_30984 (I529808,I529791,I278874);
not I_30985 (I529825,I278862);
nor I_30986 (I529842,I529808,I278868);
nor I_30987 (I529859,I529766,I529842);
DFFARX1 I_30988 (I529859,I3035,I529723,I529709,);
nor I_30989 (I529890,I278868,I278874);
nand I_30990 (I529907,I529890,I278871);
DFFARX1 I_30991 (I529907,I3035,I529723,I529712,);
nor I_30992 (I529938,I529825,I278868);
nand I_30993 (I529955,I529938,I278880);
nor I_30994 (I529972,I529749,I529955);
DFFARX1 I_30995 (I529972,I3035,I529723,I529688,);
not I_30996 (I530003,I529955);
nand I_30997 (I529700,I529766,I530003);
DFFARX1 I_30998 (I529955,I3035,I529723,I530043,);
not I_30999 (I530051,I530043);
not I_31000 (I530068,I278868);
not I_31001 (I530085,I278853);
nor I_31002 (I530102,I530085,I278862);
nor I_31003 (I529715,I530051,I530102);
nor I_31004 (I530133,I530085,I278865);
and I_31005 (I530150,I530133,I278853);
or I_31006 (I530167,I530150,I278877);
DFFARX1 I_31007 (I530167,I3035,I529723,I530193,);
nor I_31008 (I529703,I530193,I529749);
not I_31009 (I530215,I530193);
and I_31010 (I530232,I530215,I529749);
nor I_31011 (I529697,I529774,I530232);
nand I_31012 (I530263,I530215,I529825);
nor I_31013 (I529691,I530085,I530263);
nand I_31014 (I529694,I530215,I530003);
nand I_31015 (I530308,I529825,I278853);
nor I_31016 (I529706,I530068,I530308);
not I_31017 (I530369,I3042);
DFFARX1 I_31018 (I606988,I3035,I530369,I530395,);
DFFARX1 I_31019 (I606970,I3035,I530369,I530412,);
not I_31020 (I530420,I530412);
not I_31021 (I530437,I606979);
nor I_31022 (I530454,I530437,I606991);
not I_31023 (I530471,I606973);
nor I_31024 (I530488,I530454,I606982);
nor I_31025 (I530505,I530412,I530488);
DFFARX1 I_31026 (I530505,I3035,I530369,I530355,);
nor I_31027 (I530536,I606982,I606991);
nand I_31028 (I530553,I530536,I606979);
DFFARX1 I_31029 (I530553,I3035,I530369,I530358,);
nor I_31030 (I530584,I530471,I606982);
nand I_31031 (I530601,I530584,I606994);
nor I_31032 (I530618,I530395,I530601);
DFFARX1 I_31033 (I530618,I3035,I530369,I530334,);
not I_31034 (I530649,I530601);
nand I_31035 (I530346,I530412,I530649);
DFFARX1 I_31036 (I530601,I3035,I530369,I530689,);
not I_31037 (I530697,I530689);
not I_31038 (I530714,I606982);
not I_31039 (I530731,I606970);
nor I_31040 (I530748,I530731,I606973);
nor I_31041 (I530361,I530697,I530748);
nor I_31042 (I530779,I530731,I606976);
and I_31043 (I530796,I530779,I606985);
or I_31044 (I530813,I530796,I606973);
DFFARX1 I_31045 (I530813,I3035,I530369,I530839,);
nor I_31046 (I530349,I530839,I530395);
not I_31047 (I530861,I530839);
and I_31048 (I530878,I530861,I530395);
nor I_31049 (I530343,I530420,I530878);
nand I_31050 (I530909,I530861,I530471);
nor I_31051 (I530337,I530731,I530909);
nand I_31052 (I530340,I530861,I530649);
nand I_31053 (I530954,I530471,I606970);
nor I_31054 (I530352,I530714,I530954);
not I_31055 (I531015,I3042);
DFFARX1 I_31056 (I457223,I3035,I531015,I531041,);
DFFARX1 I_31057 (I457220,I3035,I531015,I531058,);
not I_31058 (I531066,I531058);
not I_31059 (I531083,I457220);
nor I_31060 (I531100,I531083,I457223);
not I_31061 (I531117,I457235);
nor I_31062 (I531134,I531100,I457229);
nor I_31063 (I531151,I531058,I531134);
DFFARX1 I_31064 (I531151,I3035,I531015,I531001,);
nor I_31065 (I531182,I457229,I457223);
nand I_31066 (I531199,I531182,I457220);
DFFARX1 I_31067 (I531199,I3035,I531015,I531004,);
nor I_31068 (I531230,I531117,I457229);
nand I_31069 (I531247,I531230,I457217);
nor I_31070 (I531264,I531041,I531247);
DFFARX1 I_31071 (I531264,I3035,I531015,I530980,);
not I_31072 (I531295,I531247);
nand I_31073 (I530992,I531058,I531295);
DFFARX1 I_31074 (I531247,I3035,I531015,I531335,);
not I_31075 (I531343,I531335);
not I_31076 (I531360,I457229);
not I_31077 (I531377,I457226);
nor I_31078 (I531394,I531377,I457235);
nor I_31079 (I531007,I531343,I531394);
nor I_31080 (I531425,I531377,I457232);
and I_31081 (I531442,I531425,I457238);
or I_31082 (I531459,I531442,I457217);
DFFARX1 I_31083 (I531459,I3035,I531015,I531485,);
nor I_31084 (I530995,I531485,I531041);
not I_31085 (I531507,I531485);
and I_31086 (I531524,I531507,I531041);
nor I_31087 (I530989,I531066,I531524);
nand I_31088 (I531555,I531507,I531117);
nor I_31089 (I530983,I531377,I531555);
nand I_31090 (I530986,I531507,I531295);
nand I_31091 (I531600,I531117,I457226);
nor I_31092 (I530998,I531360,I531600);
not I_31093 (I531661,I3042);
DFFARX1 I_31094 (I451953,I3035,I531661,I531687,);
DFFARX1 I_31095 (I451950,I3035,I531661,I531704,);
not I_31096 (I531712,I531704);
not I_31097 (I531729,I451950);
nor I_31098 (I531746,I531729,I451953);
not I_31099 (I531763,I451965);
nor I_31100 (I531780,I531746,I451959);
nor I_31101 (I531797,I531704,I531780);
DFFARX1 I_31102 (I531797,I3035,I531661,I531647,);
nor I_31103 (I531828,I451959,I451953);
nand I_31104 (I531845,I531828,I451950);
DFFARX1 I_31105 (I531845,I3035,I531661,I531650,);
nor I_31106 (I531876,I531763,I451959);
nand I_31107 (I531893,I531876,I451947);
nor I_31108 (I531910,I531687,I531893);
DFFARX1 I_31109 (I531910,I3035,I531661,I531626,);
not I_31110 (I531941,I531893);
nand I_31111 (I531638,I531704,I531941);
DFFARX1 I_31112 (I531893,I3035,I531661,I531981,);
not I_31113 (I531989,I531981);
not I_31114 (I532006,I451959);
not I_31115 (I532023,I451956);
nor I_31116 (I532040,I532023,I451965);
nor I_31117 (I531653,I531989,I532040);
nor I_31118 (I532071,I532023,I451962);
and I_31119 (I532088,I532071,I451968);
or I_31120 (I532105,I532088,I451947);
DFFARX1 I_31121 (I532105,I3035,I531661,I532131,);
nor I_31122 (I531641,I532131,I531687);
not I_31123 (I532153,I532131);
and I_31124 (I532170,I532153,I531687);
nor I_31125 (I531635,I531712,I532170);
nand I_31126 (I532201,I532153,I531763);
nor I_31127 (I531629,I532023,I532201);
nand I_31128 (I531632,I532153,I531941);
nand I_31129 (I532246,I531763,I451956);
nor I_31130 (I531644,I532006,I532246);
not I_31131 (I532307,I3042);
DFFARX1 I_31132 (I312295,I3035,I532307,I532333,);
DFFARX1 I_31133 (I312307,I3035,I532307,I532350,);
not I_31134 (I532358,I532350);
not I_31135 (I532375,I312316);
nor I_31136 (I532392,I532375,I312292);
not I_31137 (I532409,I312310);
nor I_31138 (I532426,I532392,I312304);
nor I_31139 (I532443,I532350,I532426);
DFFARX1 I_31140 (I532443,I3035,I532307,I532293,);
nor I_31141 (I532474,I312304,I312292);
nand I_31142 (I532491,I532474,I312316);
DFFARX1 I_31143 (I532491,I3035,I532307,I532296,);
nor I_31144 (I532522,I532409,I312304);
nand I_31145 (I532539,I532522,I312298);
nor I_31146 (I532556,I532333,I532539);
DFFARX1 I_31147 (I532556,I3035,I532307,I532272,);
not I_31148 (I532587,I532539);
nand I_31149 (I532284,I532350,I532587);
DFFARX1 I_31150 (I532539,I3035,I532307,I532627,);
not I_31151 (I532635,I532627);
not I_31152 (I532652,I312304);
not I_31153 (I532669,I312313);
nor I_31154 (I532686,I532669,I312310);
nor I_31155 (I532299,I532635,I532686);
nor I_31156 (I532717,I532669,I312295);
and I_31157 (I532734,I532717,I312292);
or I_31158 (I532751,I532734,I312301);
DFFARX1 I_31159 (I532751,I3035,I532307,I532777,);
nor I_31160 (I532287,I532777,I532333);
not I_31161 (I532799,I532777);
and I_31162 (I532816,I532799,I532333);
nor I_31163 (I532281,I532358,I532816);
nand I_31164 (I532847,I532799,I532409);
nor I_31165 (I532275,I532669,I532847);
nand I_31166 (I532278,I532799,I532587);
nand I_31167 (I532892,I532409,I312313);
nor I_31168 (I532290,I532652,I532892);
not I_31169 (I532953,I3042);
DFFARX1 I_31170 (I387438,I3035,I532953,I532979,);
DFFARX1 I_31171 (I387432,I3035,I532953,I532996,);
not I_31172 (I533004,I532996);
not I_31173 (I533021,I387447);
nor I_31174 (I533038,I533021,I387432);
not I_31175 (I533055,I387441);
nor I_31176 (I533072,I533038,I387450);
nor I_31177 (I533089,I532996,I533072);
DFFARX1 I_31178 (I533089,I3035,I532953,I532939,);
nor I_31179 (I533120,I387450,I387432);
nand I_31180 (I533137,I533120,I387447);
DFFARX1 I_31181 (I533137,I3035,I532953,I532942,);
nor I_31182 (I533168,I533055,I387450);
nand I_31183 (I533185,I533168,I387435);
nor I_31184 (I533202,I532979,I533185);
DFFARX1 I_31185 (I533202,I3035,I532953,I532918,);
not I_31186 (I533233,I533185);
nand I_31187 (I532930,I532996,I533233);
DFFARX1 I_31188 (I533185,I3035,I532953,I533273,);
not I_31189 (I533281,I533273);
not I_31190 (I533298,I387450);
not I_31191 (I533315,I387444);
nor I_31192 (I533332,I533315,I387441);
nor I_31193 (I532945,I533281,I533332);
nor I_31194 (I533363,I533315,I387453);
and I_31195 (I533380,I533363,I387456);
or I_31196 (I533397,I533380,I387435);
DFFARX1 I_31197 (I533397,I3035,I532953,I533423,);
nor I_31198 (I532933,I533423,I532979);
not I_31199 (I533445,I533423);
and I_31200 (I533462,I533445,I532979);
nor I_31201 (I532927,I533004,I533462);
nand I_31202 (I533493,I533445,I533055);
nor I_31203 (I532921,I533315,I533493);
nand I_31204 (I532924,I533445,I533233);
nand I_31205 (I533538,I533055,I387444);
nor I_31206 (I532936,I533298,I533538);
not I_31207 (I533599,I3042);
DFFARX1 I_31208 (I162420,I3035,I533599,I533625,);
DFFARX1 I_31209 (I162426,I3035,I533599,I533642,);
not I_31210 (I533650,I533642);
not I_31211 (I533667,I162447);
nor I_31212 (I533684,I533667,I162435);
not I_31213 (I533701,I162444);
nor I_31214 (I533718,I533684,I162429);
nor I_31215 (I533735,I533642,I533718);
DFFARX1 I_31216 (I533735,I3035,I533599,I533585,);
nor I_31217 (I533766,I162429,I162435);
nand I_31218 (I533783,I533766,I162447);
DFFARX1 I_31219 (I533783,I3035,I533599,I533588,);
nor I_31220 (I533814,I533701,I162429);
nand I_31221 (I533831,I533814,I162420);
nor I_31222 (I533848,I533625,I533831);
DFFARX1 I_31223 (I533848,I3035,I533599,I533564,);
not I_31224 (I533879,I533831);
nand I_31225 (I533576,I533642,I533879);
DFFARX1 I_31226 (I533831,I3035,I533599,I533919,);
not I_31227 (I533927,I533919);
not I_31228 (I533944,I162429);
not I_31229 (I533961,I162432);
nor I_31230 (I533978,I533961,I162444);
nor I_31231 (I533591,I533927,I533978);
nor I_31232 (I534009,I533961,I162441);
and I_31233 (I534026,I534009,I162423);
or I_31234 (I534043,I534026,I162438);
DFFARX1 I_31235 (I534043,I3035,I533599,I534069,);
nor I_31236 (I533579,I534069,I533625);
not I_31237 (I534091,I534069);
and I_31238 (I534108,I534091,I533625);
nor I_31239 (I533573,I533650,I534108);
nand I_31240 (I534139,I534091,I533701);
nor I_31241 (I533567,I533961,I534139);
nand I_31242 (I533570,I534091,I533879);
nand I_31243 (I534184,I533701,I162432);
nor I_31244 (I533582,I533944,I534184);
not I_31245 (I534245,I3042);
DFFARX1 I_31246 (I17291,I3035,I534245,I534271,);
DFFARX1 I_31247 (I17297,I3035,I534245,I534288,);
not I_31248 (I534296,I534288);
not I_31249 (I534313,I17291);
nor I_31250 (I534330,I534313,I17303);
not I_31251 (I534347,I17315);
nor I_31252 (I534364,I534330,I17309);
nor I_31253 (I534381,I534288,I534364);
DFFARX1 I_31254 (I534381,I3035,I534245,I534231,);
nor I_31255 (I534412,I17309,I17303);
nand I_31256 (I534429,I534412,I17291);
DFFARX1 I_31257 (I534429,I3035,I534245,I534234,);
nor I_31258 (I534460,I534347,I17309);
nand I_31259 (I534477,I534460,I17294);
nor I_31260 (I534494,I534271,I534477);
DFFARX1 I_31261 (I534494,I3035,I534245,I534210,);
not I_31262 (I534525,I534477);
nand I_31263 (I534222,I534288,I534525);
DFFARX1 I_31264 (I534477,I3035,I534245,I534565,);
not I_31265 (I534573,I534565);
not I_31266 (I534590,I17309);
not I_31267 (I534607,I17294);
nor I_31268 (I534624,I534607,I17315);
nor I_31269 (I534237,I534573,I534624);
nor I_31270 (I534655,I534607,I17312);
and I_31271 (I534672,I534655,I17306);
or I_31272 (I534689,I534672,I17300);
DFFARX1 I_31273 (I534689,I3035,I534245,I534715,);
nor I_31274 (I534225,I534715,I534271);
not I_31275 (I534737,I534715);
and I_31276 (I534754,I534737,I534271);
nor I_31277 (I534219,I534296,I534754);
nand I_31278 (I534785,I534737,I534347);
nor I_31279 (I534213,I534607,I534785);
nand I_31280 (I534216,I534737,I534525);
nand I_31281 (I534830,I534347,I17294);
nor I_31282 (I534228,I534590,I534830);
not I_31283 (I534891,I3042);
DFFARX1 I_31284 (I642246,I3035,I534891,I534917,);
DFFARX1 I_31285 (I642228,I3035,I534891,I534934,);
not I_31286 (I534942,I534934);
not I_31287 (I534959,I642237);
nor I_31288 (I534976,I534959,I642249);
not I_31289 (I534993,I642231);
nor I_31290 (I535010,I534976,I642240);
nor I_31291 (I535027,I534934,I535010);
DFFARX1 I_31292 (I535027,I3035,I534891,I534877,);
nor I_31293 (I535058,I642240,I642249);
nand I_31294 (I535075,I535058,I642237);
DFFARX1 I_31295 (I535075,I3035,I534891,I534880,);
nor I_31296 (I535106,I534993,I642240);
nand I_31297 (I535123,I535106,I642252);
nor I_31298 (I535140,I534917,I535123);
DFFARX1 I_31299 (I535140,I3035,I534891,I534856,);
not I_31300 (I535171,I535123);
nand I_31301 (I534868,I534934,I535171);
DFFARX1 I_31302 (I535123,I3035,I534891,I535211,);
not I_31303 (I535219,I535211);
not I_31304 (I535236,I642240);
not I_31305 (I535253,I642228);
nor I_31306 (I535270,I535253,I642231);
nor I_31307 (I534883,I535219,I535270);
nor I_31308 (I535301,I535253,I642234);
and I_31309 (I535318,I535301,I642243);
or I_31310 (I535335,I535318,I642231);
DFFARX1 I_31311 (I535335,I3035,I534891,I535361,);
nor I_31312 (I534871,I535361,I534917);
not I_31313 (I535383,I535361);
and I_31314 (I535400,I535383,I534917);
nor I_31315 (I534865,I534942,I535400);
nand I_31316 (I535431,I535383,I534993);
nor I_31317 (I534859,I535253,I535431);
nand I_31318 (I534862,I535383,I535171);
nand I_31319 (I535476,I534993,I642228);
nor I_31320 (I534874,I535236,I535476);
not I_31321 (I535537,I3042);
DFFARX1 I_31322 (I307093,I3035,I535537,I535563,);
DFFARX1 I_31323 (I307105,I3035,I535537,I535580,);
not I_31324 (I535588,I535580);
not I_31325 (I535605,I307114);
nor I_31326 (I535622,I535605,I307090);
not I_31327 (I535639,I307108);
nor I_31328 (I535656,I535622,I307102);
nor I_31329 (I535673,I535580,I535656);
DFFARX1 I_31330 (I535673,I3035,I535537,I535523,);
nor I_31331 (I535704,I307102,I307090);
nand I_31332 (I535721,I535704,I307114);
DFFARX1 I_31333 (I535721,I3035,I535537,I535526,);
nor I_31334 (I535752,I535639,I307102);
nand I_31335 (I535769,I535752,I307096);
nor I_31336 (I535786,I535563,I535769);
DFFARX1 I_31337 (I535786,I3035,I535537,I535502,);
not I_31338 (I535817,I535769);
nand I_31339 (I535514,I535580,I535817);
DFFARX1 I_31340 (I535769,I3035,I535537,I535857,);
not I_31341 (I535865,I535857);
not I_31342 (I535882,I307102);
not I_31343 (I535899,I307111);
nor I_31344 (I535916,I535899,I307108);
nor I_31345 (I535529,I535865,I535916);
nor I_31346 (I535947,I535899,I307093);
and I_31347 (I535964,I535947,I307090);
or I_31348 (I535981,I535964,I307099);
DFFARX1 I_31349 (I535981,I3035,I535537,I536007,);
nor I_31350 (I535517,I536007,I535563);
not I_31351 (I536029,I536007);
and I_31352 (I536046,I536029,I535563);
nor I_31353 (I535511,I535588,I536046);
nand I_31354 (I536077,I536029,I535639);
nor I_31355 (I535505,I535899,I536077);
nand I_31356 (I535508,I536029,I535817);
nand I_31357 (I536122,I535639,I307111);
nor I_31358 (I535520,I535882,I536122);
not I_31359 (I536183,I3042);
DFFARX1 I_31360 (I417494,I3035,I536183,I536209,);
DFFARX1 I_31361 (I417488,I3035,I536183,I536226,);
not I_31362 (I536234,I536226);
not I_31363 (I536251,I417503);
nor I_31364 (I536268,I536251,I417488);
not I_31365 (I536285,I417497);
nor I_31366 (I536302,I536268,I417506);
nor I_31367 (I536319,I536226,I536302);
DFFARX1 I_31368 (I536319,I3035,I536183,I536169,);
nor I_31369 (I536350,I417506,I417488);
nand I_31370 (I536367,I536350,I417503);
DFFARX1 I_31371 (I536367,I3035,I536183,I536172,);
nor I_31372 (I536398,I536285,I417506);
nand I_31373 (I536415,I536398,I417491);
nor I_31374 (I536432,I536209,I536415);
DFFARX1 I_31375 (I536432,I3035,I536183,I536148,);
not I_31376 (I536463,I536415);
nand I_31377 (I536160,I536226,I536463);
DFFARX1 I_31378 (I536415,I3035,I536183,I536503,);
not I_31379 (I536511,I536503);
not I_31380 (I536528,I417506);
not I_31381 (I536545,I417500);
nor I_31382 (I536562,I536545,I417497);
nor I_31383 (I536175,I536511,I536562);
nor I_31384 (I536593,I536545,I417509);
and I_31385 (I536610,I536593,I417512);
or I_31386 (I536627,I536610,I417491);
DFFARX1 I_31387 (I536627,I3035,I536183,I536653,);
nor I_31388 (I536163,I536653,I536209);
not I_31389 (I536675,I536653);
and I_31390 (I536692,I536675,I536209);
nor I_31391 (I536157,I536234,I536692);
nand I_31392 (I536723,I536675,I536285);
nor I_31393 (I536151,I536545,I536723);
nand I_31394 (I536154,I536675,I536463);
nand I_31395 (I536768,I536285,I417500);
nor I_31396 (I536166,I536528,I536768);
not I_31397 (I536829,I3042);
DFFARX1 I_31398 (I64194,I3035,I536829,I536855,);
DFFARX1 I_31399 (I64200,I3035,I536829,I536872,);
not I_31400 (I536880,I536872);
not I_31401 (I536897,I64218);
nor I_31402 (I536914,I536897,I64197);
not I_31403 (I536931,I64203);
nor I_31404 (I536948,I536914,I64209);
nor I_31405 (I536965,I536872,I536948);
DFFARX1 I_31406 (I536965,I3035,I536829,I536815,);
nor I_31407 (I536996,I64209,I64197);
nand I_31408 (I537013,I536996,I64218);
DFFARX1 I_31409 (I537013,I3035,I536829,I536818,);
nor I_31410 (I537044,I536931,I64209);
nand I_31411 (I537061,I537044,I64215);
nor I_31412 (I537078,I536855,I537061);
DFFARX1 I_31413 (I537078,I3035,I536829,I536794,);
not I_31414 (I537109,I537061);
nand I_31415 (I536806,I536872,I537109);
DFFARX1 I_31416 (I537061,I3035,I536829,I537149,);
not I_31417 (I537157,I537149);
not I_31418 (I537174,I64209);
not I_31419 (I537191,I64197);
nor I_31420 (I537208,I537191,I64203);
nor I_31421 (I536821,I537157,I537208);
nor I_31422 (I537239,I537191,I64206);
and I_31423 (I537256,I537239,I64194);
or I_31424 (I537273,I537256,I64212);
DFFARX1 I_31425 (I537273,I3035,I536829,I537299,);
nor I_31426 (I536809,I537299,I536855);
not I_31427 (I537321,I537299);
and I_31428 (I537338,I537321,I536855);
nor I_31429 (I536803,I536880,I537338);
nand I_31430 (I537369,I537321,I536931);
nor I_31431 (I536797,I537191,I537369);
nand I_31432 (I536800,I537321,I537109);
nand I_31433 (I537414,I536931,I64197);
nor I_31434 (I536812,I537174,I537414);
not I_31435 (I537475,I3042);
DFFARX1 I_31436 (I663768,I3035,I537475,I537501,);
DFFARX1 I_31437 (I663774,I3035,I537475,I537518,);
not I_31438 (I537526,I537518);
not I_31439 (I537543,I663771);
nor I_31440 (I537560,I537543,I663750);
not I_31441 (I537577,I663753);
nor I_31442 (I537594,I537560,I663759);
nor I_31443 (I537611,I537518,I537594);
DFFARX1 I_31444 (I537611,I3035,I537475,I537461,);
nor I_31445 (I537642,I663759,I663750);
nand I_31446 (I537659,I537642,I663771);
DFFARX1 I_31447 (I537659,I3035,I537475,I537464,);
nor I_31448 (I537690,I537577,I663759);
nand I_31449 (I537707,I537690,I663753);
nor I_31450 (I537724,I537501,I537707);
DFFARX1 I_31451 (I537724,I3035,I537475,I537440,);
not I_31452 (I537755,I537707);
nand I_31453 (I537452,I537518,I537755);
DFFARX1 I_31454 (I537707,I3035,I537475,I537795,);
not I_31455 (I537803,I537795);
not I_31456 (I537820,I663759);
not I_31457 (I537837,I663762);
nor I_31458 (I537854,I537837,I663753);
nor I_31459 (I537467,I537803,I537854);
nor I_31460 (I537885,I537837,I663750);
and I_31461 (I537902,I537885,I663756);
or I_31462 (I537919,I537902,I663765);
DFFARX1 I_31463 (I537919,I3035,I537475,I537945,);
nor I_31464 (I537455,I537945,I537501);
not I_31465 (I537967,I537945);
and I_31466 (I537984,I537967,I537501);
nor I_31467 (I537449,I537526,I537984);
nand I_31468 (I538015,I537967,I537577);
nor I_31469 (I537443,I537837,I538015);
nand I_31470 (I537446,I537967,I537755);
nand I_31471 (I538060,I537577,I663762);
nor I_31472 (I537458,I537820,I538060);
not I_31473 (I538121,I3042);
DFFARX1 I_31474 (I279403,I3035,I538121,I538147,);
DFFARX1 I_31475 (I279400,I3035,I538121,I538164,);
not I_31476 (I538172,I538164);
not I_31477 (I538189,I279415);
nor I_31478 (I538206,I538189,I279418);
not I_31479 (I538223,I279406);
nor I_31480 (I538240,I538206,I279412);
nor I_31481 (I538257,I538164,I538240);
DFFARX1 I_31482 (I538257,I3035,I538121,I538107,);
nor I_31483 (I538288,I279412,I279418);
nand I_31484 (I538305,I538288,I279415);
DFFARX1 I_31485 (I538305,I3035,I538121,I538110,);
nor I_31486 (I538336,I538223,I279412);
nand I_31487 (I538353,I538336,I279424);
nor I_31488 (I538370,I538147,I538353);
DFFARX1 I_31489 (I538370,I3035,I538121,I538086,);
not I_31490 (I538401,I538353);
nand I_31491 (I538098,I538164,I538401);
DFFARX1 I_31492 (I538353,I3035,I538121,I538441,);
not I_31493 (I538449,I538441);
not I_31494 (I538466,I279412);
not I_31495 (I538483,I279397);
nor I_31496 (I538500,I538483,I279406);
nor I_31497 (I538113,I538449,I538500);
nor I_31498 (I538531,I538483,I279409);
and I_31499 (I538548,I538531,I279397);
or I_31500 (I538565,I538548,I279421);
DFFARX1 I_31501 (I538565,I3035,I538121,I538591,);
nor I_31502 (I538101,I538591,I538147);
not I_31503 (I538613,I538591);
and I_31504 (I538630,I538613,I538147);
nor I_31505 (I538095,I538172,I538630);
nand I_31506 (I538661,I538613,I538223);
nor I_31507 (I538089,I538483,I538661);
nand I_31508 (I538092,I538613,I538401);
nand I_31509 (I538706,I538223,I279397);
nor I_31510 (I538104,I538466,I538706);
not I_31511 (I538767,I3042);
DFFARX1 I_31512 (I643980,I3035,I538767,I538793,);
DFFARX1 I_31513 (I643962,I3035,I538767,I538810,);
not I_31514 (I538818,I538810);
not I_31515 (I538835,I643971);
nor I_31516 (I538852,I538835,I643983);
not I_31517 (I538869,I643965);
nor I_31518 (I538886,I538852,I643974);
nor I_31519 (I538903,I538810,I538886);
DFFARX1 I_31520 (I538903,I3035,I538767,I538753,);
nor I_31521 (I538934,I643974,I643983);
nand I_31522 (I538951,I538934,I643971);
DFFARX1 I_31523 (I538951,I3035,I538767,I538756,);
nor I_31524 (I538982,I538869,I643974);
nand I_31525 (I538999,I538982,I643986);
nor I_31526 (I539016,I538793,I538999);
DFFARX1 I_31527 (I539016,I3035,I538767,I538732,);
not I_31528 (I539047,I538999);
nand I_31529 (I538744,I538810,I539047);
DFFARX1 I_31530 (I538999,I3035,I538767,I539087,);
not I_31531 (I539095,I539087);
not I_31532 (I539112,I643974);
not I_31533 (I539129,I643962);
nor I_31534 (I539146,I539129,I643965);
nor I_31535 (I538759,I539095,I539146);
nor I_31536 (I539177,I539129,I643968);
and I_31537 (I539194,I539177,I643977);
or I_31538 (I539211,I539194,I643965);
DFFARX1 I_31539 (I539211,I3035,I538767,I539237,);
nor I_31540 (I538747,I539237,I538793);
not I_31541 (I539259,I539237);
and I_31542 (I539276,I539259,I538793);
nor I_31543 (I538741,I538818,I539276);
nand I_31544 (I539307,I539259,I538869);
nor I_31545 (I538735,I539129,I539307);
nand I_31546 (I538738,I539259,I539047);
nand I_31547 (I539352,I538869,I643962);
nor I_31548 (I538750,I539112,I539352);
not I_31549 (I539413,I3042);
DFFARX1 I_31550 (I687525,I3035,I539413,I539439,);
DFFARX1 I_31551 (I687519,I3035,I539413,I539456,);
not I_31552 (I539464,I539456);
not I_31553 (I539481,I687528);
nor I_31554 (I539498,I539481,I687540);
not I_31555 (I539515,I687522);
nor I_31556 (I539532,I539498,I687519);
nor I_31557 (I539549,I539456,I539532);
DFFARX1 I_31558 (I539549,I3035,I539413,I539399,);
nor I_31559 (I539580,I687519,I687540);
nand I_31560 (I539597,I539580,I687528);
DFFARX1 I_31561 (I539597,I3035,I539413,I539402,);
nor I_31562 (I539628,I539515,I687519);
nand I_31563 (I539645,I539628,I687516);
nor I_31564 (I539662,I539439,I539645);
DFFARX1 I_31565 (I539662,I3035,I539413,I539378,);
not I_31566 (I539693,I539645);
nand I_31567 (I539390,I539456,I539693);
DFFARX1 I_31568 (I539645,I3035,I539413,I539733,);
not I_31569 (I539741,I539733);
not I_31570 (I539758,I687519);
not I_31571 (I539775,I687537);
nor I_31572 (I539792,I539775,I687522);
nor I_31573 (I539405,I539741,I539792);
nor I_31574 (I539823,I539775,I687531);
and I_31575 (I539840,I539823,I687516);
or I_31576 (I539857,I539840,I687534);
DFFARX1 I_31577 (I539857,I3035,I539413,I539883,);
nor I_31578 (I539393,I539883,I539439);
not I_31579 (I539905,I539883);
and I_31580 (I539922,I539905,I539439);
nor I_31581 (I539387,I539464,I539922);
nand I_31582 (I539953,I539905,I539515);
nor I_31583 (I539381,I539775,I539953);
nand I_31584 (I539384,I539905,I539693);
nand I_31585 (I539998,I539515,I687537);
nor I_31586 (I539396,I539758,I539998);
not I_31587 (I540059,I3042);
DFFARX1 I_31588 (I335993,I3035,I540059,I540085,);
DFFARX1 I_31589 (I336005,I3035,I540059,I540102,);
not I_31590 (I540110,I540102);
not I_31591 (I540127,I336014);
nor I_31592 (I540144,I540127,I335990);
not I_31593 (I540161,I336008);
nor I_31594 (I540178,I540144,I336002);
nor I_31595 (I540195,I540102,I540178);
DFFARX1 I_31596 (I540195,I3035,I540059,I540045,);
nor I_31597 (I540226,I336002,I335990);
nand I_31598 (I540243,I540226,I336014);
DFFARX1 I_31599 (I540243,I3035,I540059,I540048,);
nor I_31600 (I540274,I540161,I336002);
nand I_31601 (I540291,I540274,I335996);
nor I_31602 (I540308,I540085,I540291);
DFFARX1 I_31603 (I540308,I3035,I540059,I540024,);
not I_31604 (I540339,I540291);
nand I_31605 (I540036,I540102,I540339);
DFFARX1 I_31606 (I540291,I3035,I540059,I540379,);
not I_31607 (I540387,I540379);
not I_31608 (I540404,I336002);
not I_31609 (I540421,I336011);
nor I_31610 (I540438,I540421,I336008);
nor I_31611 (I540051,I540387,I540438);
nor I_31612 (I540469,I540421,I335993);
and I_31613 (I540486,I540469,I335990);
or I_31614 (I540503,I540486,I335999);
DFFARX1 I_31615 (I540503,I3035,I540059,I540529,);
nor I_31616 (I540039,I540529,I540085);
not I_31617 (I540551,I540529);
and I_31618 (I540568,I540551,I540085);
nor I_31619 (I540033,I540110,I540568);
nand I_31620 (I540599,I540551,I540161);
nor I_31621 (I540027,I540421,I540599);
nand I_31622 (I540030,I540551,I540339);
nand I_31623 (I540644,I540161,I336011);
nor I_31624 (I540042,I540404,I540644);
not I_31625 (I540705,I3042);
DFFARX1 I_31626 (I32574,I3035,I540705,I540731,);
DFFARX1 I_31627 (I32580,I3035,I540705,I540748,);
not I_31628 (I540756,I540748);
not I_31629 (I540773,I32598);
nor I_31630 (I540790,I540773,I32577);
not I_31631 (I540807,I32583);
nor I_31632 (I540824,I540790,I32589);
nor I_31633 (I540841,I540748,I540824);
DFFARX1 I_31634 (I540841,I3035,I540705,I540691,);
nor I_31635 (I540872,I32589,I32577);
nand I_31636 (I540889,I540872,I32598);
DFFARX1 I_31637 (I540889,I3035,I540705,I540694,);
nor I_31638 (I540920,I540807,I32589);
nand I_31639 (I540937,I540920,I32595);
nor I_31640 (I540954,I540731,I540937);
DFFARX1 I_31641 (I540954,I3035,I540705,I540670,);
not I_31642 (I540985,I540937);
nand I_31643 (I540682,I540748,I540985);
DFFARX1 I_31644 (I540937,I3035,I540705,I541025,);
not I_31645 (I541033,I541025);
not I_31646 (I541050,I32589);
not I_31647 (I541067,I32577);
nor I_31648 (I541084,I541067,I32583);
nor I_31649 (I540697,I541033,I541084);
nor I_31650 (I541115,I541067,I32586);
and I_31651 (I541132,I541115,I32574);
or I_31652 (I541149,I541132,I32592);
DFFARX1 I_31653 (I541149,I3035,I540705,I541175,);
nor I_31654 (I540685,I541175,I540731);
not I_31655 (I541197,I541175);
and I_31656 (I541214,I541197,I540731);
nor I_31657 (I540679,I540756,I541214);
nand I_31658 (I541245,I541197,I540807);
nor I_31659 (I540673,I541067,I541245);
nand I_31660 (I540676,I541197,I540985);
nand I_31661 (I541290,I540807,I32577);
nor I_31662 (I540688,I541050,I541290);
not I_31663 (I541351,I3042);
DFFARX1 I_31664 (I198783,I3035,I541351,I541377,);
DFFARX1 I_31665 (I198789,I3035,I541351,I541394,);
not I_31666 (I541402,I541394);
not I_31667 (I541419,I198810);
nor I_31668 (I541436,I541419,I198798);
not I_31669 (I541453,I198807);
nor I_31670 (I541470,I541436,I198792);
nor I_31671 (I541487,I541394,I541470);
DFFARX1 I_31672 (I541487,I3035,I541351,I541337,);
nor I_31673 (I541518,I198792,I198798);
nand I_31674 (I541535,I541518,I198810);
DFFARX1 I_31675 (I541535,I3035,I541351,I541340,);
nor I_31676 (I541566,I541453,I198792);
nand I_31677 (I541583,I541566,I198783);
nor I_31678 (I541600,I541377,I541583);
DFFARX1 I_31679 (I541600,I3035,I541351,I541316,);
not I_31680 (I541631,I541583);
nand I_31681 (I541328,I541394,I541631);
DFFARX1 I_31682 (I541583,I3035,I541351,I541671,);
not I_31683 (I541679,I541671);
not I_31684 (I541696,I198792);
not I_31685 (I541713,I198795);
nor I_31686 (I541730,I541713,I198807);
nor I_31687 (I541343,I541679,I541730);
nor I_31688 (I541761,I541713,I198804);
and I_31689 (I541778,I541761,I198786);
or I_31690 (I541795,I541778,I198801);
DFFARX1 I_31691 (I541795,I3035,I541351,I541821,);
nor I_31692 (I541331,I541821,I541377);
not I_31693 (I541843,I541821);
and I_31694 (I541860,I541843,I541377);
nor I_31695 (I541325,I541402,I541860);
nand I_31696 (I541891,I541843,I541453);
nor I_31697 (I541319,I541713,I541891);
nand I_31698 (I541322,I541843,I541631);
nand I_31699 (I541936,I541453,I198795);
nor I_31700 (I541334,I541696,I541936);
not I_31701 (I541997,I3042);
DFFARX1 I_31702 (I208269,I3035,I541997,I542023,);
DFFARX1 I_31703 (I208275,I3035,I541997,I542040,);
not I_31704 (I542048,I542040);
not I_31705 (I542065,I208296);
nor I_31706 (I542082,I542065,I208284);
not I_31707 (I542099,I208293);
nor I_31708 (I542116,I542082,I208278);
nor I_31709 (I542133,I542040,I542116);
DFFARX1 I_31710 (I542133,I3035,I541997,I541983,);
nor I_31711 (I542164,I208278,I208284);
nand I_31712 (I542181,I542164,I208296);
DFFARX1 I_31713 (I542181,I3035,I541997,I541986,);
nor I_31714 (I542212,I542099,I208278);
nand I_31715 (I542229,I542212,I208269);
nor I_31716 (I542246,I542023,I542229);
DFFARX1 I_31717 (I542246,I3035,I541997,I541962,);
not I_31718 (I542277,I542229);
nand I_31719 (I541974,I542040,I542277);
DFFARX1 I_31720 (I542229,I3035,I541997,I542317,);
not I_31721 (I542325,I542317);
not I_31722 (I542342,I208278);
not I_31723 (I542359,I208281);
nor I_31724 (I542376,I542359,I208293);
nor I_31725 (I541989,I542325,I542376);
nor I_31726 (I542407,I542359,I208290);
and I_31727 (I542424,I542407,I208272);
or I_31728 (I542441,I542424,I208287);
DFFARX1 I_31729 (I542441,I3035,I541997,I542467,);
nor I_31730 (I541977,I542467,I542023);
not I_31731 (I542489,I542467);
and I_31732 (I542506,I542489,I542023);
nor I_31733 (I541971,I542048,I542506);
nand I_31734 (I542537,I542489,I542099);
nor I_31735 (I541965,I542359,I542537);
nand I_31736 (I541968,I542489,I542277);
nand I_31737 (I542582,I542099,I208281);
nor I_31738 (I541980,I542342,I542582);
not I_31739 (I542643,I3042);
DFFARX1 I_31740 (I566119,I3035,I542643,I542669,);
DFFARX1 I_31741 (I566122,I3035,I542643,I542686,);
not I_31742 (I542694,I542686);
not I_31743 (I542711,I566119);
nor I_31744 (I542728,I542711,I566131);
not I_31745 (I542745,I566140);
nor I_31746 (I542762,I542728,I566128);
nor I_31747 (I542779,I542686,I542762);
DFFARX1 I_31748 (I542779,I3035,I542643,I542629,);
nor I_31749 (I542810,I566128,I566131);
nand I_31750 (I542827,I542810,I566119);
DFFARX1 I_31751 (I542827,I3035,I542643,I542632,);
nor I_31752 (I542858,I542745,I566128);
nand I_31753 (I542875,I542858,I566134);
nor I_31754 (I542892,I542669,I542875);
DFFARX1 I_31755 (I542892,I3035,I542643,I542608,);
not I_31756 (I542923,I542875);
nand I_31757 (I542620,I542686,I542923);
DFFARX1 I_31758 (I542875,I3035,I542643,I542963,);
not I_31759 (I542971,I542963);
not I_31760 (I542988,I566128);
not I_31761 (I543005,I566125);
nor I_31762 (I543022,I543005,I566140);
nor I_31763 (I542635,I542971,I543022);
nor I_31764 (I543053,I543005,I566137);
and I_31765 (I543070,I543053,I566125);
or I_31766 (I543087,I543070,I566122);
DFFARX1 I_31767 (I543087,I3035,I542643,I543113,);
nor I_31768 (I542623,I543113,I542669);
not I_31769 (I543135,I543113);
and I_31770 (I543152,I543135,I542669);
nor I_31771 (I542617,I542694,I543152);
nand I_31772 (I543183,I543135,I542745);
nor I_31773 (I542611,I543005,I543183);
nand I_31774 (I542614,I543135,I542923);
nand I_31775 (I543228,I542745,I566125);
nor I_31776 (I542626,I542988,I543228);
not I_31777 (I543289,I3042);
DFFARX1 I_31778 (I285299,I3035,I543289,I543315,);
DFFARX1 I_31779 (I285311,I3035,I543289,I543332,);
not I_31780 (I543340,I543332);
not I_31781 (I543357,I285296);
nor I_31782 (I543374,I543357,I285314);
not I_31783 (I543391,I285320);
nor I_31784 (I543408,I543374,I285302);
nor I_31785 (I543425,I543332,I543408);
DFFARX1 I_31786 (I543425,I3035,I543289,I543275,);
nor I_31787 (I543456,I285302,I285314);
nand I_31788 (I543473,I543456,I285296);
DFFARX1 I_31789 (I543473,I3035,I543289,I543278,);
nor I_31790 (I543504,I543391,I285302);
nand I_31791 (I543521,I543504,I285305);
nor I_31792 (I543538,I543315,I543521);
DFFARX1 I_31793 (I543538,I3035,I543289,I543254,);
not I_31794 (I543569,I543521);
nand I_31795 (I543266,I543332,I543569);
DFFARX1 I_31796 (I543521,I3035,I543289,I543609,);
not I_31797 (I543617,I543609);
not I_31798 (I543634,I285302);
not I_31799 (I543651,I285308);
nor I_31800 (I543668,I543651,I285320);
nor I_31801 (I543281,I543617,I543668);
nor I_31802 (I543699,I543651,I285317);
and I_31803 (I543716,I543699,I285296);
or I_31804 (I543733,I543716,I285299);
DFFARX1 I_31805 (I543733,I3035,I543289,I543759,);
nor I_31806 (I543269,I543759,I543315);
not I_31807 (I543781,I543759);
and I_31808 (I543798,I543781,I543315);
nor I_31809 (I543263,I543340,I543798);
nand I_31810 (I543829,I543781,I543391);
nor I_31811 (I543257,I543651,I543829);
nand I_31812 (I543260,I543781,I543569);
nand I_31813 (I543874,I543391,I285308);
nor I_31814 (I543272,I543634,I543874);
not I_31815 (I543935,I3042);
DFFARX1 I_31816 (I660504,I3035,I543935,I543961,);
DFFARX1 I_31817 (I660510,I3035,I543935,I543978,);
not I_31818 (I543986,I543978);
not I_31819 (I544003,I660507);
nor I_31820 (I544020,I544003,I660486);
not I_31821 (I544037,I660489);
nor I_31822 (I544054,I544020,I660495);
nor I_31823 (I544071,I543978,I544054);
DFFARX1 I_31824 (I544071,I3035,I543935,I543921,);
nor I_31825 (I544102,I660495,I660486);
nand I_31826 (I544119,I544102,I660507);
DFFARX1 I_31827 (I544119,I3035,I543935,I543924,);
nor I_31828 (I544150,I544037,I660495);
nand I_31829 (I544167,I544150,I660489);
nor I_31830 (I544184,I543961,I544167);
DFFARX1 I_31831 (I544184,I3035,I543935,I543900,);
not I_31832 (I544215,I544167);
nand I_31833 (I543912,I543978,I544215);
DFFARX1 I_31834 (I544167,I3035,I543935,I544255,);
not I_31835 (I544263,I544255);
not I_31836 (I544280,I660495);
not I_31837 (I544297,I660498);
nor I_31838 (I544314,I544297,I660489);
nor I_31839 (I543927,I544263,I544314);
nor I_31840 (I544345,I544297,I660486);
and I_31841 (I544362,I544345,I660492);
or I_31842 (I544379,I544362,I660501);
DFFARX1 I_31843 (I544379,I3035,I543935,I544405,);
nor I_31844 (I543915,I544405,I543961);
not I_31845 (I544427,I544405);
and I_31846 (I544444,I544427,I543961);
nor I_31847 (I543909,I543986,I544444);
nand I_31848 (I544475,I544427,I544037);
nor I_31849 (I543903,I544297,I544475);
nand I_31850 (I543906,I544427,I544215);
nand I_31851 (I544520,I544037,I660498);
nor I_31852 (I543918,I544280,I544520);
not I_31853 (I544581,I3042);
DFFARX1 I_31854 (I663224,I3035,I544581,I544607,);
DFFARX1 I_31855 (I663230,I3035,I544581,I544624,);
not I_31856 (I544632,I544624);
not I_31857 (I544649,I663227);
nor I_31858 (I544666,I544649,I663206);
not I_31859 (I544683,I663209);
nor I_31860 (I544700,I544666,I663215);
nor I_31861 (I544717,I544624,I544700);
DFFARX1 I_31862 (I544717,I3035,I544581,I544567,);
nor I_31863 (I544748,I663215,I663206);
nand I_31864 (I544765,I544748,I663227);
DFFARX1 I_31865 (I544765,I3035,I544581,I544570,);
nor I_31866 (I544796,I544683,I663215);
nand I_31867 (I544813,I544796,I663209);
nor I_31868 (I544830,I544607,I544813);
DFFARX1 I_31869 (I544830,I3035,I544581,I544546,);
not I_31870 (I544861,I544813);
nand I_31871 (I544558,I544624,I544861);
DFFARX1 I_31872 (I544813,I3035,I544581,I544901,);
not I_31873 (I544909,I544901);
not I_31874 (I544926,I663215);
not I_31875 (I544943,I663218);
nor I_31876 (I544960,I544943,I663209);
nor I_31877 (I544573,I544909,I544960);
nor I_31878 (I544991,I544943,I663206);
and I_31879 (I545008,I544991,I663212);
or I_31880 (I545025,I545008,I663221);
DFFARX1 I_31881 (I545025,I3035,I544581,I545051,);
nor I_31882 (I544561,I545051,I544607);
not I_31883 (I545073,I545051);
and I_31884 (I545090,I545073,I544607);
nor I_31885 (I544555,I544632,I545090);
nand I_31886 (I545121,I545073,I544683);
nor I_31887 (I544549,I544943,I545121);
nand I_31888 (I544552,I545073,I544861);
nand I_31889 (I545166,I544683,I663218);
nor I_31890 (I544564,I544926,I545166);
not I_31891 (I545227,I3042);
DFFARX1 I_31892 (I679433,I3035,I545227,I545253,);
DFFARX1 I_31893 (I679427,I3035,I545227,I545270,);
not I_31894 (I545278,I545270);
not I_31895 (I545295,I679436);
nor I_31896 (I545312,I545295,I679448);
not I_31897 (I545329,I679430);
nor I_31898 (I545346,I545312,I679427);
nor I_31899 (I545363,I545270,I545346);
DFFARX1 I_31900 (I545363,I3035,I545227,I545213,);
nor I_31901 (I545394,I679427,I679448);
nand I_31902 (I545411,I545394,I679436);
DFFARX1 I_31903 (I545411,I3035,I545227,I545216,);
nor I_31904 (I545442,I545329,I679427);
nand I_31905 (I545459,I545442,I679424);
nor I_31906 (I545476,I545253,I545459);
DFFARX1 I_31907 (I545476,I3035,I545227,I545192,);
not I_31908 (I545507,I545459);
nand I_31909 (I545204,I545270,I545507);
DFFARX1 I_31910 (I545459,I3035,I545227,I545547,);
not I_31911 (I545555,I545547);
not I_31912 (I545572,I679427);
not I_31913 (I545589,I679445);
nor I_31914 (I545606,I545589,I679430);
nor I_31915 (I545219,I545555,I545606);
nor I_31916 (I545637,I545589,I679439);
and I_31917 (I545654,I545637,I679424);
or I_31918 (I545671,I545654,I679442);
DFFARX1 I_31919 (I545671,I3035,I545227,I545697,);
nor I_31920 (I545207,I545697,I545253);
not I_31921 (I545719,I545697);
and I_31922 (I545736,I545719,I545253);
nor I_31923 (I545201,I545278,I545736);
nand I_31924 (I545767,I545719,I545329);
nor I_31925 (I545195,I545589,I545767);
nand I_31926 (I545198,I545719,I545507);
nand I_31927 (I545812,I545329,I679445);
nor I_31928 (I545210,I545572,I545812);
not I_31929 (I545873,I3042);
DFFARX1 I_31930 (I175595,I3035,I545873,I545899,);
DFFARX1 I_31931 (I175601,I3035,I545873,I545916,);
not I_31932 (I545924,I545916);
not I_31933 (I545941,I175622);
nor I_31934 (I545958,I545941,I175610);
not I_31935 (I545975,I175619);
nor I_31936 (I545992,I545958,I175604);
nor I_31937 (I546009,I545916,I545992);
DFFARX1 I_31938 (I546009,I3035,I545873,I545859,);
nor I_31939 (I546040,I175604,I175610);
nand I_31940 (I546057,I546040,I175622);
DFFARX1 I_31941 (I546057,I3035,I545873,I545862,);
nor I_31942 (I546088,I545975,I175604);
nand I_31943 (I546105,I546088,I175595);
nor I_31944 (I546122,I545899,I546105);
DFFARX1 I_31945 (I546122,I3035,I545873,I545838,);
not I_31946 (I546153,I546105);
nand I_31947 (I545850,I545916,I546153);
DFFARX1 I_31948 (I546105,I3035,I545873,I546193,);
not I_31949 (I546201,I546193);
not I_31950 (I546218,I175604);
not I_31951 (I546235,I175607);
nor I_31952 (I546252,I546235,I175619);
nor I_31953 (I545865,I546201,I546252);
nor I_31954 (I546283,I546235,I175616);
and I_31955 (I546300,I546283,I175598);
or I_31956 (I546317,I546300,I175613);
DFFARX1 I_31957 (I546317,I3035,I545873,I546343,);
nor I_31958 (I545853,I546343,I545899);
not I_31959 (I546365,I546343);
and I_31960 (I546382,I546365,I545899);
nor I_31961 (I545847,I545924,I546382);
nand I_31962 (I546413,I546365,I545975);
nor I_31963 (I545841,I546235,I546413);
nand I_31964 (I545844,I546365,I546153);
nand I_31965 (I546458,I545975,I175607);
nor I_31966 (I545856,I546218,I546458);
not I_31967 (I546513,I3042);
DFFARX1 I_31968 (I108057,I3035,I546513,I546539,);
DFFARX1 I_31969 (I546539,I3035,I546513,I546556,);
not I_31970 (I546505,I546556);
not I_31971 (I546578,I546539);
DFFARX1 I_31972 (I108072,I3035,I546513,I546604,);
nand I_31973 (I546612,I546604,I108054);
not I_31974 (I546629,I108054);
not I_31975 (I546646,I108063);
nand I_31976 (I546663,I108069,I108060);
and I_31977 (I546680,I108069,I108060);
not I_31978 (I546697,I108057);
nand I_31979 (I546714,I546697,I546646);
nor I_31980 (I546487,I546714,I546612);
nor I_31981 (I546745,I546629,I546714);
nand I_31982 (I546490,I546680,I546745);
not I_31983 (I546776,I108054);
nor I_31984 (I546793,I546776,I108069);
nor I_31985 (I546810,I546793,I108057);
nor I_31986 (I546827,I546578,I546810);
DFFARX1 I_31987 (I546827,I3035,I546513,I546499,);
not I_31988 (I546858,I546793);
DFFARX1 I_31989 (I546858,I3035,I546513,I546502,);
and I_31990 (I546496,I546604,I546793);
nor I_31991 (I546903,I546776,I108078);
and I_31992 (I546920,I546903,I108075);
or I_31993 (I546937,I546920,I108066);
DFFARX1 I_31994 (I546937,I3035,I546513,I546963,);
nor I_31995 (I546971,I546963,I546697);
DFFARX1 I_31996 (I546971,I3035,I546513,I546484,);
nand I_31997 (I547002,I546963,I546604);
nand I_31998 (I547019,I546697,I547002);
nor I_31999 (I546493,I547019,I546663);
not I_32000 (I547074,I3042);
DFFARX1 I_32001 (I232093,I3035,I547074,I547100,);
DFFARX1 I_32002 (I547100,I3035,I547074,I547117,);
not I_32003 (I547066,I547117);
not I_32004 (I547139,I547100);
DFFARX1 I_32005 (I232081,I3035,I547074,I547165,);
nand I_32006 (I547173,I547165,I232087);
not I_32007 (I547190,I232087);
not I_32008 (I547207,I232084);
nand I_32009 (I547224,I232072,I232069);
and I_32010 (I547241,I232072,I232069);
not I_32011 (I547258,I232096);
nand I_32012 (I547275,I547258,I547207);
nor I_32013 (I547048,I547275,I547173);
nor I_32014 (I547306,I547190,I547275);
nand I_32015 (I547051,I547241,I547306);
not I_32016 (I547337,I232069);
nor I_32017 (I547354,I547337,I232072);
nor I_32018 (I547371,I547354,I232096);
nor I_32019 (I547388,I547139,I547371);
DFFARX1 I_32020 (I547388,I3035,I547074,I547060,);
not I_32021 (I547419,I547354);
DFFARX1 I_32022 (I547419,I3035,I547074,I547063,);
and I_32023 (I547057,I547165,I547354);
nor I_32024 (I547464,I547337,I232078);
and I_32025 (I547481,I547464,I232075);
or I_32026 (I547498,I547481,I232090);
DFFARX1 I_32027 (I547498,I3035,I547074,I547524,);
nor I_32028 (I547532,I547524,I547258);
DFFARX1 I_32029 (I547532,I3035,I547074,I547045,);
nand I_32030 (I547563,I547524,I547165);
nand I_32031 (I547580,I547258,I547563);
nor I_32032 (I547054,I547580,I547224);
not I_32033 (I547635,I3042);
DFFARX1 I_32034 (I389747,I3035,I547635,I547661,);
DFFARX1 I_32035 (I547661,I3035,I547635,I547678,);
not I_32036 (I547627,I547678);
not I_32037 (I547700,I547661);
DFFARX1 I_32038 (I389759,I3035,I547635,I547726,);
nand I_32039 (I547734,I547726,I389768);
not I_32040 (I547751,I389768);
not I_32041 (I547768,I389750);
nand I_32042 (I547785,I389753,I389744);
and I_32043 (I547802,I389753,I389744);
not I_32044 (I547819,I389762);
nand I_32045 (I547836,I547819,I547768);
nor I_32046 (I547609,I547836,I547734);
nor I_32047 (I547867,I547751,I547836);
nand I_32048 (I547612,I547802,I547867);
not I_32049 (I547898,I389765);
nor I_32050 (I547915,I547898,I389753);
nor I_32051 (I547932,I547915,I389762);
nor I_32052 (I547949,I547700,I547932);
DFFARX1 I_32053 (I547949,I3035,I547635,I547621,);
not I_32054 (I547980,I547915);
DFFARX1 I_32055 (I547980,I3035,I547635,I547624,);
and I_32056 (I547618,I547726,I547915);
nor I_32057 (I548025,I547898,I389744);
and I_32058 (I548042,I548025,I389756);
or I_32059 (I548059,I548042,I389747);
DFFARX1 I_32060 (I548059,I3035,I547635,I548085,);
nor I_32061 (I548093,I548085,I547819);
DFFARX1 I_32062 (I548093,I3035,I547635,I547606,);
nand I_32063 (I548124,I548085,I547726);
nand I_32064 (I548141,I547819,I548124);
nor I_32065 (I547615,I548141,I547785);
not I_32066 (I548196,I3042);
DFFARX1 I_32067 (I464604,I3035,I548196,I548222,);
DFFARX1 I_32068 (I548222,I3035,I548196,I548239,);
not I_32069 (I548188,I548239);
not I_32070 (I548261,I548222);
DFFARX1 I_32071 (I464601,I3035,I548196,I548287,);
nand I_32072 (I548295,I548287,I464616);
not I_32073 (I548312,I464616);
not I_32074 (I548329,I464613);
nand I_32075 (I548346,I464610,I464598);
and I_32076 (I548363,I464610,I464598);
not I_32077 (I548380,I464595);
nand I_32078 (I548397,I548380,I548329);
nor I_32079 (I548170,I548397,I548295);
nor I_32080 (I548428,I548312,I548397);
nand I_32081 (I548173,I548363,I548428);
not I_32082 (I548459,I464601);
nor I_32083 (I548476,I548459,I464610);
nor I_32084 (I548493,I548476,I464595);
nor I_32085 (I548510,I548261,I548493);
DFFARX1 I_32086 (I548510,I3035,I548196,I548182,);
not I_32087 (I548541,I548476);
DFFARX1 I_32088 (I548541,I3035,I548196,I548185,);
and I_32089 (I548179,I548287,I548476);
nor I_32090 (I548586,I548459,I464607);
and I_32091 (I548603,I548586,I464595);
or I_32092 (I548620,I548603,I464598);
DFFARX1 I_32093 (I548620,I3035,I548196,I548646,);
nor I_32094 (I548654,I548646,I548380);
DFFARX1 I_32095 (I548654,I3035,I548196,I548167,);
nand I_32096 (I548685,I548646,I548287);
nand I_32097 (I548702,I548380,I548685);
nor I_32098 (I548176,I548702,I548346);
not I_32099 (I548757,I3042);
DFFARX1 I_32100 (I370095,I3035,I548757,I548783,);
DFFARX1 I_32101 (I548783,I3035,I548757,I548800,);
not I_32102 (I548749,I548800);
not I_32103 (I548822,I548783);
DFFARX1 I_32104 (I370107,I3035,I548757,I548848,);
nand I_32105 (I548856,I548848,I370116);
not I_32106 (I548873,I370116);
not I_32107 (I548890,I370098);
nand I_32108 (I548907,I370101,I370092);
and I_32109 (I548924,I370101,I370092);
not I_32110 (I548941,I370110);
nand I_32111 (I548958,I548941,I548890);
nor I_32112 (I548731,I548958,I548856);
nor I_32113 (I548989,I548873,I548958);
nand I_32114 (I548734,I548924,I548989);
not I_32115 (I549020,I370113);
nor I_32116 (I549037,I549020,I370101);
nor I_32117 (I549054,I549037,I370110);
nor I_32118 (I549071,I548822,I549054);
DFFARX1 I_32119 (I549071,I3035,I548757,I548743,);
not I_32120 (I549102,I549037);
DFFARX1 I_32121 (I549102,I3035,I548757,I548746,);
and I_32122 (I548740,I548848,I549037);
nor I_32123 (I549147,I549020,I370092);
and I_32124 (I549164,I549147,I370104);
or I_32125 (I549181,I549164,I370095);
DFFARX1 I_32126 (I549181,I3035,I548757,I549207,);
nor I_32127 (I549215,I549207,I548941);
DFFARX1 I_32128 (I549215,I3035,I548757,I548728,);
nand I_32129 (I549246,I549207,I548848);
nand I_32130 (I549263,I548941,I549246);
nor I_32131 (I548737,I549263,I548907);
not I_32132 (I549318,I3042);
DFFARX1 I_32133 (I338883,I3035,I549318,I549344,);
DFFARX1 I_32134 (I549344,I3035,I549318,I549361,);
not I_32135 (I549310,I549361);
not I_32136 (I549383,I549344);
DFFARX1 I_32137 (I338895,I3035,I549318,I549409,);
nand I_32138 (I549417,I549409,I338904);
not I_32139 (I549434,I338904);
not I_32140 (I549451,I338886);
nand I_32141 (I549468,I338889,I338880);
and I_32142 (I549485,I338889,I338880);
not I_32143 (I549502,I338898);
nand I_32144 (I549519,I549502,I549451);
nor I_32145 (I549292,I549519,I549417);
nor I_32146 (I549550,I549434,I549519);
nand I_32147 (I549295,I549485,I549550);
not I_32148 (I549581,I338901);
nor I_32149 (I549598,I549581,I338889);
nor I_32150 (I549615,I549598,I338898);
nor I_32151 (I549632,I549383,I549615);
DFFARX1 I_32152 (I549632,I3035,I549318,I549304,);
not I_32153 (I549663,I549598);
DFFARX1 I_32154 (I549663,I3035,I549318,I549307,);
and I_32155 (I549301,I549409,I549598);
nor I_32156 (I549708,I549581,I338880);
and I_32157 (I549725,I549708,I338892);
or I_32158 (I549742,I549725,I338883);
DFFARX1 I_32159 (I549742,I3035,I549318,I549768,);
nor I_32160 (I549776,I549768,I549502);
DFFARX1 I_32161 (I549776,I3035,I549318,I549289,);
nand I_32162 (I549807,I549768,I549409);
nand I_32163 (I549824,I549502,I549807);
nor I_32164 (I549298,I549824,I549468);
not I_32165 (I549879,I3042);
DFFARX1 I_32166 (I447740,I3035,I549879,I549905,);
DFFARX1 I_32167 (I549905,I3035,I549879,I549922,);
not I_32168 (I549871,I549922);
not I_32169 (I549944,I549905);
DFFARX1 I_32170 (I447737,I3035,I549879,I549970,);
nand I_32171 (I549978,I549970,I447752);
not I_32172 (I549995,I447752);
not I_32173 (I550012,I447749);
nand I_32174 (I550029,I447746,I447734);
and I_32175 (I550046,I447746,I447734);
not I_32176 (I550063,I447731);
nand I_32177 (I550080,I550063,I550012);
nor I_32178 (I549853,I550080,I549978);
nor I_32179 (I550111,I549995,I550080);
nand I_32180 (I549856,I550046,I550111);
not I_32181 (I550142,I447737);
nor I_32182 (I550159,I550142,I447746);
nor I_32183 (I550176,I550159,I447731);
nor I_32184 (I550193,I549944,I550176);
DFFARX1 I_32185 (I550193,I3035,I549879,I549865,);
not I_32186 (I550224,I550159);
DFFARX1 I_32187 (I550224,I3035,I549879,I549868,);
and I_32188 (I549862,I549970,I550159);
nor I_32189 (I550269,I550142,I447743);
and I_32190 (I550286,I550269,I447731);
or I_32191 (I550303,I550286,I447734);
DFFARX1 I_32192 (I550303,I3035,I549879,I550329,);
nor I_32193 (I550337,I550329,I550063);
DFFARX1 I_32194 (I550337,I3035,I549879,I549850,);
nand I_32195 (I550368,I550329,I549970);
nand I_32196 (I550385,I550063,I550368);
nor I_32197 (I549859,I550385,I550029);
not I_32198 (I550440,I3042);
DFFARX1 I_32199 (I4241,I3035,I550440,I550466,);
DFFARX1 I_32200 (I550466,I3035,I550440,I550483,);
not I_32201 (I550432,I550483);
not I_32202 (I550505,I550466);
DFFARX1 I_32203 (I4253,I3035,I550440,I550531,);
nand I_32204 (I550539,I550531,I4250);
not I_32205 (I550556,I4250);
not I_32206 (I550573,I4241);
nand I_32207 (I550590,I4235,I4235);
and I_32208 (I550607,I4235,I4235);
not I_32209 (I550624,I4256);
nand I_32210 (I550641,I550624,I550573);
nor I_32211 (I550414,I550641,I550539);
nor I_32212 (I550672,I550556,I550641);
nand I_32213 (I550417,I550607,I550672);
not I_32214 (I550703,I4247);
nor I_32215 (I550720,I550703,I4235);
nor I_32216 (I550737,I550720,I4256);
nor I_32217 (I550754,I550505,I550737);
DFFARX1 I_32218 (I550754,I3035,I550440,I550426,);
not I_32219 (I550785,I550720);
DFFARX1 I_32220 (I550785,I3035,I550440,I550429,);
and I_32221 (I550423,I550531,I550720);
nor I_32222 (I550830,I550703,I4238);
and I_32223 (I550847,I550830,I4238);
or I_32224 (I550864,I550847,I4244);
DFFARX1 I_32225 (I550864,I3035,I550440,I550890,);
nor I_32226 (I550898,I550890,I550624);
DFFARX1 I_32227 (I550898,I3035,I550440,I550411,);
nand I_32228 (I550929,I550890,I550531);
nand I_32229 (I550946,I550624,I550929);
nor I_32230 (I550420,I550946,I550590);
not I_32231 (I551001,I3042);
DFFARX1 I_32232 (I667020,I3035,I551001,I551027,);
DFFARX1 I_32233 (I551027,I3035,I551001,I551044,);
not I_32234 (I550993,I551044);
not I_32235 (I551066,I551027);
DFFARX1 I_32236 (I667026,I3035,I551001,I551092,);
nand I_32237 (I551100,I551092,I667035);
not I_32238 (I551117,I667035);
not I_32239 (I551134,I667014);
nand I_32240 (I551151,I667017,I667017);
and I_32241 (I551168,I667017,I667017);
not I_32242 (I551185,I667029);
nand I_32243 (I551202,I551185,I551134);
nor I_32244 (I550975,I551202,I551100);
nor I_32245 (I551233,I551117,I551202);
nand I_32246 (I550978,I551168,I551233);
not I_32247 (I551264,I667023);
nor I_32248 (I551281,I551264,I667017);
nor I_32249 (I551298,I551281,I667029);
nor I_32250 (I551315,I551066,I551298);
DFFARX1 I_32251 (I551315,I3035,I551001,I550987,);
not I_32252 (I551346,I551281);
DFFARX1 I_32253 (I551346,I3035,I551001,I550990,);
and I_32254 (I550984,I551092,I551281);
nor I_32255 (I551391,I551264,I667038);
and I_32256 (I551408,I551391,I667014);
or I_32257 (I551425,I551408,I667032);
DFFARX1 I_32258 (I551425,I3035,I551001,I551451,);
nor I_32259 (I551459,I551451,I551185);
DFFARX1 I_32260 (I551459,I3035,I551001,I550972,);
nand I_32261 (I551490,I551451,I551092);
nand I_32262 (I551507,I551185,I551490);
nor I_32263 (I550981,I551507,I551151);
not I_32264 (I551562,I3042);
DFFARX1 I_32265 (I524520,I3035,I551562,I551588,);
DFFARX1 I_32266 (I551588,I3035,I551562,I551605,);
not I_32267 (I551554,I551605);
not I_32268 (I551627,I551588);
DFFARX1 I_32269 (I524547,I3035,I551562,I551653,);
nand I_32270 (I551661,I551653,I524538);
not I_32271 (I551678,I524538);
not I_32272 (I551695,I524520);
nand I_32273 (I551712,I524532,I524535);
and I_32274 (I551729,I524532,I524535);
not I_32275 (I551746,I524544);
nand I_32276 (I551763,I551746,I551695);
nor I_32277 (I551536,I551763,I551661);
nor I_32278 (I551794,I551678,I551763);
nand I_32279 (I551539,I551729,I551794);
not I_32280 (I551825,I524529);
nor I_32281 (I551842,I551825,I524532);
nor I_32282 (I551859,I551842,I524544);
nor I_32283 (I551876,I551627,I551859);
DFFARX1 I_32284 (I551876,I3035,I551562,I551548,);
not I_32285 (I551907,I551842);
DFFARX1 I_32286 (I551907,I3035,I551562,I551551,);
and I_32287 (I551545,I551653,I551842);
nor I_32288 (I551952,I551825,I524523);
and I_32289 (I551969,I551952,I524526);
or I_32290 (I551986,I551969,I524541);
DFFARX1 I_32291 (I551986,I3035,I551562,I552012,);
nor I_32292 (I552020,I552012,I551746);
DFFARX1 I_32293 (I552020,I3035,I551562,I551533,);
nand I_32294 (I552051,I552012,I551653);
nand I_32295 (I552068,I551746,I552051);
nor I_32296 (I551542,I552068,I551712);
not I_32297 (I552123,I3042);
DFFARX1 I_32298 (I461969,I3035,I552123,I552149,);
DFFARX1 I_32299 (I552149,I3035,I552123,I552166,);
not I_32300 (I552115,I552166);
not I_32301 (I552188,I552149);
DFFARX1 I_32302 (I461966,I3035,I552123,I552214,);
nand I_32303 (I552222,I552214,I461981);
not I_32304 (I552239,I461981);
not I_32305 (I552256,I461978);
nand I_32306 (I552273,I461975,I461963);
and I_32307 (I552290,I461975,I461963);
not I_32308 (I552307,I461960);
nand I_32309 (I552324,I552307,I552256);
nor I_32310 (I552097,I552324,I552222);
nor I_32311 (I552355,I552239,I552324);
nand I_32312 (I552100,I552290,I552355);
not I_32313 (I552386,I461966);
nor I_32314 (I552403,I552386,I461975);
nor I_32315 (I552420,I552403,I461960);
nor I_32316 (I552437,I552188,I552420);
DFFARX1 I_32317 (I552437,I3035,I552123,I552109,);
not I_32318 (I552468,I552403);
DFFARX1 I_32319 (I552468,I3035,I552123,I552112,);
and I_32320 (I552106,I552214,I552403);
nor I_32321 (I552513,I552386,I461972);
and I_32322 (I552530,I552513,I461960);
or I_32323 (I552547,I552530,I461963);
DFFARX1 I_32324 (I552547,I3035,I552123,I552573,);
nor I_32325 (I552581,I552573,I552307);
DFFARX1 I_32326 (I552581,I3035,I552123,I552094,);
nand I_32327 (I552612,I552573,I552214);
nand I_32328 (I552629,I552307,I552612);
nor I_32329 (I552103,I552629,I552273);
not I_32330 (I552684,I3042);
DFFARX1 I_32331 (I612765,I3035,I552684,I552710,);
DFFARX1 I_32332 (I552710,I3035,I552684,I552727,);
not I_32333 (I552676,I552727);
not I_32334 (I552749,I552710);
DFFARX1 I_32335 (I612756,I3035,I552684,I552775,);
nand I_32336 (I552783,I552775,I612753);
not I_32337 (I552800,I612753);
not I_32338 (I552817,I612762);
nand I_32339 (I552834,I612771,I612753);
and I_32340 (I552851,I612771,I612753);
not I_32341 (I552868,I612750);
nand I_32342 (I552885,I552868,I552817);
nor I_32343 (I552658,I552885,I552783);
nor I_32344 (I552916,I552800,I552885);
nand I_32345 (I552661,I552851,I552916);
not I_32346 (I552947,I612759);
nor I_32347 (I552964,I552947,I612771);
nor I_32348 (I552981,I552964,I612750);
nor I_32349 (I552998,I552749,I552981);
DFFARX1 I_32350 (I552998,I3035,I552684,I552670,);
not I_32351 (I553029,I552964);
DFFARX1 I_32352 (I553029,I3035,I552684,I552673,);
and I_32353 (I552667,I552775,I552964);
nor I_32354 (I553074,I552947,I612774);
and I_32355 (I553091,I553074,I612750);
or I_32356 (I553108,I553091,I612768);
DFFARX1 I_32357 (I553108,I3035,I552684,I553134,);
nor I_32358 (I553142,I553134,I552868);
DFFARX1 I_32359 (I553142,I3035,I552684,I552655,);
nand I_32360 (I553173,I553134,I552775);
nand I_32361 (I553190,I552868,I553173);
nor I_32362 (I552664,I553190,I552834);
not I_32363 (I553245,I3042);
DFFARX1 I_32364 (I125907,I3035,I553245,I553271,);
DFFARX1 I_32365 (I553271,I3035,I553245,I553288,);
not I_32366 (I553237,I553288);
not I_32367 (I553310,I553271);
DFFARX1 I_32368 (I125922,I3035,I553245,I553336,);
nand I_32369 (I553344,I553336,I125904);
not I_32370 (I553361,I125904);
not I_32371 (I553378,I125913);
nand I_32372 (I553395,I125919,I125910);
and I_32373 (I553412,I125919,I125910);
not I_32374 (I553429,I125907);
nand I_32375 (I553446,I553429,I553378);
nor I_32376 (I553219,I553446,I553344);
nor I_32377 (I553477,I553361,I553446);
nand I_32378 (I553222,I553412,I553477);
not I_32379 (I553508,I125904);
nor I_32380 (I553525,I553508,I125919);
nor I_32381 (I553542,I553525,I125907);
nor I_32382 (I553559,I553310,I553542);
DFFARX1 I_32383 (I553559,I3035,I553245,I553231,);
not I_32384 (I553590,I553525);
DFFARX1 I_32385 (I553590,I3035,I553245,I553234,);
and I_32386 (I553228,I553336,I553525);
nor I_32387 (I553635,I553508,I125928);
and I_32388 (I553652,I553635,I125925);
or I_32389 (I553669,I553652,I125916);
DFFARX1 I_32390 (I553669,I3035,I553245,I553695,);
nor I_32391 (I553703,I553695,I553429);
DFFARX1 I_32392 (I553703,I3035,I553245,I553216,);
nand I_32393 (I553734,I553695,I553336);
nand I_32394 (I553751,I553429,I553734);
nor I_32395 (I553225,I553751,I553395);
not I_32396 (I553806,I3042);
DFFARX1 I_32397 (I103892,I3035,I553806,I553832,);
DFFARX1 I_32398 (I553832,I3035,I553806,I553849,);
not I_32399 (I553798,I553849);
not I_32400 (I553871,I553832);
DFFARX1 I_32401 (I103907,I3035,I553806,I553897,);
nand I_32402 (I553905,I553897,I103889);
not I_32403 (I553922,I103889);
not I_32404 (I553939,I103898);
nand I_32405 (I553956,I103904,I103895);
and I_32406 (I553973,I103904,I103895);
not I_32407 (I553990,I103892);
nand I_32408 (I554007,I553990,I553939);
nor I_32409 (I553780,I554007,I553905);
nor I_32410 (I554038,I553922,I554007);
nand I_32411 (I553783,I553973,I554038);
not I_32412 (I554069,I103889);
nor I_32413 (I554086,I554069,I103904);
nor I_32414 (I554103,I554086,I103892);
nor I_32415 (I554120,I553871,I554103);
DFFARX1 I_32416 (I554120,I3035,I553806,I553792,);
not I_32417 (I554151,I554086);
DFFARX1 I_32418 (I554151,I3035,I553806,I553795,);
and I_32419 (I553789,I553897,I554086);
nor I_32420 (I554196,I554069,I103913);
and I_32421 (I554213,I554196,I103910);
or I_32422 (I554230,I554213,I103901);
DFFARX1 I_32423 (I554230,I3035,I553806,I554256,);
nor I_32424 (I554264,I554256,I553990);
DFFARX1 I_32425 (I554264,I3035,I553806,I553777,);
nand I_32426 (I554295,I554256,I553897);
nand I_32427 (I554312,I553990,I554295);
nor I_32428 (I553786,I554312,I553956);
not I_32429 (I554367,I3042);
DFFARX1 I_32430 (I714493,I3035,I554367,I554393,);
DFFARX1 I_32431 (I554393,I3035,I554367,I554410,);
not I_32432 (I554359,I554410);
not I_32433 (I554432,I554393);
DFFARX1 I_32434 (I714487,I3035,I554367,I554458,);
nand I_32435 (I554466,I554458,I714478);
not I_32436 (I554483,I714478);
not I_32437 (I554500,I714505);
nand I_32438 (I554517,I714490,I714499);
and I_32439 (I554534,I714490,I714499);
not I_32440 (I554551,I714484);
nand I_32441 (I554568,I554551,I554500);
nor I_32442 (I554341,I554568,I554466);
nor I_32443 (I554599,I554483,I554568);
nand I_32444 (I554344,I554534,I554599);
not I_32445 (I554630,I714502);
nor I_32446 (I554647,I554630,I714490);
nor I_32447 (I554664,I554647,I714484);
nor I_32448 (I554681,I554432,I554664);
DFFARX1 I_32449 (I554681,I3035,I554367,I554353,);
not I_32450 (I554712,I554647);
DFFARX1 I_32451 (I554712,I3035,I554367,I554356,);
and I_32452 (I554350,I554458,I554647);
nor I_32453 (I554757,I554630,I714496);
and I_32454 (I554774,I554757,I714478);
or I_32455 (I554791,I554774,I714481);
DFFARX1 I_32456 (I554791,I3035,I554367,I554817,);
nor I_32457 (I554825,I554817,I554551);
DFFARX1 I_32458 (I554825,I3035,I554367,I554338,);
nand I_32459 (I554856,I554817,I554458);
nand I_32460 (I554873,I554551,I554856);
nor I_32461 (I554347,I554873,I554517);
not I_32462 (I554928,I3042);
DFFARX1 I_32463 (I276701,I3035,I554928,I554954,);
DFFARX1 I_32464 (I554954,I3035,I554928,I554971,);
not I_32465 (I554920,I554971);
not I_32466 (I554993,I554954);
DFFARX1 I_32467 (I276689,I3035,I554928,I555019,);
nand I_32468 (I555027,I555019,I276695);
not I_32469 (I555044,I276695);
not I_32470 (I555061,I276692);
nand I_32471 (I555078,I276680,I276677);
and I_32472 (I555095,I276680,I276677);
not I_32473 (I555112,I276704);
nand I_32474 (I555129,I555112,I555061);
nor I_32475 (I554902,I555129,I555027);
nor I_32476 (I555160,I555044,I555129);
nand I_32477 (I554905,I555095,I555160);
not I_32478 (I555191,I276677);
nor I_32479 (I555208,I555191,I276680);
nor I_32480 (I555225,I555208,I276704);
nor I_32481 (I555242,I554993,I555225);
DFFARX1 I_32482 (I555242,I3035,I554928,I554914,);
not I_32483 (I555273,I555208);
DFFARX1 I_32484 (I555273,I3035,I554928,I554917,);
and I_32485 (I554911,I555019,I555208);
nor I_32486 (I555318,I555191,I276686);
and I_32487 (I555335,I555318,I276683);
or I_32488 (I555352,I555335,I276698);
DFFARX1 I_32489 (I555352,I3035,I554928,I555378,);
nor I_32490 (I555386,I555378,I555112);
DFFARX1 I_32491 (I555386,I3035,I554928,I554899,);
nand I_32492 (I555417,I555378,I555019);
nand I_32493 (I555434,I555112,I555417);
nor I_32494 (I554908,I555434,I555078);
not I_32495 (I555489,I3042);
DFFARX1 I_32496 (I371829,I3035,I555489,I555515,);
DFFARX1 I_32497 (I555515,I3035,I555489,I555532,);
not I_32498 (I555481,I555532);
not I_32499 (I555554,I555515);
DFFARX1 I_32500 (I371841,I3035,I555489,I555580,);
nand I_32501 (I555588,I555580,I371850);
not I_32502 (I555605,I371850);
not I_32503 (I555622,I371832);
nand I_32504 (I555639,I371835,I371826);
and I_32505 (I555656,I371835,I371826);
not I_32506 (I555673,I371844);
nand I_32507 (I555690,I555673,I555622);
nor I_32508 (I555463,I555690,I555588);
nor I_32509 (I555721,I555605,I555690);
nand I_32510 (I555466,I555656,I555721);
not I_32511 (I555752,I371847);
nor I_32512 (I555769,I555752,I371835);
nor I_32513 (I555786,I555769,I371844);
nor I_32514 (I555803,I555554,I555786);
DFFARX1 I_32515 (I555803,I3035,I555489,I555475,);
not I_32516 (I555834,I555769);
DFFARX1 I_32517 (I555834,I3035,I555489,I555478,);
and I_32518 (I555472,I555580,I555769);
nor I_32519 (I555879,I555752,I371826);
and I_32520 (I555896,I555879,I371838);
or I_32521 (I555913,I555896,I371829);
DFFARX1 I_32522 (I555913,I3035,I555489,I555939,);
nor I_32523 (I555947,I555939,I555673);
DFFARX1 I_32524 (I555947,I3035,I555489,I555460,);
nand I_32525 (I555978,I555939,I555580);
nand I_32526 (I555995,I555673,I555978);
nor I_32527 (I555469,I555995,I555639);
not I_32528 (I556050,I3042);
DFFARX1 I_32529 (I645711,I3035,I556050,I556076,);
DFFARX1 I_32530 (I556076,I3035,I556050,I556093,);
not I_32531 (I556042,I556093);
not I_32532 (I556115,I556076);
DFFARX1 I_32533 (I645702,I3035,I556050,I556141,);
nand I_32534 (I556149,I556141,I645699);
not I_32535 (I556166,I645699);
not I_32536 (I556183,I645708);
nand I_32537 (I556200,I645717,I645699);
and I_32538 (I556217,I645717,I645699);
not I_32539 (I556234,I645696);
nand I_32540 (I556251,I556234,I556183);
nor I_32541 (I556024,I556251,I556149);
nor I_32542 (I556282,I556166,I556251);
nand I_32543 (I556027,I556217,I556282);
not I_32544 (I556313,I645705);
nor I_32545 (I556330,I556313,I645717);
nor I_32546 (I556347,I556330,I645696);
nor I_32547 (I556364,I556115,I556347);
DFFARX1 I_32548 (I556364,I3035,I556050,I556036,);
not I_32549 (I556395,I556330);
DFFARX1 I_32550 (I556395,I3035,I556050,I556039,);
and I_32551 (I556033,I556141,I556330);
nor I_32552 (I556440,I556313,I645720);
and I_32553 (I556457,I556440,I645696);
or I_32554 (I556474,I556457,I645714);
DFFARX1 I_32555 (I556474,I3035,I556050,I556500,);
nor I_32556 (I556508,I556500,I556234);
DFFARX1 I_32557 (I556508,I3035,I556050,I556021,);
nand I_32558 (I556539,I556500,I556141);
nand I_32559 (I556556,I556234,I556539);
nor I_32560 (I556030,I556556,I556200);
not I_32561 (I556611,I3042);
DFFARX1 I_32562 (I239165,I3035,I556611,I556637,);
DFFARX1 I_32563 (I556637,I3035,I556611,I556654,);
not I_32564 (I556603,I556654);
not I_32565 (I556676,I556637);
DFFARX1 I_32566 (I239153,I3035,I556611,I556702,);
nand I_32567 (I556710,I556702,I239159);
not I_32568 (I556727,I239159);
not I_32569 (I556744,I239156);
nand I_32570 (I556761,I239144,I239141);
and I_32571 (I556778,I239144,I239141);
not I_32572 (I556795,I239168);
nand I_32573 (I556812,I556795,I556744);
nor I_32574 (I556585,I556812,I556710);
nor I_32575 (I556843,I556727,I556812);
nand I_32576 (I556588,I556778,I556843);
not I_32577 (I556874,I239141);
nor I_32578 (I556891,I556874,I239144);
nor I_32579 (I556908,I556891,I239168);
nor I_32580 (I556925,I556676,I556908);
DFFARX1 I_32581 (I556925,I3035,I556611,I556597,);
not I_32582 (I556956,I556891);
DFFARX1 I_32583 (I556956,I3035,I556611,I556600,);
and I_32584 (I556594,I556702,I556891);
nor I_32585 (I557001,I556874,I239150);
and I_32586 (I557018,I557001,I239147);
or I_32587 (I557035,I557018,I239162);
DFFARX1 I_32588 (I557035,I3035,I556611,I557061,);
nor I_32589 (I557069,I557061,I556795);
DFFARX1 I_32590 (I557069,I3035,I556611,I556582,);
nand I_32591 (I557100,I557061,I556702);
nand I_32592 (I557117,I556795,I557100);
nor I_32593 (I556591,I557117,I556761);
not I_32594 (I557172,I3042);
DFFARX1 I_32595 (I159279,I3035,I557172,I557198,);
DFFARX1 I_32596 (I557198,I3035,I557172,I557215,);
not I_32597 (I557164,I557215);
not I_32598 (I557237,I557198);
DFFARX1 I_32599 (I159276,I3035,I557172,I557263,);
nand I_32600 (I557271,I557263,I159270);
not I_32601 (I557288,I159270);
not I_32602 (I557305,I159267);
nand I_32603 (I557322,I159261,I159258);
and I_32604 (I557339,I159261,I159258);
not I_32605 (I557356,I159273);
nand I_32606 (I557373,I557356,I557305);
nor I_32607 (I557146,I557373,I557271);
nor I_32608 (I557404,I557288,I557373);
nand I_32609 (I557149,I557339,I557404);
not I_32610 (I557435,I159285);
nor I_32611 (I557452,I557435,I159261);
nor I_32612 (I557469,I557452,I159273);
nor I_32613 (I557486,I557237,I557469);
DFFARX1 I_32614 (I557486,I3035,I557172,I557158,);
not I_32615 (I557517,I557452);
DFFARX1 I_32616 (I557517,I3035,I557172,I557161,);
and I_32617 (I557155,I557263,I557452);
nor I_32618 (I557562,I557435,I159282);
and I_32619 (I557579,I557562,I159258);
or I_32620 (I557596,I557579,I159264);
DFFARX1 I_32621 (I557596,I3035,I557172,I557622,);
nor I_32622 (I557630,I557622,I557356);
DFFARX1 I_32623 (I557630,I3035,I557172,I557143,);
nand I_32624 (I557661,I557622,I557263);
nand I_32625 (I557678,I557356,I557661);
nor I_32626 (I557152,I557678,I557322);
not I_32627 (I557733,I3042);
DFFARX1 I_32628 (I625481,I3035,I557733,I557759,);
DFFARX1 I_32629 (I557759,I3035,I557733,I557776,);
not I_32630 (I557725,I557776);
not I_32631 (I557798,I557759);
DFFARX1 I_32632 (I625472,I3035,I557733,I557824,);
nand I_32633 (I557832,I557824,I625469);
not I_32634 (I557849,I625469);
not I_32635 (I557866,I625478);
nand I_32636 (I557883,I625487,I625469);
and I_32637 (I557900,I625487,I625469);
not I_32638 (I557917,I625466);
nand I_32639 (I557934,I557917,I557866);
nor I_32640 (I557707,I557934,I557832);
nor I_32641 (I557965,I557849,I557934);
nand I_32642 (I557710,I557900,I557965);
not I_32643 (I557996,I625475);
nor I_32644 (I558013,I557996,I625487);
nor I_32645 (I558030,I558013,I625466);
nor I_32646 (I558047,I557798,I558030);
DFFARX1 I_32647 (I558047,I3035,I557733,I557719,);
not I_32648 (I558078,I558013);
DFFARX1 I_32649 (I558078,I3035,I557733,I557722,);
and I_32650 (I557716,I557824,I558013);
nor I_32651 (I558123,I557996,I625490);
and I_32652 (I558140,I558123,I625466);
or I_32653 (I558157,I558140,I625484);
DFFARX1 I_32654 (I558157,I3035,I557733,I558183,);
nor I_32655 (I558191,I558183,I557917);
DFFARX1 I_32656 (I558191,I3035,I557733,I557704,);
nand I_32657 (I558222,I558183,I557824);
nand I_32658 (I558239,I557917,I558222);
nor I_32659 (I557713,I558239,I557883);
not I_32660 (I558294,I3042);
DFFARX1 I_32661 (I273437,I3035,I558294,I558320,);
DFFARX1 I_32662 (I558320,I3035,I558294,I558337,);
not I_32663 (I558286,I558337);
not I_32664 (I558359,I558320);
DFFARX1 I_32665 (I273425,I3035,I558294,I558385,);
nand I_32666 (I558393,I558385,I273431);
not I_32667 (I558410,I273431);
not I_32668 (I558427,I273428);
nand I_32669 (I558444,I273416,I273413);
and I_32670 (I558461,I273416,I273413);
not I_32671 (I558478,I273440);
nand I_32672 (I558495,I558478,I558427);
nor I_32673 (I558268,I558495,I558393);
nor I_32674 (I558526,I558410,I558495);
nand I_32675 (I558271,I558461,I558526);
not I_32676 (I558557,I273413);
nor I_32677 (I558574,I558557,I273416);
nor I_32678 (I558591,I558574,I273440);
nor I_32679 (I558608,I558359,I558591);
DFFARX1 I_32680 (I558608,I3035,I558294,I558280,);
not I_32681 (I558639,I558574);
DFFARX1 I_32682 (I558639,I3035,I558294,I558283,);
and I_32683 (I558277,I558385,I558574);
nor I_32684 (I558684,I558557,I273422);
and I_32685 (I558701,I558684,I273419);
or I_32686 (I558718,I558701,I273434);
DFFARX1 I_32687 (I558718,I3035,I558294,I558744,);
nor I_32688 (I558752,I558744,I558478);
DFFARX1 I_32689 (I558752,I3035,I558294,I558265,);
nand I_32690 (I558783,I558744,I558385);
nand I_32691 (I558800,I558478,I558783);
nor I_32692 (I558274,I558800,I558444);
not I_32693 (I558855,I3042);
DFFARX1 I_32694 (I637619,I3035,I558855,I558881,);
DFFARX1 I_32695 (I558881,I3035,I558855,I558898,);
not I_32696 (I558847,I558898);
not I_32697 (I558920,I558881);
DFFARX1 I_32698 (I637610,I3035,I558855,I558946,);
nand I_32699 (I558954,I558946,I637607);
not I_32700 (I558971,I637607);
not I_32701 (I558988,I637616);
nand I_32702 (I559005,I637625,I637607);
and I_32703 (I559022,I637625,I637607);
not I_32704 (I559039,I637604);
nand I_32705 (I559056,I559039,I558988);
nor I_32706 (I558829,I559056,I558954);
nor I_32707 (I559087,I558971,I559056);
nand I_32708 (I558832,I559022,I559087);
not I_32709 (I559118,I637613);
nor I_32710 (I559135,I559118,I637625);
nor I_32711 (I559152,I559135,I637604);
nor I_32712 (I559169,I558920,I559152);
DFFARX1 I_32713 (I559169,I3035,I558855,I558841,);
not I_32714 (I559200,I559135);
DFFARX1 I_32715 (I559200,I3035,I558855,I558844,);
and I_32716 (I558838,I558946,I559135);
nor I_32717 (I559245,I559118,I637628);
and I_32718 (I559262,I559245,I637604);
or I_32719 (I559279,I559262,I637622);
DFFARX1 I_32720 (I559279,I3035,I558855,I559305,);
nor I_32721 (I559313,I559305,I559039);
DFFARX1 I_32722 (I559313,I3035,I558855,I558826,);
nand I_32723 (I559344,I559305,I558946);
nand I_32724 (I559361,I559039,I559344);
nor I_32725 (I558835,I559361,I559005);
not I_32726 (I559416,I3042);
DFFARX1 I_32727 (I330210,I3035,I559416,I559442,);
DFFARX1 I_32728 (I559442,I3035,I559416,I559459,);
not I_32729 (I559408,I559459);
not I_32730 (I559481,I559442);
DFFARX1 I_32731 (I330225,I3035,I559416,I559507,);
nand I_32732 (I559515,I559507,I330216);
not I_32733 (I559532,I330216);
not I_32734 (I559549,I330222);
nand I_32735 (I559566,I330219,I330228);
and I_32736 (I559583,I330219,I330228);
not I_32737 (I559600,I330213);
nand I_32738 (I559617,I559600,I559549);
nor I_32739 (I559390,I559617,I559515);
nor I_32740 (I559648,I559532,I559617);
nand I_32741 (I559393,I559583,I559648);
not I_32742 (I559679,I330210);
nor I_32743 (I559696,I559679,I330219);
nor I_32744 (I559713,I559696,I330213);
nor I_32745 (I559730,I559481,I559713);
DFFARX1 I_32746 (I559730,I3035,I559416,I559402,);
not I_32747 (I559761,I559696);
DFFARX1 I_32748 (I559761,I3035,I559416,I559405,);
and I_32749 (I559399,I559507,I559696);
nor I_32750 (I559806,I559679,I330234);
and I_32751 (I559823,I559806,I330213);
or I_32752 (I559840,I559823,I330231);
DFFARX1 I_32753 (I559840,I3035,I559416,I559866,);
nor I_32754 (I559874,I559866,I559600);
DFFARX1 I_32755 (I559874,I3035,I559416,I559387,);
nand I_32756 (I559905,I559866,I559507);
nand I_32757 (I559922,I559600,I559905);
nor I_32758 (I559396,I559922,I559566);
not I_32759 (I559977,I3042);
DFFARX1 I_32760 (I718063,I3035,I559977,I560003,);
DFFARX1 I_32761 (I560003,I3035,I559977,I560020,);
not I_32762 (I559969,I560020);
not I_32763 (I560042,I560003);
DFFARX1 I_32764 (I718057,I3035,I559977,I560068,);
nand I_32765 (I560076,I560068,I718048);
not I_32766 (I560093,I718048);
not I_32767 (I560110,I718075);
nand I_32768 (I560127,I718060,I718069);
and I_32769 (I560144,I718060,I718069);
not I_32770 (I560161,I718054);
nand I_32771 (I560178,I560161,I560110);
nor I_32772 (I559951,I560178,I560076);
nor I_32773 (I560209,I560093,I560178);
nand I_32774 (I559954,I560144,I560209);
not I_32775 (I560240,I718072);
nor I_32776 (I560257,I560240,I718060);
nor I_32777 (I560274,I560257,I718054);
nor I_32778 (I560291,I560042,I560274);
DFFARX1 I_32779 (I560291,I3035,I559977,I559963,);
not I_32780 (I560322,I560257);
DFFARX1 I_32781 (I560322,I3035,I559977,I559966,);
and I_32782 (I559960,I560068,I560257);
nor I_32783 (I560367,I560240,I718066);
and I_32784 (I560384,I560367,I718048);
or I_32785 (I560401,I560384,I718051);
DFFARX1 I_32786 (I560401,I3035,I559977,I560427,);
nor I_32787 (I560435,I560427,I560161);
DFFARX1 I_32788 (I560435,I3035,I559977,I559948,);
nand I_32789 (I560466,I560427,I560068);
nand I_32790 (I560483,I560161,I560466);
nor I_32791 (I559957,I560483,I560127);
not I_32792 (I560538,I3042);
DFFARX1 I_32793 (I198277,I3035,I560538,I560564,);
DFFARX1 I_32794 (I560564,I3035,I560538,I560581,);
not I_32795 (I560530,I560581);
not I_32796 (I560603,I560564);
DFFARX1 I_32797 (I198274,I3035,I560538,I560629,);
nand I_32798 (I560637,I560629,I198268);
not I_32799 (I560654,I198268);
not I_32800 (I560671,I198265);
nand I_32801 (I560688,I198259,I198256);
and I_32802 (I560705,I198259,I198256);
not I_32803 (I560722,I198271);
nand I_32804 (I560739,I560722,I560671);
nor I_32805 (I560512,I560739,I560637);
nor I_32806 (I560770,I560654,I560739);
nand I_32807 (I560515,I560705,I560770);
not I_32808 (I560801,I198283);
nor I_32809 (I560818,I560801,I198259);
nor I_32810 (I560835,I560818,I198271);
nor I_32811 (I560852,I560603,I560835);
DFFARX1 I_32812 (I560852,I3035,I560538,I560524,);
not I_32813 (I560883,I560818);
DFFARX1 I_32814 (I560883,I3035,I560538,I560527,);
and I_32815 (I560521,I560629,I560818);
nor I_32816 (I560928,I560801,I198280);
and I_32817 (I560945,I560928,I198256);
or I_32818 (I560962,I560945,I198262);
DFFARX1 I_32819 (I560962,I3035,I560538,I560988,);
nor I_32820 (I560996,I560988,I560722);
DFFARX1 I_32821 (I560996,I3035,I560538,I560509,);
nand I_32822 (I561027,I560988,I560629);
nand I_32823 (I561044,I560722,I561027);
nor I_32824 (I560518,I561044,I560688);
not I_32825 (I561099,I3042);
DFFARX1 I_32826 (I143162,I3035,I561099,I561125,);
DFFARX1 I_32827 (I561125,I3035,I561099,I561142,);
not I_32828 (I561091,I561142);
not I_32829 (I561164,I561125);
DFFARX1 I_32830 (I143177,I3035,I561099,I561190,);
nand I_32831 (I561198,I561190,I143159);
not I_32832 (I561215,I143159);
not I_32833 (I561232,I143168);
nand I_32834 (I561249,I143174,I143165);
and I_32835 (I561266,I143174,I143165);
not I_32836 (I561283,I143162);
nand I_32837 (I561300,I561283,I561232);
nor I_32838 (I561073,I561300,I561198);
nor I_32839 (I561331,I561215,I561300);
nand I_32840 (I561076,I561266,I561331);
not I_32841 (I561362,I143159);
nor I_32842 (I561379,I561362,I143174);
nor I_32843 (I561396,I561379,I143162);
nor I_32844 (I561413,I561164,I561396);
DFFARX1 I_32845 (I561413,I3035,I561099,I561085,);
not I_32846 (I561444,I561379);
DFFARX1 I_32847 (I561444,I3035,I561099,I561088,);
and I_32848 (I561082,I561190,I561379);
nor I_32849 (I561489,I561362,I143183);
and I_32850 (I561506,I561489,I143180);
or I_32851 (I561523,I561506,I143171);
DFFARX1 I_32852 (I561523,I3035,I561099,I561549,);
nor I_32853 (I561557,I561549,I561283);
DFFARX1 I_32854 (I561557,I3035,I561099,I561070,);
nand I_32855 (I561588,I561549,I561190);
nand I_32856 (I561605,I561283,I561588);
nor I_32857 (I561079,I561605,I561249);
not I_32858 (I561660,I3042);
DFFARX1 I_32859 (I403619,I3035,I561660,I561686,);
DFFARX1 I_32860 (I561686,I3035,I561660,I561703,);
not I_32861 (I561652,I561703);
not I_32862 (I561725,I561686);
DFFARX1 I_32863 (I403631,I3035,I561660,I561751,);
nand I_32864 (I561759,I561751,I403640);
not I_32865 (I561776,I403640);
not I_32866 (I561793,I403622);
nand I_32867 (I561810,I403625,I403616);
and I_32868 (I561827,I403625,I403616);
not I_32869 (I561844,I403634);
nand I_32870 (I561861,I561844,I561793);
nor I_32871 (I561634,I561861,I561759);
nor I_32872 (I561892,I561776,I561861);
nand I_32873 (I561637,I561827,I561892);
not I_32874 (I561923,I403637);
nor I_32875 (I561940,I561923,I403625);
nor I_32876 (I561957,I561940,I403634);
nor I_32877 (I561974,I561725,I561957);
DFFARX1 I_32878 (I561974,I3035,I561660,I561646,);
not I_32879 (I562005,I561940);
DFFARX1 I_32880 (I562005,I3035,I561660,I561649,);
and I_32881 (I561643,I561751,I561940);
nor I_32882 (I562050,I561923,I403616);
and I_32883 (I562067,I562050,I403628);
or I_32884 (I562084,I562067,I403619);
DFFARX1 I_32885 (I562084,I3035,I561660,I562110,);
nor I_32886 (I562118,I562110,I561844);
DFFARX1 I_32887 (I562118,I3035,I561660,I561631,);
nand I_32888 (I562149,I562110,I561751);
nand I_32889 (I562166,I561844,I562149);
nor I_32890 (I561640,I562166,I561810);
not I_32891 (I562221,I3042);
DFFARX1 I_32892 (I41018,I3035,I562221,I562247,);
DFFARX1 I_32893 (I562247,I3035,I562221,I562264,);
not I_32894 (I562213,I562264);
not I_32895 (I562286,I562247);
DFFARX1 I_32896 (I41006,I3035,I562221,I562312,);
nand I_32897 (I562320,I562312,I41021);
not I_32898 (I562337,I41021);
not I_32899 (I562354,I41009);
nand I_32900 (I562371,I41030,I41024);
and I_32901 (I562388,I41030,I41024);
not I_32902 (I562405,I41012);
nand I_32903 (I562422,I562405,I562354);
nor I_32904 (I562195,I562422,I562320);
nor I_32905 (I562453,I562337,I562422);
nand I_32906 (I562198,I562388,I562453);
not I_32907 (I562484,I41015);
nor I_32908 (I562501,I562484,I41030);
nor I_32909 (I562518,I562501,I41012);
nor I_32910 (I562535,I562286,I562518);
DFFARX1 I_32911 (I562535,I3035,I562221,I562207,);
not I_32912 (I562566,I562501);
DFFARX1 I_32913 (I562566,I3035,I562221,I562210,);
and I_32914 (I562204,I562312,I562501);
nor I_32915 (I562611,I562484,I41009);
and I_32916 (I562628,I562611,I41006);
or I_32917 (I562645,I562628,I41027);
DFFARX1 I_32918 (I562645,I3035,I562221,I562671,);
nor I_32919 (I562679,I562671,I562405);
DFFARX1 I_32920 (I562679,I3035,I562221,I562192,);
nand I_32921 (I562710,I562671,I562312);
nand I_32922 (I562727,I562405,I562710);
nor I_32923 (I562201,I562727,I562371);
not I_32924 (I562782,I3042);
DFFARX1 I_32925 (I27322,I3035,I562782,I562808,);
DFFARX1 I_32926 (I562808,I3035,I562782,I562825,);
not I_32927 (I562774,I562825);
not I_32928 (I562847,I562808);
DFFARX1 I_32929 (I27307,I3035,I562782,I562873,);
nand I_32930 (I562881,I562873,I27319);
not I_32931 (I562898,I27319);
not I_32932 (I562915,I27325);
nand I_32933 (I562932,I27313,I27304);
and I_32934 (I562949,I27313,I27304);
not I_32935 (I562966,I27310);
nand I_32936 (I562983,I562966,I562915);
nor I_32937 (I562756,I562983,I562881);
nor I_32938 (I563014,I562898,I562983);
nand I_32939 (I562759,I562949,I563014);
not I_32940 (I563045,I27316);
nor I_32941 (I563062,I563045,I27313);
nor I_32942 (I563079,I563062,I27310);
nor I_32943 (I563096,I562847,I563079);
DFFARX1 I_32944 (I563096,I3035,I562782,I562768,);
not I_32945 (I563127,I563062);
DFFARX1 I_32946 (I563127,I3035,I562782,I562771,);
and I_32947 (I562765,I562873,I563062);
nor I_32948 (I563172,I563045,I27304);
and I_32949 (I563189,I563172,I27328);
or I_32950 (I563206,I563189,I27307);
DFFARX1 I_32951 (I563206,I3035,I562782,I563232,);
nor I_32952 (I563240,I563232,I562966);
DFFARX1 I_32953 (I563240,I3035,I562782,I562753,);
nand I_32954 (I563271,I563232,I562873);
nand I_32955 (I563288,I562966,I563271);
nor I_32956 (I562762,I563288,I562932);
not I_32957 (I563343,I3042);
DFFARX1 I_32958 (I253309,I3035,I563343,I563369,);
DFFARX1 I_32959 (I563369,I3035,I563343,I563386,);
not I_32960 (I563335,I563386);
not I_32961 (I563408,I563369);
DFFARX1 I_32962 (I253297,I3035,I563343,I563434,);
nand I_32963 (I563442,I563434,I253303);
not I_32964 (I563459,I253303);
not I_32965 (I563476,I253300);
nand I_32966 (I563493,I253288,I253285);
and I_32967 (I563510,I253288,I253285);
not I_32968 (I563527,I253312);
nand I_32969 (I563544,I563527,I563476);
nor I_32970 (I563317,I563544,I563442);
nor I_32971 (I563575,I563459,I563544);
nand I_32972 (I563320,I563510,I563575);
not I_32973 (I563606,I253285);
nor I_32974 (I563623,I563606,I253288);
nor I_32975 (I563640,I563623,I253312);
nor I_32976 (I563657,I563408,I563640);
DFFARX1 I_32977 (I563657,I3035,I563343,I563329,);
not I_32978 (I563688,I563623);
DFFARX1 I_32979 (I563688,I3035,I563343,I563332,);
and I_32980 (I563326,I563434,I563623);
nor I_32981 (I563733,I563606,I253294);
and I_32982 (I563750,I563733,I253291);
or I_32983 (I563767,I563750,I253306);
DFFARX1 I_32984 (I563767,I3035,I563343,I563793,);
nor I_32985 (I563801,I563793,I563527);
DFFARX1 I_32986 (I563801,I3035,I563343,I563314,);
nand I_32987 (I563832,I563793,I563434);
nand I_32988 (I563849,I563527,I563832);
nor I_32989 (I563323,I563849,I563493);
not I_32990 (I563904,I3042);
DFFARX1 I_32991 (I534210,I3035,I563904,I563930,);
DFFARX1 I_32992 (I563930,I3035,I563904,I563947,);
not I_32993 (I563896,I563947);
not I_32994 (I563969,I563930);
DFFARX1 I_32995 (I534237,I3035,I563904,I563995,);
nand I_32996 (I564003,I563995,I534228);
not I_32997 (I564020,I534228);
not I_32998 (I564037,I534210);
nand I_32999 (I564054,I534222,I534225);
and I_33000 (I564071,I534222,I534225);
not I_33001 (I564088,I534234);
nand I_33002 (I564105,I564088,I564037);
nor I_33003 (I563878,I564105,I564003);
nor I_33004 (I564136,I564020,I564105);
nand I_33005 (I563881,I564071,I564136);
not I_33006 (I564167,I534219);
nor I_33007 (I564184,I564167,I534222);
nor I_33008 (I564201,I564184,I534234);
nor I_33009 (I564218,I563969,I564201);
DFFARX1 I_33010 (I564218,I3035,I563904,I563890,);
not I_33011 (I564249,I564184);
DFFARX1 I_33012 (I564249,I3035,I563904,I563893,);
and I_33013 (I563887,I563995,I564184);
nor I_33014 (I564294,I564167,I534213);
and I_33015 (I564311,I564294,I534216);
or I_33016 (I564328,I564311,I534231);
DFFARX1 I_33017 (I564328,I3035,I563904,I564354,);
nor I_33018 (I564362,I564354,I564088);
DFFARX1 I_33019 (I564362,I3035,I563904,I563875,);
nand I_33020 (I564393,I564354,I563995);
nand I_33021 (I564410,I564088,I564393);
nor I_33022 (I563884,I564410,I564054);
not I_33023 (I564465,I3042);
DFFARX1 I_33024 (I172981,I3035,I564465,I564491,);
DFFARX1 I_33025 (I564491,I3035,I564465,I564508,);
not I_33026 (I564457,I564508);
not I_33027 (I564530,I564491);
DFFARX1 I_33028 (I172978,I3035,I564465,I564556,);
nand I_33029 (I564564,I564556,I172972);
not I_33030 (I564581,I172972);
not I_33031 (I564598,I172969);
nand I_33032 (I564615,I172963,I172960);
and I_33033 (I564632,I172963,I172960);
not I_33034 (I564649,I172975);
nand I_33035 (I564666,I564649,I564598);
nor I_33036 (I564439,I564666,I564564);
nor I_33037 (I564697,I564581,I564666);
nand I_33038 (I564442,I564632,I564697);
not I_33039 (I564728,I172987);
nor I_33040 (I564745,I564728,I172963);
nor I_33041 (I564762,I564745,I172975);
nor I_33042 (I564779,I564530,I564762);
DFFARX1 I_33043 (I564779,I3035,I564465,I564451,);
not I_33044 (I564810,I564745);
DFFARX1 I_33045 (I564810,I3035,I564465,I564454,);
and I_33046 (I564448,I564556,I564745);
nor I_33047 (I564855,I564728,I172984);
and I_33048 (I564872,I564855,I172960);
or I_33049 (I564889,I564872,I172966);
DFFARX1 I_33050 (I564889,I3035,I564465,I564915,);
nor I_33051 (I564923,I564915,I564649);
DFFARX1 I_33052 (I564923,I3035,I564465,I564436,);
nand I_33053 (I564954,I564915,I564556);
nand I_33054 (I564971,I564649,I564954);
nor I_33055 (I564445,I564971,I564615);
not I_33056 (I565026,I3042);
DFFARX1 I_33057 (I702593,I3035,I565026,I565052,);
DFFARX1 I_33058 (I565052,I3035,I565026,I565069,);
not I_33059 (I565018,I565069);
not I_33060 (I565091,I565052);
DFFARX1 I_33061 (I702587,I3035,I565026,I565117,);
nand I_33062 (I565125,I565117,I702578);
not I_33063 (I565142,I702578);
not I_33064 (I565159,I702605);
nand I_33065 (I565176,I702590,I702599);
and I_33066 (I565193,I702590,I702599);
not I_33067 (I565210,I702584);
nand I_33068 (I565227,I565210,I565159);
nor I_33069 (I565000,I565227,I565125);
nor I_33070 (I565258,I565142,I565227);
nand I_33071 (I565003,I565193,I565258);
not I_33072 (I565289,I702602);
nor I_33073 (I565306,I565289,I702590);
nor I_33074 (I565323,I565306,I702584);
nor I_33075 (I565340,I565091,I565323);
DFFARX1 I_33076 (I565340,I3035,I565026,I565012,);
not I_33077 (I565371,I565306);
DFFARX1 I_33078 (I565371,I3035,I565026,I565015,);
and I_33079 (I565009,I565117,I565306);
nor I_33080 (I565416,I565289,I702596);
and I_33081 (I565433,I565416,I702578);
or I_33082 (I565450,I565433,I702581);
DFFARX1 I_33083 (I565450,I3035,I565026,I565476,);
nor I_33084 (I565484,I565476,I565210);
DFFARX1 I_33085 (I565484,I3035,I565026,I564997,);
nand I_33086 (I565515,I565476,I565117);
nand I_33087 (I565532,I565210,I565515);
nor I_33088 (I565006,I565532,I565176);
not I_33089 (I565587,I3042);
DFFARX1 I_33090 (I642821,I3035,I565587,I565613,);
DFFARX1 I_33091 (I565613,I3035,I565587,I565630,);
not I_33092 (I565579,I565630);
not I_33093 (I565652,I565613);
DFFARX1 I_33094 (I642812,I3035,I565587,I565678,);
nand I_33095 (I565686,I565678,I642809);
not I_33096 (I565703,I642809);
not I_33097 (I565720,I642818);
nand I_33098 (I565737,I642827,I642809);
and I_33099 (I565754,I642827,I642809);
not I_33100 (I565771,I642806);
nand I_33101 (I565788,I565771,I565720);
nor I_33102 (I565561,I565788,I565686);
nor I_33103 (I565819,I565703,I565788);
nand I_33104 (I565564,I565754,I565819);
not I_33105 (I565850,I642815);
nor I_33106 (I565867,I565850,I642827);
nor I_33107 (I565884,I565867,I642806);
nor I_33108 (I565901,I565652,I565884);
DFFARX1 I_33109 (I565901,I3035,I565587,I565573,);
not I_33110 (I565932,I565867);
DFFARX1 I_33111 (I565932,I3035,I565587,I565576,);
and I_33112 (I565570,I565678,I565867);
nor I_33113 (I565977,I565850,I642830);
and I_33114 (I565994,I565977,I642806);
or I_33115 (I566011,I565994,I642824);
DFFARX1 I_33116 (I566011,I3035,I565587,I566037,);
nor I_33117 (I566045,I566037,I565771);
DFFARX1 I_33118 (I566045,I3035,I565587,I565558,);
nand I_33119 (I566076,I566037,I565678);
nand I_33120 (I566093,I565771,I566076);
nor I_33121 (I565567,I566093,I565737);
not I_33122 (I566148,I3042);
DFFARX1 I_33123 (I468293,I3035,I566148,I566174,);
DFFARX1 I_33124 (I566174,I3035,I566148,I566191,);
not I_33125 (I566140,I566191);
not I_33126 (I566213,I566174);
DFFARX1 I_33127 (I468290,I3035,I566148,I566239,);
nand I_33128 (I566247,I566239,I468305);
not I_33129 (I566264,I468305);
not I_33130 (I566281,I468302);
nand I_33131 (I566298,I468299,I468287);
and I_33132 (I566315,I468299,I468287);
not I_33133 (I566332,I468284);
nand I_33134 (I566349,I566332,I566281);
nor I_33135 (I566122,I566349,I566247);
nor I_33136 (I566380,I566264,I566349);
nand I_33137 (I566125,I566315,I566380);
not I_33138 (I566411,I468290);
nor I_33139 (I566428,I566411,I468299);
nor I_33140 (I566445,I566428,I468284);
nor I_33141 (I566462,I566213,I566445);
DFFARX1 I_33142 (I566462,I3035,I566148,I566134,);
not I_33143 (I566493,I566428);
DFFARX1 I_33144 (I566493,I3035,I566148,I566137,);
and I_33145 (I566131,I566239,I566428);
nor I_33146 (I566538,I566411,I468296);
and I_33147 (I566555,I566538,I468284);
or I_33148 (I566572,I566555,I468287);
DFFARX1 I_33149 (I566572,I3035,I566148,I566598,);
nor I_33150 (I566606,I566598,I566332);
DFFARX1 I_33151 (I566606,I3035,I566148,I566119,);
nand I_33152 (I566637,I566598,I566239);
nand I_33153 (I566654,I566332,I566637);
nor I_33154 (I566128,I566654,I566298);
not I_33155 (I566709,I3042);
DFFARX1 I_33156 (I377609,I3035,I566709,I566735,);
DFFARX1 I_33157 (I566735,I3035,I566709,I566752,);
not I_33158 (I566701,I566752);
not I_33159 (I566774,I566735);
DFFARX1 I_33160 (I377621,I3035,I566709,I566800,);
nand I_33161 (I566808,I566800,I377630);
not I_33162 (I566825,I377630);
not I_33163 (I566842,I377612);
nand I_33164 (I566859,I377615,I377606);
and I_33165 (I566876,I377615,I377606);
not I_33166 (I566893,I377624);
nand I_33167 (I566910,I566893,I566842);
nor I_33168 (I566683,I566910,I566808);
nor I_33169 (I566941,I566825,I566910);
nand I_33170 (I566686,I566876,I566941);
not I_33171 (I566972,I377627);
nor I_33172 (I566989,I566972,I377615);
nor I_33173 (I567006,I566989,I377624);
nor I_33174 (I567023,I566774,I567006);
DFFARX1 I_33175 (I567023,I3035,I566709,I566695,);
not I_33176 (I567054,I566989);
DFFARX1 I_33177 (I567054,I3035,I566709,I566698,);
and I_33178 (I566692,I566800,I566989);
nor I_33179 (I567099,I566972,I377606);
and I_33180 (I567116,I567099,I377618);
or I_33181 (I567133,I567116,I377609);
DFFARX1 I_33182 (I567133,I3035,I566709,I567159,);
nor I_33183 (I567167,I567159,I566893);
DFFARX1 I_33184 (I567167,I3035,I566709,I566680,);
nand I_33185 (I567198,I567159,I566800);
nand I_33186 (I567215,I566893,I567198);
nor I_33187 (I566689,I567215,I566859);
not I_33188 (I567270,I3042);
DFFARX1 I_33189 (I350443,I3035,I567270,I567296,);
DFFARX1 I_33190 (I567296,I3035,I567270,I567313,);
not I_33191 (I567262,I567313);
not I_33192 (I567335,I567296);
DFFARX1 I_33193 (I350455,I3035,I567270,I567361,);
nand I_33194 (I567369,I567361,I350464);
not I_33195 (I567386,I350464);
not I_33196 (I567403,I350446);
nand I_33197 (I567420,I350449,I350440);
and I_33198 (I567437,I350449,I350440);
not I_33199 (I567454,I350458);
nand I_33200 (I567471,I567454,I567403);
nor I_33201 (I567244,I567471,I567369);
nor I_33202 (I567502,I567386,I567471);
nand I_33203 (I567247,I567437,I567502);
not I_33204 (I567533,I350461);
nor I_33205 (I567550,I567533,I350449);
nor I_33206 (I567567,I567550,I350458);
nor I_33207 (I567584,I567335,I567567);
DFFARX1 I_33208 (I567584,I3035,I567270,I567256,);
not I_33209 (I567615,I567550);
DFFARX1 I_33210 (I567615,I3035,I567270,I567259,);
and I_33211 (I567253,I567361,I567550);
nor I_33212 (I567660,I567533,I350440);
and I_33213 (I567677,I567660,I350452);
or I_33214 (I567694,I567677,I350443);
DFFARX1 I_33215 (I567694,I3035,I567270,I567720,);
nor I_33216 (I567728,I567720,I567454);
DFFARX1 I_33217 (I567728,I3035,I567270,I567241,);
nand I_33218 (I567759,I567720,I567361);
nand I_33219 (I567776,I567454,I567759);
nor I_33220 (I567250,I567776,I567420);
not I_33221 (I567831,I3042);
DFFARX1 I_33222 (I314026,I3035,I567831,I567857,);
DFFARX1 I_33223 (I567857,I3035,I567831,I567874,);
not I_33224 (I567823,I567874);
not I_33225 (I567896,I567857);
DFFARX1 I_33226 (I314041,I3035,I567831,I567922,);
nand I_33227 (I567930,I567922,I314032);
not I_33228 (I567947,I314032);
not I_33229 (I567964,I314038);
nand I_33230 (I567981,I314035,I314044);
and I_33231 (I567998,I314035,I314044);
not I_33232 (I568015,I314029);
nand I_33233 (I568032,I568015,I567964);
nor I_33234 (I567805,I568032,I567930);
nor I_33235 (I568063,I567947,I568032);
nand I_33236 (I567808,I567998,I568063);
not I_33237 (I568094,I314026);
nor I_33238 (I568111,I568094,I314035);
nor I_33239 (I568128,I568111,I314029);
nor I_33240 (I568145,I567896,I568128);
DFFARX1 I_33241 (I568145,I3035,I567831,I567817,);
not I_33242 (I568176,I568111);
DFFARX1 I_33243 (I568176,I3035,I567831,I567820,);
and I_33244 (I567814,I567922,I568111);
nor I_33245 (I568221,I568094,I314050);
and I_33246 (I568238,I568221,I314029);
or I_33247 (I568255,I568238,I314047);
DFFARX1 I_33248 (I568255,I3035,I567831,I568281,);
nor I_33249 (I568289,I568281,I568015);
DFFARX1 I_33250 (I568289,I3035,I567831,I567802,);
nand I_33251 (I568320,I568281,I567922);
nand I_33252 (I568337,I568015,I568320);
nor I_33253 (I567811,I568337,I567981);
not I_33254 (I568392,I3042);
DFFARX1 I_33255 (I692143,I3035,I568392,I568418,);
DFFARX1 I_33256 (I568418,I3035,I568392,I568435,);
not I_33257 (I568384,I568435);
not I_33258 (I568457,I568418);
DFFARX1 I_33259 (I692140,I3035,I568392,I568483,);
nand I_33260 (I568491,I568483,I692146);
not I_33261 (I568508,I692146);
not I_33262 (I568525,I692155);
nand I_33263 (I568542,I692149,I692143);
and I_33264 (I568559,I692149,I692143);
not I_33265 (I568576,I692161);
nand I_33266 (I568593,I568576,I568525);
nor I_33267 (I568366,I568593,I568491);
nor I_33268 (I568624,I568508,I568593);
nand I_33269 (I568369,I568559,I568624);
not I_33270 (I568655,I692158);
nor I_33271 (I568672,I568655,I692149);
nor I_33272 (I568689,I568672,I692161);
nor I_33273 (I568706,I568457,I568689);
DFFARX1 I_33274 (I568706,I3035,I568392,I568378,);
not I_33275 (I568737,I568672);
DFFARX1 I_33276 (I568737,I3035,I568392,I568381,);
and I_33277 (I568375,I568483,I568672);
nor I_33278 (I568782,I568655,I692152);
and I_33279 (I568799,I568782,I692164);
or I_33280 (I568816,I568799,I692140);
DFFARX1 I_33281 (I568816,I3035,I568392,I568842,);
nor I_33282 (I568850,I568842,I568576);
DFFARX1 I_33283 (I568850,I3035,I568392,I568363,);
nand I_33284 (I568881,I568842,I568483);
nand I_33285 (I568898,I568576,I568881);
nor I_33286 (I568372,I568898,I568542);
not I_33287 (I568953,I3042);
DFFARX1 I_33288 (I537440,I3035,I568953,I568979,);
DFFARX1 I_33289 (I568979,I3035,I568953,I568996,);
not I_33290 (I568945,I568996);
not I_33291 (I569018,I568979);
DFFARX1 I_33292 (I537467,I3035,I568953,I569044,);
nand I_33293 (I569052,I569044,I537458);
not I_33294 (I569069,I537458);
not I_33295 (I569086,I537440);
nand I_33296 (I569103,I537452,I537455);
and I_33297 (I569120,I537452,I537455);
not I_33298 (I569137,I537464);
nand I_33299 (I569154,I569137,I569086);
nor I_33300 (I568927,I569154,I569052);
nor I_33301 (I569185,I569069,I569154);
nand I_33302 (I568930,I569120,I569185);
not I_33303 (I569216,I537449);
nor I_33304 (I569233,I569216,I537452);
nor I_33305 (I569250,I569233,I537464);
nor I_33306 (I569267,I569018,I569250);
DFFARX1 I_33307 (I569267,I3035,I568953,I568939,);
not I_33308 (I569298,I569233);
DFFARX1 I_33309 (I569298,I3035,I568953,I568942,);
and I_33310 (I568936,I569044,I569233);
nor I_33311 (I569343,I569216,I537443);
and I_33312 (I569360,I569343,I537446);
or I_33313 (I569377,I569360,I537461);
DFFARX1 I_33314 (I569377,I3035,I568953,I569403,);
nor I_33315 (I569411,I569403,I569137);
DFFARX1 I_33316 (I569411,I3035,I568953,I568924,);
nand I_33317 (I569442,I569403,I569044);
nand I_33318 (I569459,I569137,I569442);
nor I_33319 (I568933,I569459,I569103);
not I_33320 (I569514,I3042);
DFFARX1 I_33321 (I160333,I3035,I569514,I569540,);
DFFARX1 I_33322 (I569540,I3035,I569514,I569557,);
not I_33323 (I569506,I569557);
not I_33324 (I569579,I569540);
DFFARX1 I_33325 (I160330,I3035,I569514,I569605,);
nand I_33326 (I569613,I569605,I160324);
not I_33327 (I569630,I160324);
not I_33328 (I569647,I160321);
nand I_33329 (I569664,I160315,I160312);
and I_33330 (I569681,I160315,I160312);
not I_33331 (I569698,I160327);
nand I_33332 (I569715,I569698,I569647);
nor I_33333 (I569488,I569715,I569613);
nor I_33334 (I569746,I569630,I569715);
nand I_33335 (I569491,I569681,I569746);
not I_33336 (I569777,I160339);
nor I_33337 (I569794,I569777,I160315);
nor I_33338 (I569811,I569794,I160327);
nor I_33339 (I569828,I569579,I569811);
DFFARX1 I_33340 (I569828,I3035,I569514,I569500,);
not I_33341 (I569859,I569794);
DFFARX1 I_33342 (I569859,I3035,I569514,I569503,);
and I_33343 (I569497,I569605,I569794);
nor I_33344 (I569904,I569777,I160336);
and I_33345 (I569921,I569904,I160312);
or I_33346 (I569938,I569921,I160318);
DFFARX1 I_33347 (I569938,I3035,I569514,I569964,);
nor I_33348 (I569972,I569964,I569698);
DFFARX1 I_33349 (I569972,I3035,I569514,I569485,);
nand I_33350 (I570003,I569964,I569605);
nand I_33351 (I570020,I569698,I570003);
nor I_33352 (I569494,I570020,I569664);
not I_33353 (I570075,I3042);
DFFARX1 I_33354 (I452483,I3035,I570075,I570101,);
DFFARX1 I_33355 (I570101,I3035,I570075,I570118,);
not I_33356 (I570067,I570118);
not I_33357 (I570140,I570101);
DFFARX1 I_33358 (I452480,I3035,I570075,I570166,);
nand I_33359 (I570174,I570166,I452495);
not I_33360 (I570191,I452495);
not I_33361 (I570208,I452492);
nand I_33362 (I570225,I452489,I452477);
and I_33363 (I570242,I452489,I452477);
not I_33364 (I570259,I452474);
nand I_33365 (I570276,I570259,I570208);
nor I_33366 (I570049,I570276,I570174);
nor I_33367 (I570307,I570191,I570276);
nand I_33368 (I570052,I570242,I570307);
not I_33369 (I570338,I452480);
nor I_33370 (I570355,I570338,I452489);
nor I_33371 (I570372,I570355,I452474);
nor I_33372 (I570389,I570140,I570372);
DFFARX1 I_33373 (I570389,I3035,I570075,I570061,);
not I_33374 (I570420,I570355);
DFFARX1 I_33375 (I570420,I3035,I570075,I570064,);
and I_33376 (I570058,I570166,I570355);
nor I_33377 (I570465,I570338,I452486);
and I_33378 (I570482,I570465,I452474);
or I_33379 (I570499,I570482,I452477);
DFFARX1 I_33380 (I570499,I3035,I570075,I570525,);
nor I_33381 (I570533,I570525,I570259);
DFFARX1 I_33382 (I570533,I3035,I570075,I570046,);
nand I_33383 (I570564,I570525,I570166);
nand I_33384 (I570581,I570259,I570564);
nor I_33385 (I570055,I570581,I570225);
not I_33386 (I570636,I3042);
DFFARX1 I_33387 (I512246,I3035,I570636,I570662,);
DFFARX1 I_33388 (I570662,I3035,I570636,I570679,);
not I_33389 (I570628,I570679);
not I_33390 (I570701,I570662);
DFFARX1 I_33391 (I512273,I3035,I570636,I570727,);
nand I_33392 (I570735,I570727,I512264);
not I_33393 (I570752,I512264);
not I_33394 (I570769,I512246);
nand I_33395 (I570786,I512258,I512261);
and I_33396 (I570803,I512258,I512261);
not I_33397 (I570820,I512270);
nand I_33398 (I570837,I570820,I570769);
nor I_33399 (I570610,I570837,I570735);
nor I_33400 (I570868,I570752,I570837);
nand I_33401 (I570613,I570803,I570868);
not I_33402 (I570899,I512255);
nor I_33403 (I570916,I570899,I512258);
nor I_33404 (I570933,I570916,I512270);
nor I_33405 (I570950,I570701,I570933);
DFFARX1 I_33406 (I570950,I3035,I570636,I570622,);
not I_33407 (I570981,I570916);
DFFARX1 I_33408 (I570981,I3035,I570636,I570625,);
and I_33409 (I570619,I570727,I570916);
nor I_33410 (I571026,I570899,I512249);
and I_33411 (I571043,I571026,I512252);
or I_33412 (I571060,I571043,I512267);
DFFARX1 I_33413 (I571060,I3035,I570636,I571086,);
nor I_33414 (I571094,I571086,I570820);
DFFARX1 I_33415 (I571094,I3035,I570636,I570607,);
nand I_33416 (I571125,I571086,I570727);
nand I_33417 (I571142,I570820,I571125);
nor I_33418 (I570616,I571142,I570786);
not I_33419 (I571197,I3042);
DFFARX1 I_33420 (I182467,I3035,I571197,I571223,);
DFFARX1 I_33421 (I571223,I3035,I571197,I571240,);
not I_33422 (I571189,I571240);
not I_33423 (I571262,I571223);
DFFARX1 I_33424 (I182464,I3035,I571197,I571288,);
nand I_33425 (I571296,I571288,I182458);
not I_33426 (I571313,I182458);
not I_33427 (I571330,I182455);
nand I_33428 (I571347,I182449,I182446);
and I_33429 (I571364,I182449,I182446);
not I_33430 (I571381,I182461);
nand I_33431 (I571398,I571381,I571330);
nor I_33432 (I571171,I571398,I571296);
nor I_33433 (I571429,I571313,I571398);
nand I_33434 (I571174,I571364,I571429);
not I_33435 (I571460,I182473);
nor I_33436 (I571477,I571460,I182449);
nor I_33437 (I571494,I571477,I182461);
nor I_33438 (I571511,I571262,I571494);
DFFARX1 I_33439 (I571511,I3035,I571197,I571183,);
not I_33440 (I571542,I571477);
DFFARX1 I_33441 (I571542,I3035,I571197,I571186,);
and I_33442 (I571180,I571288,I571477);
nor I_33443 (I571587,I571460,I182470);
and I_33444 (I571604,I571587,I182446);
or I_33445 (I571621,I571604,I182452);
DFFARX1 I_33446 (I571621,I3035,I571197,I571647,);
nor I_33447 (I571655,I571647,I571381);
DFFARX1 I_33448 (I571655,I3035,I571197,I571168,);
nand I_33449 (I571686,I571647,I571288);
nand I_33450 (I571703,I571381,I571686);
nor I_33451 (I571177,I571703,I571347);
not I_33452 (I571758,I3042);
DFFARX1 I_33453 (I103297,I3035,I571758,I571784,);
DFFARX1 I_33454 (I571784,I3035,I571758,I571801,);
not I_33455 (I571750,I571801);
not I_33456 (I571823,I571784);
DFFARX1 I_33457 (I103312,I3035,I571758,I571849,);
nand I_33458 (I571857,I571849,I103294);
not I_33459 (I571874,I103294);
not I_33460 (I571891,I103303);
nand I_33461 (I571908,I103309,I103300);
and I_33462 (I571925,I103309,I103300);
not I_33463 (I571942,I103297);
nand I_33464 (I571959,I571942,I571891);
nor I_33465 (I571732,I571959,I571857);
nor I_33466 (I571990,I571874,I571959);
nand I_33467 (I571735,I571925,I571990);
not I_33468 (I572021,I103294);
nor I_33469 (I572038,I572021,I103309);
nor I_33470 (I572055,I572038,I103297);
nor I_33471 (I572072,I571823,I572055);
DFFARX1 I_33472 (I572072,I3035,I571758,I571744,);
not I_33473 (I572103,I572038);
DFFARX1 I_33474 (I572103,I3035,I571758,I571747,);
and I_33475 (I571741,I571849,I572038);
nor I_33476 (I572148,I572021,I103318);
and I_33477 (I572165,I572148,I103315);
or I_33478 (I572182,I572165,I103306);
DFFARX1 I_33479 (I572182,I3035,I571758,I572208,);
nor I_33480 (I572216,I572208,I571942);
DFFARX1 I_33481 (I572216,I3035,I571758,I571729,);
nand I_33482 (I572247,I572208,I571849);
nand I_33483 (I572264,I571942,I572247);
nor I_33484 (I571738,I572264,I571908);
not I_33485 (I572322,I3042);
DFFARX1 I_33486 (I729380,I3035,I572322,I572348,);
and I_33487 (I572356,I572348,I729362);
DFFARX1 I_33488 (I572356,I3035,I572322,I572305,);
DFFARX1 I_33489 (I729353,I3035,I572322,I572396,);
not I_33490 (I572404,I729368);
not I_33491 (I572421,I729356);
nand I_33492 (I572438,I572421,I572404);
nor I_33493 (I572293,I572396,I572438);
DFFARX1 I_33494 (I572438,I3035,I572322,I572478,);
not I_33495 (I572314,I572478);
not I_33496 (I572500,I729365);
nand I_33497 (I572517,I572421,I572500);
DFFARX1 I_33498 (I572517,I3035,I572322,I572543,);
not I_33499 (I572551,I572543);
not I_33500 (I572568,I729374);
nand I_33501 (I572585,I572568,I729353);
and I_33502 (I572602,I572404,I572585);
nor I_33503 (I572619,I572517,I572602);
DFFARX1 I_33504 (I572619,I3035,I572322,I572290,);
DFFARX1 I_33505 (I572602,I3035,I572322,I572311,);
nor I_33506 (I572664,I729374,I729377);
nor I_33507 (I572302,I572517,I572664);
or I_33508 (I572695,I729374,I729377);
nor I_33509 (I572712,I729371,I729359);
DFFARX1 I_33510 (I572712,I3035,I572322,I572738,);
not I_33511 (I572746,I572738);
nor I_33512 (I572308,I572746,I572551);
nand I_33513 (I572777,I572746,I572396);
not I_33514 (I572794,I729371);
nand I_33515 (I572811,I572794,I572500);
nand I_33516 (I572828,I572746,I572811);
nand I_33517 (I572299,I572828,I572777);
nand I_33518 (I572296,I572811,I572695);
not I_33519 (I572900,I3042);
DFFARX1 I_33520 (I121144,I3035,I572900,I572926,);
and I_33521 (I572934,I572926,I121147);
DFFARX1 I_33522 (I572934,I3035,I572900,I572883,);
DFFARX1 I_33523 (I121147,I3035,I572900,I572974,);
not I_33524 (I572982,I121162);
not I_33525 (I572999,I121168);
nand I_33526 (I573016,I572999,I572982);
nor I_33527 (I572871,I572974,I573016);
DFFARX1 I_33528 (I573016,I3035,I572900,I573056,);
not I_33529 (I572892,I573056);
not I_33530 (I573078,I121156);
nand I_33531 (I573095,I572999,I573078);
DFFARX1 I_33532 (I573095,I3035,I572900,I573121,);
not I_33533 (I573129,I573121);
not I_33534 (I573146,I121153);
nand I_33535 (I573163,I573146,I121150);
and I_33536 (I573180,I572982,I573163);
nor I_33537 (I573197,I573095,I573180);
DFFARX1 I_33538 (I573197,I3035,I572900,I572868,);
DFFARX1 I_33539 (I573180,I3035,I572900,I572889,);
nor I_33540 (I573242,I121153,I121144);
nor I_33541 (I572880,I573095,I573242);
or I_33542 (I573273,I121153,I121144);
nor I_33543 (I573290,I121159,I121165);
DFFARX1 I_33544 (I573290,I3035,I572900,I573316,);
not I_33545 (I573324,I573316);
nor I_33546 (I572886,I573324,I573129);
nand I_33547 (I573355,I573324,I572974);
not I_33548 (I573372,I121159);
nand I_33549 (I573389,I573372,I573078);
nand I_33550 (I573406,I573324,I573389);
nand I_33551 (I572877,I573406,I573355);
nand I_33552 (I572874,I573389,I573273);
not I_33553 (I573478,I3042);
DFFARX1 I_33554 (I87229,I3035,I573478,I573504,);
and I_33555 (I573512,I573504,I87232);
DFFARX1 I_33556 (I573512,I3035,I573478,I573461,);
DFFARX1 I_33557 (I87232,I3035,I573478,I573552,);
not I_33558 (I573560,I87247);
not I_33559 (I573577,I87253);
nand I_33560 (I573594,I573577,I573560);
nor I_33561 (I573449,I573552,I573594);
DFFARX1 I_33562 (I573594,I3035,I573478,I573634,);
not I_33563 (I573470,I573634);
not I_33564 (I573656,I87241);
nand I_33565 (I573673,I573577,I573656);
DFFARX1 I_33566 (I573673,I3035,I573478,I573699,);
not I_33567 (I573707,I573699);
not I_33568 (I573724,I87238);
nand I_33569 (I573741,I573724,I87235);
and I_33570 (I573758,I573560,I573741);
nor I_33571 (I573775,I573673,I573758);
DFFARX1 I_33572 (I573775,I3035,I573478,I573446,);
DFFARX1 I_33573 (I573758,I3035,I573478,I573467,);
nor I_33574 (I573820,I87238,I87229);
nor I_33575 (I573458,I573673,I573820);
or I_33576 (I573851,I87238,I87229);
nor I_33577 (I573868,I87244,I87250);
DFFARX1 I_33578 (I573868,I3035,I573478,I573894,);
not I_33579 (I573902,I573894);
nor I_33580 (I573464,I573902,I573707);
nand I_33581 (I573933,I573902,I573552);
not I_33582 (I573950,I87244);
nand I_33583 (I573967,I573950,I573656);
nand I_33584 (I573984,I573902,I573967);
nand I_33585 (I573455,I573984,I573933);
nand I_33586 (I573452,I573967,I573851);
not I_33587 (I574056,I3042);
DFFARX1 I_33588 (I53151,I3035,I574056,I574082,);
and I_33589 (I574090,I574082,I53127);
DFFARX1 I_33590 (I574090,I3035,I574056,I574039,);
DFFARX1 I_33591 (I53145,I3035,I574056,I574130,);
not I_33592 (I574138,I53133);
not I_33593 (I574155,I53130);
nand I_33594 (I574172,I574155,I574138);
nor I_33595 (I574027,I574130,I574172);
DFFARX1 I_33596 (I574172,I3035,I574056,I574212,);
not I_33597 (I574048,I574212);
not I_33598 (I574234,I53139);
nand I_33599 (I574251,I574155,I574234);
DFFARX1 I_33600 (I574251,I3035,I574056,I574277,);
not I_33601 (I574285,I574277);
not I_33602 (I574302,I53130);
nand I_33603 (I574319,I574302,I53148);
and I_33604 (I574336,I574138,I574319);
nor I_33605 (I574353,I574251,I574336);
DFFARX1 I_33606 (I574353,I3035,I574056,I574024,);
DFFARX1 I_33607 (I574336,I3035,I574056,I574045,);
nor I_33608 (I574398,I53130,I53142);
nor I_33609 (I574036,I574251,I574398);
or I_33610 (I574429,I53130,I53142);
nor I_33611 (I574446,I53136,I53127);
DFFARX1 I_33612 (I574446,I3035,I574056,I574472,);
not I_33613 (I574480,I574472);
nor I_33614 (I574042,I574480,I574285);
nand I_33615 (I574511,I574480,I574130);
not I_33616 (I574528,I53136);
nand I_33617 (I574545,I574528,I574234);
nand I_33618 (I574562,I574480,I574545);
nand I_33619 (I574033,I574562,I574511);
nand I_33620 (I574030,I574545,I574429);
not I_33621 (I574634,I3042);
DFFARX1 I_33622 (I671387,I3035,I574634,I574660,);
and I_33623 (I574668,I574660,I671381);
DFFARX1 I_33624 (I574668,I3035,I574634,I574617,);
DFFARX1 I_33625 (I671366,I3035,I574634,I574708,);
not I_33626 (I574716,I671372);
not I_33627 (I574733,I671384);
nand I_33628 (I574750,I574733,I574716);
nor I_33629 (I574605,I574708,I574750);
DFFARX1 I_33630 (I574750,I3035,I574634,I574790,);
not I_33631 (I574626,I574790);
not I_33632 (I574812,I671366);
nand I_33633 (I574829,I574733,I574812);
DFFARX1 I_33634 (I574829,I3035,I574634,I574855,);
not I_33635 (I574863,I574855);
not I_33636 (I574880,I671390);
nand I_33637 (I574897,I574880,I671378);
and I_33638 (I574914,I574716,I574897);
nor I_33639 (I574931,I574829,I574914);
DFFARX1 I_33640 (I574931,I3035,I574634,I574602,);
DFFARX1 I_33641 (I574914,I3035,I574634,I574623,);
nor I_33642 (I574976,I671390,I671369);
nor I_33643 (I574614,I574829,I574976);
or I_33644 (I575007,I671390,I671369);
nor I_33645 (I575024,I671375,I671369);
DFFARX1 I_33646 (I575024,I3035,I574634,I575050,);
not I_33647 (I575058,I575050);
nor I_33648 (I574620,I575058,I574863);
nand I_33649 (I575089,I575058,I574708);
not I_33650 (I575106,I671375);
nand I_33651 (I575123,I575106,I574812);
nand I_33652 (I575140,I575058,I575123);
nand I_33653 (I574611,I575140,I575089);
nand I_33654 (I574608,I575123,I575007);
not I_33655 (I575212,I3042);
DFFARX1 I_33656 (I316353,I3035,I575212,I575238,);
and I_33657 (I575246,I575238,I316341);
DFFARX1 I_33658 (I575246,I3035,I575212,I575195,);
DFFARX1 I_33659 (I316356,I3035,I575212,I575286,);
not I_33660 (I575294,I316347);
not I_33661 (I575311,I316338);
nand I_33662 (I575328,I575311,I575294);
nor I_33663 (I575183,I575286,I575328);
DFFARX1 I_33664 (I575328,I3035,I575212,I575368,);
not I_33665 (I575204,I575368);
not I_33666 (I575390,I316344);
nand I_33667 (I575407,I575311,I575390);
DFFARX1 I_33668 (I575407,I3035,I575212,I575433,);
not I_33669 (I575441,I575433);
not I_33670 (I575458,I316359);
nand I_33671 (I575475,I575458,I316362);
and I_33672 (I575492,I575294,I575475);
nor I_33673 (I575509,I575407,I575492);
DFFARX1 I_33674 (I575509,I3035,I575212,I575180,);
DFFARX1 I_33675 (I575492,I3035,I575212,I575201,);
nor I_33676 (I575554,I316359,I316338);
nor I_33677 (I575192,I575407,I575554);
or I_33678 (I575585,I316359,I316338);
nor I_33679 (I575602,I316350,I316341);
DFFARX1 I_33680 (I575602,I3035,I575212,I575628,);
not I_33681 (I575636,I575628);
nor I_33682 (I575198,I575636,I575441);
nand I_33683 (I575667,I575636,I575286);
not I_33684 (I575684,I316350);
nand I_33685 (I575701,I575684,I575390);
nand I_33686 (I575718,I575636,I575701);
nand I_33687 (I575189,I575718,I575667);
nand I_33688 (I575186,I575701,I575585);
not I_33689 (I575790,I3042);
DFFARX1 I_33690 (I184054,I3035,I575790,I575816,);
and I_33691 (I575824,I575816,I184039);
DFFARX1 I_33692 (I575824,I3035,I575790,I575773,);
DFFARX1 I_33693 (I184045,I3035,I575790,I575864,);
not I_33694 (I575872,I184027);
not I_33695 (I575889,I184048);
nand I_33696 (I575906,I575889,I575872);
nor I_33697 (I575761,I575864,I575906);
DFFARX1 I_33698 (I575906,I3035,I575790,I575946,);
not I_33699 (I575782,I575946);
not I_33700 (I575968,I184051);
nand I_33701 (I575985,I575889,I575968);
DFFARX1 I_33702 (I575985,I3035,I575790,I576011,);
not I_33703 (I576019,I576011);
not I_33704 (I576036,I184042);
nand I_33705 (I576053,I576036,I184030);
and I_33706 (I576070,I575872,I576053);
nor I_33707 (I576087,I575985,I576070);
DFFARX1 I_33708 (I576087,I3035,I575790,I575758,);
DFFARX1 I_33709 (I576070,I3035,I575790,I575779,);
nor I_33710 (I576132,I184042,I184036);
nor I_33711 (I575770,I575985,I576132);
or I_33712 (I576163,I184042,I184036);
nor I_33713 (I576180,I184033,I184027);
DFFARX1 I_33714 (I576180,I3035,I575790,I576206,);
not I_33715 (I576214,I576206);
nor I_33716 (I575776,I576214,I576019);
nand I_33717 (I576245,I576214,I575864);
not I_33718 (I576262,I184033);
nand I_33719 (I576279,I576262,I575968);
nand I_33720 (I576296,I576214,I576279);
nand I_33721 (I575767,I576296,I576245);
nand I_33722 (I575764,I576279,I576163);
not I_33723 (I576368,I3042);
DFFARX1 I_33724 (I684650,I3035,I576368,I576394,);
and I_33725 (I576402,I576394,I684632);
DFFARX1 I_33726 (I576402,I3035,I576368,I576351,);
DFFARX1 I_33727 (I684641,I3035,I576368,I576442,);
not I_33728 (I576450,I684626);
not I_33729 (I576467,I684638);
nand I_33730 (I576484,I576467,I576450);
nor I_33731 (I576339,I576442,I576484);
DFFARX1 I_33732 (I576484,I3035,I576368,I576524,);
not I_33733 (I576360,I576524);
not I_33734 (I576546,I684629);
nand I_33735 (I576563,I576467,I576546);
DFFARX1 I_33736 (I576563,I3035,I576368,I576589,);
not I_33737 (I576597,I576589);
not I_33738 (I576614,I684626);
nand I_33739 (I576631,I576614,I684629);
and I_33740 (I576648,I576450,I576631);
nor I_33741 (I576665,I576563,I576648);
DFFARX1 I_33742 (I576665,I3035,I576368,I576336,);
DFFARX1 I_33743 (I576648,I3035,I576368,I576357,);
nor I_33744 (I576710,I684626,I684647);
nor I_33745 (I576348,I576563,I576710);
or I_33746 (I576741,I684626,I684647);
nor I_33747 (I576758,I684635,I684644);
DFFARX1 I_33748 (I576758,I3035,I576368,I576784,);
not I_33749 (I576792,I576784);
nor I_33750 (I576354,I576792,I576597);
nand I_33751 (I576823,I576792,I576442);
not I_33752 (I576840,I684635);
nand I_33753 (I576857,I576840,I576546);
nand I_33754 (I576874,I576792,I576857);
nand I_33755 (I576345,I576874,I576823);
nand I_33756 (I576342,I576857,I576741);
not I_33757 (I576946,I3042);
DFFARX1 I_33758 (I164555,I3035,I576946,I576972,);
and I_33759 (I576980,I576972,I164540);
DFFARX1 I_33760 (I576980,I3035,I576946,I576929,);
DFFARX1 I_33761 (I164546,I3035,I576946,I577020,);
not I_33762 (I577028,I164528);
not I_33763 (I577045,I164549);
nand I_33764 (I577062,I577045,I577028);
nor I_33765 (I576917,I577020,I577062);
DFFARX1 I_33766 (I577062,I3035,I576946,I577102,);
not I_33767 (I576938,I577102);
not I_33768 (I577124,I164552);
nand I_33769 (I577141,I577045,I577124);
DFFARX1 I_33770 (I577141,I3035,I576946,I577167,);
not I_33771 (I577175,I577167);
not I_33772 (I577192,I164543);
nand I_33773 (I577209,I577192,I164531);
and I_33774 (I577226,I577028,I577209);
nor I_33775 (I577243,I577141,I577226);
DFFARX1 I_33776 (I577243,I3035,I576946,I576914,);
DFFARX1 I_33777 (I577226,I3035,I576946,I576935,);
nor I_33778 (I577288,I164543,I164537);
nor I_33779 (I576926,I577141,I577288);
or I_33780 (I577319,I164543,I164537);
nor I_33781 (I577336,I164534,I164528);
DFFARX1 I_33782 (I577336,I3035,I576946,I577362,);
not I_33783 (I577370,I577362);
nor I_33784 (I576932,I577370,I577175);
nand I_33785 (I577401,I577370,I577020);
not I_33786 (I577418,I164534);
nand I_33787 (I577435,I577418,I577124);
nand I_33788 (I577452,I577370,I577435);
nand I_33789 (I576923,I577452,I577401);
nand I_33790 (I576920,I577435,I577319);
not I_33791 (I577524,I3042);
DFFARX1 I_33792 (I67380,I3035,I577524,I577550,);
and I_33793 (I577558,I577550,I67356);
DFFARX1 I_33794 (I577558,I3035,I577524,I577507,);
DFFARX1 I_33795 (I67374,I3035,I577524,I577598,);
not I_33796 (I577606,I67362);
not I_33797 (I577623,I67359);
nand I_33798 (I577640,I577623,I577606);
nor I_33799 (I577495,I577598,I577640);
DFFARX1 I_33800 (I577640,I3035,I577524,I577680,);
not I_33801 (I577516,I577680);
not I_33802 (I577702,I67368);
nand I_33803 (I577719,I577623,I577702);
DFFARX1 I_33804 (I577719,I3035,I577524,I577745,);
not I_33805 (I577753,I577745);
not I_33806 (I577770,I67359);
nand I_33807 (I577787,I577770,I67377);
and I_33808 (I577804,I577606,I577787);
nor I_33809 (I577821,I577719,I577804);
DFFARX1 I_33810 (I577821,I3035,I577524,I577492,);
DFFARX1 I_33811 (I577804,I3035,I577524,I577513,);
nor I_33812 (I577866,I67359,I67371);
nor I_33813 (I577504,I577719,I577866);
or I_33814 (I577897,I67359,I67371);
nor I_33815 (I577914,I67365,I67356);
DFFARX1 I_33816 (I577914,I3035,I577524,I577940,);
not I_33817 (I577948,I577940);
nor I_33818 (I577510,I577948,I577753);
nand I_33819 (I577979,I577948,I577598);
not I_33820 (I577996,I67365);
nand I_33821 (I578013,I577996,I577702);
nand I_33822 (I578030,I577948,I578013);
nand I_33823 (I577501,I578030,I577979);
nand I_33824 (I577498,I578013,I577897);
not I_33825 (I578102,I3042);
DFFARX1 I_33826 (I19399,I3035,I578102,I578128,);
and I_33827 (I578136,I578128,I19402);
DFFARX1 I_33828 (I578136,I3035,I578102,I578085,);
DFFARX1 I_33829 (I19402,I3035,I578102,I578176,);
not I_33830 (I578184,I19405);
not I_33831 (I578201,I19420);
nand I_33832 (I578218,I578201,I578184);
nor I_33833 (I578073,I578176,I578218);
DFFARX1 I_33834 (I578218,I3035,I578102,I578258,);
not I_33835 (I578094,I578258);
not I_33836 (I578280,I19414);
nand I_33837 (I578297,I578201,I578280);
DFFARX1 I_33838 (I578297,I3035,I578102,I578323,);
not I_33839 (I578331,I578323);
not I_33840 (I578348,I19417);
nand I_33841 (I578365,I578348,I19399);
and I_33842 (I578382,I578184,I578365);
nor I_33843 (I578399,I578297,I578382);
DFFARX1 I_33844 (I578399,I3035,I578102,I578070,);
DFFARX1 I_33845 (I578382,I3035,I578102,I578091,);
nor I_33846 (I578444,I19417,I19411);
nor I_33847 (I578082,I578297,I578444);
or I_33848 (I578475,I19417,I19411);
nor I_33849 (I578492,I19408,I19423);
DFFARX1 I_33850 (I578492,I3035,I578102,I578518,);
not I_33851 (I578526,I578518);
nor I_33852 (I578088,I578526,I578331);
nand I_33853 (I578557,I578526,I578176);
not I_33854 (I578574,I19408);
nand I_33855 (I578591,I578574,I578280);
nand I_33856 (I578608,I578526,I578591);
nand I_33857 (I578079,I578608,I578557);
nand I_33858 (I578076,I578591,I578475);
not I_33859 (I578680,I3042);
DFFARX1 I_33860 (I183527,I3035,I578680,I578706,);
and I_33861 (I578714,I578706,I183512);
DFFARX1 I_33862 (I578714,I3035,I578680,I578663,);
DFFARX1 I_33863 (I183518,I3035,I578680,I578754,);
not I_33864 (I578762,I183500);
not I_33865 (I578779,I183521);
nand I_33866 (I578796,I578779,I578762);
nor I_33867 (I578651,I578754,I578796);
DFFARX1 I_33868 (I578796,I3035,I578680,I578836,);
not I_33869 (I578672,I578836);
not I_33870 (I578858,I183524);
nand I_33871 (I578875,I578779,I578858);
DFFARX1 I_33872 (I578875,I3035,I578680,I578901,);
not I_33873 (I578909,I578901);
not I_33874 (I578926,I183515);
nand I_33875 (I578943,I578926,I183503);
and I_33876 (I578960,I578762,I578943);
nor I_33877 (I578977,I578875,I578960);
DFFARX1 I_33878 (I578977,I3035,I578680,I578648,);
DFFARX1 I_33879 (I578960,I3035,I578680,I578669,);
nor I_33880 (I579022,I183515,I183509);
nor I_33881 (I578660,I578875,I579022);
or I_33882 (I579053,I183515,I183509);
nor I_33883 (I579070,I183506,I183500);
DFFARX1 I_33884 (I579070,I3035,I578680,I579096,);
not I_33885 (I579104,I579096);
nor I_33886 (I578666,I579104,I578909);
nand I_33887 (I579135,I579104,I578754);
not I_33888 (I579152,I183506);
nand I_33889 (I579169,I579152,I578858);
nand I_33890 (I579186,I579104,I579169);
nand I_33891 (I578657,I579186,I579135);
nand I_33892 (I578654,I579169,I579053);
not I_33893 (I579258,I3042);
DFFARX1 I_33894 (I477368,I3035,I579258,I579284,);
and I_33895 (I579292,I579284,I477362);
DFFARX1 I_33896 (I579292,I3035,I579258,I579241,);
DFFARX1 I_33897 (I477380,I3035,I579258,I579332,);
not I_33898 (I579340,I477371);
not I_33899 (I579357,I477383);
nand I_33900 (I579374,I579357,I579340);
nor I_33901 (I579229,I579332,I579374);
DFFARX1 I_33902 (I579374,I3035,I579258,I579414,);
not I_33903 (I579250,I579414);
not I_33904 (I579436,I477389);
nand I_33905 (I579453,I579357,I579436);
DFFARX1 I_33906 (I579453,I3035,I579258,I579479,);
not I_33907 (I579487,I579479);
not I_33908 (I579504,I477365);
nand I_33909 (I579521,I579504,I477386);
and I_33910 (I579538,I579340,I579521);
nor I_33911 (I579555,I579453,I579538);
DFFARX1 I_33912 (I579555,I3035,I579258,I579226,);
DFFARX1 I_33913 (I579538,I3035,I579258,I579247,);
nor I_33914 (I579600,I477365,I477377);
nor I_33915 (I579238,I579453,I579600);
or I_33916 (I579631,I477365,I477377);
nor I_33917 (I579648,I477362,I477374);
DFFARX1 I_33918 (I579648,I3035,I579258,I579674,);
not I_33919 (I579682,I579674);
nor I_33920 (I579244,I579682,I579487);
nand I_33921 (I579713,I579682,I579332);
not I_33922 (I579730,I477362);
nand I_33923 (I579747,I579730,I579436);
nand I_33924 (I579764,I579682,I579747);
nand I_33925 (I579235,I579764,I579713);
nand I_33926 (I579232,I579747,I579631);
not I_33927 (I579836,I3042);
DFFARX1 I_33928 (I146134,I3035,I579836,I579862,);
and I_33929 (I579870,I579862,I146137);
DFFARX1 I_33930 (I579870,I3035,I579836,I579819,);
DFFARX1 I_33931 (I146137,I3035,I579836,I579910,);
not I_33932 (I579918,I146152);
not I_33933 (I579935,I146158);
nand I_33934 (I579952,I579935,I579918);
nor I_33935 (I579807,I579910,I579952);
DFFARX1 I_33936 (I579952,I3035,I579836,I579992,);
not I_33937 (I579828,I579992);
not I_33938 (I580014,I146146);
nand I_33939 (I580031,I579935,I580014);
DFFARX1 I_33940 (I580031,I3035,I579836,I580057,);
not I_33941 (I580065,I580057);
not I_33942 (I580082,I146143);
nand I_33943 (I580099,I580082,I146140);
and I_33944 (I580116,I579918,I580099);
nor I_33945 (I580133,I580031,I580116);
DFFARX1 I_33946 (I580133,I3035,I579836,I579804,);
DFFARX1 I_33947 (I580116,I3035,I579836,I579825,);
nor I_33948 (I580178,I146143,I146134);
nor I_33949 (I579816,I580031,I580178);
or I_33950 (I580209,I146143,I146134);
nor I_33951 (I580226,I146149,I146155);
DFFARX1 I_33952 (I580226,I3035,I579836,I580252,);
not I_33953 (I580260,I580252);
nor I_33954 (I579822,I580260,I580065);
nand I_33955 (I580291,I580260,I579910);
not I_33956 (I580308,I146149);
nand I_33957 (I580325,I580308,I580014);
nand I_33958 (I580342,I580260,I580325);
nand I_33959 (I579813,I580342,I580291);
nand I_33960 (I579810,I580325,I580209);
not I_33961 (I580414,I3042);
DFFARX1 I_33962 (I189324,I3035,I580414,I580440,);
and I_33963 (I580448,I580440,I189309);
DFFARX1 I_33964 (I580448,I3035,I580414,I580397,);
DFFARX1 I_33965 (I189315,I3035,I580414,I580488,);
not I_33966 (I580496,I189297);
not I_33967 (I580513,I189318);
nand I_33968 (I580530,I580513,I580496);
nor I_33969 (I580385,I580488,I580530);
DFFARX1 I_33970 (I580530,I3035,I580414,I580570,);
not I_33971 (I580406,I580570);
not I_33972 (I580592,I189321);
nand I_33973 (I580609,I580513,I580592);
DFFARX1 I_33974 (I580609,I3035,I580414,I580635,);
not I_33975 (I580643,I580635);
not I_33976 (I580660,I189312);
nand I_33977 (I580677,I580660,I189300);
and I_33978 (I580694,I580496,I580677);
nor I_33979 (I580711,I580609,I580694);
DFFARX1 I_33980 (I580711,I3035,I580414,I580382,);
DFFARX1 I_33981 (I580694,I3035,I580414,I580403,);
nor I_33982 (I580756,I189312,I189306);
nor I_33983 (I580394,I580609,I580756);
or I_33984 (I580787,I189312,I189306);
nor I_33985 (I580804,I189303,I189297);
DFFARX1 I_33986 (I580804,I3035,I580414,I580830,);
not I_33987 (I580838,I580830);
nor I_33988 (I580400,I580838,I580643);
nand I_33989 (I580869,I580838,I580488);
not I_33990 (I580886,I189303);
nand I_33991 (I580903,I580886,I580592);
nand I_33992 (I580920,I580838,I580903);
nand I_33993 (I580391,I580920,I580869);
nand I_33994 (I580388,I580903,I580787);
not I_33995 (I580992,I3042);
DFFARX1 I_33996 (I559390,I3035,I580992,I581018,);
and I_33997 (I581026,I581018,I559387);
DFFARX1 I_33998 (I581026,I3035,I580992,I580975,);
DFFARX1 I_33999 (I559393,I3035,I580992,I581066,);
not I_34000 (I581074,I559396);
not I_34001 (I581091,I559390);
nand I_34002 (I581108,I581091,I581074);
nor I_34003 (I580963,I581066,I581108);
DFFARX1 I_34004 (I581108,I3035,I580992,I581148,);
not I_34005 (I580984,I581148);
not I_34006 (I581170,I559405);
nand I_34007 (I581187,I581091,I581170);
DFFARX1 I_34008 (I581187,I3035,I580992,I581213,);
not I_34009 (I581221,I581213);
not I_34010 (I581238,I559402);
nand I_34011 (I581255,I581238,I559408);
and I_34012 (I581272,I581074,I581255);
nor I_34013 (I581289,I581187,I581272);
DFFARX1 I_34014 (I581289,I3035,I580992,I580960,);
DFFARX1 I_34015 (I581272,I3035,I580992,I580981,);
nor I_34016 (I581334,I559402,I559387);
nor I_34017 (I580972,I581187,I581334);
or I_34018 (I581365,I559402,I559387);
nor I_34019 (I581382,I559399,I559393);
DFFARX1 I_34020 (I581382,I3035,I580992,I581408,);
not I_34021 (I581416,I581408);
nor I_34022 (I580978,I581416,I581221);
nand I_34023 (I581447,I581416,I581066);
not I_34024 (I581464,I559399);
nand I_34025 (I581481,I581464,I581170);
nand I_34026 (I581498,I581416,I581481);
nand I_34027 (I580969,I581498,I581447);
nand I_34028 (I580966,I581481,I581365);
not I_34029 (I581570,I3042);
DFFARX1 I_34030 (I127689,I3035,I581570,I581596,);
and I_34031 (I581604,I581596,I127692);
DFFARX1 I_34032 (I581604,I3035,I581570,I581553,);
DFFARX1 I_34033 (I127692,I3035,I581570,I581644,);
not I_34034 (I581652,I127707);
not I_34035 (I581669,I127713);
nand I_34036 (I581686,I581669,I581652);
nor I_34037 (I581541,I581644,I581686);
DFFARX1 I_34038 (I581686,I3035,I581570,I581726,);
not I_34039 (I581562,I581726);
not I_34040 (I581748,I127701);
nand I_34041 (I581765,I581669,I581748);
DFFARX1 I_34042 (I581765,I3035,I581570,I581791,);
not I_34043 (I581799,I581791);
not I_34044 (I581816,I127698);
nand I_34045 (I581833,I581816,I127695);
and I_34046 (I581850,I581652,I581833);
nor I_34047 (I581867,I581765,I581850);
DFFARX1 I_34048 (I581867,I3035,I581570,I581538,);
DFFARX1 I_34049 (I581850,I3035,I581570,I581559,);
nor I_34050 (I581912,I127698,I127689);
nor I_34051 (I581550,I581765,I581912);
or I_34052 (I581943,I127698,I127689);
nor I_34053 (I581960,I127704,I127710);
DFFARX1 I_34054 (I581960,I3035,I581570,I581986,);
not I_34055 (I581994,I581986);
nor I_34056 (I581556,I581994,I581799);
nand I_34057 (I582025,I581994,I581644);
not I_34058 (I582042,I127704);
nand I_34059 (I582059,I582042,I581748);
nand I_34060 (I582076,I581994,I582059);
nand I_34061 (I581547,I582076,I582025);
nand I_34062 (I581544,I582059,I581943);
not I_34063 (I582148,I3042);
DFFARX1 I_34064 (I466179,I3035,I582148,I582174,);
and I_34065 (I582182,I582174,I466185);
DFFARX1 I_34066 (I582182,I3035,I582148,I582131,);
DFFARX1 I_34067 (I466191,I3035,I582148,I582222,);
not I_34068 (I582230,I466176);
not I_34069 (I582247,I466176);
nand I_34070 (I582264,I582247,I582230);
nor I_34071 (I582119,I582222,I582264);
DFFARX1 I_34072 (I582264,I3035,I582148,I582304,);
not I_34073 (I582140,I582304);
not I_34074 (I582326,I466194);
nand I_34075 (I582343,I582247,I582326);
DFFARX1 I_34076 (I582343,I3035,I582148,I582369,);
not I_34077 (I582377,I582369);
not I_34078 (I582394,I466188);
nand I_34079 (I582411,I582394,I466179);
and I_34080 (I582428,I582230,I582411);
nor I_34081 (I582445,I582343,I582428);
DFFARX1 I_34082 (I582445,I3035,I582148,I582116,);
DFFARX1 I_34083 (I582428,I3035,I582148,I582137,);
nor I_34084 (I582490,I466188,I466197);
nor I_34085 (I582128,I582343,I582490);
or I_34086 (I582521,I466188,I466197);
nor I_34087 (I582538,I466182,I466182);
DFFARX1 I_34088 (I582538,I3035,I582148,I582564,);
not I_34089 (I582572,I582564);
nor I_34090 (I582134,I582572,I582377);
nand I_34091 (I582603,I582572,I582222);
not I_34092 (I582620,I466182);
nand I_34093 (I582637,I582620,I582326);
nand I_34094 (I582654,I582572,I582637);
nand I_34095 (I582125,I582654,I582603);
nand I_34096 (I582122,I582637,I582521);
not I_34097 (I582726,I3042);
DFFARX1 I_34098 (I482536,I3035,I582726,I582752,);
and I_34099 (I582760,I582752,I482530);
DFFARX1 I_34100 (I582760,I3035,I582726,I582709,);
DFFARX1 I_34101 (I482548,I3035,I582726,I582800,);
not I_34102 (I582808,I482539);
not I_34103 (I582825,I482551);
nand I_34104 (I582842,I582825,I582808);
nor I_34105 (I582697,I582800,I582842);
DFFARX1 I_34106 (I582842,I3035,I582726,I582882,);
not I_34107 (I582718,I582882);
not I_34108 (I582904,I482557);
nand I_34109 (I582921,I582825,I582904);
DFFARX1 I_34110 (I582921,I3035,I582726,I582947,);
not I_34111 (I582955,I582947);
not I_34112 (I582972,I482533);
nand I_34113 (I582989,I582972,I482554);
and I_34114 (I583006,I582808,I582989);
nor I_34115 (I583023,I582921,I583006);
DFFARX1 I_34116 (I583023,I3035,I582726,I582694,);
DFFARX1 I_34117 (I583006,I3035,I582726,I582715,);
nor I_34118 (I583068,I482533,I482545);
nor I_34119 (I582706,I582921,I583068);
or I_34120 (I583099,I482533,I482545);
nor I_34121 (I583116,I482530,I482542);
DFFARX1 I_34122 (I583116,I3035,I582726,I583142,);
not I_34123 (I583150,I583142);
nor I_34124 (I582712,I583150,I582955);
nand I_34125 (I583181,I583150,I582800);
not I_34126 (I583198,I482530);
nand I_34127 (I583215,I583198,I582904);
nand I_34128 (I583232,I583150,I583215);
nand I_34129 (I582703,I583232,I583181);
nand I_34130 (I582700,I583215,I583099);
not I_34131 (I583304,I3042);
DFFARX1 I_34132 (I675402,I3035,I583304,I583330,);
and I_34133 (I583338,I583330,I675384);
DFFARX1 I_34134 (I583338,I3035,I583304,I583287,);
DFFARX1 I_34135 (I675393,I3035,I583304,I583378,);
not I_34136 (I583386,I675378);
not I_34137 (I583403,I675390);
nand I_34138 (I583420,I583403,I583386);
nor I_34139 (I583275,I583378,I583420);
DFFARX1 I_34140 (I583420,I3035,I583304,I583460,);
not I_34141 (I583296,I583460);
not I_34142 (I583482,I675381);
nand I_34143 (I583499,I583403,I583482);
DFFARX1 I_34144 (I583499,I3035,I583304,I583525,);
not I_34145 (I583533,I583525);
not I_34146 (I583550,I675378);
nand I_34147 (I583567,I583550,I675381);
and I_34148 (I583584,I583386,I583567);
nor I_34149 (I583601,I583499,I583584);
DFFARX1 I_34150 (I583601,I3035,I583304,I583272,);
DFFARX1 I_34151 (I583584,I3035,I583304,I583293,);
nor I_34152 (I583646,I675378,I675399);
nor I_34153 (I583284,I583499,I583646);
or I_34154 (I583677,I675378,I675399);
nor I_34155 (I583694,I675387,I675396);
DFFARX1 I_34156 (I583694,I3035,I583304,I583720,);
not I_34157 (I583728,I583720);
nor I_34158 (I583290,I583728,I583533);
nand I_34159 (I583759,I583728,I583378);
not I_34160 (I583776,I675387);
nand I_34161 (I583793,I583776,I583482);
nand I_34162 (I583810,I583728,I583793);
nand I_34163 (I583281,I583810,I583759);
nand I_34164 (I583278,I583793,I583677);
not I_34165 (I583882,I3042);
DFFARX1 I_34166 (I738305,I3035,I583882,I583908,);
and I_34167 (I583916,I583908,I738287);
DFFARX1 I_34168 (I583916,I3035,I583882,I583865,);
DFFARX1 I_34169 (I738278,I3035,I583882,I583956,);
not I_34170 (I583964,I738293);
not I_34171 (I583981,I738281);
nand I_34172 (I583998,I583981,I583964);
nor I_34173 (I583853,I583956,I583998);
DFFARX1 I_34174 (I583998,I3035,I583882,I584038,);
not I_34175 (I583874,I584038);
not I_34176 (I584060,I738290);
nand I_34177 (I584077,I583981,I584060);
DFFARX1 I_34178 (I584077,I3035,I583882,I584103,);
not I_34179 (I584111,I584103);
not I_34180 (I584128,I738299);
nand I_34181 (I584145,I584128,I738278);
and I_34182 (I584162,I583964,I584145);
nor I_34183 (I584179,I584077,I584162);
DFFARX1 I_34184 (I584179,I3035,I583882,I583850,);
DFFARX1 I_34185 (I584162,I3035,I583882,I583871,);
nor I_34186 (I584224,I738299,I738302);
nor I_34187 (I583862,I584077,I584224);
or I_34188 (I584255,I738299,I738302);
nor I_34189 (I584272,I738296,I738284);
DFFARX1 I_34190 (I584272,I3035,I583882,I584298,);
not I_34191 (I584306,I584298);
nor I_34192 (I583868,I584306,I584111);
nand I_34193 (I584337,I584306,I583956);
not I_34194 (I584354,I738296);
nand I_34195 (I584371,I584354,I584060);
nand I_34196 (I584388,I584306,I584371);
nand I_34197 (I583859,I584388,I584337);
nand I_34198 (I583856,I584371,I584255);
not I_34199 (I584460,I3042);
DFFARX1 I_34200 (I83064,I3035,I584460,I584486,);
and I_34201 (I584494,I584486,I83067);
DFFARX1 I_34202 (I584494,I3035,I584460,I584443,);
DFFARX1 I_34203 (I83067,I3035,I584460,I584534,);
not I_34204 (I584542,I83082);
not I_34205 (I584559,I83088);
nand I_34206 (I584576,I584559,I584542);
nor I_34207 (I584431,I584534,I584576);
DFFARX1 I_34208 (I584576,I3035,I584460,I584616,);
not I_34209 (I584452,I584616);
not I_34210 (I584638,I83076);
nand I_34211 (I584655,I584559,I584638);
DFFARX1 I_34212 (I584655,I3035,I584460,I584681,);
not I_34213 (I584689,I584681);
not I_34214 (I584706,I83073);
nand I_34215 (I584723,I584706,I83070);
and I_34216 (I584740,I584542,I584723);
nor I_34217 (I584757,I584655,I584740);
DFFARX1 I_34218 (I584757,I3035,I584460,I584428,);
DFFARX1 I_34219 (I584740,I3035,I584460,I584449,);
nor I_34220 (I584802,I83073,I83064);
nor I_34221 (I584440,I584655,I584802);
or I_34222 (I584833,I83073,I83064);
nor I_34223 (I584850,I83079,I83085);
DFFARX1 I_34224 (I584850,I3035,I584460,I584876,);
not I_34225 (I584884,I584876);
nor I_34226 (I584446,I584884,I584689);
nand I_34227 (I584915,I584884,I584534);
not I_34228 (I584932,I83079);
nand I_34229 (I584949,I584932,I584638);
nand I_34230 (I584966,I584884,I584949);
nand I_34231 (I584437,I584966,I584915);
nand I_34232 (I584434,I584949,I584833);
not I_34233 (I585038,I3042);
DFFARX1 I_34234 (I661595,I3035,I585038,I585064,);
and I_34235 (I585072,I585064,I661589);
DFFARX1 I_34236 (I585072,I3035,I585038,I585021,);
DFFARX1 I_34237 (I661574,I3035,I585038,I585112,);
not I_34238 (I585120,I661580);
not I_34239 (I585137,I661592);
nand I_34240 (I585154,I585137,I585120);
nor I_34241 (I585009,I585112,I585154);
DFFARX1 I_34242 (I585154,I3035,I585038,I585194,);
not I_34243 (I585030,I585194);
not I_34244 (I585216,I661574);
nand I_34245 (I585233,I585137,I585216);
DFFARX1 I_34246 (I585233,I3035,I585038,I585259,);
not I_34247 (I585267,I585259);
not I_34248 (I585284,I661598);
nand I_34249 (I585301,I585284,I661586);
and I_34250 (I585318,I585120,I585301);
nor I_34251 (I585335,I585233,I585318);
DFFARX1 I_34252 (I585335,I3035,I585038,I585006,);
DFFARX1 I_34253 (I585318,I3035,I585038,I585027,);
nor I_34254 (I585380,I661598,I661577);
nor I_34255 (I585018,I585233,I585380);
or I_34256 (I585411,I661598,I661577);
nor I_34257 (I585428,I661583,I661577);
DFFARX1 I_34258 (I585428,I3035,I585038,I585454,);
not I_34259 (I585462,I585454);
nor I_34260 (I585024,I585462,I585267);
nand I_34261 (I585493,I585462,I585112);
not I_34262 (I585510,I661583);
nand I_34263 (I585527,I585510,I585216);
nand I_34264 (I585544,I585462,I585527);
nand I_34265 (I585015,I585544,I585493);
nand I_34266 (I585012,I585527,I585411);
not I_34267 (I585616,I3042);
DFFARX1 I_34268 (I453004,I3035,I585616,I585642,);
and I_34269 (I585650,I585642,I453010);
DFFARX1 I_34270 (I585650,I3035,I585616,I585599,);
DFFARX1 I_34271 (I453016,I3035,I585616,I585690,);
not I_34272 (I585698,I453001);
not I_34273 (I585715,I453001);
nand I_34274 (I585732,I585715,I585698);
nor I_34275 (I585587,I585690,I585732);
DFFARX1 I_34276 (I585732,I3035,I585616,I585772,);
not I_34277 (I585608,I585772);
not I_34278 (I585794,I453019);
nand I_34279 (I585811,I585715,I585794);
DFFARX1 I_34280 (I585811,I3035,I585616,I585837,);
not I_34281 (I585845,I585837);
not I_34282 (I585862,I453013);
nand I_34283 (I585879,I585862,I453004);
and I_34284 (I585896,I585698,I585879);
nor I_34285 (I585913,I585811,I585896);
DFFARX1 I_34286 (I585913,I3035,I585616,I585584,);
DFFARX1 I_34287 (I585896,I3035,I585616,I585605,);
nor I_34288 (I585958,I453013,I453022);
nor I_34289 (I585596,I585811,I585958);
or I_34290 (I585989,I453013,I453022);
nor I_34291 (I586006,I453007,I453007);
DFFARX1 I_34292 (I586006,I3035,I585616,I586032,);
not I_34293 (I586040,I586032);
nor I_34294 (I585602,I586040,I585845);
nand I_34295 (I586071,I586040,I585690);
not I_34296 (I586088,I453007);
nand I_34297 (I586105,I586088,I585794);
nand I_34298 (I586122,I586040,I586105);
nand I_34299 (I585593,I586122,I586071);
nand I_34300 (I585590,I586105,I585989);
not I_34301 (I586194,I3042);
DFFARX1 I_34302 (I312885,I3035,I586194,I586220,);
and I_34303 (I586228,I586220,I312873);
DFFARX1 I_34304 (I586228,I3035,I586194,I586177,);
DFFARX1 I_34305 (I312888,I3035,I586194,I586268,);
not I_34306 (I586276,I312879);
not I_34307 (I586293,I312870);
nand I_34308 (I586310,I586293,I586276);
nor I_34309 (I586165,I586268,I586310);
DFFARX1 I_34310 (I586310,I3035,I586194,I586350,);
not I_34311 (I586186,I586350);
not I_34312 (I586372,I312876);
nand I_34313 (I586389,I586293,I586372);
DFFARX1 I_34314 (I586389,I3035,I586194,I586415,);
not I_34315 (I586423,I586415);
not I_34316 (I586440,I312891);
nand I_34317 (I586457,I586440,I312894);
and I_34318 (I586474,I586276,I586457);
nor I_34319 (I586491,I586389,I586474);
DFFARX1 I_34320 (I586491,I3035,I586194,I586162,);
DFFARX1 I_34321 (I586474,I3035,I586194,I586183,);
nor I_34322 (I586536,I312891,I312870);
nor I_34323 (I586174,I586389,I586536);
or I_34324 (I586567,I312891,I312870);
nor I_34325 (I586584,I312882,I312873);
DFFARX1 I_34326 (I586584,I3035,I586194,I586610,);
not I_34327 (I586618,I586610);
nor I_34328 (I586180,I586618,I586423);
nand I_34329 (I586649,I586618,I586268);
not I_34330 (I586666,I312882);
nand I_34331 (I586683,I586666,I586372);
nand I_34332 (I586700,I586618,I586683);
nand I_34333 (I586171,I586700,I586649);
nand I_34334 (I586168,I586683,I586567);
not I_34335 (I586772,I3042);
DFFARX1 I_34336 (I203553,I3035,I586772,I586798,);
and I_34337 (I586806,I586798,I203538);
DFFARX1 I_34338 (I586806,I3035,I586772,I586755,);
DFFARX1 I_34339 (I203544,I3035,I586772,I586846,);
not I_34340 (I586854,I203526);
not I_34341 (I586871,I203547);
nand I_34342 (I586888,I586871,I586854);
nor I_34343 (I586743,I586846,I586888);
DFFARX1 I_34344 (I586888,I3035,I586772,I586928,);
not I_34345 (I586764,I586928);
not I_34346 (I586950,I203550);
nand I_34347 (I586967,I586871,I586950);
DFFARX1 I_34348 (I586967,I3035,I586772,I586993,);
not I_34349 (I587001,I586993);
not I_34350 (I587018,I203541);
nand I_34351 (I587035,I587018,I203529);
and I_34352 (I587052,I586854,I587035);
nor I_34353 (I587069,I586967,I587052);
DFFARX1 I_34354 (I587069,I3035,I586772,I586740,);
DFFARX1 I_34355 (I587052,I3035,I586772,I586761,);
nor I_34356 (I587114,I203541,I203535);
nor I_34357 (I586752,I586967,I587114);
or I_34358 (I587145,I203541,I203535);
nor I_34359 (I587162,I203532,I203526);
DFFARX1 I_34360 (I587162,I3035,I586772,I587188,);
not I_34361 (I587196,I587188);
nor I_34362 (I586758,I587196,I587001);
nand I_34363 (I587227,I587196,I586846);
not I_34364 (I587244,I203532);
nand I_34365 (I587261,I587244,I586950);
nand I_34366 (I587278,I587196,I587261);
nand I_34367 (I586749,I587278,I587227);
nand I_34368 (I586746,I587261,I587145);
not I_34369 (I587350,I3042);
DFFARX1 I_34370 (I699035,I3035,I587350,I587376,);
and I_34371 (I587384,I587376,I699017);
DFFARX1 I_34372 (I587384,I3035,I587350,I587333,);
DFFARX1 I_34373 (I699008,I3035,I587350,I587424,);
not I_34374 (I587432,I699023);
not I_34375 (I587449,I699011);
nand I_34376 (I587466,I587449,I587432);
nor I_34377 (I587321,I587424,I587466);
DFFARX1 I_34378 (I587466,I3035,I587350,I587506,);
not I_34379 (I587342,I587506);
not I_34380 (I587528,I699020);
nand I_34381 (I587545,I587449,I587528);
DFFARX1 I_34382 (I587545,I3035,I587350,I587571,);
not I_34383 (I587579,I587571);
not I_34384 (I587596,I699029);
nand I_34385 (I587613,I587596,I699008);
and I_34386 (I587630,I587432,I587613);
nor I_34387 (I587647,I587545,I587630);
DFFARX1 I_34388 (I587647,I3035,I587350,I587318,);
DFFARX1 I_34389 (I587630,I3035,I587350,I587339,);
nor I_34390 (I587692,I699029,I699032);
nor I_34391 (I587330,I587545,I587692);
or I_34392 (I587723,I699029,I699032);
nor I_34393 (I587740,I699026,I699014);
DFFARX1 I_34394 (I587740,I3035,I587350,I587766,);
not I_34395 (I587774,I587766);
nor I_34396 (I587336,I587774,I587579);
nand I_34397 (I587805,I587774,I587424);
not I_34398 (I587822,I699026);
nand I_34399 (I587839,I587822,I587528);
nand I_34400 (I587856,I587774,I587839);
nand I_34401 (I587327,I587856,I587805);
nand I_34402 (I587324,I587839,I587723);
not I_34403 (I587928,I3042);
DFFARX1 I_34404 (I651259,I3035,I587928,I587954,);
and I_34405 (I587962,I587954,I651253);
DFFARX1 I_34406 (I587962,I3035,I587928,I587911,);
DFFARX1 I_34407 (I651238,I3035,I587928,I588002,);
not I_34408 (I588010,I651244);
not I_34409 (I588027,I651256);
nand I_34410 (I588044,I588027,I588010);
nor I_34411 (I587899,I588002,I588044);
DFFARX1 I_34412 (I588044,I3035,I587928,I588084,);
not I_34413 (I587920,I588084);
not I_34414 (I588106,I651238);
nand I_34415 (I588123,I588027,I588106);
DFFARX1 I_34416 (I588123,I3035,I587928,I588149,);
not I_34417 (I588157,I588149);
not I_34418 (I588174,I651262);
nand I_34419 (I588191,I588174,I651250);
and I_34420 (I588208,I588010,I588191);
nor I_34421 (I588225,I588123,I588208);
DFFARX1 I_34422 (I588225,I3035,I587928,I587896,);
DFFARX1 I_34423 (I588208,I3035,I587928,I587917,);
nor I_34424 (I588270,I651262,I651241);
nor I_34425 (I587908,I588123,I588270);
or I_34426 (I588301,I651262,I651241);
nor I_34427 (I588318,I651247,I651241);
DFFARX1 I_34428 (I588318,I3035,I587928,I588344,);
not I_34429 (I588352,I588344);
nor I_34430 (I587914,I588352,I588157);
nand I_34431 (I588383,I588352,I588002);
not I_34432 (I588400,I651247);
nand I_34433 (I588417,I588400,I588106);
nand I_34434 (I588434,I588352,I588417);
nand I_34435 (I587905,I588434,I588383);
nand I_34436 (I587902,I588417,I588301);
not I_34437 (I588506,I3042);
DFFARX1 I_34438 (I333115,I3035,I588506,I588532,);
and I_34439 (I588540,I588532,I333103);
DFFARX1 I_34440 (I588540,I3035,I588506,I588489,);
DFFARX1 I_34441 (I333118,I3035,I588506,I588580,);
not I_34442 (I588588,I333109);
not I_34443 (I588605,I333100);
nand I_34444 (I588622,I588605,I588588);
nor I_34445 (I588477,I588580,I588622);
DFFARX1 I_34446 (I588622,I3035,I588506,I588662,);
not I_34447 (I588498,I588662);
not I_34448 (I588684,I333106);
nand I_34449 (I588701,I588605,I588684);
DFFARX1 I_34450 (I588701,I3035,I588506,I588727,);
not I_34451 (I588735,I588727);
not I_34452 (I588752,I333121);
nand I_34453 (I588769,I588752,I333124);
and I_34454 (I588786,I588588,I588769);
nor I_34455 (I588803,I588701,I588786);
DFFARX1 I_34456 (I588803,I3035,I588506,I588474,);
DFFARX1 I_34457 (I588786,I3035,I588506,I588495,);
nor I_34458 (I588848,I333121,I333100);
nor I_34459 (I588486,I588701,I588848);
or I_34460 (I588879,I333121,I333100);
nor I_34461 (I588896,I333112,I333103);
DFFARX1 I_34462 (I588896,I3035,I588506,I588922,);
not I_34463 (I588930,I588922);
nor I_34464 (I588492,I588930,I588735);
nand I_34465 (I588961,I588930,I588580);
not I_34466 (I588978,I333112);
nand I_34467 (I588995,I588978,I588684);
nand I_34468 (I589012,I588930,I588995);
nand I_34469 (I588483,I589012,I588961);
nand I_34470 (I588480,I588995,I588879);
not I_34471 (I589084,I3042);
DFFARX1 I_34472 (I252197,I3035,I589084,I589110,);
and I_34473 (I589118,I589110,I252212);
DFFARX1 I_34474 (I589118,I3035,I589084,I589067,);
DFFARX1 I_34475 (I252215,I3035,I589084,I589158,);
not I_34476 (I589166,I252209);
not I_34477 (I589183,I252224);
nand I_34478 (I589200,I589183,I589166);
nor I_34479 (I589055,I589158,I589200);
DFFARX1 I_34480 (I589200,I3035,I589084,I589240,);
not I_34481 (I589076,I589240);
not I_34482 (I589262,I252200);
nand I_34483 (I589279,I589183,I589262);
DFFARX1 I_34484 (I589279,I3035,I589084,I589305,);
not I_34485 (I589313,I589305);
not I_34486 (I589330,I252203);
nand I_34487 (I589347,I589330,I252197);
and I_34488 (I589364,I589166,I589347);
nor I_34489 (I589381,I589279,I589364);
DFFARX1 I_34490 (I589381,I3035,I589084,I589052,);
DFFARX1 I_34491 (I589364,I3035,I589084,I589073,);
nor I_34492 (I589426,I252203,I252206);
nor I_34493 (I589064,I589279,I589426);
or I_34494 (I589457,I252203,I252206);
nor I_34495 (I589474,I252221,I252218);
DFFARX1 I_34496 (I589474,I3035,I589084,I589500,);
not I_34497 (I589508,I589500);
nor I_34498 (I589070,I589508,I589313);
nand I_34499 (I589539,I589508,I589158);
not I_34500 (I589556,I252221);
nand I_34501 (I589573,I589556,I589262);
nand I_34502 (I589590,I589508,I589573);
nand I_34503 (I589061,I589590,I589539);
nand I_34504 (I589058,I589573,I589457);
not I_34505 (I589662,I3042);
DFFARX1 I_34506 (I210931,I3035,I589662,I589688,);
and I_34507 (I589696,I589688,I210916);
DFFARX1 I_34508 (I589696,I3035,I589662,I589645,);
DFFARX1 I_34509 (I210922,I3035,I589662,I589736,);
not I_34510 (I589744,I210904);
not I_34511 (I589761,I210925);
nand I_34512 (I589778,I589761,I589744);
nor I_34513 (I589633,I589736,I589778);
DFFARX1 I_34514 (I589778,I3035,I589662,I589818,);
not I_34515 (I589654,I589818);
not I_34516 (I589840,I210928);
nand I_34517 (I589857,I589761,I589840);
DFFARX1 I_34518 (I589857,I3035,I589662,I589883,);
not I_34519 (I589891,I589883);
not I_34520 (I589908,I210919);
nand I_34521 (I589925,I589908,I210907);
and I_34522 (I589942,I589744,I589925);
nor I_34523 (I589959,I589857,I589942);
DFFARX1 I_34524 (I589959,I3035,I589662,I589630,);
DFFARX1 I_34525 (I589942,I3035,I589662,I589651,);
nor I_34526 (I590004,I210919,I210913);
nor I_34527 (I589642,I589857,I590004);
or I_34528 (I590035,I210919,I210913);
nor I_34529 (I590052,I210910,I210904);
DFFARX1 I_34530 (I590052,I3035,I589662,I590078,);
not I_34531 (I590086,I590078);
nor I_34532 (I589648,I590086,I589891);
nand I_34533 (I590117,I590086,I589736);
not I_34534 (I590134,I210910);
nand I_34535 (I590151,I590134,I589840);
nand I_34536 (I590168,I590086,I590151);
nand I_34537 (I589639,I590168,I590117);
nand I_34538 (I589636,I590151,I590035);
not I_34539 (I590240,I3042);
DFFARX1 I_34540 (I295414,I3035,I590240,I590266,);
and I_34541 (I590274,I590266,I295429);
DFFARX1 I_34542 (I590274,I3035,I590240,I590223,);
DFFARX1 I_34543 (I295420,I3035,I590240,I590314,);
not I_34544 (I590322,I295414);
not I_34545 (I590339,I295432);
nand I_34546 (I590356,I590339,I590322);
nor I_34547 (I590211,I590314,I590356);
DFFARX1 I_34548 (I590356,I3035,I590240,I590396,);
not I_34549 (I590232,I590396);
not I_34550 (I590418,I295423);
nand I_34551 (I590435,I590339,I590418);
DFFARX1 I_34552 (I590435,I3035,I590240,I590461,);
not I_34553 (I590469,I590461);
not I_34554 (I590486,I295435);
nand I_34555 (I590503,I590486,I295411);
and I_34556 (I590520,I590322,I590503);
nor I_34557 (I590537,I590435,I590520);
DFFARX1 I_34558 (I590537,I3035,I590240,I590208,);
DFFARX1 I_34559 (I590520,I3035,I590240,I590229,);
nor I_34560 (I590582,I295435,I295411);
nor I_34561 (I590220,I590435,I590582);
or I_34562 (I590613,I295435,I295411);
nor I_34563 (I590630,I295417,I295426);
DFFARX1 I_34564 (I590630,I3035,I590240,I590656,);
not I_34565 (I590664,I590656);
nor I_34566 (I590226,I590664,I590469);
nand I_34567 (I590695,I590664,I590314);
not I_34568 (I590712,I295417);
nand I_34569 (I590729,I590712,I590418);
nand I_34570 (I590746,I590664,I590729);
nand I_34571 (I590217,I590746,I590695);
nand I_34572 (I590214,I590729,I590613);
not I_34573 (I590818,I3042);
DFFARX1 I_34574 (I154542,I3035,I590818,I590844,);
and I_34575 (I590852,I590844,I154527);
DFFARX1 I_34576 (I590852,I3035,I590818,I590801,);
DFFARX1 I_34577 (I154533,I3035,I590818,I590892,);
not I_34578 (I590900,I154515);
not I_34579 (I590917,I154536);
nand I_34580 (I590934,I590917,I590900);
nor I_34581 (I590789,I590892,I590934);
DFFARX1 I_34582 (I590934,I3035,I590818,I590974,);
not I_34583 (I590810,I590974);
not I_34584 (I590996,I154539);
nand I_34585 (I591013,I590917,I590996);
DFFARX1 I_34586 (I591013,I3035,I590818,I591039,);
not I_34587 (I591047,I591039);
not I_34588 (I591064,I154530);
nand I_34589 (I591081,I591064,I154518);
and I_34590 (I591098,I590900,I591081);
nor I_34591 (I591115,I591013,I591098);
DFFARX1 I_34592 (I591115,I3035,I590818,I590786,);
DFFARX1 I_34593 (I591098,I3035,I590818,I590807,);
nor I_34594 (I591160,I154530,I154524);
nor I_34595 (I590798,I591013,I591160);
or I_34596 (I591191,I154530,I154524);
nor I_34597 (I591208,I154521,I154515);
DFFARX1 I_34598 (I591208,I3035,I590818,I591234,);
not I_34599 (I591242,I591234);
nor I_34600 (I590804,I591242,I591047);
nand I_34601 (I591273,I591242,I590892);
not I_34602 (I591290,I154521);
nand I_34603 (I591307,I591290,I590996);
nand I_34604 (I591324,I591242,I591307);
nand I_34605 (I590795,I591324,I591273);
nand I_34606 (I590792,I591307,I591191);
not I_34607 (I591396,I3042);
DFFARX1 I_34608 (I385135,I3035,I591396,I591422,);
and I_34609 (I591430,I591422,I385123);
DFFARX1 I_34610 (I591430,I3035,I591396,I591379,);
DFFARX1 I_34611 (I385126,I3035,I591396,I591470,);
not I_34612 (I591478,I385120);
not I_34613 (I591495,I385144);
nand I_34614 (I591512,I591495,I591478);
nor I_34615 (I591367,I591470,I591512);
DFFARX1 I_34616 (I591512,I3035,I591396,I591552,);
not I_34617 (I591388,I591552);
not I_34618 (I591574,I385132);
nand I_34619 (I591591,I591495,I591574);
DFFARX1 I_34620 (I591591,I3035,I591396,I591617,);
not I_34621 (I591625,I591617);
not I_34622 (I591642,I385141);
nand I_34623 (I591659,I591642,I385138);
and I_34624 (I591676,I591478,I591659);
nor I_34625 (I591693,I591591,I591676);
DFFARX1 I_34626 (I591693,I3035,I591396,I591364,);
DFFARX1 I_34627 (I591676,I3035,I591396,I591385,);
nor I_34628 (I591738,I385141,I385129);
nor I_34629 (I591376,I591591,I591738);
or I_34630 (I591769,I385141,I385129);
nor I_34631 (I591786,I385120,I385123);
DFFARX1 I_34632 (I591786,I3035,I591396,I591812,);
not I_34633 (I591820,I591812);
nor I_34634 (I591382,I591820,I591625);
nand I_34635 (I591851,I591820,I591470);
not I_34636 (I591868,I385120);
nand I_34637 (I591885,I591868,I591574);
nand I_34638 (I591902,I591820,I591885);
nand I_34639 (I591373,I591902,I591851);
nand I_34640 (I591370,I591885,I591769);
not I_34641 (I591974,I3042);
DFFARX1 I_34642 (I413457,I3035,I591974,I592000,);
and I_34643 (I592008,I592000,I413445);
DFFARX1 I_34644 (I592008,I3035,I591974,I591957,);
DFFARX1 I_34645 (I413448,I3035,I591974,I592048,);
not I_34646 (I592056,I413442);
not I_34647 (I592073,I413466);
nand I_34648 (I592090,I592073,I592056);
nor I_34649 (I591945,I592048,I592090);
DFFARX1 I_34650 (I592090,I3035,I591974,I592130,);
not I_34651 (I591966,I592130);
not I_34652 (I592152,I413454);
nand I_34653 (I592169,I592073,I592152);
DFFARX1 I_34654 (I592169,I3035,I591974,I592195,);
not I_34655 (I592203,I592195);
not I_34656 (I592220,I413463);
nand I_34657 (I592237,I592220,I413460);
and I_34658 (I592254,I592056,I592237);
nor I_34659 (I592271,I592169,I592254);
DFFARX1 I_34660 (I592271,I3035,I591974,I591942,);
DFFARX1 I_34661 (I592254,I3035,I591974,I591963,);
nor I_34662 (I592316,I413463,I413451);
nor I_34663 (I591954,I592169,I592316);
or I_34664 (I592347,I413463,I413451);
nor I_34665 (I592364,I413442,I413445);
DFFARX1 I_34666 (I592364,I3035,I591974,I592390,);
not I_34667 (I592398,I592390);
nor I_34668 (I591960,I592398,I592203);
nand I_34669 (I592429,I592398,I592048);
not I_34670 (I592446,I413442);
nand I_34671 (I592463,I592446,I592152);
nand I_34672 (I592480,I592398,I592463);
nand I_34673 (I591951,I592480,I592429);
nand I_34674 (I591948,I592463,I592347);
not I_34675 (I592552,I3042);
DFFARX1 I_34676 (I55259,I3035,I592552,I592578,);
and I_34677 (I592586,I592578,I55235);
DFFARX1 I_34678 (I592586,I3035,I592552,I592535,);
DFFARX1 I_34679 (I55253,I3035,I592552,I592626,);
not I_34680 (I592634,I55241);
not I_34681 (I592651,I55238);
nand I_34682 (I592668,I592651,I592634);
nor I_34683 (I592523,I592626,I592668);
DFFARX1 I_34684 (I592668,I3035,I592552,I592708,);
not I_34685 (I592544,I592708);
not I_34686 (I592730,I55247);
nand I_34687 (I592747,I592651,I592730);
DFFARX1 I_34688 (I592747,I3035,I592552,I592773,);
not I_34689 (I592781,I592773);
not I_34690 (I592798,I55238);
nand I_34691 (I592815,I592798,I55256);
and I_34692 (I592832,I592634,I592815);
nor I_34693 (I592849,I592747,I592832);
DFFARX1 I_34694 (I592849,I3035,I592552,I592520,);
DFFARX1 I_34695 (I592832,I3035,I592552,I592541,);
nor I_34696 (I592894,I55238,I55250);
nor I_34697 (I592532,I592747,I592894);
or I_34698 (I592925,I55238,I55250);
nor I_34699 (I592942,I55244,I55235);
DFFARX1 I_34700 (I592942,I3035,I592552,I592968,);
not I_34701 (I592976,I592968);
nor I_34702 (I592538,I592976,I592781);
nand I_34703 (I593007,I592976,I592626);
not I_34704 (I593024,I55244);
nand I_34705 (I593041,I593024,I592730);
nand I_34706 (I593058,I592976,I593041);
nand I_34707 (I592529,I593058,I593007);
nand I_34708 (I592526,I593041,I592925);
not I_34709 (I593130,I3042);
DFFARX1 I_34710 (I217782,I3035,I593130,I593156,);
and I_34711 (I593164,I593156,I217767);
DFFARX1 I_34712 (I593164,I3035,I593130,I593113,);
DFFARX1 I_34713 (I217773,I3035,I593130,I593204,);
not I_34714 (I593212,I217755);
not I_34715 (I593229,I217776);
nand I_34716 (I593246,I593229,I593212);
nor I_34717 (I593101,I593204,I593246);
DFFARX1 I_34718 (I593246,I3035,I593130,I593286,);
not I_34719 (I593122,I593286);
not I_34720 (I593308,I217779);
nand I_34721 (I593325,I593229,I593308);
DFFARX1 I_34722 (I593325,I3035,I593130,I593351,);
not I_34723 (I593359,I593351);
not I_34724 (I593376,I217770);
nand I_34725 (I593393,I593376,I217758);
and I_34726 (I593410,I593212,I593393);
nor I_34727 (I593427,I593325,I593410);
DFFARX1 I_34728 (I593427,I3035,I593130,I593098,);
DFFARX1 I_34729 (I593410,I3035,I593130,I593119,);
nor I_34730 (I593472,I217770,I217764);
nor I_34731 (I593110,I593325,I593472);
or I_34732 (I593503,I217770,I217764);
nor I_34733 (I593520,I217761,I217755);
DFFARX1 I_34734 (I593520,I3035,I593130,I593546,);
not I_34735 (I593554,I593546);
nor I_34736 (I593116,I593554,I593359);
nand I_34737 (I593585,I593554,I593204);
not I_34738 (I593602,I217761);
nand I_34739 (I593619,I593602,I593308);
nand I_34740 (I593636,I593554,I593619);
nand I_34741 (I593107,I593636,I593585);
nand I_34742 (I593104,I593619,I593503);
not I_34743 (I593708,I3042);
DFFARX1 I_34744 (I297794,I3035,I593708,I593734,);
and I_34745 (I593742,I593734,I297809);
DFFARX1 I_34746 (I593742,I3035,I593708,I593691,);
DFFARX1 I_34747 (I297800,I3035,I593708,I593782,);
not I_34748 (I593790,I297794);
not I_34749 (I593807,I297812);
nand I_34750 (I593824,I593807,I593790);
nor I_34751 (I593679,I593782,I593824);
DFFARX1 I_34752 (I593824,I3035,I593708,I593864,);
not I_34753 (I593700,I593864);
not I_34754 (I593886,I297803);
nand I_34755 (I593903,I593807,I593886);
DFFARX1 I_34756 (I593903,I3035,I593708,I593929,);
not I_34757 (I593937,I593929);
not I_34758 (I593954,I297815);
nand I_34759 (I593971,I593954,I297791);
and I_34760 (I593988,I593790,I593971);
nor I_34761 (I594005,I593903,I593988);
DFFARX1 I_34762 (I594005,I3035,I593708,I593676,);
DFFARX1 I_34763 (I593988,I3035,I593708,I593697,);
nor I_34764 (I594050,I297815,I297791);
nor I_34765 (I593688,I593903,I594050);
or I_34766 (I594081,I297815,I297791);
nor I_34767 (I594098,I297797,I297806);
DFFARX1 I_34768 (I594098,I3035,I593708,I594124,);
not I_34769 (I594132,I594124);
nor I_34770 (I593694,I594132,I593937);
nand I_34771 (I594163,I594132,I593782);
not I_34772 (I594180,I297797);
nand I_34773 (I594197,I594180,I593886);
nand I_34774 (I594214,I594132,I594197);
nand I_34775 (I593685,I594214,I594163);
nand I_34776 (I593682,I594197,I594081);
not I_34777 (I594286,I3042);
DFFARX1 I_34778 (I271237,I3035,I594286,I594312,);
and I_34779 (I594320,I594312,I271252);
DFFARX1 I_34780 (I594320,I3035,I594286,I594269,);
DFFARX1 I_34781 (I271255,I3035,I594286,I594360,);
not I_34782 (I594368,I271249);
not I_34783 (I594385,I271264);
nand I_34784 (I594402,I594385,I594368);
nor I_34785 (I594257,I594360,I594402);
DFFARX1 I_34786 (I594402,I3035,I594286,I594442,);
not I_34787 (I594278,I594442);
not I_34788 (I594464,I271240);
nand I_34789 (I594481,I594385,I594464);
DFFARX1 I_34790 (I594481,I3035,I594286,I594507,);
not I_34791 (I594515,I594507);
not I_34792 (I594532,I271243);
nand I_34793 (I594549,I594532,I271237);
and I_34794 (I594566,I594368,I594549);
nor I_34795 (I594583,I594481,I594566);
DFFARX1 I_34796 (I594583,I3035,I594286,I594254,);
DFFARX1 I_34797 (I594566,I3035,I594286,I594275,);
nor I_34798 (I594628,I271243,I271246);
nor I_34799 (I594266,I594481,I594628);
or I_34800 (I594659,I271243,I271246);
nor I_34801 (I594676,I271261,I271258);
DFFARX1 I_34802 (I594676,I3035,I594286,I594702,);
not I_34803 (I594710,I594702);
nor I_34804 (I594272,I594710,I594515);
nand I_34805 (I594741,I594710,I594360);
not I_34806 (I594758,I271261);
nand I_34807 (I594775,I594758,I594464);
nand I_34808 (I594792,I594710,I594775);
nand I_34809 (I594263,I594792,I594741);
nand I_34810 (I594260,I594775,I594659);
not I_34811 (I594864,I3042);
DFFARX1 I_34812 (I167717,I3035,I594864,I594890,);
and I_34813 (I594898,I594890,I167702);
DFFARX1 I_34814 (I594898,I3035,I594864,I594847,);
DFFARX1 I_34815 (I167708,I3035,I594864,I594938,);
not I_34816 (I594946,I167690);
not I_34817 (I594963,I167711);
nand I_34818 (I594980,I594963,I594946);
nor I_34819 (I594835,I594938,I594980);
DFFARX1 I_34820 (I594980,I3035,I594864,I595020,);
not I_34821 (I594856,I595020);
not I_34822 (I595042,I167714);
nand I_34823 (I595059,I594963,I595042);
DFFARX1 I_34824 (I595059,I3035,I594864,I595085,);
not I_34825 (I595093,I595085);
not I_34826 (I595110,I167705);
nand I_34827 (I595127,I595110,I167693);
and I_34828 (I595144,I594946,I595127);
nor I_34829 (I595161,I595059,I595144);
DFFARX1 I_34830 (I595161,I3035,I594864,I594832,);
DFFARX1 I_34831 (I595144,I3035,I594864,I594853,);
nor I_34832 (I595206,I167705,I167699);
nor I_34833 (I594844,I595059,I595206);
or I_34834 (I595237,I167705,I167699);
nor I_34835 (I595254,I167696,I167690);
DFFARX1 I_34836 (I595254,I3035,I594864,I595280,);
not I_34837 (I595288,I595280);
nor I_34838 (I594850,I595288,I595093);
nand I_34839 (I595319,I595288,I594938);
not I_34840 (I595336,I167696);
nand I_34841 (I595353,I595336,I595042);
nand I_34842 (I595370,I595288,I595353);
nand I_34843 (I594841,I595370,I595319);
nand I_34844 (I594838,I595353,I595237);
not I_34845 (I595442,I3042);
DFFARX1 I_34846 (I288274,I3035,I595442,I595468,);
and I_34847 (I595476,I595468,I288289);
DFFARX1 I_34848 (I595476,I3035,I595442,I595425,);
DFFARX1 I_34849 (I288280,I3035,I595442,I595516,);
not I_34850 (I595524,I288274);
not I_34851 (I595541,I288292);
nand I_34852 (I595558,I595541,I595524);
nor I_34853 (I595413,I595516,I595558);
DFFARX1 I_34854 (I595558,I3035,I595442,I595598,);
not I_34855 (I595434,I595598);
not I_34856 (I595620,I288283);
nand I_34857 (I595637,I595541,I595620);
DFFARX1 I_34858 (I595637,I3035,I595442,I595663,);
not I_34859 (I595671,I595663);
not I_34860 (I595688,I288295);
nand I_34861 (I595705,I595688,I288271);
and I_34862 (I595722,I595524,I595705);
nor I_34863 (I595739,I595637,I595722);
DFFARX1 I_34864 (I595739,I3035,I595442,I595410,);
DFFARX1 I_34865 (I595722,I3035,I595442,I595431,);
nor I_34866 (I595784,I288295,I288271);
nor I_34867 (I595422,I595637,I595784);
or I_34868 (I595815,I288295,I288271);
nor I_34869 (I595832,I288277,I288286);
DFFARX1 I_34870 (I595832,I3035,I595442,I595858,);
not I_34871 (I595866,I595858);
nor I_34872 (I595428,I595866,I595671);
nand I_34873 (I595897,I595866,I595516);
not I_34874 (I595914,I288277);
nand I_34875 (I595931,I595914,I595620);
nand I_34876 (I595948,I595866,I595931);
nand I_34877 (I595419,I595948,I595897);
nand I_34878 (I595416,I595931,I595815);
not I_34879 (I596020,I3042);
DFFARX1 I_34880 (I330803,I3035,I596020,I596046,);
and I_34881 (I596054,I596046,I330791);
DFFARX1 I_34882 (I596054,I3035,I596020,I596003,);
DFFARX1 I_34883 (I330806,I3035,I596020,I596094,);
not I_34884 (I596102,I330797);
not I_34885 (I596119,I330788);
nand I_34886 (I596136,I596119,I596102);
nor I_34887 (I595991,I596094,I596136);
DFFARX1 I_34888 (I596136,I3035,I596020,I596176,);
not I_34889 (I596012,I596176);
not I_34890 (I596198,I330794);
nand I_34891 (I596215,I596119,I596198);
DFFARX1 I_34892 (I596215,I3035,I596020,I596241,);
not I_34893 (I596249,I596241);
not I_34894 (I596266,I330809);
nand I_34895 (I596283,I596266,I330812);
and I_34896 (I596300,I596102,I596283);
nor I_34897 (I596317,I596215,I596300);
DFFARX1 I_34898 (I596317,I3035,I596020,I595988,);
DFFARX1 I_34899 (I596300,I3035,I596020,I596009,);
nor I_34900 (I596362,I330809,I330788);
nor I_34901 (I596000,I596215,I596362);
or I_34902 (I596393,I330809,I330788);
nor I_34903 (I596410,I330800,I330791);
DFFARX1 I_34904 (I596410,I3035,I596020,I596436,);
not I_34905 (I596444,I596436);
nor I_34906 (I596006,I596444,I596249);
nand I_34907 (I596475,I596444,I596094);
not I_34908 (I596492,I330800);
nand I_34909 (I596509,I596492,I596198);
nand I_34910 (I596526,I596444,I596509);
nand I_34911 (I595997,I596526,I596475);
nand I_34912 (I595994,I596509,I596393);
not I_34913 (I596598,I3042);
DFFARX1 I_34914 (I724025,I3035,I596598,I596624,);
and I_34915 (I596632,I596624,I724007);
DFFARX1 I_34916 (I596632,I3035,I596598,I596581,);
DFFARX1 I_34917 (I723998,I3035,I596598,I596672,);
not I_34918 (I596680,I724013);
not I_34919 (I596697,I724001);
nand I_34920 (I596714,I596697,I596680);
nor I_34921 (I596569,I596672,I596714);
DFFARX1 I_34922 (I596714,I3035,I596598,I596754,);
not I_34923 (I596590,I596754);
not I_34924 (I596776,I724010);
nand I_34925 (I596793,I596697,I596776);
DFFARX1 I_34926 (I596793,I3035,I596598,I596819,);
not I_34927 (I596827,I596819);
not I_34928 (I596844,I724019);
nand I_34929 (I596861,I596844,I723998);
and I_34930 (I596878,I596680,I596861);
nor I_34931 (I596895,I596793,I596878);
DFFARX1 I_34932 (I596895,I3035,I596598,I596566,);
DFFARX1 I_34933 (I596878,I3035,I596598,I596587,);
nor I_34934 (I596940,I724019,I724022);
nor I_34935 (I596578,I596793,I596940);
or I_34936 (I596971,I724019,I724022);
nor I_34937 (I596988,I724016,I724004);
DFFARX1 I_34938 (I596988,I3035,I596598,I597014,);
not I_34939 (I597022,I597014);
nor I_34940 (I596584,I597022,I596827);
nand I_34941 (I597053,I597022,I596672);
not I_34942 (I597070,I724016);
nand I_34943 (I597087,I597070,I596776);
nand I_34944 (I597104,I597022,I597087);
nand I_34945 (I596575,I597104,I597053);
nand I_34946 (I596572,I597087,I596971);
not I_34947 (I597176,I3042);
DFFARX1 I_34948 (I61583,I3035,I597176,I597202,);
and I_34949 (I597210,I597202,I61559);
DFFARX1 I_34950 (I597210,I3035,I597176,I597159,);
DFFARX1 I_34951 (I61577,I3035,I597176,I597250,);
not I_34952 (I597258,I61565);
not I_34953 (I597275,I61562);
nand I_34954 (I597292,I597275,I597258);
nor I_34955 (I597147,I597250,I597292);
DFFARX1 I_34956 (I597292,I3035,I597176,I597332,);
not I_34957 (I597168,I597332);
not I_34958 (I597354,I61571);
nand I_34959 (I597371,I597275,I597354);
DFFARX1 I_34960 (I597371,I3035,I597176,I597397,);
not I_34961 (I597405,I597397);
not I_34962 (I597422,I61562);
nand I_34963 (I597439,I597422,I61580);
and I_34964 (I597456,I597258,I597439);
nor I_34965 (I597473,I597371,I597456);
DFFARX1 I_34966 (I597473,I3035,I597176,I597144,);
DFFARX1 I_34967 (I597456,I3035,I597176,I597165,);
nor I_34968 (I597518,I61562,I61574);
nor I_34969 (I597156,I597371,I597518);
or I_34970 (I597549,I61562,I61574);
nor I_34971 (I597566,I61568,I61559);
DFFARX1 I_34972 (I597566,I3035,I597176,I597592,);
not I_34973 (I597600,I597592);
nor I_34974 (I597162,I597600,I597405);
nand I_34975 (I597631,I597600,I597250);
not I_34976 (I597648,I61568);
nand I_34977 (I597665,I597648,I597354);
nand I_34978 (I597682,I597600,I597665);
nand I_34979 (I597153,I597682,I597631);
nand I_34980 (I597150,I597665,I597549);
not I_34981 (I597754,I3042);
DFFARX1 I_34982 (I307683,I3035,I597754,I597780,);
and I_34983 (I597788,I597780,I307671);
DFFARX1 I_34984 (I597788,I3035,I597754,I597737,);
DFFARX1 I_34985 (I307686,I3035,I597754,I597828,);
not I_34986 (I597836,I307677);
not I_34987 (I597853,I307668);
nand I_34988 (I597870,I597853,I597836);
nor I_34989 (I597725,I597828,I597870);
DFFARX1 I_34990 (I597870,I3035,I597754,I597910,);
not I_34991 (I597746,I597910);
not I_34992 (I597932,I307674);
nand I_34993 (I597949,I597853,I597932);
DFFARX1 I_34994 (I597949,I3035,I597754,I597975,);
not I_34995 (I597983,I597975);
not I_34996 (I598000,I307689);
nand I_34997 (I598017,I598000,I307692);
and I_34998 (I598034,I597836,I598017);
nor I_34999 (I598051,I597949,I598034);
DFFARX1 I_35000 (I598051,I3035,I597754,I597722,);
DFFARX1 I_35001 (I598034,I3035,I597754,I597743,);
nor I_35002 (I598096,I307689,I307668);
nor I_35003 (I597734,I597949,I598096);
or I_35004 (I598127,I307689,I307668);
nor I_35005 (I598144,I307680,I307671);
DFFARX1 I_35006 (I598144,I3035,I597754,I598170,);
not I_35007 (I598178,I598170);
nor I_35008 (I597740,I598178,I597983);
nand I_35009 (I598209,I598178,I597828);
not I_35010 (I598226,I307680);
nand I_35011 (I598243,I598226,I597932);
nand I_35012 (I598260,I598178,I598243);
nand I_35013 (I597731,I598260,I598209);
nand I_35014 (I597728,I598243,I598127);
not I_35015 (I598332,I3042);
DFFARX1 I_35016 (I562195,I3035,I598332,I598358,);
and I_35017 (I598366,I598358,I562192);
DFFARX1 I_35018 (I598366,I3035,I598332,I598315,);
DFFARX1 I_35019 (I562198,I3035,I598332,I598406,);
not I_35020 (I598414,I562201);
not I_35021 (I598431,I562195);
nand I_35022 (I598448,I598431,I598414);
nor I_35023 (I598303,I598406,I598448);
DFFARX1 I_35024 (I598448,I3035,I598332,I598488,);
not I_35025 (I598324,I598488);
not I_35026 (I598510,I562210);
nand I_35027 (I598527,I598431,I598510);
DFFARX1 I_35028 (I598527,I3035,I598332,I598553,);
not I_35029 (I598561,I598553);
not I_35030 (I598578,I562207);
nand I_35031 (I598595,I598578,I562213);
and I_35032 (I598612,I598414,I598595);
nor I_35033 (I598629,I598527,I598612);
DFFARX1 I_35034 (I598629,I3035,I598332,I598300,);
DFFARX1 I_35035 (I598612,I3035,I598332,I598321,);
nor I_35036 (I598674,I562207,I562192);
nor I_35037 (I598312,I598527,I598674);
or I_35038 (I598705,I562207,I562192);
nor I_35039 (I598722,I562204,I562198);
DFFARX1 I_35040 (I598722,I3035,I598332,I598748,);
not I_35041 (I598756,I598748);
nor I_35042 (I598318,I598756,I598561);
nand I_35043 (I598787,I598756,I598406);
not I_35044 (I598804,I562204);
nand I_35045 (I598821,I598804,I598510);
nand I_35046 (I598838,I598756,I598821);
nand I_35047 (I598309,I598838,I598787);
nand I_35048 (I598306,I598821,I598705);
not I_35049 (I598910,I3042);
DFFARX1 I_35050 (I185635,I3035,I598910,I598936,);
and I_35051 (I598944,I598936,I185620);
DFFARX1 I_35052 (I598944,I3035,I598910,I598893,);
DFFARX1 I_35053 (I185626,I3035,I598910,I598984,);
not I_35054 (I598992,I185608);
not I_35055 (I599009,I185629);
nand I_35056 (I599026,I599009,I598992);
nor I_35057 (I598881,I598984,I599026);
DFFARX1 I_35058 (I599026,I3035,I598910,I599066,);
not I_35059 (I598902,I599066);
not I_35060 (I599088,I185632);
nand I_35061 (I599105,I599009,I599088);
DFFARX1 I_35062 (I599105,I3035,I598910,I599131,);
not I_35063 (I599139,I599131);
not I_35064 (I599156,I185623);
nand I_35065 (I599173,I599156,I185611);
and I_35066 (I599190,I598992,I599173);
nor I_35067 (I599207,I599105,I599190);
DFFARX1 I_35068 (I599207,I3035,I598910,I598878,);
DFFARX1 I_35069 (I599190,I3035,I598910,I598899,);
nor I_35070 (I599252,I185623,I185617);
nor I_35071 (I598890,I599105,I599252);
or I_35072 (I599283,I185623,I185617);
nor I_35073 (I599300,I185614,I185608);
DFFARX1 I_35074 (I599300,I3035,I598910,I599326,);
not I_35075 (I599334,I599326);
nor I_35076 (I598896,I599334,I599139);
nand I_35077 (I599365,I599334,I598984);
not I_35078 (I599382,I185614);
nand I_35079 (I599399,I599382,I599088);
nand I_35080 (I599416,I599334,I599399);
nand I_35081 (I598887,I599416,I599365);
nand I_35082 (I598884,I599399,I599283);
not I_35083 (I599488,I3042);
DFFARX1 I_35084 (I741280,I3035,I599488,I599514,);
and I_35085 (I599522,I599514,I741262);
DFFARX1 I_35086 (I599522,I3035,I599488,I599471,);
DFFARX1 I_35087 (I741253,I3035,I599488,I599562,);
not I_35088 (I599570,I741268);
not I_35089 (I599587,I741256);
nand I_35090 (I599604,I599587,I599570);
nor I_35091 (I599459,I599562,I599604);
DFFARX1 I_35092 (I599604,I3035,I599488,I599644,);
not I_35093 (I599480,I599644);
not I_35094 (I599666,I741265);
nand I_35095 (I599683,I599587,I599666);
DFFARX1 I_35096 (I599683,I3035,I599488,I599709,);
not I_35097 (I599717,I599709);
not I_35098 (I599734,I741274);
nand I_35099 (I599751,I599734,I741253);
and I_35100 (I599768,I599570,I599751);
nor I_35101 (I599785,I599683,I599768);
DFFARX1 I_35102 (I599785,I3035,I599488,I599456,);
DFFARX1 I_35103 (I599768,I3035,I599488,I599477,);
nor I_35104 (I599830,I741274,I741277);
nor I_35105 (I599468,I599683,I599830);
or I_35106 (I599861,I741274,I741277);
nor I_35107 (I599878,I741271,I741259);
DFFARX1 I_35108 (I599878,I3035,I599488,I599904,);
not I_35109 (I599912,I599904);
nor I_35110 (I599474,I599912,I599717);
nand I_35111 (I599943,I599912,I599562);
not I_35112 (I599960,I741271);
nand I_35113 (I599977,I599960,I599666);
nand I_35114 (I599994,I599912,I599977);
nand I_35115 (I599465,I599994,I599943);
nand I_35116 (I599462,I599977,I599861);
not I_35117 (I600066,I3042);
DFFARX1 I_35118 (I370685,I3035,I600066,I600092,);
and I_35119 (I600100,I600092,I370673);
DFFARX1 I_35120 (I600100,I3035,I600066,I600049,);
DFFARX1 I_35121 (I370676,I3035,I600066,I600140,);
not I_35122 (I600148,I370670);
not I_35123 (I600165,I370694);
nand I_35124 (I600182,I600165,I600148);
nor I_35125 (I600037,I600140,I600182);
DFFARX1 I_35126 (I600182,I3035,I600066,I600222,);
not I_35127 (I600058,I600222);
not I_35128 (I600244,I370682);
nand I_35129 (I600261,I600165,I600244);
DFFARX1 I_35130 (I600261,I3035,I600066,I600287,);
not I_35131 (I600295,I600287);
not I_35132 (I600312,I370691);
nand I_35133 (I600329,I600312,I370688);
and I_35134 (I600346,I600148,I600329);
nor I_35135 (I600363,I600261,I600346);
DFFARX1 I_35136 (I600363,I3035,I600066,I600034,);
DFFARX1 I_35137 (I600346,I3035,I600066,I600055,);
nor I_35138 (I600408,I370691,I370679);
nor I_35139 (I600046,I600261,I600408);
or I_35140 (I600439,I370691,I370679);
nor I_35141 (I600456,I370670,I370673);
DFFARX1 I_35142 (I600456,I3035,I600066,I600482,);
not I_35143 (I600490,I600482);
nor I_35144 (I600052,I600490,I600295);
nand I_35145 (I600521,I600490,I600140);
not I_35146 (I600538,I370670);
nand I_35147 (I600555,I600538,I600244);
nand I_35148 (I600572,I600490,I600555);
nand I_35149 (I600043,I600572,I600521);
nand I_35150 (I600040,I600555,I600439);
not I_35151 (I600644,I3042);
DFFARX1 I_35152 (I540030,I3035,I600644,I600670,);
and I_35153 (I600678,I600670,I540024);
DFFARX1 I_35154 (I600678,I3035,I600644,I600627,);
DFFARX1 I_35155 (I540042,I3035,I600644,I600718,);
not I_35156 (I600726,I540033);
not I_35157 (I600743,I540045);
nand I_35158 (I600760,I600743,I600726);
nor I_35159 (I600615,I600718,I600760);
DFFARX1 I_35160 (I600760,I3035,I600644,I600800,);
not I_35161 (I600636,I600800);
not I_35162 (I600822,I540051);
nand I_35163 (I600839,I600743,I600822);
DFFARX1 I_35164 (I600839,I3035,I600644,I600865,);
not I_35165 (I600873,I600865);
not I_35166 (I600890,I540027);
nand I_35167 (I600907,I600890,I540048);
and I_35168 (I600924,I600726,I600907);
nor I_35169 (I600941,I600839,I600924);
DFFARX1 I_35170 (I600941,I3035,I600644,I600612,);
DFFARX1 I_35171 (I600924,I3035,I600644,I600633,);
nor I_35172 (I600986,I540027,I540039);
nor I_35173 (I600624,I600839,I600986);
or I_35174 (I601017,I540027,I540039);
nor I_35175 (I601034,I540024,I540036);
DFFARX1 I_35176 (I601034,I3035,I600644,I601060,);
not I_35177 (I601068,I601060);
nor I_35178 (I600630,I601068,I600873);
nand I_35179 (I601099,I601068,I600718);
not I_35180 (I601116,I540024);
nand I_35181 (I601133,I601116,I600822);
nand I_35182 (I601150,I601068,I601133);
nand I_35183 (I600621,I601150,I601099);
nand I_35184 (I600618,I601133,I601017);
not I_35185 (I601222,I3042);
DFFARX1 I_35186 (I187743,I3035,I601222,I601248,);
and I_35187 (I601256,I601248,I187728);
DFFARX1 I_35188 (I601256,I3035,I601222,I601205,);
DFFARX1 I_35189 (I187734,I3035,I601222,I601296,);
not I_35190 (I601304,I187716);
not I_35191 (I601321,I187737);
nand I_35192 (I601338,I601321,I601304);
nor I_35193 (I601193,I601296,I601338);
DFFARX1 I_35194 (I601338,I3035,I601222,I601378,);
not I_35195 (I601214,I601378);
not I_35196 (I601400,I187740);
nand I_35197 (I601417,I601321,I601400);
DFFARX1 I_35198 (I601417,I3035,I601222,I601443,);
not I_35199 (I601451,I601443);
not I_35200 (I601468,I187731);
nand I_35201 (I601485,I601468,I187719);
and I_35202 (I601502,I601304,I601485);
nor I_35203 (I601519,I601417,I601502);
DFFARX1 I_35204 (I601519,I3035,I601222,I601190,);
DFFARX1 I_35205 (I601502,I3035,I601222,I601211,);
nor I_35206 (I601564,I187731,I187725);
nor I_35207 (I601202,I601417,I601564);
or I_35208 (I601595,I187731,I187725);
nor I_35209 (I601612,I187722,I187716);
DFFARX1 I_35210 (I601612,I3035,I601222,I601638,);
not I_35211 (I601646,I601638);
nor I_35212 (I601208,I601646,I601451);
nand I_35213 (I601677,I601646,I601296);
not I_35214 (I601694,I187722);
nand I_35215 (I601711,I601694,I601400);
nand I_35216 (I601728,I601646,I601711);
nand I_35217 (I601199,I601728,I601677);
nand I_35218 (I601196,I601711,I601595);
not I_35219 (I601800,I3042);
DFFARX1 I_35220 (I130069,I3035,I601800,I601826,);
and I_35221 (I601834,I601826,I130072);
DFFARX1 I_35222 (I601834,I3035,I601800,I601783,);
DFFARX1 I_35223 (I130072,I3035,I601800,I601874,);
not I_35224 (I601882,I130087);
not I_35225 (I601899,I130093);
nand I_35226 (I601916,I601899,I601882);
nor I_35227 (I601771,I601874,I601916);
DFFARX1 I_35228 (I601916,I3035,I601800,I601956,);
not I_35229 (I601792,I601956);
not I_35230 (I601978,I130081);
nand I_35231 (I601995,I601899,I601978);
DFFARX1 I_35232 (I601995,I3035,I601800,I602021,);
not I_35233 (I602029,I602021);
not I_35234 (I602046,I130078);
nand I_35235 (I602063,I602046,I130075);
and I_35236 (I602080,I601882,I602063);
nor I_35237 (I602097,I601995,I602080);
DFFARX1 I_35238 (I602097,I3035,I601800,I601768,);
DFFARX1 I_35239 (I602080,I3035,I601800,I601789,);
nor I_35240 (I602142,I130078,I130069);
nor I_35241 (I601780,I601995,I602142);
or I_35242 (I602173,I130078,I130069);
nor I_35243 (I602190,I130084,I130090);
DFFARX1 I_35244 (I602190,I3035,I601800,I602216,);
not I_35245 (I602224,I602216);
nor I_35246 (I601786,I602224,I602029);
nand I_35247 (I602255,I602224,I601874);
not I_35248 (I602272,I130084);
nand I_35249 (I602289,I602272,I601978);
nand I_35250 (I602306,I602224,I602289);
nand I_35251 (I601777,I602306,I602255);
nand I_35252 (I601774,I602289,I602173);
not I_35253 (I602378,I3042);
DFFARX1 I_35254 (I535508,I3035,I602378,I602404,);
and I_35255 (I602412,I602404,I535502);
DFFARX1 I_35256 (I602412,I3035,I602378,I602361,);
DFFARX1 I_35257 (I535520,I3035,I602378,I602452,);
not I_35258 (I602460,I535511);
not I_35259 (I602477,I535523);
nand I_35260 (I602494,I602477,I602460);
nor I_35261 (I602349,I602452,I602494);
DFFARX1 I_35262 (I602494,I3035,I602378,I602534,);
not I_35263 (I602370,I602534);
not I_35264 (I602556,I535529);
nand I_35265 (I602573,I602477,I602556);
DFFARX1 I_35266 (I602573,I3035,I602378,I602599,);
not I_35267 (I602607,I602599);
not I_35268 (I602624,I535505);
nand I_35269 (I602641,I602624,I535526);
and I_35270 (I602658,I602460,I602641);
nor I_35271 (I602675,I602573,I602658);
DFFARX1 I_35272 (I602675,I3035,I602378,I602346,);
DFFARX1 I_35273 (I602658,I3035,I602378,I602367,);
nor I_35274 (I602720,I535505,I535517);
nor I_35275 (I602358,I602573,I602720);
or I_35276 (I602751,I535505,I535517);
nor I_35277 (I602768,I535502,I535514);
DFFARX1 I_35278 (I602768,I3035,I602378,I602794,);
not I_35279 (I602802,I602794);
nor I_35280 (I602364,I602802,I602607);
nand I_35281 (I602833,I602802,I602452);
not I_35282 (I602850,I535502);
nand I_35283 (I602867,I602850,I602556);
nand I_35284 (I602884,I602802,I602867);
nand I_35285 (I602355,I602884,I602833);
nand I_35286 (I602352,I602867,I602751);
not I_35287 (I602956,I3042);
DFFARX1 I_35288 (I428235,I3035,I602956,I602982,);
and I_35289 (I602990,I602982,I428241);
DFFARX1 I_35290 (I602990,I3035,I602956,I602939,);
DFFARX1 I_35291 (I428247,I3035,I602956,I603030,);
not I_35292 (I603038,I428232);
not I_35293 (I603055,I428232);
nand I_35294 (I603072,I603055,I603038);
nor I_35295 (I602927,I603030,I603072);
DFFARX1 I_35296 (I603072,I3035,I602956,I603112,);
not I_35297 (I602948,I603112);
not I_35298 (I603134,I428250);
nand I_35299 (I603151,I603055,I603134);
DFFARX1 I_35300 (I603151,I3035,I602956,I603177,);
not I_35301 (I603185,I603177);
not I_35302 (I603202,I428244);
nand I_35303 (I603219,I603202,I428235);
and I_35304 (I603236,I603038,I603219);
nor I_35305 (I603253,I603151,I603236);
DFFARX1 I_35306 (I603253,I3035,I602956,I602924,);
DFFARX1 I_35307 (I603236,I3035,I602956,I602945,);
nor I_35308 (I603298,I428244,I428253);
nor I_35309 (I602936,I603151,I603298);
or I_35310 (I603329,I428244,I428253);
nor I_35311 (I603346,I428238,I428238);
DFFARX1 I_35312 (I603346,I3035,I602956,I603372,);
not I_35313 (I603380,I603372);
nor I_35314 (I602942,I603380,I603185);
nand I_35315 (I603411,I603380,I603030);
not I_35316 (I603428,I428238);
nand I_35317 (I603445,I603428,I603134);
nand I_35318 (I603462,I603380,I603445);
nand I_35319 (I602933,I603462,I603411);
nand I_35320 (I602930,I603445,I603329);
not I_35321 (I603534,I3042);
DFFARX1 I_35322 (I242949,I3035,I603534,I603560,);
and I_35323 (I603568,I603560,I242964);
DFFARX1 I_35324 (I603568,I3035,I603534,I603517,);
DFFARX1 I_35325 (I242967,I3035,I603534,I603608,);
not I_35326 (I603616,I242961);
not I_35327 (I603633,I242976);
nand I_35328 (I603650,I603633,I603616);
nor I_35329 (I603505,I603608,I603650);
DFFARX1 I_35330 (I603650,I3035,I603534,I603690,);
not I_35331 (I603526,I603690);
not I_35332 (I603712,I242952);
nand I_35333 (I603729,I603633,I603712);
DFFARX1 I_35334 (I603729,I3035,I603534,I603755,);
not I_35335 (I603763,I603755);
not I_35336 (I603780,I242955);
nand I_35337 (I603797,I603780,I242949);
and I_35338 (I603814,I603616,I603797);
nor I_35339 (I603831,I603729,I603814);
DFFARX1 I_35340 (I603831,I3035,I603534,I603502,);
DFFARX1 I_35341 (I603814,I3035,I603534,I603523,);
nor I_35342 (I603876,I242955,I242958);
nor I_35343 (I603514,I603729,I603876);
or I_35344 (I603907,I242955,I242958);
nor I_35345 (I603924,I242973,I242970);
DFFARX1 I_35346 (I603924,I3035,I603534,I603950,);
not I_35347 (I603958,I603950);
nor I_35348 (I603520,I603958,I603763);
nand I_35349 (I603989,I603958,I603608);
not I_35350 (I604006,I242973);
nand I_35351 (I604023,I604006,I603712);
nand I_35352 (I604040,I603958,I604023);
nand I_35353 (I603511,I604040,I603989);
nand I_35354 (I603508,I604023,I603907);
not I_35355 (I604112,I3042);
DFFARX1 I_35356 (I316931,I3035,I604112,I604138,);
and I_35357 (I604146,I604138,I316919);
DFFARX1 I_35358 (I604146,I3035,I604112,I604095,);
DFFARX1 I_35359 (I316934,I3035,I604112,I604186,);
not I_35360 (I604194,I316925);
not I_35361 (I604211,I316916);
nand I_35362 (I604228,I604211,I604194);
nor I_35363 (I604083,I604186,I604228);
DFFARX1 I_35364 (I604228,I3035,I604112,I604268,);
not I_35365 (I604104,I604268);
not I_35366 (I604290,I316922);
nand I_35367 (I604307,I604211,I604290);
DFFARX1 I_35368 (I604307,I3035,I604112,I604333,);
not I_35369 (I604341,I604333);
not I_35370 (I604358,I316937);
nand I_35371 (I604375,I604358,I316940);
and I_35372 (I604392,I604194,I604375);
nor I_35373 (I604409,I604307,I604392);
DFFARX1 I_35374 (I604409,I3035,I604112,I604080,);
DFFARX1 I_35375 (I604392,I3035,I604112,I604101,);
nor I_35376 (I604454,I316937,I316916);
nor I_35377 (I604092,I604307,I604454);
or I_35378 (I604485,I316937,I316916);
nor I_35379 (I604502,I316928,I316919);
DFFARX1 I_35380 (I604502,I3035,I604112,I604528,);
not I_35381 (I604536,I604528);
nor I_35382 (I604098,I604536,I604341);
nand I_35383 (I604567,I604536,I604186);
not I_35384 (I604584,I316928);
nand I_35385 (I604601,I604584,I604290);
nand I_35386 (I604618,I604536,I604601);
nand I_35387 (I604089,I604618,I604567);
nand I_35388 (I604086,I604601,I604485);
not I_35389 (I604690,I3042);
DFFARX1 I_35390 (I233701,I3035,I604690,I604716,);
and I_35391 (I604724,I604716,I233716);
DFFARX1 I_35392 (I604724,I3035,I604690,I604673,);
DFFARX1 I_35393 (I233719,I3035,I604690,I604764,);
not I_35394 (I604772,I233713);
not I_35395 (I604789,I233728);
nand I_35396 (I604806,I604789,I604772);
nor I_35397 (I604661,I604764,I604806);
DFFARX1 I_35398 (I604806,I3035,I604690,I604846,);
not I_35399 (I604682,I604846);
not I_35400 (I604868,I233704);
nand I_35401 (I604885,I604789,I604868);
DFFARX1 I_35402 (I604885,I3035,I604690,I604911,);
not I_35403 (I604919,I604911);
not I_35404 (I604936,I233707);
nand I_35405 (I604953,I604936,I233701);
and I_35406 (I604970,I604772,I604953);
nor I_35407 (I604987,I604885,I604970);
DFFARX1 I_35408 (I604987,I3035,I604690,I604658,);
DFFARX1 I_35409 (I604970,I3035,I604690,I604679,);
nor I_35410 (I605032,I233707,I233710);
nor I_35411 (I604670,I604885,I605032);
or I_35412 (I605063,I233707,I233710);
nor I_35413 (I605080,I233725,I233722);
DFFARX1 I_35414 (I605080,I3035,I604690,I605106,);
not I_35415 (I605114,I605106);
nor I_35416 (I604676,I605114,I604919);
nand I_35417 (I605145,I605114,I604764);
not I_35418 (I605162,I233725);
nand I_35419 (I605179,I605162,I604868);
nand I_35420 (I605196,I605114,I605179);
nand I_35421 (I604667,I605196,I605145);
nand I_35422 (I604664,I605179,I605063);
not I_35423 (I605268,I3042);
DFFARX1 I_35424 (I293034,I3035,I605268,I605294,);
and I_35425 (I605302,I605294,I293049);
DFFARX1 I_35426 (I605302,I3035,I605268,I605251,);
DFFARX1 I_35427 (I293040,I3035,I605268,I605342,);
not I_35428 (I605350,I293034);
not I_35429 (I605367,I293052);
nand I_35430 (I605384,I605367,I605350);
nor I_35431 (I605239,I605342,I605384);
DFFARX1 I_35432 (I605384,I3035,I605268,I605424,);
not I_35433 (I605260,I605424);
not I_35434 (I605446,I293043);
nand I_35435 (I605463,I605367,I605446);
DFFARX1 I_35436 (I605463,I3035,I605268,I605489,);
not I_35437 (I605497,I605489);
not I_35438 (I605514,I293055);
nand I_35439 (I605531,I605514,I293031);
and I_35440 (I605548,I605350,I605531);
nor I_35441 (I605565,I605463,I605548);
DFFARX1 I_35442 (I605565,I3035,I605268,I605236,);
DFFARX1 I_35443 (I605548,I3035,I605268,I605257,);
nor I_35444 (I605610,I293055,I293031);
nor I_35445 (I605248,I605463,I605610);
or I_35446 (I605641,I293055,I293031);
nor I_35447 (I605658,I293037,I293046);
DFFARX1 I_35448 (I605658,I3035,I605268,I605684,);
not I_35449 (I605692,I605684);
nor I_35450 (I605254,I605692,I605497);
nand I_35451 (I605723,I605692,I605342);
not I_35452 (I605740,I293037);
nand I_35453 (I605757,I605740,I605446);
nand I_35454 (I605774,I605692,I605757);
nand I_35455 (I605245,I605774,I605723);
nand I_35456 (I605242,I605757,I605641);
not I_35457 (I605846,I3042);
DFFARX1 I_35458 (I453531,I3035,I605846,I605872,);
and I_35459 (I605880,I605872,I453537);
DFFARX1 I_35460 (I605880,I3035,I605846,I605829,);
DFFARX1 I_35461 (I453543,I3035,I605846,I605920,);
not I_35462 (I605928,I453528);
not I_35463 (I605945,I453528);
nand I_35464 (I605962,I605945,I605928);
nor I_35465 (I605817,I605920,I605962);
DFFARX1 I_35466 (I605962,I3035,I605846,I606002,);
not I_35467 (I605838,I606002);
not I_35468 (I606024,I453546);
nand I_35469 (I606041,I605945,I606024);
DFFARX1 I_35470 (I606041,I3035,I605846,I606067,);
not I_35471 (I606075,I606067);
not I_35472 (I606092,I453540);
nand I_35473 (I606109,I606092,I453531);
and I_35474 (I606126,I605928,I606109);
nor I_35475 (I606143,I606041,I606126);
DFFARX1 I_35476 (I606143,I3035,I605846,I605814,);
DFFARX1 I_35477 (I606126,I3035,I605846,I605835,);
nor I_35478 (I606188,I453540,I453549);
nor I_35479 (I605826,I606041,I606188);
or I_35480 (I606219,I453540,I453549);
nor I_35481 (I606236,I453534,I453534);
DFFARX1 I_35482 (I606236,I3035,I605846,I606262,);
not I_35483 (I606270,I606262);
nor I_35484 (I605832,I606270,I606075);
nand I_35485 (I606301,I606270,I605920);
not I_35486 (I606318,I453534);
nand I_35487 (I606335,I606318,I606024);
nand I_35488 (I606352,I606270,I606335);
nand I_35489 (I605823,I606352,I606301);
nand I_35490 (I605820,I606335,I606219);
not I_35491 (I606424,I3042);
DFFARX1 I_35492 (I304215,I3035,I606424,I606450,);
and I_35493 (I606458,I606450,I304203);
DFFARX1 I_35494 (I606458,I3035,I606424,I606407,);
DFFARX1 I_35495 (I304218,I3035,I606424,I606498,);
not I_35496 (I606506,I304209);
not I_35497 (I606523,I304200);
nand I_35498 (I606540,I606523,I606506);
nor I_35499 (I606395,I606498,I606540);
DFFARX1 I_35500 (I606540,I3035,I606424,I606580,);
not I_35501 (I606416,I606580);
not I_35502 (I606602,I304206);
nand I_35503 (I606619,I606523,I606602);
DFFARX1 I_35504 (I606619,I3035,I606424,I606645,);
not I_35505 (I606653,I606645);
not I_35506 (I606670,I304221);
nand I_35507 (I606687,I606670,I304224);
and I_35508 (I606704,I606506,I606687);
nor I_35509 (I606721,I606619,I606704);
DFFARX1 I_35510 (I606721,I3035,I606424,I606392,);
DFFARX1 I_35511 (I606704,I3035,I606424,I606413,);
nor I_35512 (I606766,I304221,I304200);
nor I_35513 (I606404,I606619,I606766);
or I_35514 (I606797,I304221,I304200);
nor I_35515 (I606814,I304212,I304203);
DFFARX1 I_35516 (I606814,I3035,I606424,I606840,);
not I_35517 (I606848,I606840);
nor I_35518 (I606410,I606848,I606653);
nand I_35519 (I606879,I606848,I606498);
not I_35520 (I606896,I304212);
nand I_35521 (I606913,I606896,I606602);
nand I_35522 (I606930,I606848,I606913);
nand I_35523 (I606401,I606930,I606879);
nand I_35524 (I606398,I606913,I606797);
not I_35525 (I607002,I3042);
DFFARX1 I_35526 (I440356,I3035,I607002,I607028,);
and I_35527 (I607036,I607028,I440362);
DFFARX1 I_35528 (I607036,I3035,I607002,I606985,);
DFFARX1 I_35529 (I440368,I3035,I607002,I607076,);
not I_35530 (I607084,I440353);
not I_35531 (I607101,I440353);
nand I_35532 (I607118,I607101,I607084);
nor I_35533 (I606973,I607076,I607118);
DFFARX1 I_35534 (I607118,I3035,I607002,I607158,);
not I_35535 (I606994,I607158);
not I_35536 (I607180,I440371);
nand I_35537 (I607197,I607101,I607180);
DFFARX1 I_35538 (I607197,I3035,I607002,I607223,);
not I_35539 (I607231,I607223);
not I_35540 (I607248,I440365);
nand I_35541 (I607265,I607248,I440356);
and I_35542 (I607282,I607084,I607265);
nor I_35543 (I607299,I607197,I607282);
DFFARX1 I_35544 (I607299,I3035,I607002,I606970,);
DFFARX1 I_35545 (I607282,I3035,I607002,I606991,);
nor I_35546 (I607344,I440365,I440374);
nor I_35547 (I606982,I607197,I607344);
or I_35548 (I607375,I440365,I440374);
nor I_35549 (I607392,I440359,I440359);
DFFARX1 I_35550 (I607392,I3035,I607002,I607418,);
not I_35551 (I607426,I607418);
nor I_35552 (I606988,I607426,I607231);
nand I_35553 (I607457,I607426,I607076);
not I_35554 (I607474,I440359);
nand I_35555 (I607491,I607474,I607180);
nand I_35556 (I607508,I607426,I607491);
nand I_35557 (I606979,I607508,I607457);
nand I_35558 (I606976,I607491,I607375);
not I_35559 (I607580,I3042);
DFFARX1 I_35560 (I656155,I3035,I607580,I607606,);
and I_35561 (I607614,I607606,I656149);
DFFARX1 I_35562 (I607614,I3035,I607580,I607563,);
DFFARX1 I_35563 (I656134,I3035,I607580,I607654,);
not I_35564 (I607662,I656140);
not I_35565 (I607679,I656152);
nand I_35566 (I607696,I607679,I607662);
nor I_35567 (I607551,I607654,I607696);
DFFARX1 I_35568 (I607696,I3035,I607580,I607736,);
not I_35569 (I607572,I607736);
not I_35570 (I607758,I656134);
nand I_35571 (I607775,I607679,I607758);
DFFARX1 I_35572 (I607775,I3035,I607580,I607801,);
not I_35573 (I607809,I607801);
not I_35574 (I607826,I656158);
nand I_35575 (I607843,I607826,I656146);
and I_35576 (I607860,I607662,I607843);
nor I_35577 (I607877,I607775,I607860);
DFFARX1 I_35578 (I607877,I3035,I607580,I607548,);
DFFARX1 I_35579 (I607860,I3035,I607580,I607569,);
nor I_35580 (I607922,I656158,I656137);
nor I_35581 (I607560,I607775,I607922);
or I_35582 (I607953,I656158,I656137);
nor I_35583 (I607970,I656143,I656137);
DFFARX1 I_35584 (I607970,I3035,I607580,I607996,);
not I_35585 (I608004,I607996);
nor I_35586 (I607566,I608004,I607809);
nand I_35587 (I608035,I608004,I607654);
not I_35588 (I608052,I656143);
nand I_35589 (I608069,I608052,I607758);
nand I_35590 (I608086,I608004,I608069);
nand I_35591 (I607557,I608086,I608035);
nand I_35592 (I607554,I608069,I607953);
not I_35593 (I608158,I3042);
DFFARX1 I_35594 (I355079,I3035,I608158,I608184,);
and I_35595 (I608192,I608184,I355067);
DFFARX1 I_35596 (I608192,I3035,I608158,I608141,);
DFFARX1 I_35597 (I355070,I3035,I608158,I608232,);
not I_35598 (I608240,I355064);
not I_35599 (I608257,I355088);
nand I_35600 (I608274,I608257,I608240);
nor I_35601 (I608129,I608232,I608274);
DFFARX1 I_35602 (I608274,I3035,I608158,I608314,);
not I_35603 (I608150,I608314);
not I_35604 (I608336,I355076);
nand I_35605 (I608353,I608257,I608336);
DFFARX1 I_35606 (I608353,I3035,I608158,I608379,);
not I_35607 (I608387,I608379);
not I_35608 (I608404,I355085);
nand I_35609 (I608421,I608404,I355082);
and I_35610 (I608438,I608240,I608421);
nor I_35611 (I608455,I608353,I608438);
DFFARX1 I_35612 (I608455,I3035,I608158,I608126,);
DFFARX1 I_35613 (I608438,I3035,I608158,I608147,);
nor I_35614 (I608500,I355085,I355073);
nor I_35615 (I608138,I608353,I608500);
or I_35616 (I608531,I355085,I355073);
nor I_35617 (I608548,I355064,I355067);
DFFARX1 I_35618 (I608548,I3035,I608158,I608574,);
not I_35619 (I608582,I608574);
nor I_35620 (I608144,I608582,I608387);
nand I_35621 (I608613,I608582,I608232);
not I_35622 (I608630,I355064);
nand I_35623 (I608647,I608630,I608336);
nand I_35624 (I608664,I608582,I608647);
nand I_35625 (I608135,I608664,I608613);
nand I_35626 (I608132,I608647,I608531);
not I_35627 (I608736,I3042);
DFFARX1 I_35628 (I164028,I3035,I608736,I608762,);
and I_35629 (I608770,I608762,I164013);
DFFARX1 I_35630 (I608770,I3035,I608736,I608719,);
DFFARX1 I_35631 (I164019,I3035,I608736,I608810,);
not I_35632 (I608818,I164001);
not I_35633 (I608835,I164022);
nand I_35634 (I608852,I608835,I608818);
nor I_35635 (I608707,I608810,I608852);
DFFARX1 I_35636 (I608852,I3035,I608736,I608892,);
not I_35637 (I608728,I608892);
not I_35638 (I608914,I164025);
nand I_35639 (I608931,I608835,I608914);
DFFARX1 I_35640 (I608931,I3035,I608736,I608957,);
not I_35641 (I608965,I608957);
not I_35642 (I608982,I164016);
nand I_35643 (I608999,I608982,I164004);
and I_35644 (I609016,I608818,I608999);
nor I_35645 (I609033,I608931,I609016);
DFFARX1 I_35646 (I609033,I3035,I608736,I608704,);
DFFARX1 I_35647 (I609016,I3035,I608736,I608725,);
nor I_35648 (I609078,I164016,I164010);
nor I_35649 (I608716,I608931,I609078);
or I_35650 (I609109,I164016,I164010);
nor I_35651 (I609126,I164007,I164001);
DFFARX1 I_35652 (I609126,I3035,I608736,I609152,);
not I_35653 (I609160,I609152);
nor I_35654 (I608722,I609160,I608965);
nand I_35655 (I609191,I609160,I608810);
not I_35656 (I609208,I164007);
nand I_35657 (I609225,I609208,I608914);
nand I_35658 (I609242,I609160,I609225);
nand I_35659 (I608713,I609242,I609191);
nand I_35660 (I608710,I609225,I609109);
not I_35661 (I609314,I3042);
DFFARX1 I_35662 (I23615,I3035,I609314,I609340,);
and I_35663 (I609348,I609340,I23618);
DFFARX1 I_35664 (I609348,I3035,I609314,I609297,);
DFFARX1 I_35665 (I23618,I3035,I609314,I609388,);
not I_35666 (I609396,I23621);
not I_35667 (I609413,I23636);
nand I_35668 (I609430,I609413,I609396);
nor I_35669 (I609285,I609388,I609430);
DFFARX1 I_35670 (I609430,I3035,I609314,I609470,);
not I_35671 (I609306,I609470);
not I_35672 (I609492,I23630);
nand I_35673 (I609509,I609413,I609492);
DFFARX1 I_35674 (I609509,I3035,I609314,I609535,);
not I_35675 (I609543,I609535);
not I_35676 (I609560,I23633);
nand I_35677 (I609577,I609560,I23615);
and I_35678 (I609594,I609396,I609577);
nor I_35679 (I609611,I609509,I609594);
DFFARX1 I_35680 (I609611,I3035,I609314,I609282,);
DFFARX1 I_35681 (I609594,I3035,I609314,I609303,);
nor I_35682 (I609656,I23633,I23627);
nor I_35683 (I609294,I609509,I609656);
or I_35684 (I609687,I23633,I23627);
nor I_35685 (I609704,I23624,I23639);
DFFARX1 I_35686 (I609704,I3035,I609314,I609730,);
not I_35687 (I609738,I609730);
nor I_35688 (I609300,I609738,I609543);
nand I_35689 (I609769,I609738,I609388);
not I_35690 (I609786,I23624);
nand I_35691 (I609803,I609786,I609492);
nand I_35692 (I609820,I609738,I609803);
nand I_35693 (I609291,I609820,I609769);
nand I_35694 (I609288,I609803,I609687);
not I_35695 (I609892,I3042);
DFFARX1 I_35696 (I664859,I3035,I609892,I609918,);
and I_35697 (I609926,I609918,I664853);
DFFARX1 I_35698 (I609926,I3035,I609892,I609875,);
DFFARX1 I_35699 (I664838,I3035,I609892,I609966,);
not I_35700 (I609974,I664844);
not I_35701 (I609991,I664856);
nand I_35702 (I610008,I609991,I609974);
nor I_35703 (I609863,I609966,I610008);
DFFARX1 I_35704 (I610008,I3035,I609892,I610048,);
not I_35705 (I609884,I610048);
not I_35706 (I610070,I664838);
nand I_35707 (I610087,I609991,I610070);
DFFARX1 I_35708 (I610087,I3035,I609892,I610113,);
not I_35709 (I610121,I610113);
not I_35710 (I610138,I664862);
nand I_35711 (I610155,I610138,I664850);
and I_35712 (I610172,I609974,I610155);
nor I_35713 (I610189,I610087,I610172);
DFFARX1 I_35714 (I610189,I3035,I609892,I609860,);
DFFARX1 I_35715 (I610172,I3035,I609892,I609881,);
nor I_35716 (I610234,I664862,I664841);
nor I_35717 (I609872,I610087,I610234);
or I_35718 (I610265,I664862,I664841);
nor I_35719 (I610282,I664847,I664841);
DFFARX1 I_35720 (I610282,I3035,I609892,I610308,);
not I_35721 (I610316,I610308);
nor I_35722 (I609878,I610316,I610121);
nand I_35723 (I610347,I610316,I609966);
not I_35724 (I610364,I664847);
nand I_35725 (I610381,I610364,I610070);
nand I_35726 (I610398,I610316,I610381);
nand I_35727 (I609869,I610398,I610347);
nand I_35728 (I609866,I610381,I610265);
not I_35729 (I610470,I3042);
DFFARX1 I_35730 (I70015,I3035,I610470,I610496,);
and I_35731 (I610504,I610496,I69991);
DFFARX1 I_35732 (I610504,I3035,I610470,I610453,);
DFFARX1 I_35733 (I70009,I3035,I610470,I610544,);
not I_35734 (I610552,I69997);
not I_35735 (I610569,I69994);
nand I_35736 (I610586,I610569,I610552);
nor I_35737 (I610441,I610544,I610586);
DFFARX1 I_35738 (I610586,I3035,I610470,I610626,);
not I_35739 (I610462,I610626);
not I_35740 (I610648,I70003);
nand I_35741 (I610665,I610569,I610648);
DFFARX1 I_35742 (I610665,I3035,I610470,I610691,);
not I_35743 (I610699,I610691);
not I_35744 (I610716,I69994);
nand I_35745 (I610733,I610716,I70012);
and I_35746 (I610750,I610552,I610733);
nor I_35747 (I610767,I610665,I610750);
DFFARX1 I_35748 (I610767,I3035,I610470,I610438,);
DFFARX1 I_35749 (I610750,I3035,I610470,I610459,);
nor I_35750 (I610812,I69994,I70006);
nor I_35751 (I610450,I610665,I610812);
or I_35752 (I610843,I69994,I70006);
nor I_35753 (I610860,I70000,I69991);
DFFARX1 I_35754 (I610860,I3035,I610470,I610886,);
not I_35755 (I610894,I610886);
nor I_35756 (I610456,I610894,I610699);
nand I_35757 (I610925,I610894,I610544);
not I_35758 (I610942,I70000);
nand I_35759 (I610959,I610942,I610648);
nand I_35760 (I610976,I610894,I610959);
nand I_35761 (I610447,I610976,I610925);
nand I_35762 (I610444,I610959,I610843);
not I_35763 (I611048,I3042);
DFFARX1 I_35764 (I403053,I3035,I611048,I611074,);
and I_35765 (I611082,I611074,I403041);
DFFARX1 I_35766 (I611082,I3035,I611048,I611031,);
DFFARX1 I_35767 (I403044,I3035,I611048,I611122,);
not I_35768 (I611130,I403038);
not I_35769 (I611147,I403062);
nand I_35770 (I611164,I611147,I611130);
nor I_35771 (I611019,I611122,I611164);
DFFARX1 I_35772 (I611164,I3035,I611048,I611204,);
not I_35773 (I611040,I611204);
not I_35774 (I611226,I403050);
nand I_35775 (I611243,I611147,I611226);
DFFARX1 I_35776 (I611243,I3035,I611048,I611269,);
not I_35777 (I611277,I611269);
not I_35778 (I611294,I403059);
nand I_35779 (I611311,I611294,I403056);
and I_35780 (I611328,I611130,I611311);
nor I_35781 (I611345,I611243,I611328);
DFFARX1 I_35782 (I611345,I3035,I611048,I611016,);
DFFARX1 I_35783 (I611328,I3035,I611048,I611037,);
nor I_35784 (I611390,I403059,I403047);
nor I_35785 (I611028,I611243,I611390);
or I_35786 (I611421,I403059,I403047);
nor I_35787 (I611438,I403038,I403041);
DFFARX1 I_35788 (I611438,I3035,I611048,I611464,);
not I_35789 (I611472,I611464);
nor I_35790 (I611034,I611472,I611277);
nand I_35791 (I611503,I611472,I611122);
not I_35792 (I611520,I403038);
nand I_35793 (I611537,I611520,I611226);
nand I_35794 (I611554,I611472,I611537);
nand I_35795 (I611025,I611554,I611503);
nand I_35796 (I611022,I611537,I611421);
not I_35797 (I611626,I3042);
DFFARX1 I_35798 (I195121,I3035,I611626,I611652,);
and I_35799 (I611660,I611652,I195106);
DFFARX1 I_35800 (I611660,I3035,I611626,I611609,);
DFFARX1 I_35801 (I195112,I3035,I611626,I611700,);
not I_35802 (I611708,I195094);
not I_35803 (I611725,I195115);
nand I_35804 (I611742,I611725,I611708);
nor I_35805 (I611597,I611700,I611742);
DFFARX1 I_35806 (I611742,I3035,I611626,I611782,);
not I_35807 (I611618,I611782);
not I_35808 (I611804,I195118);
nand I_35809 (I611821,I611725,I611804);
DFFARX1 I_35810 (I611821,I3035,I611626,I611847,);
not I_35811 (I611855,I611847);
not I_35812 (I611872,I195109);
nand I_35813 (I611889,I611872,I195097);
and I_35814 (I611906,I611708,I611889);
nor I_35815 (I611923,I611821,I611906);
DFFARX1 I_35816 (I611923,I3035,I611626,I611594,);
DFFARX1 I_35817 (I611906,I3035,I611626,I611615,);
nor I_35818 (I611968,I195109,I195103);
nor I_35819 (I611606,I611821,I611968);
or I_35820 (I611999,I195109,I195103);
nor I_35821 (I612016,I195100,I195094);
DFFARX1 I_35822 (I612016,I3035,I611626,I612042,);
not I_35823 (I612050,I612042);
nor I_35824 (I611612,I612050,I611855);
nand I_35825 (I612081,I612050,I611700);
not I_35826 (I612098,I195100);
nand I_35827 (I612115,I612098,I611804);
nand I_35828 (I612132,I612050,I612115);
nand I_35829 (I611603,I612132,I612081);
nand I_35830 (I611600,I612115,I611999);
not I_35831 (I612204,I3042);
DFFARX1 I_35832 (I733545,I3035,I612204,I612230,);
and I_35833 (I612238,I612230,I733527);
DFFARX1 I_35834 (I612238,I3035,I612204,I612187,);
DFFARX1 I_35835 (I733518,I3035,I612204,I612278,);
not I_35836 (I612286,I733533);
not I_35837 (I612303,I733521);
nand I_35838 (I612320,I612303,I612286);
nor I_35839 (I612175,I612278,I612320);
DFFARX1 I_35840 (I612320,I3035,I612204,I612360,);
not I_35841 (I612196,I612360);
not I_35842 (I612382,I733530);
nand I_35843 (I612399,I612303,I612382);
DFFARX1 I_35844 (I612399,I3035,I612204,I612425,);
not I_35845 (I612433,I612425);
not I_35846 (I612450,I733539);
nand I_35847 (I612467,I612450,I733518);
and I_35848 (I612484,I612286,I612467);
nor I_35849 (I612501,I612399,I612484);
DFFARX1 I_35850 (I612501,I3035,I612204,I612172,);
DFFARX1 I_35851 (I612484,I3035,I612204,I612193,);
nor I_35852 (I612546,I733539,I733542);
nor I_35853 (I612184,I612399,I612546);
or I_35854 (I612577,I733539,I733542);
nor I_35855 (I612594,I733536,I733524);
DFFARX1 I_35856 (I612594,I3035,I612204,I612620,);
not I_35857 (I612628,I612620);
nor I_35858 (I612190,I612628,I612433);
nand I_35859 (I612659,I612628,I612278);
not I_35860 (I612676,I733536);
nand I_35861 (I612693,I612676,I612382);
nand I_35862 (I612710,I612628,I612693);
nand I_35863 (I612181,I612710,I612659);
nand I_35864 (I612178,I612693,I612577);
not I_35865 (I612782,I3042);
DFFARX1 I_35866 (I63164,I3035,I612782,I612808,);
and I_35867 (I612816,I612808,I63140);
DFFARX1 I_35868 (I612816,I3035,I612782,I612765,);
DFFARX1 I_35869 (I63158,I3035,I612782,I612856,);
not I_35870 (I612864,I63146);
not I_35871 (I612881,I63143);
nand I_35872 (I612898,I612881,I612864);
nor I_35873 (I612753,I612856,I612898);
DFFARX1 I_35874 (I612898,I3035,I612782,I612938,);
not I_35875 (I612774,I612938);
not I_35876 (I612960,I63152);
nand I_35877 (I612977,I612881,I612960);
DFFARX1 I_35878 (I612977,I3035,I612782,I613003,);
not I_35879 (I613011,I613003);
not I_35880 (I613028,I63143);
nand I_35881 (I613045,I613028,I63161);
and I_35882 (I613062,I612864,I613045);
nor I_35883 (I613079,I612977,I613062);
DFFARX1 I_35884 (I613079,I3035,I612782,I612750,);
DFFARX1 I_35885 (I613062,I3035,I612782,I612771,);
nor I_35886 (I613124,I63143,I63155);
nor I_35887 (I612762,I612977,I613124);
or I_35888 (I613155,I63143,I63155);
nor I_35889 (I613172,I63149,I63140);
DFFARX1 I_35890 (I613172,I3035,I612782,I613198,);
not I_35891 (I613206,I613198);
nor I_35892 (I612768,I613206,I613011);
nand I_35893 (I613237,I613206,I612856);
not I_35894 (I613254,I63149);
nand I_35895 (I613271,I613254,I612960);
nand I_35896 (I613288,I613206,I613271);
nand I_35897 (I612759,I613288,I613237);
nand I_35898 (I612756,I613271,I613155);
not I_35899 (I613360,I3042);
DFFARX1 I_35900 (I475665,I3035,I613360,I613386,);
and I_35901 (I613394,I613386,I475671);
DFFARX1 I_35902 (I613394,I3035,I613360,I613343,);
DFFARX1 I_35903 (I475677,I3035,I613360,I613434,);
not I_35904 (I613442,I475662);
not I_35905 (I613459,I475662);
nand I_35906 (I613476,I613459,I613442);
nor I_35907 (I613331,I613434,I613476);
DFFARX1 I_35908 (I613476,I3035,I613360,I613516,);
not I_35909 (I613352,I613516);
not I_35910 (I613538,I475680);
nand I_35911 (I613555,I613459,I613538);
DFFARX1 I_35912 (I613555,I3035,I613360,I613581,);
not I_35913 (I613589,I613581);
not I_35914 (I613606,I475674);
nand I_35915 (I613623,I613606,I475665);
and I_35916 (I613640,I613442,I613623);
nor I_35917 (I613657,I613555,I613640);
DFFARX1 I_35918 (I613657,I3035,I613360,I613328,);
DFFARX1 I_35919 (I613640,I3035,I613360,I613349,);
nor I_35920 (I613702,I475674,I475683);
nor I_35921 (I613340,I613555,I613702);
or I_35922 (I613733,I475674,I475683);
nor I_35923 (I613750,I475668,I475668);
DFFARX1 I_35924 (I613750,I3035,I613360,I613776,);
not I_35925 (I613784,I613776);
nor I_35926 (I613346,I613784,I613589);
nand I_35927 (I613815,I613784,I613434);
not I_35928 (I613832,I475668);
nand I_35929 (I613849,I613832,I613538);
nand I_35930 (I613866,I613784,I613849);
nand I_35931 (I613337,I613866,I613815);
nand I_35932 (I613334,I613849,I613733);
not I_35933 (I613938,I3042);
DFFARX1 I_35934 (I18345,I3035,I613938,I613964,);
and I_35935 (I613972,I613964,I18348);
DFFARX1 I_35936 (I613972,I3035,I613938,I613921,);
DFFARX1 I_35937 (I18348,I3035,I613938,I614012,);
not I_35938 (I614020,I18351);
not I_35939 (I614037,I18366);
nand I_35940 (I614054,I614037,I614020);
nor I_35941 (I613909,I614012,I614054);
DFFARX1 I_35942 (I614054,I3035,I613938,I614094,);
not I_35943 (I613930,I614094);
not I_35944 (I614116,I18360);
nand I_35945 (I614133,I614037,I614116);
DFFARX1 I_35946 (I614133,I3035,I613938,I614159,);
not I_35947 (I614167,I614159);
not I_35948 (I614184,I18363);
nand I_35949 (I614201,I614184,I18345);
and I_35950 (I614218,I614020,I614201);
nor I_35951 (I614235,I614133,I614218);
DFFARX1 I_35952 (I614235,I3035,I613938,I613906,);
DFFARX1 I_35953 (I614218,I3035,I613938,I613927,);
nor I_35954 (I614280,I18363,I18357);
nor I_35955 (I613918,I614133,I614280);
or I_35956 (I614311,I18363,I18357);
nor I_35957 (I614328,I18354,I18369);
DFFARX1 I_35958 (I614328,I3035,I613938,I614354,);
not I_35959 (I614362,I614354);
nor I_35960 (I613924,I614362,I614167);
nand I_35961 (I614393,I614362,I614012);
not I_35962 (I614410,I18354);
nand I_35963 (I614427,I614410,I614116);
nand I_35964 (I614444,I614362,I614427);
nand I_35965 (I613915,I614444,I614393);
nand I_35966 (I613912,I614427,I614311);
not I_35967 (I614516,I3042);
DFFARX1 I_35968 (I56840,I3035,I614516,I614542,);
and I_35969 (I614550,I614542,I56816);
DFFARX1 I_35970 (I614550,I3035,I614516,I614499,);
DFFARX1 I_35971 (I56834,I3035,I614516,I614590,);
not I_35972 (I614598,I56822);
not I_35973 (I614615,I56819);
nand I_35974 (I614632,I614615,I614598);
nor I_35975 (I614487,I614590,I614632);
DFFARX1 I_35976 (I614632,I3035,I614516,I614672,);
not I_35977 (I614508,I614672);
not I_35978 (I614694,I56828);
nand I_35979 (I614711,I614615,I614694);
DFFARX1 I_35980 (I614711,I3035,I614516,I614737,);
not I_35981 (I614745,I614737);
not I_35982 (I614762,I56819);
nand I_35983 (I614779,I614762,I56837);
and I_35984 (I614796,I614598,I614779);
nor I_35985 (I614813,I614711,I614796);
DFFARX1 I_35986 (I614813,I3035,I614516,I614484,);
DFFARX1 I_35987 (I614796,I3035,I614516,I614505,);
nor I_35988 (I614858,I56819,I56831);
nor I_35989 (I614496,I614711,I614858);
or I_35990 (I614889,I56819,I56831);
nor I_35991 (I614906,I56825,I56816);
DFFARX1 I_35992 (I614906,I3035,I614516,I614932,);
not I_35993 (I614940,I614932);
nor I_35994 (I614502,I614940,I614745);
nand I_35995 (I614971,I614940,I614590);
not I_35996 (I614988,I56825);
nand I_35997 (I615005,I614988,I614694);
nand I_35998 (I615022,I614940,I615005);
nand I_35999 (I614493,I615022,I614971);
nand I_36000 (I614490,I615005,I614889);
not I_36001 (I615094,I3042);
DFFARX1 I_36002 (I512898,I3035,I615094,I615120,);
and I_36003 (I615128,I615120,I512892);
DFFARX1 I_36004 (I615128,I3035,I615094,I615077,);
DFFARX1 I_36005 (I512910,I3035,I615094,I615168,);
not I_36006 (I615176,I512901);
not I_36007 (I615193,I512913);
nand I_36008 (I615210,I615193,I615176);
nor I_36009 (I615065,I615168,I615210);
DFFARX1 I_36010 (I615210,I3035,I615094,I615250,);
not I_36011 (I615086,I615250);
not I_36012 (I615272,I512919);
nand I_36013 (I615289,I615193,I615272);
DFFARX1 I_36014 (I615289,I3035,I615094,I615315,);
not I_36015 (I615323,I615315);
not I_36016 (I615340,I512895);
nand I_36017 (I615357,I615340,I512916);
and I_36018 (I615374,I615176,I615357);
nor I_36019 (I615391,I615289,I615374);
DFFARX1 I_36020 (I615391,I3035,I615094,I615062,);
DFFARX1 I_36021 (I615374,I3035,I615094,I615083,);
nor I_36022 (I615436,I512895,I512907);
nor I_36023 (I615074,I615289,I615436);
or I_36024 (I615467,I512895,I512907);
nor I_36025 (I615484,I512892,I512904);
DFFARX1 I_36026 (I615484,I3035,I615094,I615510,);
not I_36027 (I615518,I615510);
nor I_36028 (I615080,I615518,I615323);
nand I_36029 (I615549,I615518,I615168);
not I_36030 (I615566,I512892);
nand I_36031 (I615583,I615566,I615272);
nand I_36032 (I615600,I615518,I615583);
nand I_36033 (I615071,I615600,I615549);
nand I_36034 (I615068,I615583,I615467);
not I_36035 (I615672,I3042);
DFFARX1 I_36036 (I528402,I3035,I615672,I615698,);
and I_36037 (I615706,I615698,I528396);
DFFARX1 I_36038 (I615706,I3035,I615672,I615655,);
DFFARX1 I_36039 (I528414,I3035,I615672,I615746,);
not I_36040 (I615754,I528405);
not I_36041 (I615771,I528417);
nand I_36042 (I615788,I615771,I615754);
nor I_36043 (I615643,I615746,I615788);
DFFARX1 I_36044 (I615788,I3035,I615672,I615828,);
not I_36045 (I615664,I615828);
not I_36046 (I615850,I528423);
nand I_36047 (I615867,I615771,I615850);
DFFARX1 I_36048 (I615867,I3035,I615672,I615893,);
not I_36049 (I615901,I615893);
not I_36050 (I615918,I528399);
nand I_36051 (I615935,I615918,I528420);
and I_36052 (I615952,I615754,I615935);
nor I_36053 (I615969,I615867,I615952);
DFFARX1 I_36054 (I615969,I3035,I615672,I615640,);
DFFARX1 I_36055 (I615952,I3035,I615672,I615661,);
nor I_36056 (I616014,I528399,I528411);
nor I_36057 (I615652,I615867,I616014);
or I_36058 (I616045,I528399,I528411);
nor I_36059 (I616062,I528396,I528408);
DFFARX1 I_36060 (I616062,I3035,I615672,I616088,);
not I_36061 (I616096,I616088);
nor I_36062 (I615658,I616096,I615901);
nand I_36063 (I616127,I616096,I615746);
not I_36064 (I616144,I528396);
nand I_36065 (I616161,I616144,I615850);
nand I_36066 (I616178,I616096,I616161);
nand I_36067 (I615649,I616178,I616127);
nand I_36068 (I615646,I616161,I616045);
not I_36069 (I616250,I3042);
DFFARX1 I_36070 (I394961,I3035,I616250,I616276,);
and I_36071 (I616284,I616276,I394949);
DFFARX1 I_36072 (I616284,I3035,I616250,I616233,);
DFFARX1 I_36073 (I394952,I3035,I616250,I616324,);
not I_36074 (I616332,I394946);
not I_36075 (I616349,I394970);
nand I_36076 (I616366,I616349,I616332);
nor I_36077 (I616221,I616324,I616366);
DFFARX1 I_36078 (I616366,I3035,I616250,I616406,);
not I_36079 (I616242,I616406);
not I_36080 (I616428,I394958);
nand I_36081 (I616445,I616349,I616428);
DFFARX1 I_36082 (I616445,I3035,I616250,I616471,);
not I_36083 (I616479,I616471);
not I_36084 (I616496,I394967);
nand I_36085 (I616513,I616496,I394964);
and I_36086 (I616530,I616332,I616513);
nor I_36087 (I616547,I616445,I616530);
DFFARX1 I_36088 (I616547,I3035,I616250,I616218,);
DFFARX1 I_36089 (I616530,I3035,I616250,I616239,);
nor I_36090 (I616592,I394967,I394955);
nor I_36091 (I616230,I616445,I616592);
or I_36092 (I616623,I394967,I394955);
nor I_36093 (I616640,I394946,I394949);
DFFARX1 I_36094 (I616640,I3035,I616250,I616666,);
not I_36095 (I616674,I616666);
nor I_36096 (I616236,I616674,I616479);
nand I_36097 (I616705,I616674,I616324);
not I_36098 (I616722,I394946);
nand I_36099 (I616739,I616722,I616428);
nand I_36100 (I616756,I616674,I616739);
nand I_36101 (I616227,I616756,I616705);
nand I_36102 (I616224,I616739,I616623);
not I_36103 (I616828,I3042);
DFFARX1 I_36104 (I275045,I3035,I616828,I616854,);
and I_36105 (I616862,I616854,I275060);
DFFARX1 I_36106 (I616862,I3035,I616828,I616811,);
DFFARX1 I_36107 (I275063,I3035,I616828,I616902,);
not I_36108 (I616910,I275057);
not I_36109 (I616927,I275072);
nand I_36110 (I616944,I616927,I616910);
nor I_36111 (I616799,I616902,I616944);
DFFARX1 I_36112 (I616944,I3035,I616828,I616984,);
not I_36113 (I616820,I616984);
not I_36114 (I617006,I275048);
nand I_36115 (I617023,I616927,I617006);
DFFARX1 I_36116 (I617023,I3035,I616828,I617049,);
not I_36117 (I617057,I617049);
not I_36118 (I617074,I275051);
nand I_36119 (I617091,I617074,I275045);
and I_36120 (I617108,I616910,I617091);
nor I_36121 (I617125,I617023,I617108);
DFFARX1 I_36122 (I617125,I3035,I616828,I616796,);
DFFARX1 I_36123 (I617108,I3035,I616828,I616817,);
nor I_36124 (I617170,I275051,I275054);
nor I_36125 (I616808,I617023,I617170);
or I_36126 (I617201,I275051,I275054);
nor I_36127 (I617218,I275069,I275066);
DFFARX1 I_36128 (I617218,I3035,I616828,I617244,);
not I_36129 (I617252,I617244);
nor I_36130 (I616814,I617252,I617057);
nand I_36131 (I617283,I617252,I616902);
not I_36132 (I617300,I275069);
nand I_36133 (I617317,I617300,I617006);
nand I_36134 (I617334,I617252,I617317);
nand I_36135 (I616805,I617334,I617283);
nand I_36136 (I616802,I617317,I617201);
not I_36137 (I617406,I3042);
DFFARX1 I_36138 (I707960,I3035,I617406,I617432,);
and I_36139 (I617440,I617432,I707942);
DFFARX1 I_36140 (I617440,I3035,I617406,I617389,);
DFFARX1 I_36141 (I707933,I3035,I617406,I617480,);
not I_36142 (I617488,I707948);
not I_36143 (I617505,I707936);
nand I_36144 (I617522,I617505,I617488);
nor I_36145 (I617377,I617480,I617522);
DFFARX1 I_36146 (I617522,I3035,I617406,I617562,);
not I_36147 (I617398,I617562);
not I_36148 (I617584,I707945);
nand I_36149 (I617601,I617505,I617584);
DFFARX1 I_36150 (I617601,I3035,I617406,I617627,);
not I_36151 (I617635,I617627);
not I_36152 (I617652,I707954);
nand I_36153 (I617669,I617652,I707933);
and I_36154 (I617686,I617488,I617669);
nor I_36155 (I617703,I617601,I617686);
DFFARX1 I_36156 (I617703,I3035,I617406,I617374,);
DFFARX1 I_36157 (I617686,I3035,I617406,I617395,);
nor I_36158 (I617748,I707954,I707957);
nor I_36159 (I617386,I617601,I617748);
or I_36160 (I617779,I707954,I707957);
nor I_36161 (I617796,I707951,I707939);
DFFARX1 I_36162 (I617796,I3035,I617406,I617822,);
not I_36163 (I617830,I617822);
nor I_36164 (I617392,I617830,I617635);
nand I_36165 (I617861,I617830,I617480);
not I_36166 (I617878,I707951);
nand I_36167 (I617895,I617878,I617584);
nand I_36168 (I617912,I617830,I617895);
nand I_36169 (I617383,I617912,I617861);
nand I_36170 (I617380,I617895,I617779);
not I_36171 (I617984,I3042);
DFFARX1 I_36172 (I495456,I3035,I617984,I618010,);
and I_36173 (I618018,I618010,I495450);
DFFARX1 I_36174 (I618018,I3035,I617984,I617967,);
DFFARX1 I_36175 (I495468,I3035,I617984,I618058,);
not I_36176 (I618066,I495459);
not I_36177 (I618083,I495471);
nand I_36178 (I618100,I618083,I618066);
nor I_36179 (I617955,I618058,I618100);
DFFARX1 I_36180 (I618100,I3035,I617984,I618140,);
not I_36181 (I617976,I618140);
not I_36182 (I618162,I495477);
nand I_36183 (I618179,I618083,I618162);
DFFARX1 I_36184 (I618179,I3035,I617984,I618205,);
not I_36185 (I618213,I618205);
not I_36186 (I618230,I495453);
nand I_36187 (I618247,I618230,I495474);
and I_36188 (I618264,I618066,I618247);
nor I_36189 (I618281,I618179,I618264);
DFFARX1 I_36190 (I618281,I3035,I617984,I617952,);
DFFARX1 I_36191 (I618264,I3035,I617984,I617973,);
nor I_36192 (I618326,I495453,I495465);
nor I_36193 (I617964,I618179,I618326);
or I_36194 (I618357,I495453,I495465);
nor I_36195 (I618374,I495450,I495462);
DFFARX1 I_36196 (I618374,I3035,I617984,I618400,);
not I_36197 (I618408,I618400);
nor I_36198 (I617970,I618408,I618213);
nand I_36199 (I618439,I618408,I618058);
not I_36200 (I618456,I495450);
nand I_36201 (I618473,I618456,I618162);
nand I_36202 (I618490,I618408,I618473);
nand I_36203 (I617961,I618490,I618439);
nand I_36204 (I617958,I618473,I618357);
not I_36205 (I618562,I3042);
DFFARX1 I_36206 (I259813,I3035,I618562,I618588,);
and I_36207 (I618596,I618588,I259828);
DFFARX1 I_36208 (I618596,I3035,I618562,I618545,);
DFFARX1 I_36209 (I259831,I3035,I618562,I618636,);
not I_36210 (I618644,I259825);
not I_36211 (I618661,I259840);
nand I_36212 (I618678,I618661,I618644);
nor I_36213 (I618533,I618636,I618678);
DFFARX1 I_36214 (I618678,I3035,I618562,I618718,);
not I_36215 (I618554,I618718);
not I_36216 (I618740,I259816);
nand I_36217 (I618757,I618661,I618740);
DFFARX1 I_36218 (I618757,I3035,I618562,I618783,);
not I_36219 (I618791,I618783);
not I_36220 (I618808,I259819);
nand I_36221 (I618825,I618808,I259813);
and I_36222 (I618842,I618644,I618825);
nor I_36223 (I618859,I618757,I618842);
DFFARX1 I_36224 (I618859,I3035,I618562,I618530,);
DFFARX1 I_36225 (I618842,I3035,I618562,I618551,);
nor I_36226 (I618904,I259819,I259822);
nor I_36227 (I618542,I618757,I618904);
or I_36228 (I618935,I259819,I259822);
nor I_36229 (I618952,I259837,I259834);
DFFARX1 I_36230 (I618952,I3035,I618562,I618978,);
not I_36231 (I618986,I618978);
nor I_36232 (I618548,I618986,I618791);
nand I_36233 (I619017,I618986,I618636);
not I_36234 (I619034,I259837);
nand I_36235 (I619051,I619034,I618740);
nand I_36236 (I619068,I618986,I619051);
nand I_36237 (I618539,I619068,I619017);
nand I_36238 (I618536,I619051,I618935);
not I_36239 (I619140,I3042);
DFFARX1 I_36240 (I360281,I3035,I619140,I619166,);
and I_36241 (I619174,I619166,I360269);
DFFARX1 I_36242 (I619174,I3035,I619140,I619123,);
DFFARX1 I_36243 (I360272,I3035,I619140,I619214,);
not I_36244 (I619222,I360266);
not I_36245 (I619239,I360290);
nand I_36246 (I619256,I619239,I619222);
nor I_36247 (I619111,I619214,I619256);
DFFARX1 I_36248 (I619256,I3035,I619140,I619296,);
not I_36249 (I619132,I619296);
not I_36250 (I619318,I360278);
nand I_36251 (I619335,I619239,I619318);
DFFARX1 I_36252 (I619335,I3035,I619140,I619361,);
not I_36253 (I619369,I619361);
not I_36254 (I619386,I360287);
nand I_36255 (I619403,I619386,I360284);
and I_36256 (I619420,I619222,I619403);
nor I_36257 (I619437,I619335,I619420);
DFFARX1 I_36258 (I619437,I3035,I619140,I619108,);
DFFARX1 I_36259 (I619420,I3035,I619140,I619129,);
nor I_36260 (I619482,I360287,I360275);
nor I_36261 (I619120,I619335,I619482);
or I_36262 (I619513,I360287,I360275);
nor I_36263 (I619530,I360266,I360269);
DFFARX1 I_36264 (I619530,I3035,I619140,I619556,);
not I_36265 (I619564,I619556);
nor I_36266 (I619126,I619564,I619369);
nand I_36267 (I619595,I619564,I619214);
not I_36268 (I619612,I360266);
nand I_36269 (I619629,I619612,I619318);
nand I_36270 (I619646,I619564,I619629);
nand I_36271 (I619117,I619646,I619595);
nand I_36272 (I619114,I619629,I619513);
not I_36273 (I619718,I3042);
DFFARX1 I_36274 (I682338,I3035,I619718,I619744,);
and I_36275 (I619752,I619744,I682320);
DFFARX1 I_36276 (I619752,I3035,I619718,I619701,);
DFFARX1 I_36277 (I682329,I3035,I619718,I619792,);
not I_36278 (I619800,I682314);
not I_36279 (I619817,I682326);
nand I_36280 (I619834,I619817,I619800);
nor I_36281 (I619689,I619792,I619834);
DFFARX1 I_36282 (I619834,I3035,I619718,I619874,);
not I_36283 (I619710,I619874);
not I_36284 (I619896,I682317);
nand I_36285 (I619913,I619817,I619896);
DFFARX1 I_36286 (I619913,I3035,I619718,I619939,);
not I_36287 (I619947,I619939);
not I_36288 (I619964,I682314);
nand I_36289 (I619981,I619964,I682317);
and I_36290 (I619998,I619800,I619981);
nor I_36291 (I620015,I619913,I619998);
DFFARX1 I_36292 (I620015,I3035,I619718,I619686,);
DFFARX1 I_36293 (I619998,I3035,I619718,I619707,);
nor I_36294 (I620060,I682314,I682335);
nor I_36295 (I619698,I619913,I620060);
or I_36296 (I620091,I682314,I682335);
nor I_36297 (I620108,I682323,I682332);
DFFARX1 I_36298 (I620108,I3035,I619718,I620134,);
not I_36299 (I620142,I620134);
nor I_36300 (I619704,I620142,I619947);
nand I_36301 (I620173,I620142,I619792);
not I_36302 (I620190,I682323);
nand I_36303 (I620207,I620190,I619896);
nand I_36304 (I620224,I620142,I620207);
nand I_36305 (I619695,I620224,I620173);
nand I_36306 (I619692,I620207,I620091);
not I_36307 (I620296,I3042);
DFFARX1 I_36308 (I450369,I3035,I620296,I620322,);
and I_36309 (I620330,I620322,I450375);
DFFARX1 I_36310 (I620330,I3035,I620296,I620279,);
DFFARX1 I_36311 (I450381,I3035,I620296,I620370,);
not I_36312 (I620378,I450366);
not I_36313 (I620395,I450366);
nand I_36314 (I620412,I620395,I620378);
nor I_36315 (I620267,I620370,I620412);
DFFARX1 I_36316 (I620412,I3035,I620296,I620452,);
not I_36317 (I620288,I620452);
not I_36318 (I620474,I450384);
nand I_36319 (I620491,I620395,I620474);
DFFARX1 I_36320 (I620491,I3035,I620296,I620517,);
not I_36321 (I620525,I620517);
not I_36322 (I620542,I450378);
nand I_36323 (I620559,I620542,I450369);
and I_36324 (I620576,I620378,I620559);
nor I_36325 (I620593,I620491,I620576);
DFFARX1 I_36326 (I620593,I3035,I620296,I620264,);
DFFARX1 I_36327 (I620576,I3035,I620296,I620285,);
nor I_36328 (I620638,I450378,I450387);
nor I_36329 (I620276,I620491,I620638);
or I_36330 (I620669,I450378,I450387);
nor I_36331 (I620686,I450372,I450372);
DFFARX1 I_36332 (I620686,I3035,I620296,I620712,);
not I_36333 (I620720,I620712);
nor I_36334 (I620282,I620720,I620525);
nand I_36335 (I620751,I620720,I620370);
not I_36336 (I620768,I450372);
nand I_36337 (I620785,I620768,I620474);
nand I_36338 (I620802,I620720,I620785);
nand I_36339 (I620273,I620802,I620751);
nand I_36340 (I620270,I620785,I620669);
not I_36341 (I620874,I3042);
DFFARX1 I_36342 (I708555,I3035,I620874,I620900,);
and I_36343 (I620908,I620900,I708537);
DFFARX1 I_36344 (I620908,I3035,I620874,I620857,);
DFFARX1 I_36345 (I708528,I3035,I620874,I620948,);
not I_36346 (I620956,I708543);
not I_36347 (I620973,I708531);
nand I_36348 (I620990,I620973,I620956);
nor I_36349 (I620845,I620948,I620990);
DFFARX1 I_36350 (I620990,I3035,I620874,I621030,);
not I_36351 (I620866,I621030);
not I_36352 (I621052,I708540);
nand I_36353 (I621069,I620973,I621052);
DFFARX1 I_36354 (I621069,I3035,I620874,I621095,);
not I_36355 (I621103,I621095);
not I_36356 (I621120,I708549);
nand I_36357 (I621137,I621120,I708528);
and I_36358 (I621154,I620956,I621137);
nor I_36359 (I621171,I621069,I621154);
DFFARX1 I_36360 (I621171,I3035,I620874,I620842,);
DFFARX1 I_36361 (I621154,I3035,I620874,I620863,);
nor I_36362 (I621216,I708549,I708552);
nor I_36363 (I620854,I621069,I621216);
or I_36364 (I621247,I708549,I708552);
nor I_36365 (I621264,I708546,I708534);
DFFARX1 I_36366 (I621264,I3035,I620874,I621290,);
not I_36367 (I621298,I621290);
nor I_36368 (I620860,I621298,I621103);
nand I_36369 (I621329,I621298,I620948);
not I_36370 (I621346,I708546);
nand I_36371 (I621363,I621346,I621052);
nand I_36372 (I621380,I621298,I621363);
nand I_36373 (I620851,I621380,I621329);
nand I_36374 (I620848,I621363,I621247);
not I_36375 (I621452,I3042);
DFFARX1 I_36376 (I221471,I3035,I621452,I621478,);
and I_36377 (I621486,I621478,I221456);
DFFARX1 I_36378 (I621486,I3035,I621452,I621435,);
DFFARX1 I_36379 (I221462,I3035,I621452,I621526,);
not I_36380 (I621534,I221444);
not I_36381 (I621551,I221465);
nand I_36382 (I621568,I621551,I621534);
nor I_36383 (I621423,I621526,I621568);
DFFARX1 I_36384 (I621568,I3035,I621452,I621608,);
not I_36385 (I621444,I621608);
not I_36386 (I621630,I221468);
nand I_36387 (I621647,I621551,I621630);
DFFARX1 I_36388 (I621647,I3035,I621452,I621673,);
not I_36389 (I621681,I621673);
not I_36390 (I621698,I221459);
nand I_36391 (I621715,I621698,I221447);
and I_36392 (I621732,I621534,I621715);
nor I_36393 (I621749,I621647,I621732);
DFFARX1 I_36394 (I621749,I3035,I621452,I621420,);
DFFARX1 I_36395 (I621732,I3035,I621452,I621441,);
nor I_36396 (I621794,I221459,I221453);
nor I_36397 (I621432,I621647,I621794);
or I_36398 (I621825,I221459,I221453);
nor I_36399 (I621842,I221450,I221444);
DFFARX1 I_36400 (I621842,I3035,I621452,I621868,);
not I_36401 (I621876,I621868);
nor I_36402 (I621438,I621876,I621681);
nand I_36403 (I621907,I621876,I621526);
not I_36404 (I621924,I221450);
nand I_36405 (I621941,I621924,I621630);
nand I_36406 (I621958,I621876,I621941);
nand I_36407 (I621429,I621958,I621907);
nand I_36408 (I621426,I621941,I621825);
not I_36409 (I622030,I3042);
DFFARX1 I_36410 (I97344,I3035,I622030,I622056,);
and I_36411 (I622064,I622056,I97347);
DFFARX1 I_36412 (I622064,I3035,I622030,I622013,);
DFFARX1 I_36413 (I97347,I3035,I622030,I622104,);
not I_36414 (I622112,I97362);
not I_36415 (I622129,I97368);
nand I_36416 (I622146,I622129,I622112);
nor I_36417 (I622001,I622104,I622146);
DFFARX1 I_36418 (I622146,I3035,I622030,I622186,);
not I_36419 (I622022,I622186);
not I_36420 (I622208,I97356);
nand I_36421 (I622225,I622129,I622208);
DFFARX1 I_36422 (I622225,I3035,I622030,I622251,);
not I_36423 (I622259,I622251);
not I_36424 (I622276,I97353);
nand I_36425 (I622293,I622276,I97350);
and I_36426 (I622310,I622112,I622293);
nor I_36427 (I622327,I622225,I622310);
DFFARX1 I_36428 (I622327,I3035,I622030,I621998,);
DFFARX1 I_36429 (I622310,I3035,I622030,I622019,);
nor I_36430 (I622372,I97353,I97344);
nor I_36431 (I622010,I622225,I622372);
or I_36432 (I622403,I97353,I97344);
nor I_36433 (I622420,I97359,I97365);
DFFARX1 I_36434 (I622420,I3035,I622030,I622446,);
not I_36435 (I622454,I622446);
nor I_36436 (I622016,I622454,I622259);
nand I_36437 (I622485,I622454,I622104);
not I_36438 (I622502,I97359);
nand I_36439 (I622519,I622502,I622208);
nand I_36440 (I622536,I622454,I622519);
nand I_36441 (I622007,I622536,I622485);
nand I_36442 (I622004,I622519,I622403);
not I_36443 (I622608,I3042);
DFFARX1 I_36444 (I691008,I3035,I622608,I622634,);
and I_36445 (I622642,I622634,I690990);
DFFARX1 I_36446 (I622642,I3035,I622608,I622591,);
DFFARX1 I_36447 (I690999,I3035,I622608,I622682,);
not I_36448 (I622690,I690984);
not I_36449 (I622707,I690996);
nand I_36450 (I622724,I622707,I622690);
nor I_36451 (I622579,I622682,I622724);
DFFARX1 I_36452 (I622724,I3035,I622608,I622764,);
not I_36453 (I622600,I622764);
not I_36454 (I622786,I690987);
nand I_36455 (I622803,I622707,I622786);
DFFARX1 I_36456 (I622803,I3035,I622608,I622829,);
not I_36457 (I622837,I622829);
not I_36458 (I622854,I690984);
nand I_36459 (I622871,I622854,I690987);
and I_36460 (I622888,I622690,I622871);
nor I_36461 (I622905,I622803,I622888);
DFFARX1 I_36462 (I622905,I3035,I622608,I622576,);
DFFARX1 I_36463 (I622888,I3035,I622608,I622597,);
nor I_36464 (I622950,I690984,I691005);
nor I_36465 (I622588,I622803,I622950);
or I_36466 (I622981,I690984,I691005);
nor I_36467 (I622998,I690993,I691002);
DFFARX1 I_36468 (I622998,I3035,I622608,I623024,);
not I_36469 (I623032,I623024);
nor I_36470 (I622594,I623032,I622837);
nand I_36471 (I623063,I623032,I622682);
not I_36472 (I623080,I690993);
nand I_36473 (I623097,I623080,I622786);
nand I_36474 (I623114,I623032,I623097);
nand I_36475 (I622585,I623114,I623063);
nand I_36476 (I622582,I623097,I622981);
not I_36477 (I623186,I3042);
DFFARX1 I_36478 (I649083,I3035,I623186,I623212,);
and I_36479 (I623220,I623212,I649077);
DFFARX1 I_36480 (I623220,I3035,I623186,I623169,);
DFFARX1 I_36481 (I649062,I3035,I623186,I623260,);
not I_36482 (I623268,I649068);
not I_36483 (I623285,I649080);
nand I_36484 (I623302,I623285,I623268);
nor I_36485 (I623157,I623260,I623302);
DFFARX1 I_36486 (I623302,I3035,I623186,I623342,);
not I_36487 (I623178,I623342);
not I_36488 (I623364,I649062);
nand I_36489 (I623381,I623285,I623364);
DFFARX1 I_36490 (I623381,I3035,I623186,I623407,);
not I_36491 (I623415,I623407);
not I_36492 (I623432,I649086);
nand I_36493 (I623449,I623432,I649074);
and I_36494 (I623466,I623268,I623449);
nor I_36495 (I623483,I623381,I623466);
DFFARX1 I_36496 (I623483,I3035,I623186,I623154,);
DFFARX1 I_36497 (I623466,I3035,I623186,I623175,);
nor I_36498 (I623528,I649086,I649065);
nor I_36499 (I623166,I623381,I623528);
or I_36500 (I623559,I649086,I649065);
nor I_36501 (I623576,I649071,I649065);
DFFARX1 I_36502 (I623576,I3035,I623186,I623602,);
not I_36503 (I623610,I623602);
nor I_36504 (I623172,I623610,I623415);
nand I_36505 (I623641,I623610,I623260);
not I_36506 (I623658,I649071);
nand I_36507 (I623675,I623658,I623364);
nand I_36508 (I623692,I623610,I623675);
nand I_36509 (I623163,I623692,I623641);
nand I_36510 (I623160,I623675,I623559);
not I_36511 (I623764,I3042);
DFFARX1 I_36512 (I301903,I3035,I623764,I623790,);
and I_36513 (I623798,I623790,I301891);
DFFARX1 I_36514 (I623798,I3035,I623764,I623747,);
DFFARX1 I_36515 (I301906,I3035,I623764,I623838,);
not I_36516 (I623846,I301897);
not I_36517 (I623863,I301888);
nand I_36518 (I623880,I623863,I623846);
nor I_36519 (I623735,I623838,I623880);
DFFARX1 I_36520 (I623880,I3035,I623764,I623920,);
not I_36521 (I623756,I623920);
not I_36522 (I623942,I301894);
nand I_36523 (I623959,I623863,I623942);
DFFARX1 I_36524 (I623959,I3035,I623764,I623985,);
not I_36525 (I623993,I623985);
not I_36526 (I624010,I301909);
nand I_36527 (I624027,I624010,I301912);
and I_36528 (I624044,I623846,I624027);
nor I_36529 (I624061,I623959,I624044);
DFFARX1 I_36530 (I624061,I3035,I623764,I623732,);
DFFARX1 I_36531 (I624044,I3035,I623764,I623753,);
nor I_36532 (I624106,I301909,I301888);
nor I_36533 (I623744,I623959,I624106);
or I_36534 (I624137,I301909,I301888);
nor I_36535 (I624154,I301900,I301891);
DFFARX1 I_36536 (I624154,I3035,I623764,I624180,);
not I_36537 (I624188,I624180);
nor I_36538 (I623750,I624188,I623993);
nand I_36539 (I624219,I624188,I623838);
not I_36540 (I624236,I301900);
nand I_36541 (I624253,I624236,I623942);
nand I_36542 (I624270,I624188,I624253);
nand I_36543 (I623741,I624270,I624219);
nand I_36544 (I623738,I624253,I624137);
not I_36545 (I624342,I3042);
DFFARX1 I_36546 (I73704,I3035,I624342,I624368,);
and I_36547 (I624376,I624368,I73680);
DFFARX1 I_36548 (I624376,I3035,I624342,I624325,);
DFFARX1 I_36549 (I73698,I3035,I624342,I624416,);
not I_36550 (I624424,I73686);
not I_36551 (I624441,I73683);
nand I_36552 (I624458,I624441,I624424);
nor I_36553 (I624313,I624416,I624458);
DFFARX1 I_36554 (I624458,I3035,I624342,I624498,);
not I_36555 (I624334,I624498);
not I_36556 (I624520,I73692);
nand I_36557 (I624537,I624441,I624520);
DFFARX1 I_36558 (I624537,I3035,I624342,I624563,);
not I_36559 (I624571,I624563);
not I_36560 (I624588,I73683);
nand I_36561 (I624605,I624588,I73701);
and I_36562 (I624622,I624424,I624605);
nor I_36563 (I624639,I624537,I624622);
DFFARX1 I_36564 (I624639,I3035,I624342,I624310,);
DFFARX1 I_36565 (I624622,I3035,I624342,I624331,);
nor I_36566 (I624684,I73683,I73695);
nor I_36567 (I624322,I624537,I624684);
or I_36568 (I624715,I73683,I73695);
nor I_36569 (I624732,I73689,I73680);
DFFARX1 I_36570 (I624732,I3035,I624342,I624758,);
not I_36571 (I624766,I624758);
nor I_36572 (I624328,I624766,I624571);
nand I_36573 (I624797,I624766,I624416);
not I_36574 (I624814,I73689);
nand I_36575 (I624831,I624814,I624520);
nand I_36576 (I624848,I624766,I624831);
nand I_36577 (I624319,I624848,I624797);
nand I_36578 (I624316,I624831,I624715);
not I_36579 (I624920,I3042);
DFFARX1 I_36580 (I446680,I3035,I624920,I624946,);
and I_36581 (I624954,I624946,I446686);
DFFARX1 I_36582 (I624954,I3035,I624920,I624903,);
DFFARX1 I_36583 (I446692,I3035,I624920,I624994,);
not I_36584 (I625002,I446677);
not I_36585 (I625019,I446677);
nand I_36586 (I625036,I625019,I625002);
nor I_36587 (I624891,I624994,I625036);
DFFARX1 I_36588 (I625036,I3035,I624920,I625076,);
not I_36589 (I624912,I625076);
not I_36590 (I625098,I446695);
nand I_36591 (I625115,I625019,I625098);
DFFARX1 I_36592 (I625115,I3035,I624920,I625141,);
not I_36593 (I625149,I625141);
not I_36594 (I625166,I446689);
nand I_36595 (I625183,I625166,I446680);
and I_36596 (I625200,I625002,I625183);
nor I_36597 (I625217,I625115,I625200);
DFFARX1 I_36598 (I625217,I3035,I624920,I624888,);
DFFARX1 I_36599 (I625200,I3035,I624920,I624909,);
nor I_36600 (I625262,I446689,I446698);
nor I_36601 (I624900,I625115,I625262);
or I_36602 (I625293,I446689,I446698);
nor I_36603 (I625310,I446683,I446683);
DFFARX1 I_36604 (I625310,I3035,I624920,I625336,);
not I_36605 (I625344,I625336);
nor I_36606 (I624906,I625344,I625149);
nand I_36607 (I625375,I625344,I624994);
not I_36608 (I625392,I446683);
nand I_36609 (I625409,I625392,I625098);
nand I_36610 (I625426,I625344,I625409);
nand I_36611 (I624897,I625426,I625375);
nand I_36612 (I624894,I625409,I625293);
not I_36613 (I625498,I3042);
DFFARX1 I_36614 (I99129,I3035,I625498,I625524,);
and I_36615 (I625532,I625524,I99132);
DFFARX1 I_36616 (I625532,I3035,I625498,I625481,);
DFFARX1 I_36617 (I99132,I3035,I625498,I625572,);
not I_36618 (I625580,I99147);
not I_36619 (I625597,I99153);
nand I_36620 (I625614,I625597,I625580);
nor I_36621 (I625469,I625572,I625614);
DFFARX1 I_36622 (I625614,I3035,I625498,I625654,);
not I_36623 (I625490,I625654);
not I_36624 (I625676,I99141);
nand I_36625 (I625693,I625597,I625676);
DFFARX1 I_36626 (I625693,I3035,I625498,I625719,);
not I_36627 (I625727,I625719);
not I_36628 (I625744,I99138);
nand I_36629 (I625761,I625744,I99135);
and I_36630 (I625778,I625580,I625761);
nor I_36631 (I625795,I625693,I625778);
DFFARX1 I_36632 (I625795,I3035,I625498,I625466,);
DFFARX1 I_36633 (I625778,I3035,I625498,I625487,);
nor I_36634 (I625840,I99138,I99129);
nor I_36635 (I625478,I625693,I625840);
or I_36636 (I625871,I99138,I99129);
nor I_36637 (I625888,I99144,I99150);
DFFARX1 I_36638 (I625888,I3035,I625498,I625914,);
not I_36639 (I625922,I625914);
nor I_36640 (I625484,I625922,I625727);
nand I_36641 (I625953,I625922,I625572);
not I_36642 (I625970,I99144);
nand I_36643 (I625987,I625970,I625676);
nand I_36644 (I626004,I625922,I625987);
nand I_36645 (I625475,I626004,I625953);
nand I_36646 (I625472,I625987,I625871);
not I_36647 (I626076,I3042);
DFFARX1 I_36648 (I565561,I3035,I626076,I626102,);
and I_36649 (I626110,I626102,I565558);
DFFARX1 I_36650 (I626110,I3035,I626076,I626059,);
DFFARX1 I_36651 (I565564,I3035,I626076,I626150,);
not I_36652 (I626158,I565567);
not I_36653 (I626175,I565561);
nand I_36654 (I626192,I626175,I626158);
nor I_36655 (I626047,I626150,I626192);
DFFARX1 I_36656 (I626192,I3035,I626076,I626232,);
not I_36657 (I626068,I626232);
not I_36658 (I626254,I565576);
nand I_36659 (I626271,I626175,I626254);
DFFARX1 I_36660 (I626271,I3035,I626076,I626297,);
not I_36661 (I626305,I626297);
not I_36662 (I626322,I565573);
nand I_36663 (I626339,I626322,I565579);
and I_36664 (I626356,I626158,I626339);
nor I_36665 (I626373,I626271,I626356);
DFFARX1 I_36666 (I626373,I3035,I626076,I626044,);
DFFARX1 I_36667 (I626356,I3035,I626076,I626065,);
nor I_36668 (I626418,I565573,I565558);
nor I_36669 (I626056,I626271,I626418);
or I_36670 (I626449,I565573,I565558);
nor I_36671 (I626466,I565570,I565564);
DFFARX1 I_36672 (I626466,I3035,I626076,I626492,);
not I_36673 (I626500,I626492);
nor I_36674 (I626062,I626500,I626305);
nand I_36675 (I626531,I626500,I626150);
not I_36676 (I626548,I565570);
nand I_36677 (I626565,I626548,I626254);
nand I_36678 (I626582,I626500,I626565);
nand I_36679 (I626053,I626582,I626531);
nand I_36680 (I626050,I626565,I626449);
not I_36681 (I626654,I3042);
DFFARX1 I_36682 (I433505,I3035,I626654,I626680,);
and I_36683 (I626688,I626680,I433511);
DFFARX1 I_36684 (I626688,I3035,I626654,I626637,);
DFFARX1 I_36685 (I433517,I3035,I626654,I626728,);
not I_36686 (I626736,I433502);
not I_36687 (I626753,I433502);
nand I_36688 (I626770,I626753,I626736);
nor I_36689 (I626625,I626728,I626770);
DFFARX1 I_36690 (I626770,I3035,I626654,I626810,);
not I_36691 (I626646,I626810);
not I_36692 (I626832,I433520);
nand I_36693 (I626849,I626753,I626832);
DFFARX1 I_36694 (I626849,I3035,I626654,I626875,);
not I_36695 (I626883,I626875);
not I_36696 (I626900,I433514);
nand I_36697 (I626917,I626900,I433505);
and I_36698 (I626934,I626736,I626917);
nor I_36699 (I626951,I626849,I626934);
DFFARX1 I_36700 (I626951,I3035,I626654,I626622,);
DFFARX1 I_36701 (I626934,I3035,I626654,I626643,);
nor I_36702 (I626996,I433514,I433523);
nor I_36703 (I626634,I626849,I626996);
or I_36704 (I627027,I433514,I433523);
nor I_36705 (I627044,I433508,I433508);
DFFARX1 I_36706 (I627044,I3035,I626654,I627070,);
not I_36707 (I627078,I627070);
nor I_36708 (I626640,I627078,I626883);
nand I_36709 (I627109,I627078,I626728);
not I_36710 (I627126,I433508);
nand I_36711 (I627143,I627126,I626832);
nand I_36712 (I627160,I627078,I627143);
nand I_36713 (I626631,I627160,I627109);
nand I_36714 (I626628,I627143,I627027);
not I_36715 (I627232,I3042);
DFFARX1 I_36716 (I340629,I3035,I627232,I627258,);
and I_36717 (I627266,I627258,I340617);
DFFARX1 I_36718 (I627266,I3035,I627232,I627215,);
DFFARX1 I_36719 (I340620,I3035,I627232,I627306,);
not I_36720 (I627314,I340614);
not I_36721 (I627331,I340638);
nand I_36722 (I627348,I627331,I627314);
nor I_36723 (I627203,I627306,I627348);
DFFARX1 I_36724 (I627348,I3035,I627232,I627388,);
not I_36725 (I627224,I627388);
not I_36726 (I627410,I340626);
nand I_36727 (I627427,I627331,I627410);
DFFARX1 I_36728 (I627427,I3035,I627232,I627453,);
not I_36729 (I627461,I627453);
not I_36730 (I627478,I340635);
nand I_36731 (I627495,I627478,I340632);
and I_36732 (I627512,I627314,I627495);
nor I_36733 (I627529,I627427,I627512);
DFFARX1 I_36734 (I627529,I3035,I627232,I627200,);
DFFARX1 I_36735 (I627512,I3035,I627232,I627221,);
nor I_36736 (I627574,I340635,I340623);
nor I_36737 (I627212,I627427,I627574);
or I_36738 (I627605,I340635,I340623);
nor I_36739 (I627622,I340614,I340617);
DFFARX1 I_36740 (I627622,I3035,I627232,I627648,);
not I_36741 (I627656,I627648);
nor I_36742 (I627218,I627656,I627461);
nand I_36743 (I627687,I627656,I627306);
not I_36744 (I627704,I340614);
nand I_36745 (I627721,I627704,I627410);
nand I_36746 (I627738,I627656,I627721);
nand I_36747 (I627209,I627738,I627687);
nand I_36748 (I627206,I627721,I627605);
not I_36749 (I627810,I3042);
DFFARX1 I_36750 (I455112,I3035,I627810,I627836,);
and I_36751 (I627844,I627836,I455118);
DFFARX1 I_36752 (I627844,I3035,I627810,I627793,);
DFFARX1 I_36753 (I455124,I3035,I627810,I627884,);
not I_36754 (I627892,I455109);
not I_36755 (I627909,I455109);
nand I_36756 (I627926,I627909,I627892);
nor I_36757 (I627781,I627884,I627926);
DFFARX1 I_36758 (I627926,I3035,I627810,I627966,);
not I_36759 (I627802,I627966);
not I_36760 (I627988,I455127);
nand I_36761 (I628005,I627909,I627988);
DFFARX1 I_36762 (I628005,I3035,I627810,I628031,);
not I_36763 (I628039,I628031);
not I_36764 (I628056,I455121);
nand I_36765 (I628073,I628056,I455112);
and I_36766 (I628090,I627892,I628073);
nor I_36767 (I628107,I628005,I628090);
DFFARX1 I_36768 (I628107,I3035,I627810,I627778,);
DFFARX1 I_36769 (I628090,I3035,I627810,I627799,);
nor I_36770 (I628152,I455121,I455130);
nor I_36771 (I627790,I628005,I628152);
or I_36772 (I628183,I455121,I455130);
nor I_36773 (I628200,I455115,I455115);
DFFARX1 I_36774 (I628200,I3035,I627810,I628226,);
not I_36775 (I628234,I628226);
nor I_36776 (I627796,I628234,I628039);
nand I_36777 (I628265,I628234,I627884);
not I_36778 (I628282,I455115);
nand I_36779 (I628299,I628282,I627988);
nand I_36780 (I628316,I628234,I628299);
nand I_36781 (I627787,I628316,I628265);
nand I_36782 (I627784,I628299,I628183);
not I_36783 (I628388,I3042);
DFFARX1 I_36784 (I662139,I3035,I628388,I628414,);
and I_36785 (I628422,I628414,I662133);
DFFARX1 I_36786 (I628422,I3035,I628388,I628371,);
DFFARX1 I_36787 (I662118,I3035,I628388,I628462,);
not I_36788 (I628470,I662124);
not I_36789 (I628487,I662136);
nand I_36790 (I628504,I628487,I628470);
nor I_36791 (I628359,I628462,I628504);
DFFARX1 I_36792 (I628504,I3035,I628388,I628544,);
not I_36793 (I628380,I628544);
not I_36794 (I628566,I662118);
nand I_36795 (I628583,I628487,I628566);
DFFARX1 I_36796 (I628583,I3035,I628388,I628609,);
not I_36797 (I628617,I628609);
not I_36798 (I628634,I662142);
nand I_36799 (I628651,I628634,I662130);
and I_36800 (I628668,I628470,I628651);
nor I_36801 (I628685,I628583,I628668);
DFFARX1 I_36802 (I628685,I3035,I628388,I628356,);
DFFARX1 I_36803 (I628668,I3035,I628388,I628377,);
nor I_36804 (I628730,I662142,I662121);
nor I_36805 (I628368,I628583,I628730);
or I_36806 (I628761,I662142,I662121);
nor I_36807 (I628778,I662127,I662121);
DFFARX1 I_36808 (I628778,I3035,I628388,I628804,);
not I_36809 (I628812,I628804);
nor I_36810 (I628374,I628812,I628617);
nand I_36811 (I628843,I628812,I628462);
not I_36812 (I628860,I662127);
nand I_36813 (I628877,I628860,I628566);
nand I_36814 (I628894,I628812,I628877);
nand I_36815 (I628365,I628894,I628843);
nand I_36816 (I628362,I628877,I628761);
not I_36817 (I628966,I3042);
DFFARX1 I_36818 (I26250,I3035,I628966,I628992,);
and I_36819 (I629000,I628992,I26253);
DFFARX1 I_36820 (I629000,I3035,I628966,I628949,);
DFFARX1 I_36821 (I26253,I3035,I628966,I629040,);
not I_36822 (I629048,I26256);
not I_36823 (I629065,I26271);
nand I_36824 (I629082,I629065,I629048);
nor I_36825 (I628937,I629040,I629082);
DFFARX1 I_36826 (I629082,I3035,I628966,I629122,);
not I_36827 (I628958,I629122);
not I_36828 (I629144,I26265);
nand I_36829 (I629161,I629065,I629144);
DFFARX1 I_36830 (I629161,I3035,I628966,I629187,);
not I_36831 (I629195,I629187);
not I_36832 (I629212,I26268);
nand I_36833 (I629229,I629212,I26250);
and I_36834 (I629246,I629048,I629229);
nor I_36835 (I629263,I629161,I629246);
DFFARX1 I_36836 (I629263,I3035,I628966,I628934,);
DFFARX1 I_36837 (I629246,I3035,I628966,I628955,);
nor I_36838 (I629308,I26268,I26262);
nor I_36839 (I628946,I629161,I629308);
or I_36840 (I629339,I26268,I26262);
nor I_36841 (I629356,I26259,I26274);
DFFARX1 I_36842 (I629356,I3035,I628966,I629382,);
not I_36843 (I629390,I629382);
nor I_36844 (I628952,I629390,I629195);
nand I_36845 (I629421,I629390,I629040);
not I_36846 (I629438,I26259);
nand I_36847 (I629455,I629438,I629144);
nand I_36848 (I629472,I629390,I629455);
nand I_36849 (I628943,I629472,I629421);
nand I_36850 (I628940,I629455,I629339);
not I_36851 (I629544,I3042);
DFFARX1 I_36852 (I2404,I3035,I629544,I629570,);
and I_36853 (I629578,I629570,I1740);
DFFARX1 I_36854 (I629578,I3035,I629544,I629527,);
DFFARX1 I_36855 (I2236,I3035,I629544,I629618,);
not I_36856 (I629626,I1372);
not I_36857 (I629643,I2044);
nand I_36858 (I629660,I629643,I629626);
nor I_36859 (I629515,I629618,I629660);
DFFARX1 I_36860 (I629660,I3035,I629544,I629700,);
not I_36861 (I629536,I629700);
not I_36862 (I629722,I2836);
nand I_36863 (I629739,I629643,I629722);
DFFARX1 I_36864 (I629739,I3035,I629544,I629765,);
not I_36865 (I629773,I629765);
not I_36866 (I629790,I2300);
nand I_36867 (I629807,I629790,I2900);
and I_36868 (I629824,I629626,I629807);
nor I_36869 (I629841,I629739,I629824);
DFFARX1 I_36870 (I629841,I3035,I629544,I629512,);
DFFARX1 I_36871 (I629824,I3035,I629544,I629533,);
nor I_36872 (I629886,I2300,I2684);
nor I_36873 (I629524,I629739,I629886);
or I_36874 (I629917,I2300,I2684);
nor I_36875 (I629934,I2980,I2676);
DFFARX1 I_36876 (I629934,I3035,I629544,I629960,);
not I_36877 (I629968,I629960);
nor I_36878 (I629530,I629968,I629773);
nand I_36879 (I629999,I629968,I629618);
not I_36880 (I630016,I2980);
nand I_36881 (I630033,I630016,I629722);
nand I_36882 (I630050,I629968,I630033);
nand I_36883 (I629521,I630050,I629999);
nand I_36884 (I629518,I630033,I629917);
not I_36885 (I630122,I3042);
DFFARX1 I_36886 (I404209,I3035,I630122,I630148,);
and I_36887 (I630156,I630148,I404197);
DFFARX1 I_36888 (I630156,I3035,I630122,I630105,);
DFFARX1 I_36889 (I404200,I3035,I630122,I630196,);
not I_36890 (I630204,I404194);
not I_36891 (I630221,I404218);
nand I_36892 (I630238,I630221,I630204);
nor I_36893 (I630093,I630196,I630238);
DFFARX1 I_36894 (I630238,I3035,I630122,I630278,);
not I_36895 (I630114,I630278);
not I_36896 (I630300,I404206);
nand I_36897 (I630317,I630221,I630300);
DFFARX1 I_36898 (I630317,I3035,I630122,I630343,);
not I_36899 (I630351,I630343);
not I_36900 (I630368,I404215);
nand I_36901 (I630385,I630368,I404212);
and I_36902 (I630402,I630204,I630385);
nor I_36903 (I630419,I630317,I630402);
DFFARX1 I_36904 (I630419,I3035,I630122,I630090,);
DFFARX1 I_36905 (I630402,I3035,I630122,I630111,);
nor I_36906 (I630464,I404215,I404203);
nor I_36907 (I630102,I630317,I630464);
or I_36908 (I630495,I404215,I404203);
nor I_36909 (I630512,I404194,I404197);
DFFARX1 I_36910 (I630512,I3035,I630122,I630538,);
not I_36911 (I630546,I630538);
nor I_36912 (I630108,I630546,I630351);
nand I_36913 (I630577,I630546,I630196);
not I_36914 (I630594,I404194);
nand I_36915 (I630611,I630594,I630300);
nand I_36916 (I630628,I630546,I630611);
nand I_36917 (I630099,I630628,I630577);
nand I_36918 (I630096,I630611,I630495);
not I_36919 (I630700,I3042);
DFFARX1 I_36920 (I518066,I3035,I630700,I630726,);
and I_36921 (I630734,I630726,I518060);
DFFARX1 I_36922 (I630734,I3035,I630700,I630683,);
DFFARX1 I_36923 (I518078,I3035,I630700,I630774,);
not I_36924 (I630782,I518069);
not I_36925 (I630799,I518081);
nand I_36926 (I630816,I630799,I630782);
nor I_36927 (I630671,I630774,I630816);
DFFARX1 I_36928 (I630816,I3035,I630700,I630856,);
not I_36929 (I630692,I630856);
not I_36930 (I630878,I518087);
nand I_36931 (I630895,I630799,I630878);
DFFARX1 I_36932 (I630895,I3035,I630700,I630921,);
not I_36933 (I630929,I630921);
not I_36934 (I630946,I518063);
nand I_36935 (I630963,I630946,I518084);
and I_36936 (I630980,I630782,I630963);
nor I_36937 (I630997,I630895,I630980);
DFFARX1 I_36938 (I630997,I3035,I630700,I630668,);
DFFARX1 I_36939 (I630980,I3035,I630700,I630689,);
nor I_36940 (I631042,I518063,I518075);
nor I_36941 (I630680,I630895,I631042);
or I_36942 (I631073,I518063,I518075);
nor I_36943 (I631090,I518060,I518072);
DFFARX1 I_36944 (I631090,I3035,I630700,I631116,);
not I_36945 (I631124,I631116);
nor I_36946 (I630686,I631124,I630929);
nand I_36947 (I631155,I631124,I630774);
not I_36948 (I631172,I518060);
nand I_36949 (I631189,I631172,I630878);
nand I_36950 (I631206,I631124,I631189);
nand I_36951 (I630677,I631206,I631155);
nand I_36952 (I630674,I631189,I631073);
not I_36953 (I631278,I3042);
DFFARX1 I_36954 (I510314,I3035,I631278,I631304,);
and I_36955 (I631312,I631304,I510308);
DFFARX1 I_36956 (I631312,I3035,I631278,I631261,);
DFFARX1 I_36957 (I510326,I3035,I631278,I631352,);
not I_36958 (I631360,I510317);
not I_36959 (I631377,I510329);
nand I_36960 (I631394,I631377,I631360);
nor I_36961 (I631249,I631352,I631394);
DFFARX1 I_36962 (I631394,I3035,I631278,I631434,);
not I_36963 (I631270,I631434);
not I_36964 (I631456,I510335);
nand I_36965 (I631473,I631377,I631456);
DFFARX1 I_36966 (I631473,I3035,I631278,I631499,);
not I_36967 (I631507,I631499);
not I_36968 (I631524,I510311);
nand I_36969 (I631541,I631524,I510332);
and I_36970 (I631558,I631360,I631541);
nor I_36971 (I631575,I631473,I631558);
DFFARX1 I_36972 (I631575,I3035,I631278,I631246,);
DFFARX1 I_36973 (I631558,I3035,I631278,I631267,);
nor I_36974 (I631620,I510311,I510323);
nor I_36975 (I631258,I631473,I631620);
or I_36976 (I631651,I510311,I510323);
nor I_36977 (I631668,I510308,I510320);
DFFARX1 I_36978 (I631668,I3035,I631278,I631694,);
not I_36979 (I631702,I631694);
nor I_36980 (I631264,I631702,I631507);
nand I_36981 (I631733,I631702,I631352);
not I_36982 (I631750,I510308);
nand I_36983 (I631767,I631750,I631456);
nand I_36984 (I631784,I631702,I631767);
nand I_36985 (I631255,I631784,I631733);
nand I_36986 (I631252,I631767,I631651);
not I_36987 (I631856,I3042);
DFFARX1 I_36988 (I678870,I3035,I631856,I631882,);
and I_36989 (I631890,I631882,I678852);
DFFARX1 I_36990 (I631890,I3035,I631856,I631839,);
DFFARX1 I_36991 (I678861,I3035,I631856,I631930,);
not I_36992 (I631938,I678846);
not I_36993 (I631955,I678858);
nand I_36994 (I631972,I631955,I631938);
nor I_36995 (I631827,I631930,I631972);
DFFARX1 I_36996 (I631972,I3035,I631856,I632012,);
not I_36997 (I631848,I632012);
not I_36998 (I632034,I678849);
nand I_36999 (I632051,I631955,I632034);
DFFARX1 I_37000 (I632051,I3035,I631856,I632077,);
not I_37001 (I632085,I632077);
not I_37002 (I632102,I678846);
nand I_37003 (I632119,I632102,I678849);
and I_37004 (I632136,I631938,I632119);
nor I_37005 (I632153,I632051,I632136);
DFFARX1 I_37006 (I632153,I3035,I631856,I631824,);
DFFARX1 I_37007 (I632136,I3035,I631856,I631845,);
nor I_37008 (I632198,I678846,I678867);
nor I_37009 (I631836,I632051,I632198);
or I_37010 (I632229,I678846,I678867);
nor I_37011 (I632246,I678855,I678864);
DFFARX1 I_37012 (I632246,I3035,I631856,I632272,);
not I_37013 (I632280,I632272);
nor I_37014 (I631842,I632280,I632085);
nand I_37015 (I632311,I632280,I631930);
not I_37016 (I632328,I678855);
nand I_37017 (I632345,I632328,I632034);
nand I_37018 (I632362,I632280,I632345);
nand I_37019 (I631833,I632362,I632311);
nand I_37020 (I631830,I632345,I632229);
not I_37021 (I632434,I3042);
DFFARX1 I_37022 (I399585,I3035,I632434,I632460,);
and I_37023 (I632468,I632460,I399573);
DFFARX1 I_37024 (I632468,I3035,I632434,I632417,);
DFFARX1 I_37025 (I399576,I3035,I632434,I632508,);
not I_37026 (I632516,I399570);
not I_37027 (I632533,I399594);
nand I_37028 (I632550,I632533,I632516);
nor I_37029 (I632405,I632508,I632550);
DFFARX1 I_37030 (I632550,I3035,I632434,I632590,);
not I_37031 (I632426,I632590);
not I_37032 (I632612,I399582);
nand I_37033 (I632629,I632533,I632612);
DFFARX1 I_37034 (I632629,I3035,I632434,I632655,);
not I_37035 (I632663,I632655);
not I_37036 (I632680,I399591);
nand I_37037 (I632697,I632680,I399588);
and I_37038 (I632714,I632516,I632697);
nor I_37039 (I632731,I632629,I632714);
DFFARX1 I_37040 (I632731,I3035,I632434,I632402,);
DFFARX1 I_37041 (I632714,I3035,I632434,I632423,);
nor I_37042 (I632776,I399591,I399579);
nor I_37043 (I632414,I632629,I632776);
or I_37044 (I632807,I399591,I399579);
nor I_37045 (I632824,I399570,I399573);
DFFARX1 I_37046 (I632824,I3035,I632434,I632850,);
not I_37047 (I632858,I632850);
nor I_37048 (I632420,I632858,I632663);
nand I_37049 (I632889,I632858,I632508);
not I_37050 (I632906,I399570);
nand I_37051 (I632923,I632906,I632612);
nand I_37052 (I632940,I632858,I632923);
nand I_37053 (I632411,I632940,I632889);
nand I_37054 (I632408,I632923,I632807);
not I_37055 (I633012,I3042);
DFFARX1 I_37056 (I411145,I3035,I633012,I633038,);
and I_37057 (I633046,I633038,I411133);
DFFARX1 I_37058 (I633046,I3035,I633012,I632995,);
DFFARX1 I_37059 (I411136,I3035,I633012,I633086,);
not I_37060 (I633094,I411130);
not I_37061 (I633111,I411154);
nand I_37062 (I633128,I633111,I633094);
nor I_37063 (I632983,I633086,I633128);
DFFARX1 I_37064 (I633128,I3035,I633012,I633168,);
not I_37065 (I633004,I633168);
not I_37066 (I633190,I411142);
nand I_37067 (I633207,I633111,I633190);
DFFARX1 I_37068 (I633207,I3035,I633012,I633233,);
not I_37069 (I633241,I633233);
not I_37070 (I633258,I411151);
nand I_37071 (I633275,I633258,I411148);
and I_37072 (I633292,I633094,I633275);
nor I_37073 (I633309,I633207,I633292);
DFFARX1 I_37074 (I633309,I3035,I633012,I632980,);
DFFARX1 I_37075 (I633292,I3035,I633012,I633001,);
nor I_37076 (I633354,I411151,I411139);
nor I_37077 (I632992,I633207,I633354);
or I_37078 (I633385,I411151,I411139);
nor I_37079 (I633402,I411130,I411133);
DFFARX1 I_37080 (I633402,I3035,I633012,I633428,);
not I_37081 (I633436,I633428);
nor I_37082 (I632998,I633436,I633241);
nand I_37083 (I633467,I633436,I633086);
not I_37084 (I633484,I411130);
nand I_37085 (I633501,I633484,I633190);
nand I_37086 (I633518,I633436,I633501);
nand I_37087 (I632989,I633518,I633467);
nand I_37088 (I632986,I633501,I633385);
not I_37089 (I633590,I3042);
DFFARX1 I_37090 (I374731,I3035,I633590,I633616,);
and I_37091 (I633624,I633616,I374719);
DFFARX1 I_37092 (I633624,I3035,I633590,I633573,);
DFFARX1 I_37093 (I374722,I3035,I633590,I633664,);
not I_37094 (I633672,I374716);
not I_37095 (I633689,I374740);
nand I_37096 (I633706,I633689,I633672);
nor I_37097 (I633561,I633664,I633706);
DFFARX1 I_37098 (I633706,I3035,I633590,I633746,);
not I_37099 (I633582,I633746);
not I_37100 (I633768,I374728);
nand I_37101 (I633785,I633689,I633768);
DFFARX1 I_37102 (I633785,I3035,I633590,I633811,);
not I_37103 (I633819,I633811);
not I_37104 (I633836,I374737);
nand I_37105 (I633853,I633836,I374734);
and I_37106 (I633870,I633672,I633853);
nor I_37107 (I633887,I633785,I633870);
DFFARX1 I_37108 (I633887,I3035,I633590,I633558,);
DFFARX1 I_37109 (I633870,I3035,I633590,I633579,);
nor I_37110 (I633932,I374737,I374725);
nor I_37111 (I633570,I633785,I633932);
or I_37112 (I633963,I374737,I374725);
nor I_37113 (I633980,I374716,I374719);
DFFARX1 I_37114 (I633980,I3035,I633590,I634006,);
not I_37115 (I634014,I634006);
nor I_37116 (I633576,I634014,I633819);
nand I_37117 (I634045,I634014,I633664);
not I_37118 (I634062,I374716);
nand I_37119 (I634079,I634062,I633768);
nand I_37120 (I634096,I634014,I634079);
nand I_37121 (I633567,I634096,I634045);
nand I_37122 (I633564,I634079,I633963);
not I_37123 (I634168,I3042);
DFFARX1 I_37124 (I207769,I3035,I634168,I634194,);
and I_37125 (I634202,I634194,I207754);
DFFARX1 I_37126 (I634202,I3035,I634168,I634151,);
DFFARX1 I_37127 (I207760,I3035,I634168,I634242,);
not I_37128 (I634250,I207742);
not I_37129 (I634267,I207763);
nand I_37130 (I634284,I634267,I634250);
nor I_37131 (I634139,I634242,I634284);
DFFARX1 I_37132 (I634284,I3035,I634168,I634324,);
not I_37133 (I634160,I634324);
not I_37134 (I634346,I207766);
nand I_37135 (I634363,I634267,I634346);
DFFARX1 I_37136 (I634363,I3035,I634168,I634389,);
not I_37137 (I634397,I634389);
not I_37138 (I634414,I207757);
nand I_37139 (I634431,I634414,I207745);
and I_37140 (I634448,I634250,I634431);
nor I_37141 (I634465,I634363,I634448);
DFFARX1 I_37142 (I634465,I3035,I634168,I634136,);
DFFARX1 I_37143 (I634448,I3035,I634168,I634157,);
nor I_37144 (I634510,I207757,I207751);
nor I_37145 (I634148,I634363,I634510);
or I_37146 (I634541,I207757,I207751);
nor I_37147 (I634558,I207748,I207742);
DFFARX1 I_37148 (I634558,I3035,I634168,I634584,);
not I_37149 (I634592,I634584);
nor I_37150 (I634154,I634592,I634397);
nand I_37151 (I634623,I634592,I634242);
not I_37152 (I634640,I207748);
nand I_37153 (I634657,I634640,I634346);
nand I_37154 (I634674,I634592,I634657);
nand I_37155 (I634145,I634674,I634623);
nand I_37156 (I634142,I634657,I634541);
not I_37157 (I634746,I3042);
DFFARX1 I_37158 (I351033,I3035,I634746,I634772,);
and I_37159 (I634780,I634772,I351021);
DFFARX1 I_37160 (I634780,I3035,I634746,I634729,);
DFFARX1 I_37161 (I351024,I3035,I634746,I634820,);
not I_37162 (I634828,I351018);
not I_37163 (I634845,I351042);
nand I_37164 (I634862,I634845,I634828);
nor I_37165 (I634717,I634820,I634862);
DFFARX1 I_37166 (I634862,I3035,I634746,I634902,);
not I_37167 (I634738,I634902);
not I_37168 (I634924,I351030);
nand I_37169 (I634941,I634845,I634924);
DFFARX1 I_37170 (I634941,I3035,I634746,I634967,);
not I_37171 (I634975,I634967);
not I_37172 (I634992,I351039);
nand I_37173 (I635009,I634992,I351036);
and I_37174 (I635026,I634828,I635009);
nor I_37175 (I635043,I634941,I635026);
DFFARX1 I_37176 (I635043,I3035,I634746,I634714,);
DFFARX1 I_37177 (I635026,I3035,I634746,I634735,);
nor I_37178 (I635088,I351039,I351027);
nor I_37179 (I634726,I634941,I635088);
or I_37180 (I635119,I351039,I351027);
nor I_37181 (I635136,I351018,I351021);
DFFARX1 I_37182 (I635136,I3035,I634746,I635162,);
not I_37183 (I635170,I635162);
nor I_37184 (I634732,I635170,I634975);
nand I_37185 (I635201,I635170,I634820);
not I_37186 (I635218,I351018);
nand I_37187 (I635235,I635218,I634924);
nand I_37188 (I635252,I635170,I635235);
nand I_37189 (I634723,I635252,I635201);
nand I_37190 (I634720,I635235,I635119);
not I_37191 (I635324,I3042);
DFFARX1 I_37192 (I253829,I3035,I635324,I635350,);
and I_37193 (I635358,I635350,I253844);
DFFARX1 I_37194 (I635358,I3035,I635324,I635307,);
DFFARX1 I_37195 (I253847,I3035,I635324,I635398,);
not I_37196 (I635406,I253841);
not I_37197 (I635423,I253856);
nand I_37198 (I635440,I635423,I635406);
nor I_37199 (I635295,I635398,I635440);
DFFARX1 I_37200 (I635440,I3035,I635324,I635480,);
not I_37201 (I635316,I635480);
not I_37202 (I635502,I253832);
nand I_37203 (I635519,I635423,I635502);
DFFARX1 I_37204 (I635519,I3035,I635324,I635545,);
not I_37205 (I635553,I635545);
not I_37206 (I635570,I253835);
nand I_37207 (I635587,I635570,I253829);
and I_37208 (I635604,I635406,I635587);
nor I_37209 (I635621,I635519,I635604);
DFFARX1 I_37210 (I635621,I3035,I635324,I635292,);
DFFARX1 I_37211 (I635604,I3035,I635324,I635313,);
nor I_37212 (I635666,I253835,I253838);
nor I_37213 (I635304,I635519,I635666);
or I_37214 (I635697,I253835,I253838);
nor I_37215 (I635714,I253853,I253850);
DFFARX1 I_37216 (I635714,I3035,I635324,I635740,);
not I_37217 (I635748,I635740);
nor I_37218 (I635310,I635748,I635553);
nand I_37219 (I635779,I635748,I635398);
not I_37220 (I635796,I253853);
nand I_37221 (I635813,I635796,I635502);
nand I_37222 (I635830,I635748,I635813);
nand I_37223 (I635301,I635830,I635779);
nand I_37224 (I635298,I635813,I635697);
not I_37225 (I635902,I3042);
DFFARX1 I_37226 (I377043,I3035,I635902,I635928,);
and I_37227 (I635936,I635928,I377031);
DFFARX1 I_37228 (I635936,I3035,I635902,I635885,);
DFFARX1 I_37229 (I377034,I3035,I635902,I635976,);
not I_37230 (I635984,I377028);
not I_37231 (I636001,I377052);
nand I_37232 (I636018,I636001,I635984);
nor I_37233 (I635873,I635976,I636018);
DFFARX1 I_37234 (I636018,I3035,I635902,I636058,);
not I_37235 (I635894,I636058);
not I_37236 (I636080,I377040);
nand I_37237 (I636097,I636001,I636080);
DFFARX1 I_37238 (I636097,I3035,I635902,I636123,);
not I_37239 (I636131,I636123);
not I_37240 (I636148,I377049);
nand I_37241 (I636165,I636148,I377046);
and I_37242 (I636182,I635984,I636165);
nor I_37243 (I636199,I636097,I636182);
DFFARX1 I_37244 (I636199,I3035,I635902,I635870,);
DFFARX1 I_37245 (I636182,I3035,I635902,I635891,);
nor I_37246 (I636244,I377049,I377037);
nor I_37247 (I635882,I636097,I636244);
or I_37248 (I636275,I377049,I377037);
nor I_37249 (I636292,I377028,I377031);
DFFARX1 I_37250 (I636292,I3035,I635902,I636318,);
not I_37251 (I636326,I636318);
nor I_37252 (I635888,I636326,I636131);
nand I_37253 (I636357,I636326,I635976);
not I_37254 (I636374,I377028);
nand I_37255 (I636391,I636374,I636080);
nand I_37256 (I636408,I636326,I636391);
nand I_37257 (I635879,I636408,I636357);
nand I_37258 (I635876,I636391,I636275);
not I_37259 (I636480,I3042);
DFFARX1 I_37260 (I386869,I3035,I636480,I636506,);
and I_37261 (I636514,I636506,I386857);
DFFARX1 I_37262 (I636514,I3035,I636480,I636463,);
DFFARX1 I_37263 (I386860,I3035,I636480,I636554,);
not I_37264 (I636562,I386854);
not I_37265 (I636579,I386878);
nand I_37266 (I636596,I636579,I636562);
nor I_37267 (I636451,I636554,I636596);
DFFARX1 I_37268 (I636596,I3035,I636480,I636636,);
not I_37269 (I636472,I636636);
not I_37270 (I636658,I386866);
nand I_37271 (I636675,I636579,I636658);
DFFARX1 I_37272 (I636675,I3035,I636480,I636701,);
not I_37273 (I636709,I636701);
not I_37274 (I636726,I386875);
nand I_37275 (I636743,I636726,I386872);
and I_37276 (I636760,I636562,I636743);
nor I_37277 (I636777,I636675,I636760);
DFFARX1 I_37278 (I636777,I3035,I636480,I636448,);
DFFARX1 I_37279 (I636760,I3035,I636480,I636469,);
nor I_37280 (I636822,I386875,I386863);
nor I_37281 (I636460,I636675,I636822);
or I_37282 (I636853,I386875,I386863);
nor I_37283 (I636870,I386854,I386857);
DFFARX1 I_37284 (I636870,I3035,I636480,I636896,);
not I_37285 (I636904,I636896);
nor I_37286 (I636466,I636904,I636709);
nand I_37287 (I636935,I636904,I636554);
not I_37288 (I636952,I386854);
nand I_37289 (I636969,I636952,I636658);
nand I_37290 (I636986,I636904,I636969);
nand I_37291 (I636457,I636986,I636935);
nand I_37292 (I636454,I636969,I636853);
not I_37293 (I637058,I3042);
DFFARX1 I_37294 (I177203,I3035,I637058,I637084,);
and I_37295 (I637092,I637084,I177188);
DFFARX1 I_37296 (I637092,I3035,I637058,I637041,);
DFFARX1 I_37297 (I177194,I3035,I637058,I637132,);
not I_37298 (I637140,I177176);
not I_37299 (I637157,I177197);
nand I_37300 (I637174,I637157,I637140);
nor I_37301 (I637029,I637132,I637174);
DFFARX1 I_37302 (I637174,I3035,I637058,I637214,);
not I_37303 (I637050,I637214);
not I_37304 (I637236,I177200);
nand I_37305 (I637253,I637157,I637236);
DFFARX1 I_37306 (I637253,I3035,I637058,I637279,);
not I_37307 (I637287,I637279);
not I_37308 (I637304,I177191);
nand I_37309 (I637321,I637304,I177179);
and I_37310 (I637338,I637140,I637321);
nor I_37311 (I637355,I637253,I637338);
DFFARX1 I_37312 (I637355,I3035,I637058,I637026,);
DFFARX1 I_37313 (I637338,I3035,I637058,I637047,);
nor I_37314 (I637400,I177191,I177185);
nor I_37315 (I637038,I637253,I637400);
or I_37316 (I637431,I177191,I177185);
nor I_37317 (I637448,I177182,I177176);
DFFARX1 I_37318 (I637448,I3035,I637058,I637474,);
not I_37319 (I637482,I637474);
nor I_37320 (I637044,I637482,I637287);
nand I_37321 (I637513,I637482,I637132);
not I_37322 (I637530,I177182);
nand I_37323 (I637547,I637530,I637236);
nand I_37324 (I637564,I637482,I637547);
nand I_37325 (I637035,I637564,I637513);
nand I_37326 (I637032,I637547,I637431);
not I_37327 (I637636,I3042);
DFFARX1 I_37328 (I419803,I3035,I637636,I637662,);
and I_37329 (I637670,I637662,I419809);
DFFARX1 I_37330 (I637670,I3035,I637636,I637619,);
DFFARX1 I_37331 (I419815,I3035,I637636,I637710,);
not I_37332 (I637718,I419800);
not I_37333 (I637735,I419800);
nand I_37334 (I637752,I637735,I637718);
nor I_37335 (I637607,I637710,I637752);
DFFARX1 I_37336 (I637752,I3035,I637636,I637792,);
not I_37337 (I637628,I637792);
not I_37338 (I637814,I419818);
nand I_37339 (I637831,I637735,I637814);
DFFARX1 I_37340 (I637831,I3035,I637636,I637857,);
not I_37341 (I637865,I637857);
not I_37342 (I637882,I419812);
nand I_37343 (I637899,I637882,I419803);
and I_37344 (I637916,I637718,I637899);
nor I_37345 (I637933,I637831,I637916);
DFFARX1 I_37346 (I637933,I3035,I637636,I637604,);
DFFARX1 I_37347 (I637916,I3035,I637636,I637625,);
nor I_37348 (I637978,I419812,I419821);
nor I_37349 (I637616,I637831,I637978);
or I_37350 (I638009,I419812,I419821);
nor I_37351 (I638026,I419806,I419806);
DFFARX1 I_37352 (I638026,I3035,I637636,I638052,);
not I_37353 (I638060,I638052);
nor I_37354 (I637622,I638060,I637865);
nand I_37355 (I638091,I638060,I637710);
not I_37356 (I638108,I419806);
nand I_37357 (I638125,I638108,I637814);
nand I_37358 (I638142,I638060,I638125);
nand I_37359 (I637613,I638142,I638091);
nand I_37360 (I637610,I638125,I638009);
not I_37361 (I638214,I3042);
DFFARX1 I_37362 (I196702,I3035,I638214,I638240,);
and I_37363 (I638248,I638240,I196687);
DFFARX1 I_37364 (I638248,I3035,I638214,I638197,);
DFFARX1 I_37365 (I196693,I3035,I638214,I638288,);
not I_37366 (I638296,I196675);
not I_37367 (I638313,I196696);
nand I_37368 (I638330,I638313,I638296);
nor I_37369 (I638185,I638288,I638330);
DFFARX1 I_37370 (I638330,I3035,I638214,I638370,);
not I_37371 (I638206,I638370);
not I_37372 (I638392,I196699);
nand I_37373 (I638409,I638313,I638392);
DFFARX1 I_37374 (I638409,I3035,I638214,I638435,);
not I_37375 (I638443,I638435);
not I_37376 (I638460,I196690);
nand I_37377 (I638477,I638460,I196678);
and I_37378 (I638494,I638296,I638477);
nor I_37379 (I638511,I638409,I638494);
DFFARX1 I_37380 (I638511,I3035,I638214,I638182,);
DFFARX1 I_37381 (I638494,I3035,I638214,I638203,);
nor I_37382 (I638556,I196690,I196684);
nor I_37383 (I638194,I638409,I638556);
or I_37384 (I638587,I196690,I196684);
nor I_37385 (I638604,I196681,I196675);
DFFARX1 I_37386 (I638604,I3035,I638214,I638630,);
not I_37387 (I638638,I638630);
nor I_37388 (I638200,I638638,I638443);
nand I_37389 (I638669,I638638,I638288);
not I_37390 (I638686,I196681);
nand I_37391 (I638703,I638686,I638392);
nand I_37392 (I638720,I638638,I638703);
nand I_37393 (I638191,I638720,I638669);
nand I_37394 (I638188,I638703,I638587);
not I_37395 (I638792,I3042);
DFFARX1 I_37396 (I170352,I3035,I638792,I638818,);
and I_37397 (I638826,I638818,I170337);
DFFARX1 I_37398 (I638826,I3035,I638792,I638775,);
DFFARX1 I_37399 (I170343,I3035,I638792,I638866,);
not I_37400 (I638874,I170325);
not I_37401 (I638891,I170346);
nand I_37402 (I638908,I638891,I638874);
nor I_37403 (I638763,I638866,I638908);
DFFARX1 I_37404 (I638908,I3035,I638792,I638948,);
not I_37405 (I638784,I638948);
not I_37406 (I638970,I170349);
nand I_37407 (I638987,I638891,I638970);
DFFARX1 I_37408 (I638987,I3035,I638792,I639013,);
not I_37409 (I639021,I639013);
not I_37410 (I639038,I170340);
nand I_37411 (I639055,I639038,I170328);
and I_37412 (I639072,I638874,I639055);
nor I_37413 (I639089,I638987,I639072);
DFFARX1 I_37414 (I639089,I3035,I638792,I638760,);
DFFARX1 I_37415 (I639072,I3035,I638792,I638781,);
nor I_37416 (I639134,I170340,I170334);
nor I_37417 (I638772,I638987,I639134);
or I_37418 (I639165,I170340,I170334);
nor I_37419 (I639182,I170331,I170325);
DFFARX1 I_37420 (I639182,I3035,I638792,I639208,);
not I_37421 (I639216,I639208);
nor I_37422 (I638778,I639216,I639021);
nand I_37423 (I639247,I639216,I638866);
not I_37424 (I639264,I170331);
nand I_37425 (I639281,I639264,I638970);
nand I_37426 (I639298,I639216,I639281);
nand I_37427 (I638769,I639298,I639247);
nand I_37428 (I638766,I639281,I639165);
not I_37429 (I639370,I3042);
DFFARX1 I_37430 (I171406,I3035,I639370,I639396,);
and I_37431 (I639404,I639396,I171391);
DFFARX1 I_37432 (I639404,I3035,I639370,I639353,);
DFFARX1 I_37433 (I171397,I3035,I639370,I639444,);
not I_37434 (I639452,I171379);
not I_37435 (I639469,I171400);
nand I_37436 (I639486,I639469,I639452);
nor I_37437 (I639341,I639444,I639486);
DFFARX1 I_37438 (I639486,I3035,I639370,I639526,);
not I_37439 (I639362,I639526);
not I_37440 (I639548,I171403);
nand I_37441 (I639565,I639469,I639548);
DFFARX1 I_37442 (I639565,I3035,I639370,I639591,);
not I_37443 (I639599,I639591);
not I_37444 (I639616,I171394);
nand I_37445 (I639633,I639616,I171382);
and I_37446 (I639650,I639452,I639633);
nor I_37447 (I639667,I639565,I639650);
DFFARX1 I_37448 (I639667,I3035,I639370,I639338,);
DFFARX1 I_37449 (I639650,I3035,I639370,I639359,);
nor I_37450 (I639712,I171394,I171388);
nor I_37451 (I639350,I639565,I639712);
or I_37452 (I639743,I171394,I171388);
nor I_37453 (I639760,I171385,I171379);
DFFARX1 I_37454 (I639760,I3035,I639370,I639786,);
not I_37455 (I639794,I639786);
nor I_37456 (I639356,I639794,I639599);
nand I_37457 (I639825,I639794,I639444);
not I_37458 (I639842,I171385);
nand I_37459 (I639859,I639842,I639548);
nand I_37460 (I639876,I639794,I639859);
nand I_37461 (I639347,I639876,I639825);
nand I_37462 (I639344,I639859,I639743);
not I_37463 (I639948,I3042);
DFFARX1 I_37464 (I366061,I3035,I639948,I639974,);
and I_37465 (I639982,I639974,I366049);
DFFARX1 I_37466 (I639982,I3035,I639948,I639931,);
DFFARX1 I_37467 (I366052,I3035,I639948,I640022,);
not I_37468 (I640030,I366046);
not I_37469 (I640047,I366070);
nand I_37470 (I640064,I640047,I640030);
nor I_37471 (I639919,I640022,I640064);
DFFARX1 I_37472 (I640064,I3035,I639948,I640104,);
not I_37473 (I639940,I640104);
not I_37474 (I640126,I366058);
nand I_37475 (I640143,I640047,I640126);
DFFARX1 I_37476 (I640143,I3035,I639948,I640169,);
not I_37477 (I640177,I640169);
not I_37478 (I640194,I366067);
nand I_37479 (I640211,I640194,I366064);
and I_37480 (I640228,I640030,I640211);
nor I_37481 (I640245,I640143,I640228);
DFFARX1 I_37482 (I640245,I3035,I639948,I639916,);
DFFARX1 I_37483 (I640228,I3035,I639948,I639937,);
nor I_37484 (I640290,I366067,I366055);
nor I_37485 (I639928,I640143,I640290);
or I_37486 (I640321,I366067,I366055);
nor I_37487 (I640338,I366046,I366049);
DFFARX1 I_37488 (I640338,I3035,I639948,I640364,);
not I_37489 (I640372,I640364);
nor I_37490 (I639934,I640372,I640177);
nand I_37491 (I640403,I640372,I640022);
not I_37492 (I640420,I366046);
nand I_37493 (I640437,I640420,I640126);
nand I_37494 (I640454,I640372,I640437);
nand I_37495 (I639925,I640454,I640403);
nand I_37496 (I639922,I640437,I640321);
not I_37497 (I640526,I3042);
DFFARX1 I_37498 (I282324,I3035,I640526,I640552,);
and I_37499 (I640560,I640552,I282339);
DFFARX1 I_37500 (I640560,I3035,I640526,I640509,);
DFFARX1 I_37501 (I282330,I3035,I640526,I640600,);
not I_37502 (I640608,I282324);
not I_37503 (I640625,I282342);
nand I_37504 (I640642,I640625,I640608);
nor I_37505 (I640497,I640600,I640642);
DFFARX1 I_37506 (I640642,I3035,I640526,I640682,);
not I_37507 (I640518,I640682);
not I_37508 (I640704,I282333);
nand I_37509 (I640721,I640625,I640704);
DFFARX1 I_37510 (I640721,I3035,I640526,I640747,);
not I_37511 (I640755,I640747);
not I_37512 (I640772,I282345);
nand I_37513 (I640789,I640772,I282321);
and I_37514 (I640806,I640608,I640789);
nor I_37515 (I640823,I640721,I640806);
DFFARX1 I_37516 (I640823,I3035,I640526,I640494,);
DFFARX1 I_37517 (I640806,I3035,I640526,I640515,);
nor I_37518 (I640868,I282345,I282321);
nor I_37519 (I640506,I640721,I640868);
or I_37520 (I640899,I282345,I282321);
nor I_37521 (I640916,I282327,I282336);
DFFARX1 I_37522 (I640916,I3035,I640526,I640942,);
not I_37523 (I640950,I640942);
nor I_37524 (I640512,I640950,I640755);
nand I_37525 (I640981,I640950,I640600);
not I_37526 (I640998,I282327);
nand I_37527 (I641015,I640998,I640704);
nand I_37528 (I641032,I640950,I641015);
nand I_37529 (I640503,I641032,I640981);
nand I_37530 (I640500,I641015,I640899);
not I_37531 (I641104,I3042);
DFFARX1 I_37532 (I245125,I3035,I641104,I641130,);
and I_37533 (I641138,I641130,I245140);
DFFARX1 I_37534 (I641138,I3035,I641104,I641087,);
DFFARX1 I_37535 (I245143,I3035,I641104,I641178,);
not I_37536 (I641186,I245137);
not I_37537 (I641203,I245152);
nand I_37538 (I641220,I641203,I641186);
nor I_37539 (I641075,I641178,I641220);
DFFARX1 I_37540 (I641220,I3035,I641104,I641260,);
not I_37541 (I641096,I641260);
not I_37542 (I641282,I245128);
nand I_37543 (I641299,I641203,I641282);
DFFARX1 I_37544 (I641299,I3035,I641104,I641325,);
not I_37545 (I641333,I641325);
not I_37546 (I641350,I245131);
nand I_37547 (I641367,I641350,I245125);
and I_37548 (I641384,I641186,I641367);
nor I_37549 (I641401,I641299,I641384);
DFFARX1 I_37550 (I641401,I3035,I641104,I641072,);
DFFARX1 I_37551 (I641384,I3035,I641104,I641093,);
nor I_37552 (I641446,I245131,I245134);
nor I_37553 (I641084,I641299,I641446);
or I_37554 (I641477,I245131,I245134);
nor I_37555 (I641494,I245149,I245146);
DFFARX1 I_37556 (I641494,I3035,I641104,I641520,);
not I_37557 (I641528,I641520);
nor I_37558 (I641090,I641528,I641333);
nand I_37559 (I641559,I641528,I641178);
not I_37560 (I641576,I245149);
nand I_37561 (I641593,I641576,I641282);
nand I_37562 (I641610,I641528,I641593);
nand I_37563 (I641081,I641610,I641559);
nand I_37564 (I641078,I641593,I641477);
not I_37565 (I641682,I3042);
DFFARX1 I_37566 (I181419,I3035,I641682,I641708,);
and I_37567 (I641716,I641708,I181404);
DFFARX1 I_37568 (I641716,I3035,I641682,I641665,);
DFFARX1 I_37569 (I181410,I3035,I641682,I641756,);
not I_37570 (I641764,I181392);
not I_37571 (I641781,I181413);
nand I_37572 (I641798,I641781,I641764);
nor I_37573 (I641653,I641756,I641798);
DFFARX1 I_37574 (I641798,I3035,I641682,I641838,);
not I_37575 (I641674,I641838);
not I_37576 (I641860,I181416);
nand I_37577 (I641877,I641781,I641860);
DFFARX1 I_37578 (I641877,I3035,I641682,I641903,);
not I_37579 (I641911,I641903);
not I_37580 (I641928,I181407);
nand I_37581 (I641945,I641928,I181395);
and I_37582 (I641962,I641764,I641945);
nor I_37583 (I641979,I641877,I641962);
DFFARX1 I_37584 (I641979,I3035,I641682,I641650,);
DFFARX1 I_37585 (I641962,I3035,I641682,I641671,);
nor I_37586 (I642024,I181407,I181401);
nor I_37587 (I641662,I641877,I642024);
or I_37588 (I642055,I181407,I181401);
nor I_37589 (I642072,I181398,I181392);
DFFARX1 I_37590 (I642072,I3035,I641682,I642098,);
not I_37591 (I642106,I642098);
nor I_37592 (I641668,I642106,I641911);
nand I_37593 (I642137,I642106,I641756);
not I_37594 (I642154,I181398);
nand I_37595 (I642171,I642154,I641860);
nand I_37596 (I642188,I642106,I642171);
nand I_37597 (I641659,I642188,I642137);
nand I_37598 (I641656,I642171,I642055);
not I_37599 (I642260,I3042);
DFFARX1 I_37600 (I556585,I3035,I642260,I642286,);
and I_37601 (I642294,I642286,I556582);
DFFARX1 I_37602 (I642294,I3035,I642260,I642243,);
DFFARX1 I_37603 (I556588,I3035,I642260,I642334,);
not I_37604 (I642342,I556591);
not I_37605 (I642359,I556585);
nand I_37606 (I642376,I642359,I642342);
nor I_37607 (I642231,I642334,I642376);
DFFARX1 I_37608 (I642376,I3035,I642260,I642416,);
not I_37609 (I642252,I642416);
not I_37610 (I642438,I556600);
nand I_37611 (I642455,I642359,I642438);
DFFARX1 I_37612 (I642455,I3035,I642260,I642481,);
not I_37613 (I642489,I642481);
not I_37614 (I642506,I556597);
nand I_37615 (I642523,I642506,I556603);
and I_37616 (I642540,I642342,I642523);
nor I_37617 (I642557,I642455,I642540);
DFFARX1 I_37618 (I642557,I3035,I642260,I642228,);
DFFARX1 I_37619 (I642540,I3035,I642260,I642249,);
nor I_37620 (I642602,I556597,I556582);
nor I_37621 (I642240,I642455,I642602);
or I_37622 (I642633,I556597,I556582);
nor I_37623 (I642650,I556594,I556588);
DFFARX1 I_37624 (I642650,I3035,I642260,I642676,);
not I_37625 (I642684,I642676);
nor I_37626 (I642246,I642684,I642489);
nand I_37627 (I642715,I642684,I642334);
not I_37628 (I642732,I556594);
nand I_37629 (I642749,I642732,I642438);
nand I_37630 (I642766,I642684,I642749);
nand I_37631 (I642237,I642766,I642715);
nand I_37632 (I642234,I642749,I642633);
not I_37633 (I642838,I3042);
DFFARX1 I_37634 (I141969,I3035,I642838,I642864,);
and I_37635 (I642872,I642864,I141972);
DFFARX1 I_37636 (I642872,I3035,I642838,I642821,);
DFFARX1 I_37637 (I141972,I3035,I642838,I642912,);
not I_37638 (I642920,I141987);
not I_37639 (I642937,I141993);
nand I_37640 (I642954,I642937,I642920);
nor I_37641 (I642809,I642912,I642954);
DFFARX1 I_37642 (I642954,I3035,I642838,I642994,);
not I_37643 (I642830,I642994);
not I_37644 (I643016,I141981);
nand I_37645 (I643033,I642937,I643016);
DFFARX1 I_37646 (I643033,I3035,I642838,I643059,);
not I_37647 (I643067,I643059);
not I_37648 (I643084,I141978);
nand I_37649 (I643101,I643084,I141975);
and I_37650 (I643118,I642920,I643101);
nor I_37651 (I643135,I643033,I643118);
DFFARX1 I_37652 (I643135,I3035,I642838,I642806,);
DFFARX1 I_37653 (I643118,I3035,I642838,I642827,);
nor I_37654 (I643180,I141978,I141969);
nor I_37655 (I642818,I643033,I643180);
or I_37656 (I643211,I141978,I141969);
nor I_37657 (I643228,I141984,I141990);
DFFARX1 I_37658 (I643228,I3035,I642838,I643254,);
not I_37659 (I643262,I643254);
nor I_37660 (I642824,I643262,I643067);
nand I_37661 (I643293,I643262,I642912);
not I_37662 (I643310,I141984);
nand I_37663 (I643327,I643310,I643016);
nand I_37664 (I643344,I643262,I643327);
nand I_37665 (I642815,I643344,I643293);
nand I_37666 (I642812,I643327,I643211);
not I_37667 (I643416,I3042);
DFFARX1 I_37668 (I314619,I3035,I643416,I643442,);
and I_37669 (I643450,I643442,I314607);
DFFARX1 I_37670 (I643450,I3035,I643416,I643399,);
DFFARX1 I_37671 (I314622,I3035,I643416,I643490,);
not I_37672 (I643498,I314613);
not I_37673 (I643515,I314604);
nand I_37674 (I643532,I643515,I643498);
nor I_37675 (I643387,I643490,I643532);
DFFARX1 I_37676 (I643532,I3035,I643416,I643572,);
not I_37677 (I643408,I643572);
not I_37678 (I643594,I314610);
nand I_37679 (I643611,I643515,I643594);
DFFARX1 I_37680 (I643611,I3035,I643416,I643637,);
not I_37681 (I643645,I643637);
not I_37682 (I643662,I314625);
nand I_37683 (I643679,I643662,I314628);
and I_37684 (I643696,I643498,I643679);
nor I_37685 (I643713,I643611,I643696);
DFFARX1 I_37686 (I643713,I3035,I643416,I643384,);
DFFARX1 I_37687 (I643696,I3035,I643416,I643405,);
nor I_37688 (I643758,I314625,I314604);
nor I_37689 (I643396,I643611,I643758);
or I_37690 (I643789,I314625,I314604);
nor I_37691 (I643806,I314616,I314607);
DFFARX1 I_37692 (I643806,I3035,I643416,I643832,);
not I_37693 (I643840,I643832);
nor I_37694 (I643402,I643840,I643645);
nand I_37695 (I643871,I643840,I643490);
not I_37696 (I643888,I314616);
nand I_37697 (I643905,I643888,I643594);
nand I_37698 (I643922,I643840,I643905);
nand I_37699 (I643393,I643922,I643871);
nand I_37700 (I643390,I643905,I643789);
not I_37701 (I643994,I3042);
DFFARX1 I_37702 (I492226,I3035,I643994,I644020,);
and I_37703 (I644028,I644020,I492220);
DFFARX1 I_37704 (I644028,I3035,I643994,I643977,);
DFFARX1 I_37705 (I492238,I3035,I643994,I644068,);
not I_37706 (I644076,I492229);
not I_37707 (I644093,I492241);
nand I_37708 (I644110,I644093,I644076);
nor I_37709 (I643965,I644068,I644110);
DFFARX1 I_37710 (I644110,I3035,I643994,I644150,);
not I_37711 (I643986,I644150);
not I_37712 (I644172,I492247);
nand I_37713 (I644189,I644093,I644172);
DFFARX1 I_37714 (I644189,I3035,I643994,I644215,);
not I_37715 (I644223,I644215);
not I_37716 (I644240,I492223);
nand I_37717 (I644257,I644240,I492244);
and I_37718 (I644274,I644076,I644257);
nor I_37719 (I644291,I644189,I644274);
DFFARX1 I_37720 (I644291,I3035,I643994,I643962,);
DFFARX1 I_37721 (I644274,I3035,I643994,I643983,);
nor I_37722 (I644336,I492223,I492235);
nor I_37723 (I643974,I644189,I644336);
or I_37724 (I644367,I492223,I492235);
nor I_37725 (I644384,I492220,I492232);
DFFARX1 I_37726 (I644384,I3035,I643994,I644410,);
not I_37727 (I644418,I644410);
nor I_37728 (I643980,I644418,I644223);
nand I_37729 (I644449,I644418,I644068);
not I_37730 (I644466,I492220);
nand I_37731 (I644483,I644466,I644172);
nand I_37732 (I644500,I644418,I644483);
nand I_37733 (I643971,I644500,I644449);
nand I_37734 (I643968,I644483,I644367);
not I_37735 (I644572,I3042);
DFFARX1 I_37736 (I229349,I3035,I644572,I644598,);
and I_37737 (I644606,I644598,I229364);
DFFARX1 I_37738 (I644606,I3035,I644572,I644555,);
DFFARX1 I_37739 (I229367,I3035,I644572,I644646,);
not I_37740 (I644654,I229361);
not I_37741 (I644671,I229376);
nand I_37742 (I644688,I644671,I644654);
nor I_37743 (I644543,I644646,I644688);
DFFARX1 I_37744 (I644688,I3035,I644572,I644728,);
not I_37745 (I644564,I644728);
not I_37746 (I644750,I229352);
nand I_37747 (I644767,I644671,I644750);
DFFARX1 I_37748 (I644767,I3035,I644572,I644793,);
not I_37749 (I644801,I644793);
not I_37750 (I644818,I229355);
nand I_37751 (I644835,I644818,I229349);
and I_37752 (I644852,I644654,I644835);
nor I_37753 (I644869,I644767,I644852);
DFFARX1 I_37754 (I644869,I3035,I644572,I644540,);
DFFARX1 I_37755 (I644852,I3035,I644572,I644561,);
nor I_37756 (I644914,I229355,I229358);
nor I_37757 (I644552,I644767,I644914);
or I_37758 (I644945,I229355,I229358);
nor I_37759 (I644962,I229373,I229370);
DFFARX1 I_37760 (I644962,I3035,I644572,I644988,);
not I_37761 (I644996,I644988);
nor I_37762 (I644558,I644996,I644801);
nand I_37763 (I645027,I644996,I644646);
not I_37764 (I645044,I229373);
nand I_37765 (I645061,I645044,I644750);
nand I_37766 (I645078,I644996,I645061);
nand I_37767 (I644549,I645078,I645027);
nand I_37768 (I644546,I645061,I644945);
not I_37769 (I645150,I3042);
DFFARX1 I_37770 (I91394,I3035,I645150,I645176,);
and I_37771 (I645184,I645176,I91397);
DFFARX1 I_37772 (I645184,I3035,I645150,I645133,);
DFFARX1 I_37773 (I91397,I3035,I645150,I645224,);
not I_37774 (I645232,I91412);
not I_37775 (I645249,I91418);
nand I_37776 (I645266,I645249,I645232);
nor I_37777 (I645121,I645224,I645266);
DFFARX1 I_37778 (I645266,I3035,I645150,I645306,);
not I_37779 (I645142,I645306);
not I_37780 (I645328,I91406);
nand I_37781 (I645345,I645249,I645328);
DFFARX1 I_37782 (I645345,I3035,I645150,I645371,);
not I_37783 (I645379,I645371);
not I_37784 (I645396,I91403);
nand I_37785 (I645413,I645396,I91400);
and I_37786 (I645430,I645232,I645413);
nor I_37787 (I645447,I645345,I645430);
DFFARX1 I_37788 (I645447,I3035,I645150,I645118,);
DFFARX1 I_37789 (I645430,I3035,I645150,I645139,);
nor I_37790 (I645492,I91403,I91394);
nor I_37791 (I645130,I645345,I645492);
or I_37792 (I645523,I91403,I91394);
nor I_37793 (I645540,I91409,I91415);
DFFARX1 I_37794 (I645540,I3035,I645150,I645566,);
not I_37795 (I645574,I645566);
nor I_37796 (I645136,I645574,I645379);
nand I_37797 (I645605,I645574,I645224);
not I_37798 (I645622,I91409);
nand I_37799 (I645639,I645622,I645328);
nand I_37800 (I645656,I645574,I645639);
nand I_37801 (I645127,I645656,I645605);
nand I_37802 (I645124,I645639,I645523);
not I_37803 (I645728,I3042);
DFFARX1 I_37804 (I464071,I3035,I645728,I645754,);
and I_37805 (I645762,I645754,I464077);
DFFARX1 I_37806 (I645762,I3035,I645728,I645711,);
DFFARX1 I_37807 (I464083,I3035,I645728,I645802,);
not I_37808 (I645810,I464068);
not I_37809 (I645827,I464068);
nand I_37810 (I645844,I645827,I645810);
nor I_37811 (I645699,I645802,I645844);
DFFARX1 I_37812 (I645844,I3035,I645728,I645884,);
not I_37813 (I645720,I645884);
not I_37814 (I645906,I464086);
nand I_37815 (I645923,I645827,I645906);
DFFARX1 I_37816 (I645923,I3035,I645728,I645949,);
not I_37817 (I645957,I645949);
not I_37818 (I645974,I464080);
nand I_37819 (I645991,I645974,I464071);
and I_37820 (I646008,I645810,I645991);
nor I_37821 (I646025,I645923,I646008);
DFFARX1 I_37822 (I646025,I3035,I645728,I645696,);
DFFARX1 I_37823 (I646008,I3035,I645728,I645717,);
nor I_37824 (I646070,I464080,I464089);
nor I_37825 (I645708,I645923,I646070);
or I_37826 (I646101,I464080,I464089);
nor I_37827 (I646118,I464074,I464074);
DFFARX1 I_37828 (I646118,I3035,I645728,I646144,);
not I_37829 (I646152,I646144);
nor I_37830 (I645714,I646152,I645957);
nand I_37831 (I646183,I646152,I645802);
not I_37832 (I646200,I464074);
nand I_37833 (I646217,I646200,I645906);
nand I_37834 (I646234,I646152,I646217);
nand I_37835 (I645705,I646234,I646183);
nand I_37836 (I645702,I646217,I646101);
not I_37837 (I646306,I3042);
DFFARX1 I_37838 (I218309,I3035,I646306,I646332,);
and I_37839 (I646340,I646332,I218294);
DFFARX1 I_37840 (I646340,I3035,I646306,I646289,);
DFFARX1 I_37841 (I218300,I3035,I646306,I646380,);
not I_37842 (I646388,I218282);
not I_37843 (I646405,I218303);
nand I_37844 (I646422,I646405,I646388);
nor I_37845 (I646277,I646380,I646422);
DFFARX1 I_37846 (I646422,I3035,I646306,I646462,);
not I_37847 (I646298,I646462);
not I_37848 (I646484,I218306);
nand I_37849 (I646501,I646405,I646484);
DFFARX1 I_37850 (I646501,I3035,I646306,I646527,);
not I_37851 (I646535,I646527);
not I_37852 (I646552,I218297);
nand I_37853 (I646569,I646552,I218285);
and I_37854 (I646586,I646388,I646569);
nor I_37855 (I646603,I646501,I646586);
DFFARX1 I_37856 (I646603,I3035,I646306,I646274,);
DFFARX1 I_37857 (I646586,I3035,I646306,I646295,);
nor I_37858 (I646648,I218297,I218291);
nor I_37859 (I646286,I646501,I646648);
or I_37860 (I646679,I218297,I218291);
nor I_37861 (I646696,I218288,I218282);
DFFARX1 I_37862 (I646696,I3035,I646306,I646722,);
not I_37863 (I646730,I646722);
nor I_37864 (I646292,I646730,I646535);
nand I_37865 (I646761,I646730,I646380);
not I_37866 (I646778,I218288);
nand I_37867 (I646795,I646778,I646484);
nand I_37868 (I646812,I646730,I646795);
nand I_37869 (I646283,I646812,I646761);
nand I_37870 (I646280,I646795,I646679);
not I_37871 (I646884,I3042);
DFFARX1 I_37872 (I706175,I3035,I646884,I646910,);
and I_37873 (I646918,I646910,I706157);
DFFARX1 I_37874 (I646918,I3035,I646884,I646867,);
DFFARX1 I_37875 (I706148,I3035,I646884,I646958,);
not I_37876 (I646966,I706163);
not I_37877 (I646983,I706151);
nand I_37878 (I647000,I646983,I646966);
nor I_37879 (I646855,I646958,I647000);
DFFARX1 I_37880 (I647000,I3035,I646884,I647040,);
not I_37881 (I646876,I647040);
not I_37882 (I647062,I706160);
nand I_37883 (I647079,I646983,I647062);
DFFARX1 I_37884 (I647079,I3035,I646884,I647105,);
not I_37885 (I647113,I647105);
not I_37886 (I647130,I706169);
nand I_37887 (I647147,I647130,I706148);
and I_37888 (I647164,I646966,I647147);
nor I_37889 (I647181,I647079,I647164);
DFFARX1 I_37890 (I647181,I3035,I646884,I646852,);
DFFARX1 I_37891 (I647164,I3035,I646884,I646873,);
nor I_37892 (I647226,I706169,I706172);
nor I_37893 (I646864,I647079,I647226);
or I_37894 (I647257,I706169,I706172);
nor I_37895 (I647274,I706166,I706154);
DFFARX1 I_37896 (I647274,I3035,I646884,I647300,);
not I_37897 (I647308,I647300);
nor I_37898 (I646870,I647308,I647113);
nand I_37899 (I647339,I647308,I646958);
not I_37900 (I647356,I706166);
nand I_37901 (I647373,I647356,I647062);
nand I_37902 (I647390,I647308,I647373);
nand I_37903 (I646861,I647390,I647339);
nand I_37904 (I646858,I647373,I647257);
not I_37905 (I647462,I3042);
DFFARX1 I_37906 (I211970,I3035,I647462,I647488,);
nand I_37907 (I647496,I647488,I211973);
DFFARX1 I_37908 (I211967,I3035,I647462,I647522,);
DFFARX1 I_37909 (I647522,I3035,I647462,I647539,);
not I_37910 (I647454,I647539);
not I_37911 (I647561,I211976);
nor I_37912 (I647578,I211976,I211961);
not I_37913 (I647595,I211985);
nand I_37914 (I647612,I647561,I647595);
nor I_37915 (I647629,I211985,I211976);
and I_37916 (I647433,I647629,I647496);
not I_37917 (I647660,I211964);
nand I_37918 (I647677,I647660,I211982);
nor I_37919 (I647694,I211964,I211958);
not I_37920 (I647711,I647694);
nand I_37921 (I647436,I647578,I647711);
DFFARX1 I_37922 (I647694,I3035,I647462,I647451,);
nor I_37923 (I647756,I211979,I211985);
nor I_37924 (I647773,I647756,I211961);
and I_37925 (I647790,I647773,I647677);
DFFARX1 I_37926 (I647790,I3035,I647462,I647448,);
nor I_37927 (I647445,I647756,I647612);
or I_37928 (I647442,I647694,I647756);
nor I_37929 (I647849,I211979,I211958);
DFFARX1 I_37930 (I647849,I3035,I647462,I647875,);
not I_37931 (I647883,I647875);
nand I_37932 (I647900,I647883,I647561);
nor I_37933 (I647917,I647900,I211961);
DFFARX1 I_37934 (I647917,I3035,I647462,I647430,);
nor I_37935 (I647948,I647883,I647612);
nor I_37936 (I647439,I647756,I647948);
not I_37937 (I648006,I3042);
DFFARX1 I_37938 (I157162,I3035,I648006,I648032,);
nand I_37939 (I648040,I648032,I157165);
DFFARX1 I_37940 (I157159,I3035,I648006,I648066,);
DFFARX1 I_37941 (I648066,I3035,I648006,I648083,);
not I_37942 (I647998,I648083);
not I_37943 (I648105,I157168);
nor I_37944 (I648122,I157168,I157153);
not I_37945 (I648139,I157177);
nand I_37946 (I648156,I648105,I648139);
nor I_37947 (I648173,I157177,I157168);
and I_37948 (I647977,I648173,I648040);
not I_37949 (I648204,I157156);
nand I_37950 (I648221,I648204,I157174);
nor I_37951 (I648238,I157156,I157150);
not I_37952 (I648255,I648238);
nand I_37953 (I647980,I648122,I648255);
DFFARX1 I_37954 (I648238,I3035,I648006,I647995,);
nor I_37955 (I648300,I157171,I157177);
nor I_37956 (I648317,I648300,I157153);
and I_37957 (I648334,I648317,I648221);
DFFARX1 I_37958 (I648334,I3035,I648006,I647992,);
nor I_37959 (I647989,I648300,I648156);
or I_37960 (I647986,I648238,I648300);
nor I_37961 (I648393,I157171,I157150);
DFFARX1 I_37962 (I648393,I3035,I648006,I648419,);
not I_37963 (I648427,I648419);
nand I_37964 (I648444,I648427,I648105);
nor I_37965 (I648461,I648444,I157153);
DFFARX1 I_37966 (I648461,I3035,I648006,I647974,);
nor I_37967 (I648492,I648427,I648156);
nor I_37968 (I647983,I648300,I648492);
not I_37969 (I648550,I3042);
DFFARX1 I_37970 (I223037,I3035,I648550,I648576,);
nand I_37971 (I648584,I648576,I223040);
DFFARX1 I_37972 (I223034,I3035,I648550,I648610,);
DFFARX1 I_37973 (I648610,I3035,I648550,I648627,);
not I_37974 (I648542,I648627);
not I_37975 (I648649,I223043);
nor I_37976 (I648666,I223043,I223028);
not I_37977 (I648683,I223052);
nand I_37978 (I648700,I648649,I648683);
nor I_37979 (I648717,I223052,I223043);
and I_37980 (I648521,I648717,I648584);
not I_37981 (I648748,I223031);
nand I_37982 (I648765,I648748,I223049);
nor I_37983 (I648782,I223031,I223025);
not I_37984 (I648799,I648782);
nand I_37985 (I648524,I648666,I648799);
DFFARX1 I_37986 (I648782,I3035,I648550,I648539,);
nor I_37987 (I648844,I223046,I223052);
nor I_37988 (I648861,I648844,I223028);
and I_37989 (I648878,I648861,I648765);
DFFARX1 I_37990 (I648878,I3035,I648550,I648536,);
nor I_37991 (I648533,I648844,I648700);
or I_37992 (I648530,I648782,I648844);
nor I_37993 (I648937,I223046,I223025);
DFFARX1 I_37994 (I648937,I3035,I648550,I648963,);
not I_37995 (I648971,I648963);
nand I_37996 (I648988,I648971,I648649);
nor I_37997 (I649005,I648988,I223028);
DFFARX1 I_37998 (I649005,I3035,I648550,I648518,);
nor I_37999 (I649036,I648971,I648700);
nor I_38000 (I648527,I648844,I649036);
not I_38001 (I649094,I3042);
DFFARX1 I_38002 (I541316,I3035,I649094,I649120,);
nand I_38003 (I649128,I649120,I541316);
DFFARX1 I_38004 (I541328,I3035,I649094,I649154,);
DFFARX1 I_38005 (I649154,I3035,I649094,I649171,);
not I_38006 (I649086,I649171);
not I_38007 (I649193,I541322);
nor I_38008 (I649210,I541322,I541343);
not I_38009 (I649227,I541331);
nand I_38010 (I649244,I649193,I649227);
nor I_38011 (I649261,I541331,I541322);
and I_38012 (I649065,I649261,I649128);
not I_38013 (I649292,I541325);
nand I_38014 (I649309,I649292,I541340);
nor I_38015 (I649326,I541325,I541334);
not I_38016 (I649343,I649326);
nand I_38017 (I649068,I649210,I649343);
DFFARX1 I_38018 (I649326,I3035,I649094,I649083,);
nor I_38019 (I649388,I541337,I541331);
nor I_38020 (I649405,I649388,I541343);
and I_38021 (I649422,I649405,I649309);
DFFARX1 I_38022 (I649422,I3035,I649094,I649080,);
nor I_38023 (I649077,I649388,I649244);
or I_38024 (I649074,I649326,I649388);
nor I_38025 (I649481,I541337,I541319);
DFFARX1 I_38026 (I649481,I3035,I649094,I649507,);
not I_38027 (I649515,I649507);
nand I_38028 (I649532,I649515,I649193);
nor I_38029 (I649549,I649532,I541343);
DFFARX1 I_38030 (I649549,I3035,I649094,I649062,);
nor I_38031 (I649580,I649515,I649244);
nor I_38032 (I649071,I649388,I649580);
not I_38033 (I649638,I3042);
DFFARX1 I_38034 (I39973,I3035,I649638,I649664,);
nand I_38035 (I649672,I649664,I39955);
DFFARX1 I_38036 (I39952,I3035,I649638,I649698,);
DFFARX1 I_38037 (I649698,I3035,I649638,I649715,);
not I_38038 (I649630,I649715);
not I_38039 (I649737,I39970);
nor I_38040 (I649754,I39970,I39964);
not I_38041 (I649771,I39952);
nand I_38042 (I649788,I649737,I649771);
nor I_38043 (I649805,I39952,I39970);
and I_38044 (I649609,I649805,I649672);
not I_38045 (I649836,I39961);
nand I_38046 (I649853,I649836,I39967);
nor I_38047 (I649870,I39961,I39955);
not I_38048 (I649887,I649870);
nand I_38049 (I649612,I649754,I649887);
DFFARX1 I_38050 (I649870,I3035,I649638,I649627,);
nor I_38051 (I649932,I39958,I39952);
nor I_38052 (I649949,I649932,I39964);
and I_38053 (I649966,I649949,I649853);
DFFARX1 I_38054 (I649966,I3035,I649638,I649624,);
nor I_38055 (I649621,I649932,I649788);
or I_38056 (I649618,I649870,I649932);
nor I_38057 (I650025,I39958,I39976);
DFFARX1 I_38058 (I650025,I3035,I649638,I650051,);
not I_38059 (I650059,I650051);
nand I_38060 (I650076,I650059,I649737);
nor I_38061 (I650093,I650076,I39964);
DFFARX1 I_38062 (I650093,I3035,I649638,I649606,);
nor I_38063 (I650124,I650059,I649788);
nor I_38064 (I649615,I649932,I650124);
not I_38065 (I650182,I3042);
DFFARX1 I_38066 (I328497,I3035,I650182,I650208,);
nand I_38067 (I650216,I650208,I328485);
DFFARX1 I_38068 (I328491,I3035,I650182,I650242,);
DFFARX1 I_38069 (I650242,I3035,I650182,I650259,);
not I_38070 (I650174,I650259);
not I_38071 (I650281,I328476);
nor I_38072 (I650298,I328476,I328488);
not I_38073 (I650315,I328479);
nand I_38074 (I650332,I650281,I650315);
nor I_38075 (I650349,I328479,I328476);
and I_38076 (I650153,I650349,I650216);
not I_38077 (I650380,I328494);
nand I_38078 (I650397,I650380,I328476);
nor I_38079 (I650414,I328494,I328500);
not I_38080 (I650431,I650414);
nand I_38081 (I650156,I650298,I650431);
DFFARX1 I_38082 (I650414,I3035,I650182,I650171,);
nor I_38083 (I650476,I328482,I328479);
nor I_38084 (I650493,I650476,I328488);
and I_38085 (I650510,I650493,I650397);
DFFARX1 I_38086 (I650510,I3035,I650182,I650168,);
nor I_38087 (I650165,I650476,I650332);
or I_38088 (I650162,I650414,I650476);
nor I_38089 (I650569,I328482,I328479);
DFFARX1 I_38090 (I650569,I3035,I650182,I650595,);
not I_38091 (I650603,I650595);
nand I_38092 (I650620,I650603,I650281);
nor I_38093 (I650637,I650620,I328488);
DFFARX1 I_38094 (I650637,I3035,I650182,I650150,);
nor I_38095 (I650668,I650603,I650332);
nor I_38096 (I650159,I650476,I650668);
not I_38097 (I650726,I3042);
DFFARX1 I_38098 (I677121,I3035,I650726,I650752,);
nand I_38099 (I650760,I650752,I677130);
DFFARX1 I_38100 (I677133,I3035,I650726,I650786,);
DFFARX1 I_38101 (I650786,I3035,I650726,I650803,);
not I_38102 (I650718,I650803);
not I_38103 (I650825,I677127);
nor I_38104 (I650842,I677127,I677124);
not I_38105 (I650859,I677118);
nand I_38106 (I650876,I650825,I650859);
nor I_38107 (I650893,I677118,I677127);
and I_38108 (I650697,I650893,I650760);
not I_38109 (I650924,I677115);
nand I_38110 (I650941,I650924,I677112);
nor I_38111 (I650958,I677115,I677112);
not I_38112 (I650975,I650958);
nand I_38113 (I650700,I650842,I650975);
DFFARX1 I_38114 (I650958,I3035,I650726,I650715,);
nor I_38115 (I651020,I677115,I677118);
nor I_38116 (I651037,I651020,I677124);
and I_38117 (I651054,I651037,I650941);
DFFARX1 I_38118 (I651054,I3035,I650726,I650712,);
nor I_38119 (I650709,I651020,I650876);
or I_38120 (I650706,I650958,I651020);
nor I_38121 (I651113,I677115,I677136);
DFFARX1 I_38122 (I651113,I3035,I650726,I651139,);
not I_38123 (I651147,I651139);
nand I_38124 (I651164,I651147,I650825);
nor I_38125 (I651181,I651164,I677124);
DFFARX1 I_38126 (I651181,I3035,I650726,I650694,);
nor I_38127 (I651212,I651147,I650876);
nor I_38128 (I650703,I651020,I651212);
not I_38129 (I651270,I3042);
DFFARX1 I_38130 (I609884,I3035,I651270,I651296,);
nand I_38131 (I651304,I651296,I609863);
DFFARX1 I_38132 (I609860,I3035,I651270,I651330,);
DFFARX1 I_38133 (I651330,I3035,I651270,I651347,);
not I_38134 (I651262,I651347);
not I_38135 (I651369,I609872);
nor I_38136 (I651386,I609872,I609881);
not I_38137 (I651403,I609869);
nand I_38138 (I651420,I651369,I651403);
nor I_38139 (I651437,I609869,I609872);
and I_38140 (I651241,I651437,I651304);
not I_38141 (I651468,I609878);
nand I_38142 (I651485,I651468,I609875);
nor I_38143 (I651502,I609878,I609860);
not I_38144 (I651519,I651502);
nand I_38145 (I651244,I651386,I651519);
DFFARX1 I_38146 (I651502,I3035,I651270,I651259,);
nor I_38147 (I651564,I609863,I609869);
nor I_38148 (I651581,I651564,I609881);
and I_38149 (I651598,I651581,I651485);
DFFARX1 I_38150 (I651598,I3035,I651270,I651256,);
nor I_38151 (I651253,I651564,I651420);
or I_38152 (I651250,I651502,I651564);
nor I_38153 (I651657,I609863,I609866);
DFFARX1 I_38154 (I651657,I3035,I651270,I651683,);
not I_38155 (I651691,I651683);
nand I_38156 (I651708,I651691,I651369);
nor I_38157 (I651725,I651708,I609881);
DFFARX1 I_38158 (I651725,I3035,I651270,I651238,);
nor I_38159 (I651756,I651691,I651420);
nor I_38160 (I651247,I651564,I651756);
not I_38161 (I651814,I3042);
DFFARX1 I_38162 (I484468,I3035,I651814,I651840,);
nand I_38163 (I651848,I651840,I484468);
DFFARX1 I_38164 (I484480,I3035,I651814,I651874,);
DFFARX1 I_38165 (I651874,I3035,I651814,I651891,);
not I_38166 (I651806,I651891);
not I_38167 (I651913,I484474);
nor I_38168 (I651930,I484474,I484495);
not I_38169 (I651947,I484483);
nand I_38170 (I651964,I651913,I651947);
nor I_38171 (I651981,I484483,I484474);
and I_38172 (I651785,I651981,I651848);
not I_38173 (I652012,I484477);
nand I_38174 (I652029,I652012,I484492);
nor I_38175 (I652046,I484477,I484486);
not I_38176 (I652063,I652046);
nand I_38177 (I651788,I651930,I652063);
DFFARX1 I_38178 (I652046,I3035,I651814,I651803,);
nor I_38179 (I652108,I484489,I484483);
nor I_38180 (I652125,I652108,I484495);
and I_38181 (I652142,I652125,I652029);
DFFARX1 I_38182 (I652142,I3035,I651814,I651800,);
nor I_38183 (I651797,I652108,I651964);
or I_38184 (I651794,I652046,I652108);
nor I_38185 (I652201,I484489,I484471);
DFFARX1 I_38186 (I652201,I3035,I651814,I652227,);
not I_38187 (I652235,I652227);
nand I_38188 (I652252,I652235,I651913);
nor I_38189 (I652269,I652252,I484495);
DFFARX1 I_38190 (I652269,I3035,I651814,I651782,);
nor I_38191 (I652300,I652235,I651964);
nor I_38192 (I651791,I652108,I652300);
not I_38193 (I652358,I3042);
DFFARX1 I_38194 (I229917,I3035,I652358,I652384,);
nand I_38195 (I652392,I652384,I229914);
DFFARX1 I_38196 (I229893,I3035,I652358,I652418,);
DFFARX1 I_38197 (I652418,I3035,I652358,I652435,);
not I_38198 (I652350,I652435);
not I_38199 (I652457,I229908);
nor I_38200 (I652474,I229908,I229911);
not I_38201 (I652491,I229902);
nand I_38202 (I652508,I652457,I652491);
nor I_38203 (I652525,I229902,I229908);
and I_38204 (I652329,I652525,I652392);
not I_38205 (I652556,I229899);
nand I_38206 (I652573,I652556,I229920);
nor I_38207 (I652590,I229899,I229896);
not I_38208 (I652607,I652590);
nand I_38209 (I652332,I652474,I652607);
DFFARX1 I_38210 (I652590,I3035,I652358,I652347,);
nor I_38211 (I652652,I229905,I229902);
nor I_38212 (I652669,I652652,I229911);
and I_38213 (I652686,I652669,I652573);
DFFARX1 I_38214 (I652686,I3035,I652358,I652344,);
nor I_38215 (I652341,I652652,I652508);
or I_38216 (I652338,I652590,I652652);
nor I_38217 (I652745,I229905,I229893);
DFFARX1 I_38218 (I652745,I3035,I652358,I652771,);
not I_38219 (I652779,I652771);
nand I_38220 (I652796,I652779,I652457);
nor I_38221 (I652813,I652796,I229911);
DFFARX1 I_38222 (I652813,I3035,I652358,I652326,);
nor I_38223 (I652844,I652779,I652508);
nor I_38224 (I652335,I652652,I652844);
not I_38225 (I652902,I3042);
DFFARX1 I_38226 (I78331,I3035,I652902,I652928,);
nand I_38227 (I652936,I652928,I78304);
DFFARX1 I_38228 (I78322,I3035,I652902,I652962,);
DFFARX1 I_38229 (I652962,I3035,I652902,I652979,);
not I_38230 (I652894,I652979);
not I_38231 (I653001,I78316);
nor I_38232 (I653018,I78316,I78304);
not I_38233 (I653035,I78319);
nand I_38234 (I653052,I653001,I653035);
nor I_38235 (I653069,I78319,I78316);
and I_38236 (I652873,I653069,I652936);
not I_38237 (I653100,I78307);
nand I_38238 (I653117,I653100,I78325);
nor I_38239 (I653134,I78307,I78328);
not I_38240 (I653151,I653134);
nand I_38241 (I652876,I653018,I653151);
DFFARX1 I_38242 (I653134,I3035,I652902,I652891,);
nor I_38243 (I653196,I78310,I78319);
nor I_38244 (I653213,I653196,I78304);
and I_38245 (I653230,I653213,I653117);
DFFARX1 I_38246 (I653230,I3035,I652902,I652888,);
nor I_38247 (I652885,I653196,I653052);
or I_38248 (I652882,I653134,I653196);
nor I_38249 (I653289,I78310,I78313);
DFFARX1 I_38250 (I653289,I3035,I652902,I653315,);
not I_38251 (I653323,I653315);
nand I_38252 (I653340,I653323,I653001);
nor I_38253 (I653357,I653340,I78304);
DFFARX1 I_38254 (I653357,I3035,I652902,I652870,);
nor I_38255 (I653388,I653323,I653052);
nor I_38256 (I652879,I653196,I653388);
not I_38257 (I653446,I3042);
DFFARX1 I_38258 (I621444,I3035,I653446,I653472,);
nand I_38259 (I653480,I653472,I621423);
DFFARX1 I_38260 (I621420,I3035,I653446,I653506,);
DFFARX1 I_38261 (I653506,I3035,I653446,I653523,);
not I_38262 (I653438,I653523);
not I_38263 (I653545,I621432);
nor I_38264 (I653562,I621432,I621441);
not I_38265 (I653579,I621429);
nand I_38266 (I653596,I653545,I653579);
nor I_38267 (I653613,I621429,I621432);
and I_38268 (I653417,I653613,I653480);
not I_38269 (I653644,I621438);
nand I_38270 (I653661,I653644,I621435);
nor I_38271 (I653678,I621438,I621420);
not I_38272 (I653695,I653678);
nand I_38273 (I653420,I653562,I653695);
DFFARX1 I_38274 (I653678,I3035,I653446,I653435,);
nor I_38275 (I653740,I621423,I621429);
nor I_38276 (I653757,I653740,I621441);
and I_38277 (I653774,I653757,I653661);
DFFARX1 I_38278 (I653774,I3035,I653446,I653432,);
nor I_38279 (I653429,I653740,I653596);
or I_38280 (I653426,I653678,I653740);
nor I_38281 (I653833,I621423,I621426);
DFFARX1 I_38282 (I653833,I3035,I653446,I653859,);
not I_38283 (I653867,I653859);
nand I_38284 (I653884,I653867,I653545);
nor I_38285 (I653901,I653884,I621441);
DFFARX1 I_38286 (I653901,I3035,I653446,I653414,);
nor I_38287 (I653932,I653867,I653596);
nor I_38288 (I653423,I653740,I653932);
not I_38289 (I653990,I3042);
DFFARX1 I_38290 (I233181,I3035,I653990,I654016,);
nand I_38291 (I654024,I654016,I233178);
DFFARX1 I_38292 (I233157,I3035,I653990,I654050,);
DFFARX1 I_38293 (I654050,I3035,I653990,I654067,);
not I_38294 (I653982,I654067);
not I_38295 (I654089,I233172);
nor I_38296 (I654106,I233172,I233175);
not I_38297 (I654123,I233166);
nand I_38298 (I654140,I654089,I654123);
nor I_38299 (I654157,I233166,I233172);
and I_38300 (I653961,I654157,I654024);
not I_38301 (I654188,I233163);
nand I_38302 (I654205,I654188,I233184);
nor I_38303 (I654222,I233163,I233160);
not I_38304 (I654239,I654222);
nand I_38305 (I653964,I654106,I654239);
DFFARX1 I_38306 (I654222,I3035,I653990,I653979,);
nor I_38307 (I654284,I233169,I233166);
nor I_38308 (I654301,I654284,I233175);
and I_38309 (I654318,I654301,I654205);
DFFARX1 I_38310 (I654318,I3035,I653990,I653976,);
nor I_38311 (I653973,I654284,I654140);
or I_38312 (I653970,I654222,I654284);
nor I_38313 (I654377,I233169,I233157);
DFFARX1 I_38314 (I654377,I3035,I653990,I654403,);
not I_38315 (I654411,I654403);
nand I_38316 (I654428,I654411,I654089);
nor I_38317 (I654445,I654428,I233175);
DFFARX1 I_38318 (I654445,I3035,I653990,I653958,);
nor I_38319 (I654476,I654411,I654140);
nor I_38320 (I653967,I654284,I654476);
not I_38321 (I654534,I3042);
DFFARX1 I_38322 (I677699,I3035,I654534,I654560,);
nand I_38323 (I654568,I654560,I677708);
DFFARX1 I_38324 (I677711,I3035,I654534,I654594,);
DFFARX1 I_38325 (I654594,I3035,I654534,I654611,);
not I_38326 (I654526,I654611);
not I_38327 (I654633,I677705);
nor I_38328 (I654650,I677705,I677702);
not I_38329 (I654667,I677696);
nand I_38330 (I654684,I654633,I654667);
nor I_38331 (I654701,I677696,I677705);
and I_38332 (I654505,I654701,I654568);
not I_38333 (I654732,I677693);
nand I_38334 (I654749,I654732,I677690);
nor I_38335 (I654766,I677693,I677690);
not I_38336 (I654783,I654766);
nand I_38337 (I654508,I654650,I654783);
DFFARX1 I_38338 (I654766,I3035,I654534,I654523,);
nor I_38339 (I654828,I677693,I677696);
nor I_38340 (I654845,I654828,I677702);
and I_38341 (I654862,I654845,I654749);
DFFARX1 I_38342 (I654862,I3035,I654534,I654520,);
nor I_38343 (I654517,I654828,I654684);
or I_38344 (I654514,I654766,I654828);
nor I_38345 (I654921,I677693,I677714);
DFFARX1 I_38346 (I654921,I3035,I654534,I654947,);
not I_38347 (I654955,I654947);
nand I_38348 (I654972,I654955,I654633);
nor I_38349 (I654989,I654972,I677702);
DFFARX1 I_38350 (I654989,I3035,I654534,I654502,);
nor I_38351 (I655020,I654955,I654684);
nor I_38352 (I654511,I654828,I655020);
not I_38353 (I655078,I3042);
DFFARX1 I_38354 (I673075,I3035,I655078,I655104,);
nand I_38355 (I655112,I655104,I673084);
DFFARX1 I_38356 (I673087,I3035,I655078,I655138,);
DFFARX1 I_38357 (I655138,I3035,I655078,I655155,);
not I_38358 (I655070,I655155);
not I_38359 (I655177,I673081);
nor I_38360 (I655194,I673081,I673078);
not I_38361 (I655211,I673072);
nand I_38362 (I655228,I655177,I655211);
nor I_38363 (I655245,I673072,I673081);
and I_38364 (I655049,I655245,I655112);
not I_38365 (I655276,I673069);
nand I_38366 (I655293,I655276,I673066);
nor I_38367 (I655310,I673069,I673066);
not I_38368 (I655327,I655310);
nand I_38369 (I655052,I655194,I655327);
DFFARX1 I_38370 (I655310,I3035,I655078,I655067,);
nor I_38371 (I655372,I673069,I673072);
nor I_38372 (I655389,I655372,I673078);
and I_38373 (I655406,I655389,I655293);
DFFARX1 I_38374 (I655406,I3035,I655078,I655064,);
nor I_38375 (I655061,I655372,I655228);
or I_38376 (I655058,I655310,I655372);
nor I_38377 (I655465,I673069,I673090);
DFFARX1 I_38378 (I655465,I3035,I655078,I655491,);
not I_38379 (I655499,I655491);
nand I_38380 (I655516,I655499,I655177);
nor I_38381 (I655533,I655516,I673078);
DFFARX1 I_38382 (I655533,I3035,I655078,I655046,);
nor I_38383 (I655564,I655499,I655228);
nor I_38384 (I655055,I655372,I655564);
not I_38385 (I655622,I3042);
DFFARX1 I_38386 (I92593,I3035,I655622,I655648,);
nand I_38387 (I655656,I655648,I92608);
DFFARX1 I_38388 (I92605,I3035,I655622,I655682,);
DFFARX1 I_38389 (I655682,I3035,I655622,I655699,);
not I_38390 (I655614,I655699);
not I_38391 (I655721,I92584);
nor I_38392 (I655738,I92584,I92590);
not I_38393 (I655755,I92596);
nand I_38394 (I655772,I655721,I655755);
nor I_38395 (I655789,I92596,I92584);
and I_38396 (I655593,I655789,I655656);
not I_38397 (I655820,I92602);
nand I_38398 (I655837,I655820,I92584);
nor I_38399 (I655854,I92602,I92587);
not I_38400 (I655871,I655854);
nand I_38401 (I655596,I655738,I655871);
DFFARX1 I_38402 (I655854,I3035,I655622,I655611,);
nor I_38403 (I655916,I92587,I92596);
nor I_38404 (I655933,I655916,I92590);
and I_38405 (I655950,I655933,I655837);
DFFARX1 I_38406 (I655950,I3035,I655622,I655608,);
nor I_38407 (I655605,I655916,I655772);
or I_38408 (I655602,I655854,I655916);
nor I_38409 (I656009,I92587,I92599);
DFFARX1 I_38410 (I656009,I3035,I655622,I656035,);
not I_38411 (I656043,I656035);
nand I_38412 (I656060,I656043,I655721);
nor I_38413 (I656077,I656060,I92590);
DFFARX1 I_38414 (I656077,I3035,I655622,I655590,);
nor I_38415 (I656108,I656043,I655772);
nor I_38416 (I655599,I655916,I656108);
not I_38417 (I656166,I3042);
DFFARX1 I_38418 (I430346,I3035,I656166,I656192,);
nand I_38419 (I656200,I656192,I430340);
DFFARX1 I_38420 (I430343,I3035,I656166,I656226,);
DFFARX1 I_38421 (I656226,I3035,I656166,I656243,);
not I_38422 (I656158,I656243);
not I_38423 (I656265,I430349);
nor I_38424 (I656282,I430349,I430343);
not I_38425 (I656299,I430352);
nand I_38426 (I656316,I656265,I656299);
nor I_38427 (I656333,I430352,I430349);
and I_38428 (I656137,I656333,I656200);
not I_38429 (I656364,I430361);
nand I_38430 (I656381,I656364,I430355);
nor I_38431 (I656398,I430361,I430358);
not I_38432 (I656415,I656398);
nand I_38433 (I656140,I656282,I656415);
DFFARX1 I_38434 (I656398,I3035,I656166,I656155,);
nor I_38435 (I656460,I430340,I430352);
nor I_38436 (I656477,I656460,I430343);
and I_38437 (I656494,I656477,I656381);
DFFARX1 I_38438 (I656494,I3035,I656166,I656152,);
nor I_38439 (I656149,I656460,I656316);
or I_38440 (I656146,I656398,I656460);
nor I_38441 (I656553,I430340,I430346);
DFFARX1 I_38442 (I656553,I3035,I656166,I656579,);
not I_38443 (I656587,I656579);
nand I_38444 (I656604,I656587,I656265);
nor I_38445 (I656621,I656604,I430343);
DFFARX1 I_38446 (I656621,I3035,I656166,I656134,);
nor I_38447 (I656652,I656587,I656316);
nor I_38448 (I656143,I656460,I656652);
not I_38449 (I656710,I3042);
DFFARX1 I_38450 (I151892,I3035,I656710,I656736,);
nand I_38451 (I656744,I656736,I151895);
DFFARX1 I_38452 (I151889,I3035,I656710,I656770,);
DFFARX1 I_38453 (I656770,I3035,I656710,I656787,);
not I_38454 (I656702,I656787);
not I_38455 (I656809,I151898);
nor I_38456 (I656826,I151898,I151883);
not I_38457 (I656843,I151907);
nand I_38458 (I656860,I656809,I656843);
nor I_38459 (I656877,I151907,I151898);
and I_38460 (I656681,I656877,I656744);
not I_38461 (I656908,I151886);
nand I_38462 (I656925,I656908,I151904);
nor I_38463 (I656942,I151886,I151880);
not I_38464 (I656959,I656942);
nand I_38465 (I656684,I656826,I656959);
DFFARX1 I_38466 (I656942,I3035,I656710,I656699,);
nor I_38467 (I657004,I151901,I151907);
nor I_38468 (I657021,I657004,I151883);
and I_38469 (I657038,I657021,I656925);
DFFARX1 I_38470 (I657038,I3035,I656710,I656696,);
nor I_38471 (I656693,I657004,I656860);
or I_38472 (I656690,I656942,I657004);
nor I_38473 (I657097,I151901,I151880);
DFFARX1 I_38474 (I657097,I3035,I656710,I657123,);
not I_38475 (I657131,I657123);
nand I_38476 (I657148,I657131,I656809);
nor I_38477 (I657165,I657148,I151883);
DFFARX1 I_38478 (I657165,I3035,I656710,I656678,);
nor I_38479 (I657196,I657131,I656860);
nor I_38480 (I656687,I657004,I657196);
not I_38481 (I657254,I3042);
DFFARX1 I_38482 (I591388,I3035,I657254,I657280,);
nand I_38483 (I657288,I657280,I591367);
DFFARX1 I_38484 (I591364,I3035,I657254,I657314,);
DFFARX1 I_38485 (I657314,I3035,I657254,I657331,);
not I_38486 (I657246,I657331);
not I_38487 (I657353,I591376);
nor I_38488 (I657370,I591376,I591385);
not I_38489 (I657387,I591373);
nand I_38490 (I657404,I657353,I657387);
nor I_38491 (I657421,I591373,I591376);
and I_38492 (I657225,I657421,I657288);
not I_38493 (I657452,I591382);
nand I_38494 (I657469,I657452,I591379);
nor I_38495 (I657486,I591382,I591364);
not I_38496 (I657503,I657486);
nand I_38497 (I657228,I657370,I657503);
DFFARX1 I_38498 (I657486,I3035,I657254,I657243,);
nor I_38499 (I657548,I591367,I591373);
nor I_38500 (I657565,I657548,I591385);
and I_38501 (I657582,I657565,I657469);
DFFARX1 I_38502 (I657582,I3035,I657254,I657240,);
nor I_38503 (I657237,I657548,I657404);
or I_38504 (I657234,I657486,I657548);
nor I_38505 (I657641,I591367,I591370);
DFFARX1 I_38506 (I657641,I3035,I657254,I657667,);
not I_38507 (I657675,I657667);
nand I_38508 (I657692,I657675,I657353);
nor I_38509 (I657709,I657692,I591385);
DFFARX1 I_38510 (I657709,I3035,I657254,I657222,);
nor I_38511 (I657740,I657675,I657404);
nor I_38512 (I657231,I657548,I657740);
not I_38513 (I657798,I3042);
DFFARX1 I_38514 (I691571,I3035,I657798,I657824,);
nand I_38515 (I657832,I657824,I691580);
DFFARX1 I_38516 (I691583,I3035,I657798,I657858,);
DFFARX1 I_38517 (I657858,I3035,I657798,I657875,);
not I_38518 (I657790,I657875);
not I_38519 (I657897,I691577);
nor I_38520 (I657914,I691577,I691574);
not I_38521 (I657931,I691568);
nand I_38522 (I657948,I657897,I657931);
nor I_38523 (I657965,I691568,I691577);
and I_38524 (I657769,I657965,I657832);
not I_38525 (I657996,I691565);
nand I_38526 (I658013,I657996,I691562);
nor I_38527 (I658030,I691565,I691562);
not I_38528 (I658047,I658030);
nand I_38529 (I657772,I657914,I658047);
DFFARX1 I_38530 (I658030,I3035,I657798,I657787,);
nor I_38531 (I658092,I691565,I691568);
nor I_38532 (I658109,I658092,I691574);
and I_38533 (I658126,I658109,I658013);
DFFARX1 I_38534 (I658126,I3035,I657798,I657784,);
nor I_38535 (I657781,I658092,I657948);
or I_38536 (I657778,I658030,I658092);
nor I_38537 (I658185,I691565,I691586);
DFFARX1 I_38538 (I658185,I3035,I657798,I658211,);
not I_38539 (I658219,I658211);
nand I_38540 (I658236,I658219,I657897);
nor I_38541 (I658253,I658236,I691574);
DFFARX1 I_38542 (I658253,I3035,I657798,I657766,);
nor I_38543 (I658284,I658219,I657948);
nor I_38544 (I657775,I658092,I658284);
not I_38545 (I658342,I3042);
DFFARX1 I_38546 (I440886,I3035,I658342,I658368,);
nand I_38547 (I658376,I658368,I440880);
DFFARX1 I_38548 (I440883,I3035,I658342,I658402,);
DFFARX1 I_38549 (I658402,I3035,I658342,I658419,);
not I_38550 (I658334,I658419);
not I_38551 (I658441,I440889);
nor I_38552 (I658458,I440889,I440883);
not I_38553 (I658475,I440892);
nand I_38554 (I658492,I658441,I658475);
nor I_38555 (I658509,I440892,I440889);
and I_38556 (I658313,I658509,I658376);
not I_38557 (I658540,I440901);
nand I_38558 (I658557,I658540,I440895);
nor I_38559 (I658574,I440901,I440898);
not I_38560 (I658591,I658574);
nand I_38561 (I658316,I658458,I658591);
DFFARX1 I_38562 (I658574,I3035,I658342,I658331,);
nor I_38563 (I658636,I440880,I440892);
nor I_38564 (I658653,I658636,I440883);
and I_38565 (I658670,I658653,I658557);
DFFARX1 I_38566 (I658670,I3035,I658342,I658328,);
nor I_38567 (I658325,I658636,I658492);
or I_38568 (I658322,I658574,I658636);
nor I_38569 (I658729,I440880,I440886);
DFFARX1 I_38570 (I658729,I3035,I658342,I658755,);
not I_38571 (I658763,I658755);
nand I_38572 (I658780,I658763,I658441);
nor I_38573 (I658797,I658780,I440883);
DFFARX1 I_38574 (I658797,I3035,I658342,I658310,);
nor I_38575 (I658828,I658763,I658492);
nor I_38576 (I658319,I658636,I658828);
not I_38577 (I658886,I3042);
DFFARX1 I_38578 (I400151,I3035,I658886,I658912,);
nand I_38579 (I658920,I658912,I400166);
DFFARX1 I_38580 (I400160,I3035,I658886,I658946,);
DFFARX1 I_38581 (I658946,I3035,I658886,I658963,);
not I_38582 (I658878,I658963);
not I_38583 (I658985,I400163);
nor I_38584 (I659002,I400163,I400169);
not I_38585 (I659019,I400151);
nand I_38586 (I659036,I658985,I659019);
nor I_38587 (I659053,I400151,I400163);
and I_38588 (I658857,I659053,I658920);
not I_38589 (I659084,I400148);
nand I_38590 (I659101,I659084,I400154);
nor I_38591 (I659118,I400148,I400148);
not I_38592 (I659135,I659118);
nand I_38593 (I658860,I659002,I659135);
DFFARX1 I_38594 (I659118,I3035,I658886,I658875,);
nor I_38595 (I659180,I400157,I400151);
nor I_38596 (I659197,I659180,I400169);
and I_38597 (I659214,I659197,I659101);
DFFARX1 I_38598 (I659214,I3035,I658886,I658872,);
nor I_38599 (I658869,I659180,I659036);
or I_38600 (I658866,I659118,I659180);
nor I_38601 (I659273,I400157,I400172);
DFFARX1 I_38602 (I659273,I3035,I658886,I659299,);
not I_38603 (I659307,I659299);
nand I_38604 (I659324,I659307,I658985);
nor I_38605 (I659341,I659324,I400169);
DFFARX1 I_38606 (I659341,I3035,I658886,I658854,);
nor I_38607 (I659372,I659307,I659036);
nor I_38608 (I658863,I659180,I659372);
not I_38609 (I659430,I3042);
DFFARX1 I_38610 (I169810,I3035,I659430,I659456,);
nand I_38611 (I659464,I659456,I169813);
DFFARX1 I_38612 (I169807,I3035,I659430,I659490,);
DFFARX1 I_38613 (I659490,I3035,I659430,I659507,);
not I_38614 (I659422,I659507);
not I_38615 (I659529,I169816);
nor I_38616 (I659546,I169816,I169801);
not I_38617 (I659563,I169825);
nand I_38618 (I659580,I659529,I659563);
nor I_38619 (I659597,I169825,I169816);
and I_38620 (I659401,I659597,I659464);
not I_38621 (I659628,I169804);
nand I_38622 (I659645,I659628,I169822);
nor I_38623 (I659662,I169804,I169798);
not I_38624 (I659679,I659662);
nand I_38625 (I659404,I659546,I659679);
DFFARX1 I_38626 (I659662,I3035,I659430,I659419,);
nor I_38627 (I659724,I169819,I169825);
nor I_38628 (I659741,I659724,I169801);
and I_38629 (I659758,I659741,I659645);
DFFARX1 I_38630 (I659758,I3035,I659430,I659416,);
nor I_38631 (I659413,I659724,I659580);
or I_38632 (I659410,I659662,I659724);
nor I_38633 (I659817,I169819,I169798);
DFFARX1 I_38634 (I659817,I3035,I659430,I659843,);
not I_38635 (I659851,I659843);
nand I_38636 (I659868,I659851,I659529);
nor I_38637 (I659885,I659868,I169801);
DFFARX1 I_38638 (I659885,I3035,I659430,I659398,);
nor I_38639 (I659916,I659851,I659580);
nor I_38640 (I659407,I659724,I659916);
not I_38641 (I659974,I3042);
DFFARX1 I_38642 (I49986,I3035,I659974,I660000,);
nand I_38643 (I660008,I660000,I49968);
DFFARX1 I_38644 (I49965,I3035,I659974,I660034,);
DFFARX1 I_38645 (I660034,I3035,I659974,I660051,);
not I_38646 (I659966,I660051);
not I_38647 (I660073,I49983);
nor I_38648 (I660090,I49983,I49977);
not I_38649 (I660107,I49965);
nand I_38650 (I660124,I660073,I660107);
nor I_38651 (I660141,I49965,I49983);
and I_38652 (I659945,I660141,I660008);
not I_38653 (I660172,I49974);
nand I_38654 (I660189,I660172,I49980);
nor I_38655 (I660206,I49974,I49968);
not I_38656 (I660223,I660206);
nand I_38657 (I659948,I660090,I660223);
DFFARX1 I_38658 (I660206,I3035,I659974,I659963,);
nor I_38659 (I660268,I49971,I49965);
nor I_38660 (I660285,I660268,I49977);
and I_38661 (I660302,I660285,I660189);
DFFARX1 I_38662 (I660302,I3035,I659974,I659960,);
nor I_38663 (I659957,I660268,I660124);
or I_38664 (I659954,I660206,I660268);
nor I_38665 (I660361,I49971,I49989);
DFFARX1 I_38666 (I660361,I3035,I659974,I660387,);
not I_38667 (I660395,I660387);
nand I_38668 (I660412,I660395,I660073);
nor I_38669 (I660429,I660412,I49977);
DFFARX1 I_38670 (I660429,I3035,I659974,I659942,);
nor I_38671 (I660460,I660395,I660124);
nor I_38672 (I659951,I660268,I660460);
not I_38673 (I660518,I3042);
DFFARX1 I_38674 (I410555,I3035,I660518,I660544,);
nand I_38675 (I660552,I660544,I410570);
DFFARX1 I_38676 (I410564,I3035,I660518,I660578,);
DFFARX1 I_38677 (I660578,I3035,I660518,I660595,);
not I_38678 (I660510,I660595);
not I_38679 (I660617,I410567);
nor I_38680 (I660634,I410567,I410573);
not I_38681 (I660651,I410555);
nand I_38682 (I660668,I660617,I660651);
nor I_38683 (I660685,I410555,I410567);
and I_38684 (I660489,I660685,I660552);
not I_38685 (I660716,I410552);
nand I_38686 (I660733,I660716,I410558);
nor I_38687 (I660750,I410552,I410552);
not I_38688 (I660767,I660750);
nand I_38689 (I660492,I660634,I660767);
DFFARX1 I_38690 (I660750,I3035,I660518,I660507,);
nor I_38691 (I660812,I410561,I410555);
nor I_38692 (I660829,I660812,I410573);
and I_38693 (I660846,I660829,I660733);
DFFARX1 I_38694 (I660846,I3035,I660518,I660504,);
nor I_38695 (I660501,I660812,I660668);
or I_38696 (I660498,I660750,I660812);
nor I_38697 (I660905,I410561,I410576);
DFFARX1 I_38698 (I660905,I3035,I660518,I660931,);
not I_38699 (I660939,I660931);
nand I_38700 (I660956,I660939,I660617);
nor I_38701 (I660973,I660956,I410573);
DFFARX1 I_38702 (I660973,I3035,I660518,I660486,);
nor I_38703 (I661004,I660939,I660668);
nor I_38704 (I660495,I660812,I661004);
not I_38705 (I661062,I3042);
DFFARX1 I_38706 (I46824,I3035,I661062,I661088,);
nand I_38707 (I661096,I661088,I46806);
DFFARX1 I_38708 (I46803,I3035,I661062,I661122,);
DFFARX1 I_38709 (I661122,I3035,I661062,I661139,);
not I_38710 (I661054,I661139);
not I_38711 (I661161,I46821);
nor I_38712 (I661178,I46821,I46815);
not I_38713 (I661195,I46803);
nand I_38714 (I661212,I661161,I661195);
nor I_38715 (I661229,I46803,I46821);
and I_38716 (I661033,I661229,I661096);
not I_38717 (I661260,I46812);
nand I_38718 (I661277,I661260,I46818);
nor I_38719 (I661294,I46812,I46806);
not I_38720 (I661311,I661294);
nand I_38721 (I661036,I661178,I661311);
DFFARX1 I_38722 (I661294,I3035,I661062,I661051,);
nor I_38723 (I661356,I46809,I46803);
nor I_38724 (I661373,I661356,I46815);
and I_38725 (I661390,I661373,I661277);
DFFARX1 I_38726 (I661390,I3035,I661062,I661048,);
nor I_38727 (I661045,I661356,I661212);
or I_38728 (I661042,I661294,I661356);
nor I_38729 (I661449,I46809,I46827);
DFFARX1 I_38730 (I661449,I3035,I661062,I661475,);
not I_38731 (I661483,I661475);
nand I_38732 (I661500,I661483,I661161);
nor I_38733 (I661517,I661500,I46815);
DFFARX1 I_38734 (I661517,I3035,I661062,I661030,);
nor I_38735 (I661548,I661483,I661212);
nor I_38736 (I661039,I661356,I661548);
not I_38737 (I661606,I3042);
DFFARX1 I_38738 (I363737,I3035,I661606,I661632,);
nand I_38739 (I661640,I661632,I363752);
DFFARX1 I_38740 (I363746,I3035,I661606,I661666,);
DFFARX1 I_38741 (I661666,I3035,I661606,I661683,);
not I_38742 (I661598,I661683);
not I_38743 (I661705,I363749);
nor I_38744 (I661722,I363749,I363755);
not I_38745 (I661739,I363737);
nand I_38746 (I661756,I661705,I661739);
nor I_38747 (I661773,I363737,I363749);
and I_38748 (I661577,I661773,I661640);
not I_38749 (I661804,I363734);
nand I_38750 (I661821,I661804,I363740);
nor I_38751 (I661838,I363734,I363734);
not I_38752 (I661855,I661838);
nand I_38753 (I661580,I661722,I661855);
DFFARX1 I_38754 (I661838,I3035,I661606,I661595,);
nor I_38755 (I661900,I363743,I363737);
nor I_38756 (I661917,I661900,I363755);
and I_38757 (I661934,I661917,I661821);
DFFARX1 I_38758 (I661934,I3035,I661606,I661592,);
nor I_38759 (I661589,I661900,I661756);
or I_38760 (I661586,I661838,I661900);
nor I_38761 (I661993,I363743,I363758);
DFFARX1 I_38762 (I661993,I3035,I661606,I662019,);
not I_38763 (I662027,I662019);
nand I_38764 (I662044,I662027,I661705);
nor I_38765 (I662061,I662044,I363755);
DFFARX1 I_38766 (I662061,I3035,I661606,I661574,);
nor I_38767 (I662092,I662027,I661756);
nor I_38768 (I661583,I661900,I662092);
not I_38769 (I662150,I3042);
DFFARX1 I_38770 (I429819,I3035,I662150,I662176,);
nand I_38771 (I662184,I662176,I429813);
DFFARX1 I_38772 (I429816,I3035,I662150,I662210,);
DFFARX1 I_38773 (I662210,I3035,I662150,I662227,);
not I_38774 (I662142,I662227);
not I_38775 (I662249,I429822);
nor I_38776 (I662266,I429822,I429816);
not I_38777 (I662283,I429825);
nand I_38778 (I662300,I662249,I662283);
nor I_38779 (I662317,I429825,I429822);
and I_38780 (I662121,I662317,I662184);
not I_38781 (I662348,I429834);
nand I_38782 (I662365,I662348,I429828);
nor I_38783 (I662382,I429834,I429831);
not I_38784 (I662399,I662382);
nand I_38785 (I662124,I662266,I662399);
DFFARX1 I_38786 (I662382,I3035,I662150,I662139,);
nor I_38787 (I662444,I429813,I429825);
nor I_38788 (I662461,I662444,I429816);
and I_38789 (I662478,I662461,I662365);
DFFARX1 I_38790 (I662478,I3035,I662150,I662136,);
nor I_38791 (I662133,I662444,I662300);
or I_38792 (I662130,I662382,I662444);
nor I_38793 (I662537,I429813,I429819);
DFFARX1 I_38794 (I662537,I3035,I662150,I662563,);
not I_38795 (I662571,I662563);
nand I_38796 (I662588,I662571,I662249);
nor I_38797 (I662605,I662588,I429816);
DFFARX1 I_38798 (I662605,I3035,I662150,I662118,);
nor I_38799 (I662636,I662571,I662300);
nor I_38800 (I662127,I662444,I662636);
not I_38801 (I662694,I3042);
DFFARX1 I_38802 (I138408,I3035,I662694,I662720,);
nand I_38803 (I662728,I662720,I138423);
DFFARX1 I_38804 (I138420,I3035,I662694,I662754,);
DFFARX1 I_38805 (I662754,I3035,I662694,I662771,);
not I_38806 (I662686,I662771);
not I_38807 (I662793,I138399);
nor I_38808 (I662810,I138399,I138405);
not I_38809 (I662827,I138411);
nand I_38810 (I662844,I662793,I662827);
nor I_38811 (I662861,I138411,I138399);
and I_38812 (I662665,I662861,I662728);
not I_38813 (I662892,I138417);
nand I_38814 (I662909,I662892,I138399);
nor I_38815 (I662926,I138417,I138402);
not I_38816 (I662943,I662926);
nand I_38817 (I662668,I662810,I662943);
DFFARX1 I_38818 (I662926,I3035,I662694,I662683,);
nor I_38819 (I662988,I138402,I138411);
nor I_38820 (I663005,I662988,I138405);
and I_38821 (I663022,I663005,I662909);
DFFARX1 I_38822 (I663022,I3035,I662694,I662680,);
nor I_38823 (I662677,I662988,I662844);
or I_38824 (I662674,I662926,I662988);
nor I_38825 (I663081,I138402,I138414);
DFFARX1 I_38826 (I663081,I3035,I662694,I663107,);
not I_38827 (I663115,I663107);
nand I_38828 (I663132,I663115,I662793);
nor I_38829 (I663149,I663132,I138405);
DFFARX1 I_38830 (I663149,I3035,I662694,I662662,);
nor I_38831 (I663180,I663115,I662844);
nor I_38832 (I662671,I662988,I663180);
not I_38833 (I663238,I3042);
DFFARX1 I_38834 (I704985,I3035,I663238,I663264,);
nand I_38835 (I663272,I663264,I704970);
DFFARX1 I_38836 (I704964,I3035,I663238,I663298,);
DFFARX1 I_38837 (I663298,I3035,I663238,I663315,);
not I_38838 (I663230,I663315);
not I_38839 (I663337,I704958);
nor I_38840 (I663354,I704958,I704979);
not I_38841 (I663371,I704967);
nand I_38842 (I663388,I663337,I663371);
nor I_38843 (I663405,I704967,I704958);
and I_38844 (I663209,I663405,I663272);
not I_38845 (I663436,I704976);
nand I_38846 (I663453,I663436,I704982);
nor I_38847 (I663470,I704976,I704973);
not I_38848 (I663487,I663470);
nand I_38849 (I663212,I663354,I663487);
DFFARX1 I_38850 (I663470,I3035,I663238,I663227,);
nor I_38851 (I663532,I704961,I704967);
nor I_38852 (I663549,I663532,I704979);
and I_38853 (I663566,I663549,I663453);
DFFARX1 I_38854 (I663566,I3035,I663238,I663224,);
nor I_38855 (I663221,I663532,I663388);
or I_38856 (I663218,I663470,I663532);
nor I_38857 (I663625,I704961,I704958);
DFFARX1 I_38858 (I663625,I3035,I663238,I663651,);
not I_38859 (I663659,I663651);
nand I_38860 (I663676,I663659,I663337);
nor I_38861 (I663693,I663676,I704979);
DFFARX1 I_38862 (I663693,I3035,I663238,I663206,);
nor I_38863 (I663724,I663659,I663388);
nor I_38864 (I663215,I663532,I663724);
not I_38865 (I663782,I3042);
DFFARX1 I_38866 (I31541,I3035,I663782,I663808,);
nand I_38867 (I663816,I663808,I31523);
DFFARX1 I_38868 (I31520,I3035,I663782,I663842,);
DFFARX1 I_38869 (I663842,I3035,I663782,I663859,);
not I_38870 (I663774,I663859);
not I_38871 (I663881,I31538);
nor I_38872 (I663898,I31538,I31532);
not I_38873 (I663915,I31520);
nand I_38874 (I663932,I663881,I663915);
nor I_38875 (I663949,I31520,I31538);
and I_38876 (I663753,I663949,I663816);
not I_38877 (I663980,I31529);
nand I_38878 (I663997,I663980,I31535);
nor I_38879 (I664014,I31529,I31523);
not I_38880 (I664031,I664014);
nand I_38881 (I663756,I663898,I664031);
DFFARX1 I_38882 (I664014,I3035,I663782,I663771,);
nor I_38883 (I664076,I31526,I31520);
nor I_38884 (I664093,I664076,I31532);
and I_38885 (I664110,I664093,I663997);
DFFARX1 I_38886 (I664110,I3035,I663782,I663768,);
nor I_38887 (I663765,I664076,I663932);
or I_38888 (I663762,I664014,I664076);
nor I_38889 (I664169,I31526,I31544);
DFFARX1 I_38890 (I664169,I3035,I663782,I664195,);
not I_38891 (I664203,I664195);
nand I_38892 (I664220,I664203,I663881);
nor I_38893 (I664237,I664220,I31532);
DFFARX1 I_38894 (I664237,I3035,I663782,I663750,);
nor I_38895 (I664268,I664203,I663932);
nor I_38896 (I663759,I664076,I664268);
not I_38897 (I664326,I3042);
DFFARX1 I_38898 (I200903,I3035,I664326,I664352,);
nand I_38899 (I664360,I664352,I200906);
DFFARX1 I_38900 (I200900,I3035,I664326,I664386,);
DFFARX1 I_38901 (I664386,I3035,I664326,I664403,);
not I_38902 (I664318,I664403);
not I_38903 (I664425,I200909);
nor I_38904 (I664442,I200909,I200894);
not I_38905 (I664459,I200918);
nand I_38906 (I664476,I664425,I664459);
nor I_38907 (I664493,I200918,I200909);
and I_38908 (I664297,I664493,I664360);
not I_38909 (I664524,I200897);
nand I_38910 (I664541,I664524,I200915);
nor I_38911 (I664558,I200897,I200891);
not I_38912 (I664575,I664558);
nand I_38913 (I664300,I664442,I664575);
DFFARX1 I_38914 (I664558,I3035,I664326,I664315,);
nor I_38915 (I664620,I200912,I200918);
nor I_38916 (I664637,I664620,I200894);
and I_38917 (I664654,I664637,I664541);
DFFARX1 I_38918 (I664654,I3035,I664326,I664312,);
nor I_38919 (I664309,I664620,I664476);
or I_38920 (I664306,I664558,I664620);
nor I_38921 (I664713,I200912,I200891);
DFFARX1 I_38922 (I664713,I3035,I664326,I664739,);
not I_38923 (I664747,I664739);
nand I_38924 (I664764,I664747,I664425);
nor I_38925 (I664781,I664764,I200894);
DFFARX1 I_38926 (I664781,I3035,I664326,I664294,);
nor I_38927 (I664812,I664747,I664476);
nor I_38928 (I664303,I664620,I664812);
not I_38929 (I664870,I3042);
DFFARX1 I_38930 (I458277,I3035,I664870,I664896,);
nand I_38931 (I664904,I664896,I458271);
DFFARX1 I_38932 (I458274,I3035,I664870,I664930,);
DFFARX1 I_38933 (I664930,I3035,I664870,I664947,);
not I_38934 (I664862,I664947);
not I_38935 (I664969,I458280);
nor I_38936 (I664986,I458280,I458274);
not I_38937 (I665003,I458283);
nand I_38938 (I665020,I664969,I665003);
nor I_38939 (I665037,I458283,I458280);
and I_38940 (I664841,I665037,I664904);
not I_38941 (I665068,I458292);
nand I_38942 (I665085,I665068,I458286);
nor I_38943 (I665102,I458292,I458289);
not I_38944 (I665119,I665102);
nand I_38945 (I664844,I664986,I665119);
DFFARX1 I_38946 (I665102,I3035,I664870,I664859,);
nor I_38947 (I665164,I458271,I458283);
nor I_38948 (I665181,I665164,I458274);
and I_38949 (I665198,I665181,I665085);
DFFARX1 I_38950 (I665198,I3035,I664870,I664856,);
nor I_38951 (I664853,I665164,I665020);
or I_38952 (I664850,I665102,I665164);
nor I_38953 (I665257,I458271,I458277);
DFFARX1 I_38954 (I665257,I3035,I664870,I665283,);
not I_38955 (I665291,I665283);
nand I_38956 (I665308,I665291,I664969);
nor I_38957 (I665325,I665308,I458274);
DFFARX1 I_38958 (I665325,I3035,I664870,I664838,);
nor I_38959 (I665356,I665291,I665020);
nor I_38960 (I664847,I665164,I665356);
not I_38961 (I665414,I3042);
DFFARX1 I_38962 (I732355,I3035,I665414,I665440,);
nand I_38963 (I665448,I665440,I732340);
DFFARX1 I_38964 (I732334,I3035,I665414,I665474,);
DFFARX1 I_38965 (I665474,I3035,I665414,I665491,);
not I_38966 (I665406,I665491);
not I_38967 (I665513,I732328);
nor I_38968 (I665530,I732328,I732349);
not I_38969 (I665547,I732337);
nand I_38970 (I665564,I665513,I665547);
nor I_38971 (I665581,I732337,I732328);
and I_38972 (I665385,I665581,I665448);
not I_38973 (I665612,I732346);
nand I_38974 (I665629,I665612,I732352);
nor I_38975 (I665646,I732346,I732343);
not I_38976 (I665663,I665646);
nand I_38977 (I665388,I665530,I665663);
DFFARX1 I_38978 (I665646,I3035,I665414,I665403,);
nor I_38979 (I665708,I732331,I732337);
nor I_38980 (I665725,I665708,I732349);
and I_38981 (I665742,I665725,I665629);
DFFARX1 I_38982 (I665742,I3035,I665414,I665400,);
nor I_38983 (I665397,I665708,I665564);
or I_38984 (I665394,I665646,I665708);
nor I_38985 (I665801,I732331,I732328);
DFFARX1 I_38986 (I665801,I3035,I665414,I665827,);
not I_38987 (I665835,I665827);
nand I_38988 (I665852,I665835,I665513);
nor I_38989 (I665869,I665852,I732349);
DFFARX1 I_38990 (I665869,I3035,I665414,I665382,);
nor I_38991 (I665900,I665835,I665564);
nor I_38992 (I665391,I665708,I665900);
not I_38993 (I665958,I3042);
DFFARX1 I_38994 (I225145,I3035,I665958,I665984,);
nand I_38995 (I665992,I665984,I225148);
DFFARX1 I_38996 (I225142,I3035,I665958,I666018,);
DFFARX1 I_38997 (I666018,I3035,I665958,I666035,);
not I_38998 (I665950,I666035);
not I_38999 (I666057,I225151);
nor I_39000 (I666074,I225151,I225136);
not I_39001 (I666091,I225160);
nand I_39002 (I666108,I666057,I666091);
nor I_39003 (I666125,I225160,I225151);
and I_39004 (I665929,I666125,I665992);
not I_39005 (I666156,I225139);
nand I_39006 (I666173,I666156,I225157);
nor I_39007 (I666190,I225139,I225133);
not I_39008 (I666207,I666190);
nand I_39009 (I665932,I666074,I666207);
DFFARX1 I_39010 (I666190,I3035,I665958,I665947,);
nor I_39011 (I666252,I225154,I225160);
nor I_39012 (I666269,I666252,I225136);
and I_39013 (I666286,I666269,I666173);
DFFARX1 I_39014 (I666286,I3035,I665958,I665944,);
nor I_39015 (I665941,I666252,I666108);
or I_39016 (I665938,I666190,I666252);
nor I_39017 (I666345,I225154,I225133);
DFFARX1 I_39018 (I666345,I3035,I665958,I666371,);
not I_39019 (I666379,I666371);
nand I_39020 (I666396,I666379,I666057);
nor I_39021 (I666413,I666396,I225136);
DFFARX1 I_39022 (I666413,I3035,I665958,I665926,);
nor I_39023 (I666444,I666379,I666108);
nor I_39024 (I665935,I666252,I666444);
not I_39025 (I666502,I3042);
DFFARX1 I_39026 (I526458,I3035,I666502,I666528,);
nand I_39027 (I666536,I666528,I526458);
DFFARX1 I_39028 (I526470,I3035,I666502,I666562,);
DFFARX1 I_39029 (I666562,I3035,I666502,I666579,);
not I_39030 (I666494,I666579);
not I_39031 (I666601,I526464);
nor I_39032 (I666618,I526464,I526485);
not I_39033 (I666635,I526473);
nand I_39034 (I666652,I666601,I666635);
nor I_39035 (I666669,I526473,I526464);
and I_39036 (I666473,I666669,I666536);
not I_39037 (I666700,I526467);
nand I_39038 (I666717,I666700,I526482);
nor I_39039 (I666734,I526467,I526476);
not I_39040 (I666751,I666734);
nand I_39041 (I666476,I666618,I666751);
DFFARX1 I_39042 (I666734,I3035,I666502,I666491,);
nor I_39043 (I666796,I526479,I526473);
nor I_39044 (I666813,I666796,I526485);
and I_39045 (I666830,I666813,I666717);
DFFARX1 I_39046 (I666830,I3035,I666502,I666488,);
nor I_39047 (I666485,I666796,I666652);
or I_39048 (I666482,I666734,I666796);
nor I_39049 (I666889,I526479,I526461);
DFFARX1 I_39050 (I666889,I3035,I666502,I666915,);
not I_39051 (I666923,I666915);
nand I_39052 (I666940,I666923,I666601);
nor I_39053 (I666957,I666940,I526485);
DFFARX1 I_39054 (I666957,I3035,I666502,I666470,);
nor I_39055 (I666988,I666923,I666652);
nor I_39056 (I666479,I666796,I666988);
not I_39057 (I667046,I3042);
DFFARX1 I_39058 (I725215,I3035,I667046,I667072,);
nand I_39059 (I667080,I667072,I725200);
DFFARX1 I_39060 (I725194,I3035,I667046,I667106,);
DFFARX1 I_39061 (I667106,I3035,I667046,I667123,);
not I_39062 (I667038,I667123);
not I_39063 (I667145,I725188);
nor I_39064 (I667162,I725188,I725209);
not I_39065 (I667179,I725197);
nand I_39066 (I667196,I667145,I667179);
nor I_39067 (I667213,I725197,I725188);
and I_39068 (I667017,I667213,I667080);
not I_39069 (I667244,I725206);
nand I_39070 (I667261,I667244,I725212);
nor I_39071 (I667278,I725206,I725203);
not I_39072 (I667295,I667278);
nand I_39073 (I667020,I667162,I667295);
DFFARX1 I_39074 (I667278,I3035,I667046,I667035,);
nor I_39075 (I667340,I725191,I725197);
nor I_39076 (I667357,I667340,I725209);
and I_39077 (I667374,I667357,I667261);
DFFARX1 I_39078 (I667374,I3035,I667046,I667032,);
nor I_39079 (I667029,I667340,I667196);
or I_39080 (I667026,I667278,I667340);
nor I_39081 (I667433,I725191,I725188);
DFFARX1 I_39082 (I667433,I3035,I667046,I667459,);
not I_39083 (I667467,I667459);
nand I_39084 (I667484,I667467,I667145);
nor I_39085 (I667501,I667484,I725209);
DFFARX1 I_39086 (I667501,I3035,I667046,I667014,);
nor I_39087 (I667532,I667467,I667196);
nor I_39088 (I667023,I667340,I667532);
not I_39089 (I667590,I3042);
DFFARX1 I_39090 (I90808,I3035,I667590,I667616,);
nand I_39091 (I667624,I667616,I90823);
DFFARX1 I_39092 (I90820,I3035,I667590,I667650,);
DFFARX1 I_39093 (I667650,I3035,I667590,I667667,);
not I_39094 (I667582,I667667);
not I_39095 (I667689,I90799);
nor I_39096 (I667706,I90799,I90805);
not I_39097 (I667723,I90811);
nand I_39098 (I667740,I667689,I667723);
nor I_39099 (I667757,I90811,I90799);
and I_39100 (I667561,I667757,I667624);
not I_39101 (I667788,I90817);
nand I_39102 (I667805,I667788,I90799);
nor I_39103 (I667822,I90817,I90802);
not I_39104 (I667839,I667822);
nand I_39105 (I667564,I667706,I667839);
DFFARX1 I_39106 (I667822,I3035,I667590,I667579,);
nor I_39107 (I667884,I90802,I90811);
nor I_39108 (I667901,I667884,I90805);
and I_39109 (I667918,I667901,I667805);
DFFARX1 I_39110 (I667918,I3035,I667590,I667576,);
nor I_39111 (I667573,I667884,I667740);
or I_39112 (I667570,I667822,I667884);
nor I_39113 (I667977,I90802,I90814);
DFFARX1 I_39114 (I667977,I3035,I667590,I668003,);
not I_39115 (I668011,I668003);
nand I_39116 (I668028,I668011,I667689);
nor I_39117 (I668045,I668028,I90805);
DFFARX1 I_39118 (I668045,I3035,I667590,I667558,);
nor I_39119 (I668076,I668011,I667740);
nor I_39120 (I667567,I667884,I668076);
not I_39121 (I668134,I3042);
DFFARX1 I_39122 (I202484,I3035,I668134,I668160,);
nand I_39123 (I668168,I668160,I202487);
DFFARX1 I_39124 (I202481,I3035,I668134,I668194,);
DFFARX1 I_39125 (I668194,I3035,I668134,I668211,);
not I_39126 (I668126,I668211);
not I_39127 (I668233,I202490);
nor I_39128 (I668250,I202490,I202475);
not I_39129 (I668267,I202499);
nand I_39130 (I668284,I668233,I668267);
nor I_39131 (I668301,I202499,I202490);
and I_39132 (I668105,I668301,I668168);
not I_39133 (I668332,I202478);
nand I_39134 (I668349,I668332,I202496);
nor I_39135 (I668366,I202478,I202472);
not I_39136 (I668383,I668366);
nand I_39137 (I668108,I668250,I668383);
DFFARX1 I_39138 (I668366,I3035,I668134,I668123,);
nor I_39139 (I668428,I202493,I202499);
nor I_39140 (I668445,I668428,I202475);
and I_39141 (I668462,I668445,I668349);
DFFARX1 I_39142 (I668462,I3035,I668134,I668120,);
nor I_39143 (I668117,I668428,I668284);
or I_39144 (I668114,I668366,I668428);
nor I_39145 (I668521,I202493,I202472);
DFFARX1 I_39146 (I668521,I3035,I668134,I668547,);
not I_39147 (I668555,I668547);
nand I_39148 (I668572,I668555,I668233);
nor I_39149 (I668589,I668572,I202475);
DFFARX1 I_39150 (I668589,I3035,I668134,I668102,);
nor I_39151 (I668620,I668555,I668284);
nor I_39152 (I668111,I668428,I668620);
not I_39153 (I668678,I3042);
DFFARX1 I_39154 (I434035,I3035,I668678,I668704,);
nand I_39155 (I668712,I668704,I434029);
DFFARX1 I_39156 (I434032,I3035,I668678,I668738,);
DFFARX1 I_39157 (I668738,I3035,I668678,I668755,);
not I_39158 (I668670,I668755);
not I_39159 (I668777,I434038);
nor I_39160 (I668794,I434038,I434032);
not I_39161 (I668811,I434041);
nand I_39162 (I668828,I668777,I668811);
nor I_39163 (I668845,I434041,I434038);
and I_39164 (I668649,I668845,I668712);
not I_39165 (I668876,I434050);
nand I_39166 (I668893,I668876,I434044);
nor I_39167 (I668910,I434050,I434047);
not I_39168 (I668927,I668910);
nand I_39169 (I668652,I668794,I668927);
DFFARX1 I_39170 (I668910,I3035,I668678,I668667,);
nor I_39171 (I668972,I434029,I434041);
nor I_39172 (I668989,I668972,I434032);
and I_39173 (I669006,I668989,I668893);
DFFARX1 I_39174 (I669006,I3035,I668678,I668664,);
nor I_39175 (I668661,I668972,I668828);
or I_39176 (I668658,I668910,I668972);
nor I_39177 (I669065,I434029,I434035);
DFFARX1 I_39178 (I669065,I3035,I668678,I669091,);
not I_39179 (I669099,I669091);
nand I_39180 (I669116,I669099,I668777);
nor I_39181 (I669133,I669116,I434032);
DFFARX1 I_39182 (I669133,I3035,I668678,I668646,);
nor I_39183 (I669164,I669099,I668828);
nor I_39184 (I668655,I668972,I669164);
not I_39185 (I669222,I3042);
DFFARX1 I_39186 (I283511,I3035,I669222,I669248,);
nand I_39187 (I669256,I669248,I283535);
DFFARX1 I_39188 (I283514,I3035,I669222,I669282,);
DFFARX1 I_39189 (I669282,I3035,I669222,I669299,);
not I_39190 (I669214,I669299);
not I_39191 (I669321,I283517);
nor I_39192 (I669338,I283517,I283532);
not I_39193 (I669355,I283523);
nand I_39194 (I669372,I669321,I669355);
nor I_39195 (I669389,I283523,I283517);
and I_39196 (I669193,I669389,I669256);
not I_39197 (I669420,I283520);
nand I_39198 (I669437,I669420,I283514);
nor I_39199 (I669454,I283520,I283529);
not I_39200 (I669471,I669454);
nand I_39201 (I669196,I669338,I669471);
DFFARX1 I_39202 (I669454,I3035,I669222,I669211,);
nor I_39203 (I669516,I283526,I283523);
nor I_39204 (I669533,I669516,I283532);
and I_39205 (I669550,I669533,I669437);
DFFARX1 I_39206 (I669550,I3035,I669222,I669208,);
nor I_39207 (I669205,I669516,I669372);
or I_39208 (I669202,I669454,I669516);
nor I_39209 (I669609,I283526,I283511);
DFFARX1 I_39210 (I669609,I3035,I669222,I669635,);
not I_39211 (I669643,I669635);
nand I_39212 (I669660,I669643,I669321);
nor I_39213 (I669677,I669660,I283532);
DFFARX1 I_39214 (I669677,I3035,I669222,I669190,);
nor I_39215 (I669708,I669643,I669372);
nor I_39216 (I669199,I669516,I669708);
not I_39217 (I669766,I3042);
DFFARX1 I_39218 (I735925,I3035,I669766,I669792,);
nand I_39219 (I669800,I669792,I735910);
DFFARX1 I_39220 (I735904,I3035,I669766,I669826,);
DFFARX1 I_39221 (I669826,I3035,I669766,I669843,);
not I_39222 (I669758,I669843);
not I_39223 (I669865,I735898);
nor I_39224 (I669882,I735898,I735919);
not I_39225 (I669899,I735907);
nand I_39226 (I669916,I669865,I669899);
nor I_39227 (I669933,I735907,I735898);
and I_39228 (I669737,I669933,I669800);
not I_39229 (I669964,I735916);
nand I_39230 (I669981,I669964,I735922);
nor I_39231 (I669998,I735916,I735913);
not I_39232 (I670015,I669998);
nand I_39233 (I669740,I669882,I670015);
DFFARX1 I_39234 (I669998,I3035,I669766,I669755,);
nor I_39235 (I670060,I735901,I735907);
nor I_39236 (I670077,I670060,I735919);
and I_39237 (I670094,I670077,I669981);
DFFARX1 I_39238 (I670094,I3035,I669766,I669752,);
nor I_39239 (I669749,I670060,I669916);
or I_39240 (I669746,I669998,I670060);
nor I_39241 (I670153,I735901,I735898);
DFFARX1 I_39242 (I670153,I3035,I669766,I670179,);
not I_39243 (I670187,I670179);
nand I_39244 (I670204,I670187,I669865);
nor I_39245 (I670221,I670204,I735919);
DFFARX1 I_39246 (I670221,I3035,I669766,I669734,);
nor I_39247 (I670252,I670187,I669916);
nor I_39248 (I669743,I670060,I670252);
not I_39249 (I670310,I3042);
DFFARX1 I_39250 (I222510,I3035,I670310,I670336,);
nand I_39251 (I670344,I670336,I222513);
DFFARX1 I_39252 (I222507,I3035,I670310,I670370,);
DFFARX1 I_39253 (I670370,I3035,I670310,I670387,);
not I_39254 (I670302,I670387);
not I_39255 (I670409,I222516);
nor I_39256 (I670426,I222516,I222501);
not I_39257 (I670443,I222525);
nand I_39258 (I670460,I670409,I670443);
nor I_39259 (I670477,I222525,I222516);
and I_39260 (I670281,I670477,I670344);
not I_39261 (I670508,I222504);
nand I_39262 (I670525,I670508,I222522);
nor I_39263 (I670542,I222504,I222498);
not I_39264 (I670559,I670542);
nand I_39265 (I670284,I670426,I670559);
DFFARX1 I_39266 (I670542,I3035,I670310,I670299,);
nor I_39267 (I670604,I222519,I222525);
nor I_39268 (I670621,I670604,I222501);
and I_39269 (I670638,I670621,I670525);
DFFARX1 I_39270 (I670638,I3035,I670310,I670296,);
nor I_39271 (I670293,I670604,I670460);
or I_39272 (I670290,I670542,I670604);
nor I_39273 (I670697,I222519,I222498);
DFFARX1 I_39274 (I670697,I3035,I670310,I670723,);
not I_39275 (I670731,I670723);
nand I_39276 (I670748,I670731,I670409);
nor I_39277 (I670765,I670748,I222501);
DFFARX1 I_39278 (I670765,I3035,I670310,I670278,);
nor I_39279 (I670796,I670731,I670460);
nor I_39280 (I670287,I670604,I670796);
not I_39281 (I670854,I3042);
DFFARX1 I_39282 (I470398,I3035,I670854,I670880,);
nand I_39283 (I670888,I670880,I470392);
DFFARX1 I_39284 (I470395,I3035,I670854,I670914,);
DFFARX1 I_39285 (I670914,I3035,I670854,I670931,);
not I_39286 (I670846,I670931);
not I_39287 (I670953,I470401);
nor I_39288 (I670970,I470401,I470395);
not I_39289 (I670987,I470404);
nand I_39290 (I671004,I670953,I670987);
nor I_39291 (I671021,I470404,I470401);
and I_39292 (I670825,I671021,I670888);
not I_39293 (I671052,I470413);
nand I_39294 (I671069,I671052,I470407);
nor I_39295 (I671086,I470413,I470410);
not I_39296 (I671103,I671086);
nand I_39297 (I670828,I670970,I671103);
DFFARX1 I_39298 (I671086,I3035,I670854,I670843,);
nor I_39299 (I671148,I470392,I470404);
nor I_39300 (I671165,I671148,I470395);
and I_39301 (I671182,I671165,I671069);
DFFARX1 I_39302 (I671182,I3035,I670854,I670840,);
nor I_39303 (I670837,I671148,I671004);
or I_39304 (I670834,I671086,I671148);
nor I_39305 (I671241,I470392,I470398);
DFFARX1 I_39306 (I671241,I3035,I670854,I671267,);
not I_39307 (I671275,I671267);
nand I_39308 (I671292,I671275,I670953);
nor I_39309 (I671309,I671292,I470395);
DFFARX1 I_39310 (I671309,I3035,I670854,I670822,);
nor I_39311 (I671340,I671275,I671004);
nor I_39312 (I670831,I671148,I671340);
not I_39313 (I671398,I3042);
DFFARX1 I_39314 (I82478,I3035,I671398,I671424,);
nand I_39315 (I671432,I671424,I82493);
DFFARX1 I_39316 (I82490,I3035,I671398,I671458,);
DFFARX1 I_39317 (I671458,I3035,I671398,I671475,);
not I_39318 (I671390,I671475);
not I_39319 (I671497,I82469);
nor I_39320 (I671514,I82469,I82475);
not I_39321 (I671531,I82481);
nand I_39322 (I671548,I671497,I671531);
nor I_39323 (I671565,I82481,I82469);
and I_39324 (I671369,I671565,I671432);
not I_39325 (I671596,I82487);
nand I_39326 (I671613,I671596,I82469);
nor I_39327 (I671630,I82487,I82472);
not I_39328 (I671647,I671630);
nand I_39329 (I671372,I671514,I671647);
DFFARX1 I_39330 (I671630,I3035,I671398,I671387,);
nor I_39331 (I671692,I82472,I82481);
nor I_39332 (I671709,I671692,I82475);
and I_39333 (I671726,I671709,I671613);
DFFARX1 I_39334 (I671726,I3035,I671398,I671384,);
nor I_39335 (I671381,I671692,I671548);
or I_39336 (I671378,I671630,I671692);
nor I_39337 (I671785,I82472,I82484);
DFFARX1 I_39338 (I671785,I3035,I671398,I671811,);
not I_39339 (I671819,I671811);
nand I_39340 (I671836,I671819,I671497);
nor I_39341 (I671853,I671836,I82475);
DFFARX1 I_39342 (I671853,I3035,I671398,I671366,);
nor I_39343 (I671884,I671819,I671548);
nor I_39344 (I671375,I671692,I671884);
not I_39345 (I671942,I3042);
DFFARX1 I_39346 (I362000,I3035,I671942,I671968,);
nand I_39347 (I671976,I671968,I362003);
not I_39348 (I671993,I671976);
DFFARX1 I_39349 (I362015,I3035,I671942,I672019,);
not I_39350 (I672027,I672019);
not I_39351 (I672044,I362000);
or I_39352 (I672061,I362009,I362000);
nor I_39353 (I672078,I362009,I362000);
or I_39354 (I672095,I362018,I362009);
DFFARX1 I_39355 (I672095,I3035,I671942,I671934,);
not I_39356 (I672126,I362021);
nand I_39357 (I672143,I672126,I362003);
nand I_39358 (I672160,I672044,I672143);
and I_39359 (I671913,I672027,I672160);
nor I_39360 (I672191,I362021,I362006);
and I_39361 (I672208,I672027,I672191);
nor I_39362 (I671919,I671993,I672208);
DFFARX1 I_39363 (I672191,I3035,I671942,I672248,);
not I_39364 (I672256,I672248);
nor I_39365 (I671928,I672027,I672256);
or I_39366 (I672287,I672095,I362012);
nor I_39367 (I672304,I362012,I362018);
nand I_39368 (I672321,I672160,I672304);
nand I_39369 (I672338,I672287,I672321);
DFFARX1 I_39370 (I672338,I3035,I671942,I671931,);
nor I_39371 (I672369,I672304,I672061);
DFFARX1 I_39372 (I672369,I3035,I671942,I671910,);
nor I_39373 (I672400,I362012,I362024);
DFFARX1 I_39374 (I672400,I3035,I671942,I672426,);
DFFARX1 I_39375 (I672426,I3035,I671942,I671925,);
not I_39376 (I672448,I672426);
nand I_39377 (I671922,I672448,I671976);
nand I_39378 (I671916,I672448,I672078);
not I_39379 (I672520,I3042);
DFFARX1 I_39380 (I407084,I3035,I672520,I672546,);
nand I_39381 (I672554,I672546,I407087);
not I_39382 (I672571,I672554);
DFFARX1 I_39383 (I407099,I3035,I672520,I672597,);
not I_39384 (I672605,I672597);
not I_39385 (I672622,I407084);
or I_39386 (I672639,I407093,I407084);
nor I_39387 (I672656,I407093,I407084);
or I_39388 (I672673,I407102,I407093);
DFFARX1 I_39389 (I672673,I3035,I672520,I672512,);
not I_39390 (I672704,I407105);
nand I_39391 (I672721,I672704,I407087);
nand I_39392 (I672738,I672622,I672721);
and I_39393 (I672491,I672605,I672738);
nor I_39394 (I672769,I407105,I407090);
and I_39395 (I672786,I672605,I672769);
nor I_39396 (I672497,I672571,I672786);
DFFARX1 I_39397 (I672769,I3035,I672520,I672826,);
not I_39398 (I672834,I672826);
nor I_39399 (I672506,I672605,I672834);
or I_39400 (I672865,I672673,I407096);
nor I_39401 (I672882,I407096,I407102);
nand I_39402 (I672899,I672738,I672882);
nand I_39403 (I672916,I672865,I672899);
DFFARX1 I_39404 (I672916,I3035,I672520,I672509,);
nor I_39405 (I672947,I672882,I672639);
DFFARX1 I_39406 (I672947,I3035,I672520,I672488,);
nor I_39407 (I672978,I407096,I407108);
DFFARX1 I_39408 (I672978,I3035,I672520,I673004,);
DFFARX1 I_39409 (I673004,I3035,I672520,I672503,);
not I_39410 (I673026,I673004);
nand I_39411 (I672500,I673026,I672554);
nand I_39412 (I672494,I673026,I672656);
not I_39413 (I673098,I3042);
DFFARX1 I_39414 (I538092,I3035,I673098,I673124,);
nand I_39415 (I673132,I673124,I538113);
not I_39416 (I673149,I673132);
DFFARX1 I_39417 (I538086,I3035,I673098,I673175,);
not I_39418 (I673183,I673175);
not I_39419 (I673200,I538107);
or I_39420 (I673217,I538098,I538107);
nor I_39421 (I673234,I538098,I538107);
or I_39422 (I673251,I538101,I538098);
DFFARX1 I_39423 (I673251,I3035,I673098,I673090,);
not I_39424 (I673282,I538089);
nand I_39425 (I673299,I673282,I538104);
nand I_39426 (I673316,I673200,I673299);
and I_39427 (I673069,I673183,I673316);
nor I_39428 (I673347,I538089,I538086);
and I_39429 (I673364,I673183,I673347);
nor I_39430 (I673075,I673149,I673364);
DFFARX1 I_39431 (I673347,I3035,I673098,I673404,);
not I_39432 (I673412,I673404);
nor I_39433 (I673084,I673183,I673412);
or I_39434 (I673443,I673251,I538110);
nor I_39435 (I673460,I538110,I538101);
nand I_39436 (I673477,I673316,I673460);
nand I_39437 (I673494,I673443,I673477);
DFFARX1 I_39438 (I673494,I3035,I673098,I673087,);
nor I_39439 (I673525,I673460,I673217);
DFFARX1 I_39440 (I673525,I3035,I673098,I673066,);
nor I_39441 (I673556,I538110,I538095);
DFFARX1 I_39442 (I673556,I3035,I673098,I673582,);
DFFARX1 I_39443 (I673582,I3035,I673098,I673081,);
not I_39444 (I673604,I673582);
nand I_39445 (I673078,I673604,I673132);
nand I_39446 (I673072,I673604,I673234);
not I_39447 (I673676,I3042);
DFFARX1 I_39448 (I427708,I3035,I673676,I673702,);
nand I_39449 (I673710,I673702,I427708);
not I_39450 (I673727,I673710);
DFFARX1 I_39451 (I427714,I3035,I673676,I673753,);
not I_39452 (I673761,I673753);
not I_39453 (I673778,I427726);
or I_39454 (I673795,I427711,I427726);
nor I_39455 (I673812,I427711,I427726);
or I_39456 (I673829,I427705,I427711);
DFFARX1 I_39457 (I673829,I3035,I673676,I673668,);
not I_39458 (I673860,I427723);
nand I_39459 (I673877,I673860,I427717);
nand I_39460 (I673894,I673778,I673877);
and I_39461 (I673647,I673761,I673894);
nor I_39462 (I673925,I427723,I427705);
and I_39463 (I673942,I673761,I673925);
nor I_39464 (I673653,I673727,I673942);
DFFARX1 I_39465 (I673925,I3035,I673676,I673982,);
not I_39466 (I673990,I673982);
nor I_39467 (I673662,I673761,I673990);
or I_39468 (I674021,I673829,I427720);
nor I_39469 (I674038,I427720,I427705);
nand I_39470 (I674055,I673894,I674038);
nand I_39471 (I674072,I674021,I674055);
DFFARX1 I_39472 (I674072,I3035,I673676,I673665,);
nor I_39473 (I674103,I674038,I673795);
DFFARX1 I_39474 (I674103,I3035,I673676,I673644,);
nor I_39475 (I674134,I427720,I427711);
DFFARX1 I_39476 (I674134,I3035,I673676,I674160,);
DFFARX1 I_39477 (I674160,I3035,I673676,I673659,);
not I_39478 (I674182,I674160);
nand I_39479 (I673656,I674182,I673710);
nand I_39480 (I673650,I674182,I673812);
not I_39481 (I674254,I3042);
DFFARX1 I_39482 (I210383,I3035,I674254,I674280,);
nand I_39483 (I674288,I674280,I210404);
not I_39484 (I674305,I674288);
DFFARX1 I_39485 (I210398,I3035,I674254,I674331,);
not I_39486 (I674339,I674331);
not I_39487 (I674356,I210386);
or I_39488 (I674373,I210401,I210386);
nor I_39489 (I674390,I210401,I210386);
or I_39490 (I674407,I210392,I210401);
DFFARX1 I_39491 (I674407,I3035,I674254,I674246,);
not I_39492 (I674438,I210380);
nand I_39493 (I674455,I674438,I210377);
nand I_39494 (I674472,I674356,I674455);
and I_39495 (I674225,I674339,I674472);
nor I_39496 (I674503,I210380,I210389);
and I_39497 (I674520,I674339,I674503);
nor I_39498 (I674231,I674305,I674520);
DFFARX1 I_39499 (I674503,I3035,I674254,I674560,);
not I_39500 (I674568,I674560);
nor I_39501 (I674240,I674339,I674568);
or I_39502 (I674599,I674407,I210395);
nor I_39503 (I674616,I210395,I210392);
nand I_39504 (I674633,I674472,I674616);
nand I_39505 (I674650,I674599,I674633);
DFFARX1 I_39506 (I674650,I3035,I674254,I674243,);
nor I_39507 (I674681,I674616,I674373);
DFFARX1 I_39508 (I674681,I3035,I674254,I674222,);
nor I_39509 (I674712,I210395,I210377);
DFFARX1 I_39510 (I674712,I3035,I674254,I674738,);
DFFARX1 I_39511 (I674738,I3035,I674254,I674237,);
not I_39512 (I674760,I674738);
nand I_39513 (I674234,I674760,I674288);
nand I_39514 (I674228,I674760,I674390);
not I_39515 (I674832,I3042);
DFFARX1 I_39516 (I40491,I3035,I674832,I674858,);
nand I_39517 (I674866,I674858,I40482);
not I_39518 (I674883,I674866);
DFFARX1 I_39519 (I40479,I3035,I674832,I674909,);
not I_39520 (I674917,I674909);
not I_39521 (I674934,I40488);
or I_39522 (I674951,I40479,I40488);
nor I_39523 (I674968,I40479,I40488);
or I_39524 (I674985,I40485,I40479);
DFFARX1 I_39525 (I674985,I3035,I674832,I674824,);
not I_39526 (I675016,I40494);
nand I_39527 (I675033,I675016,I40503);
nand I_39528 (I675050,I674934,I675033);
and I_39529 (I674803,I674917,I675050);
nor I_39530 (I675081,I40494,I40497);
and I_39531 (I675098,I674917,I675081);
nor I_39532 (I674809,I674883,I675098);
DFFARX1 I_39533 (I675081,I3035,I674832,I675138,);
not I_39534 (I675146,I675138);
nor I_39535 (I674818,I674917,I675146);
or I_39536 (I675177,I674985,I40482);
nor I_39537 (I675194,I40482,I40485);
nand I_39538 (I675211,I675050,I675194);
nand I_39539 (I675228,I675177,I675211);
DFFARX1 I_39540 (I675228,I3035,I674832,I674821,);
nor I_39541 (I675259,I675194,I674951);
DFFARX1 I_39542 (I675259,I3035,I674832,I674800,);
nor I_39543 (I675290,I40482,I40500);
DFFARX1 I_39544 (I675290,I3035,I674832,I675316,);
DFFARX1 I_39545 (I675316,I3035,I674832,I674815,);
not I_39546 (I675338,I675316);
nand I_39547 (I674812,I675338,I674866);
nand I_39548 (I674806,I675338,I674968);
not I_39549 (I675410,I3042);
DFFARX1 I_39550 (I296601,I3035,I675410,I675436,);
nand I_39551 (I675444,I675436,I296610);
not I_39552 (I675461,I675444);
DFFARX1 I_39553 (I296622,I3035,I675410,I675487,);
not I_39554 (I675495,I675487);
not I_39555 (I675512,I296613);
or I_39556 (I675529,I296607,I296613);
nor I_39557 (I675546,I296607,I296613);
or I_39558 (I675563,I296601,I296607);
DFFARX1 I_39559 (I675563,I3035,I675410,I675402,);
not I_39560 (I675594,I296604);
nand I_39561 (I675611,I675594,I296616);
nand I_39562 (I675628,I675512,I675611);
and I_39563 (I675381,I675495,I675628);
nor I_39564 (I675659,I296604,I296625);
and I_39565 (I675676,I675495,I675659);
nor I_39566 (I675387,I675461,I675676);
DFFARX1 I_39567 (I675659,I3035,I675410,I675716,);
not I_39568 (I675724,I675716);
nor I_39569 (I675396,I675495,I675724);
or I_39570 (I675755,I675563,I296619);
nor I_39571 (I675772,I296619,I296601);
nand I_39572 (I675789,I675628,I675772);
nand I_39573 (I675806,I675755,I675789);
DFFARX1 I_39574 (I675806,I3035,I675410,I675399,);
nor I_39575 (I675837,I675772,I675529);
DFFARX1 I_39576 (I675837,I3035,I675410,I675378,);
nor I_39577 (I675868,I296619,I296604);
DFFARX1 I_39578 (I675868,I3035,I675410,I675894,);
DFFARX1 I_39579 (I675894,I3035,I675410,I675393,);
not I_39580 (I675916,I675894);
nand I_39581 (I675390,I675916,I675444);
nand I_39582 (I675384,I675916,I675546);
not I_39583 (I675988,I3042);
DFFARX1 I_39584 (I346972,I3035,I675988,I676014,);
nand I_39585 (I676022,I676014,I346975);
not I_39586 (I676039,I676022);
DFFARX1 I_39587 (I346987,I3035,I675988,I676065,);
not I_39588 (I676073,I676065);
not I_39589 (I676090,I346972);
or I_39590 (I676107,I346981,I346972);
nor I_39591 (I676124,I346981,I346972);
or I_39592 (I676141,I346990,I346981);
DFFARX1 I_39593 (I676141,I3035,I675988,I675980,);
not I_39594 (I676172,I346993);
nand I_39595 (I676189,I676172,I346975);
nand I_39596 (I676206,I676090,I676189);
and I_39597 (I675959,I676073,I676206);
nor I_39598 (I676237,I346993,I346978);
and I_39599 (I676254,I676073,I676237);
nor I_39600 (I675965,I676039,I676254);
DFFARX1 I_39601 (I676237,I3035,I675988,I676294,);
not I_39602 (I676302,I676294);
nor I_39603 (I675974,I676073,I676302);
or I_39604 (I676333,I676141,I346984);
nor I_39605 (I676350,I346984,I346990);
nand I_39606 (I676367,I676206,I676350);
nand I_39607 (I676384,I676333,I676367);
DFFARX1 I_39608 (I676384,I3035,I675988,I675977,);
nor I_39609 (I676415,I676350,I676107);
DFFARX1 I_39610 (I676415,I3035,I675988,I675956,);
nor I_39611 (I676446,I346984,I346996);
DFFARX1 I_39612 (I676446,I3035,I675988,I676472,);
DFFARX1 I_39613 (I676472,I3035,I675988,I675971,);
not I_39614 (I676494,I676472);
nand I_39615 (I675968,I676494,I676022);
nand I_39616 (I675962,I676494,I676124);
not I_39617 (I676566,I3042);
DFFARX1 I_39618 (I420330,I3035,I676566,I676592,);
nand I_39619 (I676600,I676592,I420330);
not I_39620 (I676617,I676600);
DFFARX1 I_39621 (I420336,I3035,I676566,I676643,);
not I_39622 (I676651,I676643);
not I_39623 (I676668,I420348);
or I_39624 (I676685,I420333,I420348);
nor I_39625 (I676702,I420333,I420348);
or I_39626 (I676719,I420327,I420333);
DFFARX1 I_39627 (I676719,I3035,I676566,I676558,);
not I_39628 (I676750,I420345);
nand I_39629 (I676767,I676750,I420339);
nand I_39630 (I676784,I676668,I676767);
and I_39631 (I676537,I676651,I676784);
nor I_39632 (I676815,I420345,I420327);
and I_39633 (I676832,I676651,I676815);
nor I_39634 (I676543,I676617,I676832);
DFFARX1 I_39635 (I676815,I3035,I676566,I676872,);
not I_39636 (I676880,I676872);
nor I_39637 (I676552,I676651,I676880);
or I_39638 (I676911,I676719,I420342);
nor I_39639 (I676928,I420342,I420327);
nand I_39640 (I676945,I676784,I676928);
nand I_39641 (I676962,I676911,I676945);
DFFARX1 I_39642 (I676962,I3035,I676566,I676555,);
nor I_39643 (I676993,I676928,I676685);
DFFARX1 I_39644 (I676993,I3035,I676566,I676534,);
nor I_39645 (I677024,I420342,I420333);
DFFARX1 I_39646 (I677024,I3035,I676566,I677050,);
DFFARX1 I_39647 (I677050,I3035,I676566,I676549,);
not I_39648 (I677072,I677050);
nand I_39649 (I676546,I677072,I676600);
nand I_39650 (I676540,I677072,I676702);
not I_39651 (I677144,I3042);
DFFARX1 I_39652 (I442991,I3035,I677144,I677170,);
nand I_39653 (I677178,I677170,I442991);
not I_39654 (I677195,I677178);
DFFARX1 I_39655 (I442997,I3035,I677144,I677221,);
not I_39656 (I677229,I677221);
not I_39657 (I677246,I443009);
or I_39658 (I677263,I442994,I443009);
nor I_39659 (I677280,I442994,I443009);
or I_39660 (I677297,I442988,I442994);
DFFARX1 I_39661 (I677297,I3035,I677144,I677136,);
not I_39662 (I677328,I443006);
nand I_39663 (I677345,I677328,I443000);
nand I_39664 (I677362,I677246,I677345);
and I_39665 (I677115,I677229,I677362);
nor I_39666 (I677393,I443006,I442988);
and I_39667 (I677410,I677229,I677393);
nor I_39668 (I677121,I677195,I677410);
DFFARX1 I_39669 (I677393,I3035,I677144,I677450,);
not I_39670 (I677458,I677450);
nor I_39671 (I677130,I677229,I677458);
or I_39672 (I677489,I677297,I443003);
nor I_39673 (I677506,I443003,I442988);
nand I_39674 (I677523,I677362,I677506);
nand I_39675 (I677540,I677489,I677523);
DFFARX1 I_39676 (I677540,I3035,I677144,I677133,);
nor I_39677 (I677571,I677506,I677263);
DFFARX1 I_39678 (I677571,I3035,I677144,I677112,);
nor I_39679 (I677602,I443003,I442994);
DFFARX1 I_39680 (I677602,I3035,I677144,I677628,);
DFFARX1 I_39681 (I677628,I3035,I677144,I677127,);
not I_39682 (I677650,I677628);
nand I_39683 (I677124,I677650,I677178);
nand I_39684 (I677118,I677650,I677280);
not I_39685 (I677722,I3042);
DFFARX1 I_39686 (I45761,I3035,I677722,I677748,);
nand I_39687 (I677756,I677748,I45752);
not I_39688 (I677773,I677756);
DFFARX1 I_39689 (I45749,I3035,I677722,I677799,);
not I_39690 (I677807,I677799);
not I_39691 (I677824,I45758);
or I_39692 (I677841,I45749,I45758);
nor I_39693 (I677858,I45749,I45758);
or I_39694 (I677875,I45755,I45749);
DFFARX1 I_39695 (I677875,I3035,I677722,I677714,);
not I_39696 (I677906,I45764);
nand I_39697 (I677923,I677906,I45773);
nand I_39698 (I677940,I677824,I677923);
and I_39699 (I677693,I677807,I677940);
nor I_39700 (I677971,I45764,I45767);
and I_39701 (I677988,I677807,I677971);
nor I_39702 (I677699,I677773,I677988);
DFFARX1 I_39703 (I677971,I3035,I677722,I678028,);
not I_39704 (I678036,I678028);
nor I_39705 (I677708,I677807,I678036);
or I_39706 (I678067,I677875,I45752);
nor I_39707 (I678084,I45752,I45755);
nand I_39708 (I678101,I677940,I678084);
nand I_39709 (I678118,I678067,I678101);
DFFARX1 I_39710 (I678118,I3035,I677722,I677711,);
nor I_39711 (I678149,I678084,I677841);
DFFARX1 I_39712 (I678149,I3035,I677722,I677690,);
nor I_39713 (I678180,I45752,I45770);
DFFARX1 I_39714 (I678180,I3035,I677722,I678206,);
DFFARX1 I_39715 (I678206,I3035,I677722,I677705,);
not I_39716 (I678228,I678206);
nand I_39717 (I677702,I678228,I677756);
nand I_39718 (I677696,I678228,I677858);
not I_39719 (I678300,I3042);
DFFARX1 I_39720 (I228828,I3035,I678300,I678326,);
nand I_39721 (I678334,I678326,I228849);
not I_39722 (I678351,I678334);
DFFARX1 I_39723 (I228843,I3035,I678300,I678377,);
not I_39724 (I678385,I678377);
not I_39725 (I678402,I228831);
or I_39726 (I678419,I228846,I228831);
nor I_39727 (I678436,I228846,I228831);
or I_39728 (I678453,I228837,I228846);
DFFARX1 I_39729 (I678453,I3035,I678300,I678292,);
not I_39730 (I678484,I228825);
nand I_39731 (I678501,I678484,I228822);
nand I_39732 (I678518,I678402,I678501);
and I_39733 (I678271,I678385,I678518);
nor I_39734 (I678549,I228825,I228834);
and I_39735 (I678566,I678385,I678549);
nor I_39736 (I678277,I678351,I678566);
DFFARX1 I_39737 (I678549,I3035,I678300,I678606,);
not I_39738 (I678614,I678606);
nor I_39739 (I678286,I678385,I678614);
or I_39740 (I678645,I678453,I228840);
nor I_39741 (I678662,I228840,I228837);
nand I_39742 (I678679,I678518,I678662);
nand I_39743 (I678696,I678645,I678679);
DFFARX1 I_39744 (I678696,I3035,I678300,I678289,);
nor I_39745 (I678727,I678662,I678419);
DFFARX1 I_39746 (I678727,I3035,I678300,I678268,);
nor I_39747 (I678758,I228840,I228822);
DFFARX1 I_39748 (I678758,I3035,I678300,I678784,);
DFFARX1 I_39749 (I678784,I3035,I678300,I678283,);
not I_39750 (I678806,I678784);
nand I_39751 (I678280,I678806,I678334);
nand I_39752 (I678274,I678806,I678436);
not I_39753 (I678878,I3042);
DFFARX1 I_39754 (I448788,I3035,I678878,I678904,);
nand I_39755 (I678912,I678904,I448788);
not I_39756 (I678929,I678912);
DFFARX1 I_39757 (I448794,I3035,I678878,I678955,);
not I_39758 (I678963,I678955);
not I_39759 (I678980,I448806);
or I_39760 (I678997,I448791,I448806);
nor I_39761 (I679014,I448791,I448806);
or I_39762 (I679031,I448785,I448791);
DFFARX1 I_39763 (I679031,I3035,I678878,I678870,);
not I_39764 (I679062,I448803);
nand I_39765 (I679079,I679062,I448797);
nand I_39766 (I679096,I678980,I679079);
and I_39767 (I678849,I678963,I679096);
nor I_39768 (I679127,I448803,I448785);
and I_39769 (I679144,I678963,I679127);
nor I_39770 (I678855,I678929,I679144);
DFFARX1 I_39771 (I679127,I3035,I678878,I679184,);
not I_39772 (I679192,I679184);
nor I_39773 (I678864,I678963,I679192);
or I_39774 (I679223,I679031,I448800);
nor I_39775 (I679240,I448800,I448785);
nand I_39776 (I679257,I679096,I679240);
nand I_39777 (I679274,I679223,I679257);
DFFARX1 I_39778 (I679274,I3035,I678878,I678867,);
nor I_39779 (I679305,I679240,I678997);
DFFARX1 I_39780 (I679305,I3035,I678878,I678846,);
nor I_39781 (I679336,I448800,I448791);
DFFARX1 I_39782 (I679336,I3035,I678878,I679362,);
DFFARX1 I_39783 (I679362,I3035,I678878,I678861,);
not I_39784 (I679384,I679362);
nand I_39785 (I678858,I679384,I678912);
nand I_39786 (I678852,I679384,I679014);
not I_39787 (I679456,I3042);
DFFARX1 I_39788 (I709147,I3035,I679456,I679482,);
nand I_39789 (I679490,I679482,I709138);
not I_39790 (I679507,I679490);
DFFARX1 I_39791 (I709123,I3035,I679456,I679533,);
not I_39792 (I679541,I679533);
not I_39793 (I679558,I709126);
or I_39794 (I679575,I709135,I709126);
nor I_39795 (I679592,I709135,I709126);
or I_39796 (I679609,I709132,I709135);
DFFARX1 I_39797 (I679609,I3035,I679456,I679448,);
not I_39798 (I679640,I709144);
nand I_39799 (I679657,I679640,I709123);
nand I_39800 (I679674,I679558,I679657);
and I_39801 (I679427,I679541,I679674);
nor I_39802 (I679705,I709144,I709129);
and I_39803 (I679722,I679541,I679705);
nor I_39804 (I679433,I679507,I679722);
DFFARX1 I_39805 (I679705,I3035,I679456,I679762,);
not I_39806 (I679770,I679762);
nor I_39807 (I679442,I679541,I679770);
or I_39808 (I679801,I679609,I709150);
nor I_39809 (I679818,I709150,I709132);
nand I_39810 (I679835,I679674,I679818);
nand I_39811 (I679852,I679801,I679835);
DFFARX1 I_39812 (I679852,I3035,I679456,I679445,);
nor I_39813 (I679883,I679818,I679575);
DFFARX1 I_39814 (I679883,I3035,I679456,I679424,);
nor I_39815 (I679914,I709150,I709141);
DFFARX1 I_39816 (I679914,I3035,I679456,I679940,);
DFFARX1 I_39817 (I679940,I3035,I679456,I679439,);
not I_39818 (I679962,I679940);
nand I_39819 (I679436,I679962,I679490);
nand I_39820 (I679430,I679962,I679592);
not I_39821 (I680034,I3042);
DFFARX1 I_39822 (I43653,I3035,I680034,I680060,);
nand I_39823 (I680068,I680060,I43644);
not I_39824 (I680085,I680068);
DFFARX1 I_39825 (I43641,I3035,I680034,I680111,);
not I_39826 (I680119,I680111);
not I_39827 (I680136,I43650);
or I_39828 (I680153,I43641,I43650);
nor I_39829 (I680170,I43641,I43650);
or I_39830 (I680187,I43647,I43641);
DFFARX1 I_39831 (I680187,I3035,I680034,I680026,);
not I_39832 (I680218,I43656);
nand I_39833 (I680235,I680218,I43665);
nand I_39834 (I680252,I680136,I680235);
and I_39835 (I680005,I680119,I680252);
nor I_39836 (I680283,I43656,I43659);
and I_39837 (I680300,I680119,I680283);
nor I_39838 (I680011,I680085,I680300);
DFFARX1 I_39839 (I680283,I3035,I680034,I680340,);
not I_39840 (I680348,I680340);
nor I_39841 (I680020,I680119,I680348);
or I_39842 (I680379,I680187,I43644);
nor I_39843 (I680396,I43644,I43647);
nand I_39844 (I680413,I680252,I680396);
nand I_39845 (I680430,I680379,I680413);
DFFARX1 I_39846 (I680430,I3035,I680034,I680023,);
nor I_39847 (I680461,I680396,I680153);
DFFARX1 I_39848 (I680461,I3035,I680034,I680002,);
nor I_39849 (I680492,I43644,I43662);
DFFARX1 I_39850 (I680492,I3035,I680034,I680518,);
DFFARX1 I_39851 (I680518,I3035,I680034,I680017,);
not I_39852 (I680540,I680518);
nand I_39853 (I680014,I680540,I680068);
nand I_39854 (I680008,I680540,I680170);
not I_39855 (I680612,I3042);
DFFARX1 I_39856 (I639356,I3035,I680612,I680638,);
nand I_39857 (I680646,I680638,I639341);
not I_39858 (I680663,I680646);
DFFARX1 I_39859 (I639344,I3035,I680612,I680689,);
not I_39860 (I680697,I680689);
not I_39861 (I680714,I639359);
or I_39862 (I680731,I639362,I639359);
nor I_39863 (I680748,I639362,I639359);
or I_39864 (I680765,I639338,I639362);
DFFARX1 I_39865 (I680765,I3035,I680612,I680604,);
not I_39866 (I680796,I639350);
nand I_39867 (I680813,I680796,I639353);
nand I_39868 (I680830,I680714,I680813);
and I_39869 (I680583,I680697,I680830);
nor I_39870 (I680861,I639350,I639347);
and I_39871 (I680878,I680697,I680861);
nor I_39872 (I680589,I680663,I680878);
DFFARX1 I_39873 (I680861,I3035,I680612,I680918,);
not I_39874 (I680926,I680918);
nor I_39875 (I680598,I680697,I680926);
or I_39876 (I680957,I680765,I639338);
nor I_39877 (I680974,I639338,I639338);
nand I_39878 (I680991,I680830,I680974);
nand I_39879 (I681008,I680957,I680991);
DFFARX1 I_39880 (I681008,I3035,I680612,I680601,);
nor I_39881 (I681039,I680974,I680731);
DFFARX1 I_39882 (I681039,I3035,I680612,I680580,);
nor I_39883 (I681070,I639338,I639341);
DFFARX1 I_39884 (I681070,I3035,I680612,I681096,);
DFFARX1 I_39885 (I681096,I3035,I680612,I680595,);
not I_39886 (I681118,I681096);
nand I_39887 (I680592,I681118,I680646);
nand I_39888 (I680586,I681118,I680748);
not I_39889 (I681190,I3042);
DFFARX1 I_39890 (I599474,I3035,I681190,I681216,);
nand I_39891 (I681224,I681216,I599459);
not I_39892 (I681241,I681224);
DFFARX1 I_39893 (I599462,I3035,I681190,I681267,);
not I_39894 (I681275,I681267);
not I_39895 (I681292,I599477);
or I_39896 (I681309,I599480,I599477);
nor I_39897 (I681326,I599480,I599477);
or I_39898 (I681343,I599456,I599480);
DFFARX1 I_39899 (I681343,I3035,I681190,I681182,);
not I_39900 (I681374,I599468);
nand I_39901 (I681391,I681374,I599471);
nand I_39902 (I681408,I681292,I681391);
and I_39903 (I681161,I681275,I681408);
nor I_39904 (I681439,I599468,I599465);
and I_39905 (I681456,I681275,I681439);
nor I_39906 (I681167,I681241,I681456);
DFFARX1 I_39907 (I681439,I3035,I681190,I681496,);
not I_39908 (I681504,I681496);
nor I_39909 (I681176,I681275,I681504);
or I_39910 (I681535,I681343,I599456);
nor I_39911 (I681552,I599456,I599456);
nand I_39912 (I681569,I681408,I681552);
nand I_39913 (I681586,I681535,I681569);
DFFARX1 I_39914 (I681586,I3035,I681190,I681179,);
nor I_39915 (I681617,I681552,I681309);
DFFARX1 I_39916 (I681617,I3035,I681190,I681158,);
nor I_39917 (I681648,I599456,I599459);
DFFARX1 I_39918 (I681648,I3035,I681190,I681674,);
DFFARX1 I_39919 (I681674,I3035,I681190,I681173,);
not I_39920 (I681696,I681674);
nand I_39921 (I681170,I681696,I681224);
nand I_39922 (I681164,I681696,I681326);
not I_39923 (I681768,I3042);
DFFARX1 I_39924 (I257096,I3035,I681768,I681794,);
nand I_39925 (I681802,I681794,I257105);
not I_39926 (I681819,I681802);
DFFARX1 I_39927 (I257093,I3035,I681768,I681845,);
not I_39928 (I681853,I681845);
not I_39929 (I681870,I257099);
or I_39930 (I681887,I257093,I257099);
nor I_39931 (I681904,I257093,I257099);
or I_39932 (I681921,I257108,I257093);
DFFARX1 I_39933 (I681921,I3035,I681768,I681760,);
not I_39934 (I681952,I257102);
nand I_39935 (I681969,I681952,I257117);
nand I_39936 (I681986,I681870,I681969);
and I_39937 (I681739,I681853,I681986);
nor I_39938 (I682017,I257102,I257120);
and I_39939 (I682034,I681853,I682017);
nor I_39940 (I681745,I681819,I682034);
DFFARX1 I_39941 (I682017,I3035,I681768,I682074,);
not I_39942 (I682082,I682074);
nor I_39943 (I681754,I681853,I682082);
or I_39944 (I682113,I681921,I257111);
nor I_39945 (I682130,I257111,I257108);
nand I_39946 (I682147,I681986,I682130);
nand I_39947 (I682164,I682113,I682147);
DFFARX1 I_39948 (I682164,I3035,I681768,I681757,);
nor I_39949 (I682195,I682130,I681887);
DFFARX1 I_39950 (I682195,I3035,I681768,I681736,);
nor I_39951 (I682226,I257111,I257114);
DFFARX1 I_39952 (I682226,I3035,I681768,I682252,);
DFFARX1 I_39953 (I682252,I3035,I681768,I681751,);
not I_39954 (I682274,I682252);
nand I_39955 (I681748,I682274,I681802);
nand I_39956 (I681742,I682274,I681904);
not I_39957 (I682346,I3042);
DFFARX1 I_39958 (I173493,I3035,I682346,I682372,);
nand I_39959 (I682380,I682372,I173514);
not I_39960 (I682397,I682380);
DFFARX1 I_39961 (I173508,I3035,I682346,I682423,);
not I_39962 (I682431,I682423);
not I_39963 (I682448,I173496);
or I_39964 (I682465,I173511,I173496);
nor I_39965 (I682482,I173511,I173496);
or I_39966 (I682499,I173502,I173511);
DFFARX1 I_39967 (I682499,I3035,I682346,I682338,);
not I_39968 (I682530,I173490);
nand I_39969 (I682547,I682530,I173487);
nand I_39970 (I682564,I682448,I682547);
and I_39971 (I682317,I682431,I682564);
nor I_39972 (I682595,I173490,I173499);
and I_39973 (I682612,I682431,I682595);
nor I_39974 (I682323,I682397,I682612);
DFFARX1 I_39975 (I682595,I3035,I682346,I682652,);
not I_39976 (I682660,I682652);
nor I_39977 (I682332,I682431,I682660);
or I_39978 (I682691,I682499,I173505);
nor I_39979 (I682708,I173505,I173502);
nand I_39980 (I682725,I682564,I682708);
nand I_39981 (I682742,I682691,I682725);
DFFARX1 I_39982 (I682742,I3035,I682346,I682335,);
nor I_39983 (I682773,I682708,I682465);
DFFARX1 I_39984 (I682773,I3035,I682346,I682314,);
nor I_39985 (I682804,I173505,I173487);
DFFARX1 I_39986 (I682804,I3035,I682346,I682830,);
DFFARX1 I_39987 (I682830,I3035,I682346,I682329,);
not I_39988 (I682852,I682830);
nand I_39989 (I682326,I682852,I682380);
nand I_39990 (I682320,I682852,I682482);
not I_39991 (I682924,I3042);
DFFARX1 I_39992 (I226193,I3035,I682924,I682950,);
nand I_39993 (I682958,I682950,I226214);
not I_39994 (I682975,I682958);
DFFARX1 I_39995 (I226208,I3035,I682924,I683001,);
not I_39996 (I683009,I683001);
not I_39997 (I683026,I226196);
or I_39998 (I683043,I226211,I226196);
nor I_39999 (I683060,I226211,I226196);
or I_40000 (I683077,I226202,I226211);
DFFARX1 I_40001 (I683077,I3035,I682924,I682916,);
not I_40002 (I683108,I226190);
nand I_40003 (I683125,I683108,I226187);
nand I_40004 (I683142,I683026,I683125);
and I_40005 (I682895,I683009,I683142);
nor I_40006 (I683173,I226190,I226199);
and I_40007 (I683190,I683009,I683173);
nor I_40008 (I682901,I682975,I683190);
DFFARX1 I_40009 (I683173,I3035,I682924,I683230,);
not I_40010 (I683238,I683230);
nor I_40011 (I682910,I683009,I683238);
or I_40012 (I683269,I683077,I226205);
nor I_40013 (I683286,I226205,I226202);
nand I_40014 (I683303,I683142,I683286);
nand I_40015 (I683320,I683269,I683303);
DFFARX1 I_40016 (I683320,I3035,I682924,I682913,);
nor I_40017 (I683351,I683286,I683043);
DFFARX1 I_40018 (I683351,I3035,I682924,I682892,);
nor I_40019 (I683382,I226205,I226187);
DFFARX1 I_40020 (I683382,I3035,I682924,I683408,);
DFFARX1 I_40021 (I683408,I3035,I682924,I682907,);
not I_40022 (I683430,I683408);
nand I_40023 (I682904,I683430,I682958);
nand I_40024 (I682898,I683430,I683060);
not I_40025 (I683502,I3042);
DFFARX1 I_40026 (I571177,I3035,I683502,I683528,);
nand I_40027 (I683536,I683528,I571174);
not I_40028 (I683553,I683536);
DFFARX1 I_40029 (I571174,I3035,I683502,I683579,);
not I_40030 (I683587,I683579);
not I_40031 (I683604,I571171);
or I_40032 (I683621,I571180,I571171);
nor I_40033 (I683638,I571180,I571171);
or I_40034 (I683655,I571183,I571180);
DFFARX1 I_40035 (I683655,I3035,I683502,I683494,);
not I_40036 (I683686,I571171);
nand I_40037 (I683703,I683686,I571168);
nand I_40038 (I683720,I683604,I683703);
and I_40039 (I683473,I683587,I683720);
nor I_40040 (I683751,I571171,I571186);
and I_40041 (I683768,I683587,I683751);
nor I_40042 (I683479,I683553,I683768);
DFFARX1 I_40043 (I683751,I3035,I683502,I683808,);
not I_40044 (I683816,I683808);
nor I_40045 (I683488,I683587,I683816);
or I_40046 (I683847,I683655,I571189);
nor I_40047 (I683864,I571189,I571183);
nand I_40048 (I683881,I683720,I683864);
nand I_40049 (I683898,I683847,I683881);
DFFARX1 I_40050 (I683898,I3035,I683502,I683491,);
nor I_40051 (I683929,I683864,I683621);
DFFARX1 I_40052 (I683929,I3035,I683502,I683470,);
nor I_40053 (I683960,I571189,I571168);
DFFARX1 I_40054 (I683960,I3035,I683502,I683986,);
DFFARX1 I_40055 (I683986,I3035,I683502,I683485,);
not I_40056 (I684008,I683986);
nand I_40057 (I683482,I684008,I683536);
nand I_40058 (I683476,I684008,I683638);
not I_40059 (I684080,I3042);
DFFARX1 I_40060 (I300735,I3035,I684080,I684106,);
nand I_40061 (I684114,I684106,I300750);
not I_40062 (I684131,I684114);
DFFARX1 I_40063 (I300732,I3035,I684080,I684157,);
not I_40064 (I684165,I684157);
not I_40065 (I684182,I300741);
or I_40066 (I684199,I300735,I300741);
nor I_40067 (I684216,I300735,I300741);
or I_40068 (I684233,I300732,I300735);
DFFARX1 I_40069 (I684233,I3035,I684080,I684072,);
not I_40070 (I684264,I300753);
nand I_40071 (I684281,I684264,I300756);
nand I_40072 (I684298,I684182,I684281);
and I_40073 (I684051,I684165,I684298);
nor I_40074 (I684329,I300753,I300738);
and I_40075 (I684346,I684165,I684329);
nor I_40076 (I684057,I684131,I684346);
DFFARX1 I_40077 (I684329,I3035,I684080,I684386,);
not I_40078 (I684394,I684386);
nor I_40079 (I684066,I684165,I684394);
or I_40080 (I684425,I684233,I300744);
nor I_40081 (I684442,I300744,I300732);
nand I_40082 (I684459,I684298,I684442);
nand I_40083 (I684476,I684425,I684459);
DFFARX1 I_40084 (I684476,I3035,I684080,I684069,);
nor I_40085 (I684507,I684442,I684199);
DFFARX1 I_40086 (I684507,I3035,I684080,I684048,);
nor I_40087 (I684538,I300744,I300747);
DFFARX1 I_40088 (I684538,I3035,I684080,I684564,);
DFFARX1 I_40089 (I684564,I3035,I684080,I684063,);
not I_40090 (I684586,I684564);
nand I_40091 (I684060,I684586,I684114);
nand I_40092 (I684054,I684586,I684216);
not I_40093 (I684658,I3042);
DFFARX1 I_40094 (I28364,I3035,I684658,I684684,);
nand I_40095 (I684692,I684684,I28358);
not I_40096 (I684709,I684692);
DFFARX1 I_40097 (I28376,I3035,I684658,I684735,);
not I_40098 (I684743,I684735);
not I_40099 (I684760,I28379);
or I_40100 (I684777,I28382,I28379);
nor I_40101 (I684794,I28382,I28379);
or I_40102 (I684811,I28367,I28382);
DFFARX1 I_40103 (I684811,I3035,I684658,I684650,);
not I_40104 (I684842,I28370);
nand I_40105 (I684859,I684842,I28373);
nand I_40106 (I684876,I684760,I684859);
and I_40107 (I684629,I684743,I684876);
nor I_40108 (I684907,I28370,I28361);
and I_40109 (I684924,I684743,I684907);
nor I_40110 (I684635,I684709,I684924);
DFFARX1 I_40111 (I684907,I3035,I684658,I684964,);
not I_40112 (I684972,I684964);
nor I_40113 (I684644,I684743,I684972);
or I_40114 (I685003,I684811,I28361);
nor I_40115 (I685020,I28361,I28367);
nand I_40116 (I685037,I684876,I685020);
nand I_40117 (I685054,I685003,I685037);
DFFARX1 I_40118 (I685054,I3035,I684658,I684647,);
nor I_40119 (I685085,I685020,I684777);
DFFARX1 I_40120 (I685085,I3035,I684658,I684626,);
nor I_40121 (I685116,I28361,I28358);
DFFARX1 I_40122 (I685116,I3035,I684658,I685142,);
DFFARX1 I_40123 (I685142,I3035,I684658,I684641,);
not I_40124 (I685164,I685142);
nand I_40125 (I684638,I685164,I684692);
nand I_40126 (I684632,I685164,I684794);
not I_40127 (I685236,I3042);
DFFARX1 I_40128 (I570616,I3035,I685236,I685262,);
nand I_40129 (I685270,I685262,I570613);
not I_40130 (I685287,I685270);
DFFARX1 I_40131 (I570613,I3035,I685236,I685313,);
not I_40132 (I685321,I685313);
not I_40133 (I685338,I570610);
or I_40134 (I685355,I570619,I570610);
nor I_40135 (I685372,I570619,I570610);
or I_40136 (I685389,I570622,I570619);
DFFARX1 I_40137 (I685389,I3035,I685236,I685228,);
not I_40138 (I685420,I570610);
nand I_40139 (I685437,I685420,I570607);
nand I_40140 (I685454,I685338,I685437);
and I_40141 (I685207,I685321,I685454);
nor I_40142 (I685485,I570610,I570625);
and I_40143 (I685502,I685321,I685485);
nor I_40144 (I685213,I685287,I685502);
DFFARX1 I_40145 (I685485,I3035,I685236,I685542,);
not I_40146 (I685550,I685542);
nor I_40147 (I685222,I685321,I685550);
or I_40148 (I685581,I685389,I570628);
nor I_40149 (I685598,I570628,I570622);
nand I_40150 (I685615,I685454,I685598);
nand I_40151 (I685632,I685581,I685615);
DFFARX1 I_40152 (I685632,I3035,I685236,I685225,);
nor I_40153 (I685663,I685598,I685355);
DFFARX1 I_40154 (I685663,I3035,I685236,I685204,);
nor I_40155 (I685694,I570628,I570607);
DFFARX1 I_40156 (I685694,I3035,I685236,I685720,);
DFFARX1 I_40157 (I685720,I3035,I685236,I685219,);
not I_40158 (I685742,I685720);
nand I_40159 (I685216,I685742,I685270);
nand I_40160 (I685210,I685742,I685372);
not I_40161 (I685814,I3042);
DFFARX1 I_40162 (I591960,I3035,I685814,I685840,);
nand I_40163 (I685848,I685840,I591945);
not I_40164 (I685865,I685848);
DFFARX1 I_40165 (I591948,I3035,I685814,I685891,);
not I_40166 (I685899,I685891);
not I_40167 (I685916,I591963);
or I_40168 (I685933,I591966,I591963);
nor I_40169 (I685950,I591966,I591963);
or I_40170 (I685967,I591942,I591966);
DFFARX1 I_40171 (I685967,I3035,I685814,I685806,);
not I_40172 (I685998,I591954);
nand I_40173 (I686015,I685998,I591957);
nand I_40174 (I686032,I685916,I686015);
and I_40175 (I685785,I685899,I686032);
nor I_40176 (I686063,I591954,I591951);
and I_40177 (I686080,I685899,I686063);
nor I_40178 (I685791,I685865,I686080);
DFFARX1 I_40179 (I686063,I3035,I685814,I686120,);
not I_40180 (I686128,I686120);
nor I_40181 (I685800,I685899,I686128);
or I_40182 (I686159,I685967,I591942);
nor I_40183 (I686176,I591942,I591942);
nand I_40184 (I686193,I686032,I686176);
nand I_40185 (I686210,I686159,I686193);
DFFARX1 I_40186 (I686210,I3035,I685814,I685803,);
nor I_40187 (I686241,I686176,I685933);
DFFARX1 I_40188 (I686241,I3035,I685814,I685782,);
nor I_40189 (I686272,I591942,I591945);
DFFARX1 I_40190 (I686272,I3035,I685814,I686298,);
DFFARX1 I_40191 (I686298,I3035,I685814,I685797,);
not I_40192 (I686320,I686298);
nand I_40193 (I685794,I686320,I685848);
nand I_40194 (I685788,I686320,I685950);
not I_40195 (I686392,I3042);
DFFARX1 I_40196 (I501916,I3035,I686392,I686418,);
nand I_40197 (I686426,I686418,I501937);
not I_40198 (I686443,I686426);
DFFARX1 I_40199 (I501910,I3035,I686392,I686469,);
not I_40200 (I686477,I686469);
not I_40201 (I686494,I501931);
or I_40202 (I686511,I501922,I501931);
nor I_40203 (I686528,I501922,I501931);
or I_40204 (I686545,I501925,I501922);
DFFARX1 I_40205 (I686545,I3035,I686392,I686384,);
not I_40206 (I686576,I501913);
nand I_40207 (I686593,I686576,I501928);
nand I_40208 (I686610,I686494,I686593);
and I_40209 (I686363,I686477,I686610);
nor I_40210 (I686641,I501913,I501910);
and I_40211 (I686658,I686477,I686641);
nor I_40212 (I686369,I686443,I686658);
DFFARX1 I_40213 (I686641,I3035,I686392,I686698,);
not I_40214 (I686706,I686698);
nor I_40215 (I686378,I686477,I686706);
or I_40216 (I686737,I686545,I501934);
nor I_40217 (I686754,I501934,I501925);
nand I_40218 (I686771,I686610,I686754);
nand I_40219 (I686788,I686737,I686771);
DFFARX1 I_40220 (I686788,I3035,I686392,I686381,);
nor I_40221 (I686819,I686754,I686511);
DFFARX1 I_40222 (I686819,I3035,I686392,I686360,);
nor I_40223 (I686850,I501934,I501919);
DFFARX1 I_40224 (I686850,I3035,I686392,I686876,);
DFFARX1 I_40225 (I686876,I3035,I686392,I686375,);
not I_40226 (I686898,I686876);
nand I_40227 (I686372,I686898,I686426);
nand I_40228 (I686366,I686898,I686528);
not I_40229 (I686970,I3042);
DFFARX1 I_40230 (I265800,I3035,I686970,I686996,);
nand I_40231 (I687004,I686996,I265809);
not I_40232 (I687021,I687004);
DFFARX1 I_40233 (I265797,I3035,I686970,I687047,);
not I_40234 (I687055,I687047);
not I_40235 (I687072,I265803);
or I_40236 (I687089,I265797,I265803);
nor I_40237 (I687106,I265797,I265803);
or I_40238 (I687123,I265812,I265797);
DFFARX1 I_40239 (I687123,I3035,I686970,I686962,);
not I_40240 (I687154,I265806);
nand I_40241 (I687171,I687154,I265821);
nand I_40242 (I687188,I687072,I687171);
and I_40243 (I686941,I687055,I687188);
nor I_40244 (I687219,I265806,I265824);
and I_40245 (I687236,I687055,I687219);
nor I_40246 (I686947,I687021,I687236);
DFFARX1 I_40247 (I687219,I3035,I686970,I687276,);
not I_40248 (I687284,I687276);
nor I_40249 (I686956,I687055,I687284);
or I_40250 (I687315,I687123,I265815);
nor I_40251 (I687332,I265815,I265812);
nand I_40252 (I687349,I687188,I687332);
nand I_40253 (I687366,I687315,I687349);
DFFARX1 I_40254 (I687366,I3035,I686970,I686959,);
nor I_40255 (I687397,I687332,I687089);
DFFARX1 I_40256 (I687397,I3035,I686970,I686938,);
nor I_40257 (I687428,I265815,I265818);
DFFARX1 I_40258 (I687428,I3035,I686970,I687454,);
DFFARX1 I_40259 (I687454,I3035,I686970,I686953,);
not I_40260 (I687476,I687454);
nand I_40261 (I686950,I687476,I687004);
nand I_40262 (I686944,I687476,I687106);
not I_40263 (I687548,I3042);
DFFARX1 I_40264 (I732947,I3035,I687548,I687574,);
nand I_40265 (I687582,I687574,I732938);
not I_40266 (I687599,I687582);
DFFARX1 I_40267 (I732923,I3035,I687548,I687625,);
not I_40268 (I687633,I687625);
not I_40269 (I687650,I732926);
or I_40270 (I687667,I732935,I732926);
nor I_40271 (I687684,I732935,I732926);
or I_40272 (I687701,I732932,I732935);
DFFARX1 I_40273 (I687701,I3035,I687548,I687540,);
not I_40274 (I687732,I732944);
nand I_40275 (I687749,I687732,I732923);
nand I_40276 (I687766,I687650,I687749);
and I_40277 (I687519,I687633,I687766);
nor I_40278 (I687797,I732944,I732929);
and I_40279 (I687814,I687633,I687797);
nor I_40280 (I687525,I687599,I687814);
DFFARX1 I_40281 (I687797,I3035,I687548,I687854,);
not I_40282 (I687862,I687854);
nor I_40283 (I687534,I687633,I687862);
or I_40284 (I687893,I687701,I732950);
nor I_40285 (I687910,I732950,I732932);
nand I_40286 (I687927,I687766,I687910);
nand I_40287 (I687944,I687893,I687927);
DFFARX1 I_40288 (I687944,I3035,I687548,I687537,);
nor I_40289 (I687975,I687910,I687667);
DFFARX1 I_40290 (I687975,I3035,I687548,I687516,);
nor I_40291 (I688006,I732950,I732941);
DFFARX1 I_40292 (I688006,I3035,I687548,I688032,);
DFFARX1 I_40293 (I688032,I3035,I687548,I687531,);
not I_40294 (I688054,I688032);
nand I_40295 (I687528,I688054,I687582);
nand I_40296 (I687522,I688054,I687684);
not I_40297 (I688126,I3042);
DFFARX1 I_40298 (I213545,I3035,I688126,I688152,);
nand I_40299 (I688160,I688152,I213566);
not I_40300 (I688177,I688160);
DFFARX1 I_40301 (I213560,I3035,I688126,I688203,);
not I_40302 (I688211,I688203);
not I_40303 (I688228,I213548);
or I_40304 (I688245,I213563,I213548);
nor I_40305 (I688262,I213563,I213548);
or I_40306 (I688279,I213554,I213563);
DFFARX1 I_40307 (I688279,I3035,I688126,I688118,);
not I_40308 (I688310,I213542);
nand I_40309 (I688327,I688310,I213539);
nand I_40310 (I688344,I688228,I688327);
and I_40311 (I688097,I688211,I688344);
nor I_40312 (I688375,I213542,I213551);
and I_40313 (I688392,I688211,I688375);
nor I_40314 (I688103,I688177,I688392);
DFFARX1 I_40315 (I688375,I3035,I688126,I688432,);
not I_40316 (I688440,I688432);
nor I_40317 (I688112,I688211,I688440);
or I_40318 (I688471,I688279,I213557);
nor I_40319 (I688488,I213557,I213554);
nand I_40320 (I688505,I688344,I688488);
nand I_40321 (I688522,I688471,I688505);
DFFARX1 I_40322 (I688522,I3035,I688126,I688115,);
nor I_40323 (I688553,I688488,I688245);
DFFARX1 I_40324 (I688553,I3035,I688126,I688094,);
nor I_40325 (I688584,I213557,I213539);
DFFARX1 I_40326 (I688584,I3035,I688126,I688610,);
DFFARX1 I_40327 (I688610,I3035,I688126,I688109,);
not I_40328 (I688632,I688610);
nand I_40329 (I688106,I688632,I688160);
nand I_40330 (I688100,I688632,I688262);
not I_40331 (I688704,I3042);
DFFARX1 I_40332 (I471976,I3035,I688704,I688730,);
nand I_40333 (I688738,I688730,I471976);
not I_40334 (I688755,I688738);
DFFARX1 I_40335 (I471982,I3035,I688704,I688781,);
not I_40336 (I688789,I688781);
not I_40337 (I688806,I471994);
or I_40338 (I688823,I471979,I471994);
nor I_40339 (I688840,I471979,I471994);
or I_40340 (I688857,I471973,I471979);
DFFARX1 I_40341 (I688857,I3035,I688704,I688696,);
not I_40342 (I688888,I471991);
nand I_40343 (I688905,I688888,I471985);
nand I_40344 (I688922,I688806,I688905);
and I_40345 (I688675,I688789,I688922);
nor I_40346 (I688953,I471991,I471973);
and I_40347 (I688970,I688789,I688953);
nor I_40348 (I688681,I688755,I688970);
DFFARX1 I_40349 (I688953,I3035,I688704,I689010,);
not I_40350 (I689018,I689010);
nor I_40351 (I688690,I688789,I689018);
or I_40352 (I689049,I688857,I471988);
nor I_40353 (I689066,I471988,I471973);
nand I_40354 (I689083,I688922,I689066);
nand I_40355 (I689100,I689049,I689083);
DFFARX1 I_40356 (I689100,I3035,I688704,I688693,);
nor I_40357 (I689131,I689066,I688823);
DFFARX1 I_40358 (I689131,I3035,I688704,I688672,);
nor I_40359 (I689162,I471988,I471979);
DFFARX1 I_40360 (I689162,I3035,I688704,I689188,);
DFFARX1 I_40361 (I689188,I3035,I688704,I688687,);
not I_40362 (I689210,I689188);
nand I_40363 (I688684,I689210,I688738);
nand I_40364 (I688678,I689210,I688840);
not I_40365 (I689282,I3042);
DFFARX1 I_40366 (I26783,I3035,I689282,I689308,);
nand I_40367 (I689316,I689308,I26777);
not I_40368 (I689333,I689316);
DFFARX1 I_40369 (I26795,I3035,I689282,I689359,);
not I_40370 (I689367,I689359);
not I_40371 (I689384,I26798);
or I_40372 (I689401,I26801,I26798);
nor I_40373 (I689418,I26801,I26798);
or I_40374 (I689435,I26786,I26801);
DFFARX1 I_40375 (I689435,I3035,I689282,I689274,);
not I_40376 (I689466,I26789);
nand I_40377 (I689483,I689466,I26792);
nand I_40378 (I689500,I689384,I689483);
and I_40379 (I689253,I689367,I689500);
nor I_40380 (I689531,I26789,I26780);
and I_40381 (I689548,I689367,I689531);
nor I_40382 (I689259,I689333,I689548);
DFFARX1 I_40383 (I689531,I3035,I689282,I689588,);
not I_40384 (I689596,I689588);
nor I_40385 (I689268,I689367,I689596);
or I_40386 (I689627,I689435,I26780);
nor I_40387 (I689644,I26780,I26786);
nand I_40388 (I689661,I689500,I689644);
nand I_40389 (I689678,I689627,I689661);
DFFARX1 I_40390 (I689678,I3035,I689282,I689271,);
nor I_40391 (I689709,I689644,I689401);
DFFARX1 I_40392 (I689709,I3035,I689282,I689250,);
nor I_40393 (I689740,I26780,I26777);
DFFARX1 I_40394 (I689740,I3035,I689282,I689766,);
DFFARX1 I_40395 (I689766,I3035,I689282,I689265,);
not I_40396 (I689788,I689766);
nand I_40397 (I689262,I689788,I689316);
nand I_40398 (I689256,I689788,I689418);
not I_40399 (I689860,I3042);
DFFARX1 I_40400 (I115194,I3035,I689860,I689886,);
nand I_40401 (I689894,I689886,I115197);
not I_40402 (I689911,I689894);
DFFARX1 I_40403 (I115206,I3035,I689860,I689937,);
not I_40404 (I689945,I689937);
not I_40405 (I689962,I115209);
or I_40406 (I689979,I115200,I115209);
nor I_40407 (I689996,I115200,I115209);
or I_40408 (I690013,I115212,I115200);
DFFARX1 I_40409 (I690013,I3035,I689860,I689852,);
not I_40410 (I690044,I115197);
nand I_40411 (I690061,I690044,I115203);
nand I_40412 (I690078,I689962,I690061);
and I_40413 (I689831,I689945,I690078);
nor I_40414 (I690109,I115197,I115215);
and I_40415 (I690126,I689945,I690109);
nor I_40416 (I689837,I689911,I690126);
DFFARX1 I_40417 (I690109,I3035,I689860,I690166,);
not I_40418 (I690174,I690166);
nor I_40419 (I689846,I689945,I690174);
or I_40420 (I690205,I690013,I115194);
nor I_40421 (I690222,I115194,I115212);
nand I_40422 (I690239,I690078,I690222);
nand I_40423 (I690256,I690205,I690239);
DFFARX1 I_40424 (I690256,I3035,I689860,I689849,);
nor I_40425 (I690287,I690222,I689979);
DFFARX1 I_40426 (I690287,I3035,I689860,I689828,);
nor I_40427 (I690318,I115194,I115218);
DFFARX1 I_40428 (I690318,I3035,I689860,I690344,);
DFFARX1 I_40429 (I690344,I3035,I689860,I689843,);
not I_40430 (I690366,I690344);
nand I_40431 (I689840,I690366,I689894);
nand I_40432 (I689834,I690366,I689996);
not I_40433 (I690438,I3042);
DFFARX1 I_40434 (I311139,I3035,I690438,I690464,);
nand I_40435 (I690472,I690464,I311154);
not I_40436 (I690489,I690472);
DFFARX1 I_40437 (I311136,I3035,I690438,I690515,);
not I_40438 (I690523,I690515);
not I_40439 (I690540,I311145);
or I_40440 (I690557,I311139,I311145);
nor I_40441 (I690574,I311139,I311145);
or I_40442 (I690591,I311136,I311139);
DFFARX1 I_40443 (I690591,I3035,I690438,I690430,);
not I_40444 (I690622,I311157);
nand I_40445 (I690639,I690622,I311160);
nand I_40446 (I690656,I690540,I690639);
and I_40447 (I690409,I690523,I690656);
nor I_40448 (I690687,I311157,I311142);
and I_40449 (I690704,I690523,I690687);
nor I_40450 (I690415,I690489,I690704);
DFFARX1 I_40451 (I690687,I3035,I690438,I690744,);
not I_40452 (I690752,I690744);
nor I_40453 (I690424,I690523,I690752);
or I_40454 (I690783,I690591,I311148);
nor I_40455 (I690800,I311148,I311136);
nand I_40456 (I690817,I690656,I690800);
nand I_40457 (I690834,I690783,I690817);
DFFARX1 I_40458 (I690834,I3035,I690438,I690427,);
nor I_40459 (I690865,I690800,I690557);
DFFARX1 I_40460 (I690865,I3035,I690438,I690406,);
nor I_40461 (I690896,I311148,I311151);
DFFARX1 I_40462 (I690896,I3035,I690438,I690922,);
DFFARX1 I_40463 (I690922,I3035,I690438,I690421,);
not I_40464 (I690944,I690922);
nand I_40465 (I690418,I690944,I690472);
nand I_40466 (I690412,I690944,I690574);
not I_40467 (I691016,I3042);
DFFARX1 I_40468 (I114599,I3035,I691016,I691042,);
nand I_40469 (I691050,I691042,I114602);
not I_40470 (I691067,I691050);
DFFARX1 I_40471 (I114611,I3035,I691016,I691093,);
not I_40472 (I691101,I691093);
not I_40473 (I691118,I114614);
or I_40474 (I691135,I114605,I114614);
nor I_40475 (I691152,I114605,I114614);
or I_40476 (I691169,I114617,I114605);
DFFARX1 I_40477 (I691169,I3035,I691016,I691008,);
not I_40478 (I691200,I114602);
nand I_40479 (I691217,I691200,I114608);
nand I_40480 (I691234,I691118,I691217);
and I_40481 (I690987,I691101,I691234);
nor I_40482 (I691265,I114602,I114620);
and I_40483 (I691282,I691101,I691265);
nor I_40484 (I690993,I691067,I691282);
DFFARX1 I_40485 (I691265,I3035,I691016,I691322,);
not I_40486 (I691330,I691322);
nor I_40487 (I691002,I691101,I691330);
or I_40488 (I691361,I691169,I114599);
nor I_40489 (I691378,I114599,I114617);
nand I_40490 (I691395,I691234,I691378);
nand I_40491 (I691412,I691361,I691395);
DFFARX1 I_40492 (I691412,I3035,I691016,I691005,);
nor I_40493 (I691443,I691378,I691135);
DFFARX1 I_40494 (I691443,I3035,I691016,I690984,);
nor I_40495 (I691474,I114599,I114623);
DFFARX1 I_40496 (I691474,I3035,I691016,I691500,);
DFFARX1 I_40497 (I691500,I3035,I691016,I690999,);
not I_40498 (I691522,I691500);
nand I_40499 (I690996,I691522,I691050);
nand I_40500 (I690990,I691522,I691152);
not I_40501 (I691594,I3042);
DFFARX1 I_40502 (I579822,I3035,I691594,I691620,);
nand I_40503 (I691628,I691620,I579807);
not I_40504 (I691645,I691628);
DFFARX1 I_40505 (I579810,I3035,I691594,I691671,);
not I_40506 (I691679,I691671);
not I_40507 (I691696,I579825);
or I_40508 (I691713,I579828,I579825);
nor I_40509 (I691730,I579828,I579825);
or I_40510 (I691747,I579804,I579828);
DFFARX1 I_40511 (I691747,I3035,I691594,I691586,);
not I_40512 (I691778,I579816);
nand I_40513 (I691795,I691778,I579819);
nand I_40514 (I691812,I691696,I691795);
and I_40515 (I691565,I691679,I691812);
nor I_40516 (I691843,I579816,I579813);
and I_40517 (I691860,I691679,I691843);
nor I_40518 (I691571,I691645,I691860);
DFFARX1 I_40519 (I691843,I3035,I691594,I691900,);
not I_40520 (I691908,I691900);
nor I_40521 (I691580,I691679,I691908);
or I_40522 (I691939,I691747,I579804);
nor I_40523 (I691956,I579804,I579804);
nand I_40524 (I691973,I691812,I691956);
nand I_40525 (I691990,I691939,I691973);
DFFARX1 I_40526 (I691990,I3035,I691594,I691583,);
nor I_40527 (I692021,I691956,I691713);
DFFARX1 I_40528 (I692021,I3035,I691594,I691562,);
nor I_40529 (I692052,I579804,I579807);
DFFARX1 I_40530 (I692052,I3035,I691594,I692078,);
DFFARX1 I_40531 (I692078,I3035,I691594,I691577,);
not I_40532 (I692100,I692078);
nand I_40533 (I691574,I692100,I691628);
nand I_40534 (I691568,I692100,I691730);
not I_40535 (I692172,I3042);
DFFARX1 I_40536 (I509022,I3035,I692172,I692198,);
nand I_40537 (I692206,I692198,I509043);
not I_40538 (I692223,I692206);
DFFARX1 I_40539 (I509016,I3035,I692172,I692249,);
not I_40540 (I692257,I692249);
not I_40541 (I692274,I509037);
or I_40542 (I692291,I509028,I509037);
nor I_40543 (I692308,I509028,I509037);
or I_40544 (I692325,I509031,I509028);
DFFARX1 I_40545 (I692325,I3035,I692172,I692164,);
not I_40546 (I692356,I509019);
nand I_40547 (I692373,I692356,I509034);
nand I_40548 (I692390,I692274,I692373);
and I_40549 (I692143,I692257,I692390);
nor I_40550 (I692421,I509019,I509016);
and I_40551 (I692438,I692257,I692421);
nor I_40552 (I692149,I692223,I692438);
DFFARX1 I_40553 (I692421,I3035,I692172,I692478,);
not I_40554 (I692486,I692478);
nor I_40555 (I692158,I692257,I692486);
or I_40556 (I692517,I692325,I509040);
nor I_40557 (I692534,I509040,I509031);
nand I_40558 (I692551,I692390,I692534);
nand I_40559 (I692568,I692517,I692551);
DFFARX1 I_40560 (I692568,I3035,I692172,I692161,);
nor I_40561 (I692599,I692534,I692291);
DFFARX1 I_40562 (I692599,I3035,I692172,I692140,);
nor I_40563 (I692630,I509040,I509025);
DFFARX1 I_40564 (I692630,I3035,I692172,I692656,);
DFFARX1 I_40565 (I692656,I3035,I692172,I692155,);
not I_40566 (I692678,I692656);
nand I_40567 (I692152,I692678,I692206);
nand I_40568 (I692146,I692678,I692308);
not I_40569 (I692750,I3042);
DFFARX1 I_40570 (I355642,I3035,I692750,I692776,);
nand I_40571 (I692784,I692776,I355645);
not I_40572 (I692801,I692784);
DFFARX1 I_40573 (I355657,I3035,I692750,I692827,);
not I_40574 (I692835,I692827);
not I_40575 (I692852,I355642);
or I_40576 (I692869,I355651,I355642);
nor I_40577 (I692886,I355651,I355642);
or I_40578 (I692903,I355660,I355651);
DFFARX1 I_40579 (I692903,I3035,I692750,I692742,);
not I_40580 (I692934,I355663);
nand I_40581 (I692951,I692934,I355645);
nand I_40582 (I692968,I692852,I692951);
and I_40583 (I692721,I692835,I692968);
nor I_40584 (I692999,I355663,I355648);
and I_40585 (I693016,I692835,I692999);
nor I_40586 (I692727,I692801,I693016);
DFFARX1 I_40587 (I692999,I3035,I692750,I693056,);
not I_40588 (I693064,I693056);
nor I_40589 (I692736,I692835,I693064);
or I_40590 (I693095,I692903,I355654);
nor I_40591 (I693112,I355654,I355660);
nand I_40592 (I693129,I692968,I693112);
nand I_40593 (I693146,I693095,I693129);
DFFARX1 I_40594 (I693146,I3035,I692750,I692739,);
nor I_40595 (I693177,I693112,I692869);
DFFARX1 I_40596 (I693177,I3035,I692750,I692718,);
nor I_40597 (I693208,I355654,I355666);
DFFARX1 I_40598 (I693208,I3035,I692750,I693234,);
DFFARX1 I_40599 (I693234,I3035,I692750,I692733,);
not I_40600 (I693256,I693234);
nand I_40601 (I692730,I693256,I692784);
nand I_40602 (I692724,I693256,I692886);
not I_40603 (I693331,I3042);
DFFARX1 I_40604 (I602927,I3035,I693331,I693357,);
nand I_40605 (I693365,I693357,I602924);
not I_40606 (I693382,I693365);
DFFARX1 I_40607 (I602927,I3035,I693331,I693408,);
not I_40608 (I693416,I693408);
nor I_40609 (I693433,I602945,I602939);
not I_40610 (I693450,I693433);
DFFARX1 I_40611 (I693450,I3035,I693331,I693317,);
or I_40612 (I693481,I602948,I602945);
DFFARX1 I_40613 (I693481,I3035,I693331,I693320,);
not I_40614 (I693512,I602936);
nor I_40615 (I693529,I693512,I602933);
nor I_40616 (I693546,I693529,I602939);
nor I_40617 (I693563,I602933,I602924);
nor I_40618 (I693580,I693416,I693563);
nor I_40619 (I693305,I693382,I693580);
not I_40620 (I693611,I693563);
nand I_40621 (I693308,I693611,I693365);
nand I_40622 (I693302,I693611,I693433);
nor I_40623 (I693299,I693563,I693546);
nor I_40624 (I693670,I602930,I602948);
not I_40625 (I693687,I693670);
DFFARX1 I_40626 (I693670,I3035,I693331,I693713,);
not I_40627 (I693323,I693713);
nor I_40628 (I693735,I602930,I602942);
DFFARX1 I_40629 (I693735,I3035,I693331,I693761,);
and I_40630 (I693769,I693761,I602945);
nor I_40631 (I693786,I693769,I693687);
DFFARX1 I_40632 (I693786,I3035,I693331,I693314,);
nor I_40633 (I693817,I693761,I693546);
DFFARX1 I_40634 (I693817,I3035,I693331,I693296,);
nor I_40635 (I693311,I693761,I693450);
not I_40636 (I693892,I3042);
DFFARX1 I_40637 (I251674,I3035,I693892,I693918,);
nand I_40638 (I693926,I693918,I251656);
not I_40639 (I693943,I693926);
DFFARX1 I_40640 (I251653,I3035,I693892,I693969,);
not I_40641 (I693977,I693969);
nor I_40642 (I693994,I251659,I251653);
not I_40643 (I694011,I693994);
DFFARX1 I_40644 (I694011,I3035,I693892,I693878,);
or I_40645 (I694042,I251662,I251659);
DFFARX1 I_40646 (I694042,I3035,I693892,I693881,);
not I_40647 (I694073,I251668);
nor I_40648 (I694090,I694073,I251680);
nor I_40649 (I694107,I694090,I251653);
nor I_40650 (I694124,I251680,I251665);
nor I_40651 (I694141,I693977,I694124);
nor I_40652 (I693866,I693943,I694141);
not I_40653 (I694172,I694124);
nand I_40654 (I693869,I694172,I693926);
nand I_40655 (I693863,I694172,I693994);
nor I_40656 (I693860,I694124,I694107);
nor I_40657 (I694231,I251671,I251662);
not I_40658 (I694248,I694231);
DFFARX1 I_40659 (I694231,I3035,I693892,I694274,);
not I_40660 (I693884,I694274);
nor I_40661 (I694296,I251671,I251677);
DFFARX1 I_40662 (I694296,I3035,I693892,I694322,);
and I_40663 (I694330,I694322,I251659);
nor I_40664 (I694347,I694330,I694248);
DFFARX1 I_40665 (I694347,I3035,I693892,I693875,);
nor I_40666 (I694378,I694322,I694107);
DFFARX1 I_40667 (I694378,I3035,I693892,I693857,);
nor I_40668 (I693872,I694322,I694011);
not I_40669 (I694453,I3042);
DFFARX1 I_40670 (I574027,I3035,I694453,I694479,);
nand I_40671 (I694487,I694479,I574024);
not I_40672 (I694504,I694487);
DFFARX1 I_40673 (I574027,I3035,I694453,I694530,);
not I_40674 (I694538,I694530);
nor I_40675 (I694555,I574045,I574039);
not I_40676 (I694572,I694555);
DFFARX1 I_40677 (I694572,I3035,I694453,I694439,);
or I_40678 (I694603,I574048,I574045);
DFFARX1 I_40679 (I694603,I3035,I694453,I694442,);
not I_40680 (I694634,I574036);
nor I_40681 (I694651,I694634,I574033);
nor I_40682 (I694668,I694651,I574039);
nor I_40683 (I694685,I574033,I574024);
nor I_40684 (I694702,I694538,I694685);
nor I_40685 (I694427,I694504,I694702);
not I_40686 (I694733,I694685);
nand I_40687 (I694430,I694733,I694487);
nand I_40688 (I694424,I694733,I694555);
nor I_40689 (I694421,I694685,I694668);
nor I_40690 (I694792,I574030,I574048);
not I_40691 (I694809,I694792);
DFFARX1 I_40692 (I694792,I3035,I694453,I694835,);
not I_40693 (I694445,I694835);
nor I_40694 (I694857,I574030,I574042);
DFFARX1 I_40695 (I694857,I3035,I694453,I694883,);
and I_40696 (I694891,I694883,I574045);
nor I_40697 (I694908,I694891,I694809);
DFFARX1 I_40698 (I694908,I3035,I694453,I694436,);
nor I_40699 (I694939,I694883,I694668);
DFFARX1 I_40700 (I694939,I3035,I694453,I694418,);
nor I_40701 (I694433,I694883,I694572);
not I_40702 (I695014,I3042);
DFFARX1 I_40703 (I6621,I3035,I695014,I695040,);
nand I_40704 (I695048,I695040,I6618);
not I_40705 (I695065,I695048);
DFFARX1 I_40706 (I6618,I3035,I695014,I695091,);
not I_40707 (I695099,I695091);
nor I_40708 (I695116,I6636,I6630);
not I_40709 (I695133,I695116);
DFFARX1 I_40710 (I695133,I3035,I695014,I695000,);
or I_40711 (I695164,I6633,I6636);
DFFARX1 I_40712 (I695164,I3035,I695014,I695003,);
not I_40713 (I695195,I6621);
nor I_40714 (I695212,I695195,I6615);
nor I_40715 (I695229,I695212,I6630);
nor I_40716 (I695246,I6615,I6627);
nor I_40717 (I695263,I695099,I695246);
nor I_40718 (I694988,I695065,I695263);
not I_40719 (I695294,I695246);
nand I_40720 (I694991,I695294,I695048);
nand I_40721 (I694985,I695294,I695116);
nor I_40722 (I694982,I695246,I695229);
nor I_40723 (I695353,I6624,I6633);
not I_40724 (I695370,I695353);
DFFARX1 I_40725 (I695353,I3035,I695014,I695396,);
not I_40726 (I695006,I695396);
nor I_40727 (I695418,I6624,I6615);
DFFARX1 I_40728 (I695418,I3035,I695014,I695444,);
and I_40729 (I695452,I695444,I6636);
nor I_40730 (I695469,I695452,I695370);
DFFARX1 I_40731 (I695469,I3035,I695014,I694997,);
nor I_40732 (I695500,I695444,I695229);
DFFARX1 I_40733 (I695500,I3035,I695014,I694979,);
nor I_40734 (I694994,I695444,I695133);
not I_40735 (I695575,I3042);
DFFARX1 I_40736 (I565009,I3035,I695575,I695601,);
nand I_40737 (I695609,I695601,I565012);
not I_40738 (I695626,I695609);
DFFARX1 I_40739 (I565000,I3035,I695575,I695652,);
not I_40740 (I695660,I695652);
nor I_40741 (I695677,I565018,I565015);
not I_40742 (I695694,I695677);
DFFARX1 I_40743 (I695694,I3035,I695575,I695561,);
or I_40744 (I695725,I564997,I565018);
DFFARX1 I_40745 (I695725,I3035,I695575,I695564,);
not I_40746 (I695756,I564997);
nor I_40747 (I695773,I695756,I565000);
nor I_40748 (I695790,I695773,I565015);
nor I_40749 (I695807,I565000,I565003);
nor I_40750 (I695824,I695660,I695807);
nor I_40751 (I695549,I695626,I695824);
not I_40752 (I695855,I695807);
nand I_40753 (I695552,I695855,I695609);
nand I_40754 (I695546,I695855,I695677);
nor I_40755 (I695543,I695807,I695790);
nor I_40756 (I695914,I565006,I564997);
not I_40757 (I695931,I695914);
DFFARX1 I_40758 (I695914,I3035,I695575,I695957,);
not I_40759 (I695567,I695957);
nor I_40760 (I695979,I565006,I565003);
DFFARX1 I_40761 (I695979,I3035,I695575,I696005,);
and I_40762 (I696013,I696005,I565018);
nor I_40763 (I696030,I696013,I695931);
DFFARX1 I_40764 (I696030,I3035,I695575,I695558,);
nor I_40765 (I696061,I696005,I695790);
DFFARX1 I_40766 (I696061,I3035,I695575,I695540,);
nor I_40767 (I695555,I696005,I695694);
not I_40768 (I696136,I3042);
DFFARX1 I_40769 (I594835,I3035,I696136,I696162,);
nand I_40770 (I696170,I696162,I594832);
not I_40771 (I696187,I696170);
DFFARX1 I_40772 (I594835,I3035,I696136,I696213,);
not I_40773 (I696221,I696213);
nor I_40774 (I696238,I594853,I594847);
not I_40775 (I696255,I696238);
DFFARX1 I_40776 (I696255,I3035,I696136,I696122,);
or I_40777 (I696286,I594856,I594853);
DFFARX1 I_40778 (I696286,I3035,I696136,I696125,);
not I_40779 (I696317,I594844);
nor I_40780 (I696334,I696317,I594841);
nor I_40781 (I696351,I696334,I594847);
nor I_40782 (I696368,I594841,I594832);
nor I_40783 (I696385,I696221,I696368);
nor I_40784 (I696110,I696187,I696385);
not I_40785 (I696416,I696368);
nand I_40786 (I696113,I696416,I696170);
nand I_40787 (I696107,I696416,I696238);
nor I_40788 (I696104,I696368,I696351);
nor I_40789 (I696475,I594838,I594856);
not I_40790 (I696492,I696475);
DFFARX1 I_40791 (I696475,I3035,I696136,I696518,);
not I_40792 (I696128,I696518);
nor I_40793 (I696540,I594838,I594850);
DFFARX1 I_40794 (I696540,I3035,I696136,I696566,);
and I_40795 (I696574,I696566,I594853);
nor I_40796 (I696591,I696574,I696492);
DFFARX1 I_40797 (I696591,I3035,I696136,I696119,);
nor I_40798 (I696622,I696566,I696351);
DFFARX1 I_40799 (I696622,I3035,I696136,I696101,);
nor I_40800 (I696116,I696566,I696255);
not I_40801 (I696697,I3042);
DFFARX1 I_40802 (I397276,I3035,I696697,I696723,);
nand I_40803 (I696731,I696723,I397261);
not I_40804 (I696748,I696731);
DFFARX1 I_40805 (I397279,I3035,I696697,I696774,);
not I_40806 (I696782,I696774);
nor I_40807 (I696799,I397258,I397273);
not I_40808 (I696816,I696799);
DFFARX1 I_40809 (I696816,I3035,I696697,I696683,);
or I_40810 (I696847,I397270,I397258);
DFFARX1 I_40811 (I696847,I3035,I696697,I696686,);
not I_40812 (I696878,I397258);
nor I_40813 (I696895,I696878,I397267);
nor I_40814 (I696912,I696895,I397273);
nor I_40815 (I696929,I397267,I397261);
nor I_40816 (I696946,I696782,I696929);
nor I_40817 (I696671,I696748,I696946);
not I_40818 (I696977,I696929);
nand I_40819 (I696674,I696977,I696731);
nand I_40820 (I696668,I696977,I696799);
nor I_40821 (I696665,I696929,I696912);
nor I_40822 (I697036,I397264,I397270);
not I_40823 (I697053,I697036);
DFFARX1 I_40824 (I697036,I3035,I696697,I697079,);
not I_40825 (I696689,I697079);
nor I_40826 (I697101,I397264,I397282);
DFFARX1 I_40827 (I697101,I3035,I696697,I697127,);
and I_40828 (I697135,I697127,I397258);
nor I_40829 (I697152,I697135,I697053);
DFFARX1 I_40830 (I697152,I3035,I696697,I696680,);
nor I_40831 (I697183,I697127,I696912);
DFFARX1 I_40832 (I697183,I3035,I696697,I696662,);
nor I_40833 (I696677,I697127,I696816);
not I_40834 (I697258,I3042);
DFFARX1 I_40835 (I149704,I3035,I697258,I697284,);
DFFARX1 I_40836 (I149707,I3035,I697258,I697301,);
not I_40837 (I697309,I697301);
nor I_40838 (I697226,I697284,I697309);
DFFARX1 I_40839 (I697309,I3035,I697258,I697241,);
nor I_40840 (I697354,I149713,I149707);
and I_40841 (I697371,I697354,I149710);
nor I_40842 (I697388,I697371,I149713);
not I_40843 (I697405,I149713);
and I_40844 (I697422,I697405,I149704);
nand I_40845 (I697439,I697422,I149722);
nor I_40846 (I697456,I697405,I697439);
DFFARX1 I_40847 (I697456,I3035,I697258,I697223,);
not I_40848 (I697487,I697439);
nand I_40849 (I697504,I697309,I697487);
nand I_40850 (I697235,I697371,I697487);
DFFARX1 I_40851 (I697405,I3035,I697258,I697250,);
not I_40852 (I697549,I149716);
nor I_40853 (I697566,I697549,I149704);
nor I_40854 (I697583,I697566,I697388);
DFFARX1 I_40855 (I697583,I3035,I697258,I697247,);
not I_40856 (I697614,I697566);
DFFARX1 I_40857 (I697614,I3035,I697258,I697640,);
not I_40858 (I697648,I697640);
nor I_40859 (I697244,I697648,I697566);
nor I_40860 (I697679,I697549,I149719);
and I_40861 (I697696,I697679,I149725);
or I_40862 (I697713,I697696,I149728);
DFFARX1 I_40863 (I697713,I3035,I697258,I697739,);
not I_40864 (I697747,I697739);
nand I_40865 (I697764,I697747,I697487);
not I_40866 (I697238,I697764);
nand I_40867 (I697232,I697764,I697504);
nand I_40868 (I697229,I697747,I697371);
not I_40869 (I697853,I3042);
DFFARX1 I_40870 (I305377,I3035,I697853,I697879,);
DFFARX1 I_40871 (I305371,I3035,I697853,I697896,);
not I_40872 (I697904,I697896);
nor I_40873 (I697821,I697879,I697904);
DFFARX1 I_40874 (I697904,I3035,I697853,I697836,);
nor I_40875 (I697949,I305368,I305359);
and I_40876 (I697966,I697949,I305356);
nor I_40877 (I697983,I697966,I305368);
not I_40878 (I698000,I305368);
and I_40879 (I698017,I698000,I305362);
nand I_40880 (I698034,I698017,I305374);
nor I_40881 (I698051,I698000,I698034);
DFFARX1 I_40882 (I698051,I3035,I697853,I697818,);
not I_40883 (I698082,I698034);
nand I_40884 (I698099,I697904,I698082);
nand I_40885 (I697830,I697966,I698082);
DFFARX1 I_40886 (I698000,I3035,I697853,I697845,);
not I_40887 (I698144,I305380);
nor I_40888 (I698161,I698144,I305362);
nor I_40889 (I698178,I698161,I697983);
DFFARX1 I_40890 (I698178,I3035,I697853,I697842,);
not I_40891 (I698209,I698161);
DFFARX1 I_40892 (I698209,I3035,I697853,I698235,);
not I_40893 (I698243,I698235);
nor I_40894 (I697839,I698243,I698161);
nor I_40895 (I698274,I698144,I305359);
and I_40896 (I698291,I698274,I305365);
or I_40897 (I698308,I698291,I305356);
DFFARX1 I_40898 (I698308,I3035,I697853,I698334,);
not I_40899 (I698342,I698334);
nand I_40900 (I698359,I698342,I698082);
not I_40901 (I697833,I698359);
nand I_40902 (I697827,I698359,I698099);
nand I_40903 (I697824,I698342,I697966);
not I_40904 (I698448,I3042);
DFFARX1 I_40905 (I467766,I3035,I698448,I698474,);
DFFARX1 I_40906 (I467763,I3035,I698448,I698491,);
not I_40907 (I698499,I698491);
nor I_40908 (I698416,I698474,I698499);
DFFARX1 I_40909 (I698499,I3035,I698448,I698431,);
nor I_40910 (I698544,I467778,I467760);
and I_40911 (I698561,I698544,I467757);
nor I_40912 (I698578,I698561,I467778);
not I_40913 (I698595,I467778);
and I_40914 (I698612,I698595,I467763);
nand I_40915 (I698629,I698612,I467775);
nor I_40916 (I698646,I698595,I698629);
DFFARX1 I_40917 (I698646,I3035,I698448,I698413,);
not I_40918 (I698677,I698629);
nand I_40919 (I698694,I698499,I698677);
nand I_40920 (I698425,I698561,I698677);
DFFARX1 I_40921 (I698595,I3035,I698448,I698440,);
not I_40922 (I698739,I467769);
nor I_40923 (I698756,I698739,I467763);
nor I_40924 (I698773,I698756,I698578);
DFFARX1 I_40925 (I698773,I3035,I698448,I698437,);
not I_40926 (I698804,I698756);
DFFARX1 I_40927 (I698804,I3035,I698448,I698830,);
not I_40928 (I698838,I698830);
nor I_40929 (I698434,I698838,I698756);
nor I_40930 (I698869,I698739,I467757);
and I_40931 (I698886,I698869,I467772);
or I_40932 (I698903,I698886,I467760);
DFFARX1 I_40933 (I698903,I3035,I698448,I698929,);
not I_40934 (I698937,I698929);
nand I_40935 (I698954,I698937,I698677);
not I_40936 (I698428,I698954);
nand I_40937 (I698422,I698954,I698694);
nand I_40938 (I698419,I698937,I698561);
not I_40939 (I699043,I3042);
DFFARX1 I_40940 (I689268,I3035,I699043,I699069,);
DFFARX1 I_40941 (I689259,I3035,I699043,I699086,);
not I_40942 (I699094,I699086);
nor I_40943 (I699011,I699069,I699094);
DFFARX1 I_40944 (I699094,I3035,I699043,I699026,);
nor I_40945 (I699139,I689250,I689265);
and I_40946 (I699156,I699139,I689253);
nor I_40947 (I699173,I699156,I689250);
not I_40948 (I699190,I689250);
and I_40949 (I699207,I699190,I689256);
nand I_40950 (I699224,I699207,I689274);
nor I_40951 (I699241,I699190,I699224);
DFFARX1 I_40952 (I699241,I3035,I699043,I699008,);
not I_40953 (I699272,I699224);
nand I_40954 (I699289,I699094,I699272);
nand I_40955 (I699020,I699156,I699272);
DFFARX1 I_40956 (I699190,I3035,I699043,I699035,);
not I_40957 (I699334,I689250);
nor I_40958 (I699351,I699334,I689256);
nor I_40959 (I699368,I699351,I699173);
DFFARX1 I_40960 (I699368,I3035,I699043,I699032,);
not I_40961 (I699399,I699351);
DFFARX1 I_40962 (I699399,I3035,I699043,I699425,);
not I_40963 (I699433,I699425);
nor I_40964 (I699029,I699433,I699351);
nor I_40965 (I699464,I699334,I689253);
and I_40966 (I699481,I699464,I689262);
or I_40967 (I699498,I699481,I689271);
DFFARX1 I_40968 (I699498,I3035,I699043,I699524,);
not I_40969 (I699532,I699524);
nand I_40970 (I699549,I699532,I699272);
not I_40971 (I699023,I699549);
nand I_40972 (I699017,I699549,I699289);
nand I_40973 (I699014,I699532,I699156);
not I_40974 (I699638,I3042);
DFFARX1 I_40975 (I201439,I3035,I699638,I699664,);
DFFARX1 I_40976 (I201433,I3035,I699638,I699681,);
not I_40977 (I699689,I699681);
nor I_40978 (I699606,I699664,I699689);
DFFARX1 I_40979 (I699689,I3035,I699638,I699621,);
nor I_40980 (I699734,I201421,I201442);
and I_40981 (I699751,I699734,I201436);
nor I_40982 (I699768,I699751,I201421);
not I_40983 (I699785,I201421);
and I_40984 (I699802,I699785,I201418);
nand I_40985 (I699819,I699802,I201430);
nor I_40986 (I699836,I699785,I699819);
DFFARX1 I_40987 (I699836,I3035,I699638,I699603,);
not I_40988 (I699867,I699819);
nand I_40989 (I699884,I699689,I699867);
nand I_40990 (I699615,I699751,I699867);
DFFARX1 I_40991 (I699785,I3035,I699638,I699630,);
not I_40992 (I699929,I201445);
nor I_40993 (I699946,I699929,I201418);
nor I_40994 (I699963,I699946,I699768);
DFFARX1 I_40995 (I699963,I3035,I699638,I699627,);
not I_40996 (I699994,I699946);
DFFARX1 I_40997 (I699994,I3035,I699638,I700020,);
not I_40998 (I700028,I700020);
nor I_40999 (I699624,I700028,I699946);
nor I_41000 (I700059,I699929,I201427);
and I_41001 (I700076,I700059,I201424);
or I_41002 (I700093,I700076,I201418);
DFFARX1 I_41003 (I700093,I3035,I699638,I700119,);
not I_41004 (I700127,I700119);
nand I_41005 (I700144,I700127,I699867);
not I_41006 (I699618,I700144);
nand I_41007 (I699612,I700144,I699884);
nand I_41008 (I699609,I700127,I699751);
not I_41009 (I700233,I3042);
DFFARX1 I_41010 (I15728,I3035,I700233,I700259,);
DFFARX1 I_41011 (I15710,I3035,I700233,I700276,);
not I_41012 (I700284,I700276);
nor I_41013 (I700201,I700259,I700284);
DFFARX1 I_41014 (I700284,I3035,I700233,I700216,);
nor I_41015 (I700329,I15710,I15725);
and I_41016 (I700346,I700329,I15719);
nor I_41017 (I700363,I700346,I15710);
not I_41018 (I700380,I15710);
and I_41019 (I700397,I700380,I15713);
nand I_41020 (I700414,I700397,I15716);
nor I_41021 (I700431,I700380,I700414);
DFFARX1 I_41022 (I700431,I3035,I700233,I700198,);
not I_41023 (I700462,I700414);
nand I_41024 (I700479,I700284,I700462);
nand I_41025 (I700210,I700346,I700462);
DFFARX1 I_41026 (I700380,I3035,I700233,I700225,);
not I_41027 (I700524,I15722);
nor I_41028 (I700541,I700524,I15713);
nor I_41029 (I700558,I700541,I700363);
DFFARX1 I_41030 (I700558,I3035,I700233,I700222,);
not I_41031 (I700589,I700541);
DFFARX1 I_41032 (I700589,I3035,I700233,I700615,);
not I_41033 (I700623,I700615);
nor I_41034 (I700219,I700623,I700541);
nor I_41035 (I700654,I700524,I15734);
and I_41036 (I700671,I700654,I15731);
or I_41037 (I700688,I700671,I15713);
DFFARX1 I_41038 (I700688,I3035,I700233,I700714,);
not I_41039 (I700722,I700714);
nand I_41040 (I700739,I700722,I700462);
not I_41041 (I700213,I700739);
nand I_41042 (I700207,I700739,I700479);
nand I_41043 (I700204,I700722,I700346);
not I_41044 (I700828,I3042);
DFFARX1 I_41045 (I266885,I3035,I700828,I700854,);
DFFARX1 I_41046 (I266891,I3035,I700828,I700871,);
not I_41047 (I700879,I700871);
nor I_41048 (I700796,I700854,I700879);
DFFARX1 I_41049 (I700879,I3035,I700828,I700811,);
nor I_41050 (I700924,I266900,I266885);
and I_41051 (I700941,I700924,I266912);
nor I_41052 (I700958,I700941,I266900);
not I_41053 (I700975,I266900);
and I_41054 (I700992,I700975,I266888);
nand I_41055 (I701009,I700992,I266909);
nor I_41056 (I701026,I700975,I701009);
DFFARX1 I_41057 (I701026,I3035,I700828,I700793,);
not I_41058 (I701057,I701009);
nand I_41059 (I701074,I700879,I701057);
nand I_41060 (I700805,I700941,I701057);
DFFARX1 I_41061 (I700975,I3035,I700828,I700820,);
not I_41062 (I701119,I266897);
nor I_41063 (I701136,I701119,I266888);
nor I_41064 (I701153,I701136,I700958);
DFFARX1 I_41065 (I701153,I3035,I700828,I700817,);
not I_41066 (I701184,I701136);
DFFARX1 I_41067 (I701184,I3035,I700828,I701210,);
not I_41068 (I701218,I701210);
nor I_41069 (I700814,I701218,I701136);
nor I_41070 (I701249,I701119,I266894);
and I_41071 (I701266,I701249,I266906);
or I_41072 (I701283,I701266,I266903);
DFFARX1 I_41073 (I701283,I3035,I700828,I701309,);
not I_41074 (I701317,I701309);
nand I_41075 (I701334,I701317,I701057);
not I_41076 (I700808,I701334);
nand I_41077 (I700802,I701334,I701074);
nand I_41078 (I700799,I701317,I700941);
not I_41079 (I701423,I3042);
DFFARX1 I_41080 (I191953,I3035,I701423,I701449,);
DFFARX1 I_41081 (I191947,I3035,I701423,I701466,);
not I_41082 (I701474,I701466);
nor I_41083 (I701391,I701449,I701474);
DFFARX1 I_41084 (I701474,I3035,I701423,I701406,);
nor I_41085 (I701519,I191935,I191956);
and I_41086 (I701536,I701519,I191950);
nor I_41087 (I701553,I701536,I191935);
not I_41088 (I701570,I191935);
and I_41089 (I701587,I701570,I191932);
nand I_41090 (I701604,I701587,I191944);
nor I_41091 (I701621,I701570,I701604);
DFFARX1 I_41092 (I701621,I3035,I701423,I701388,);
not I_41093 (I701652,I701604);
nand I_41094 (I701669,I701474,I701652);
nand I_41095 (I701400,I701536,I701652);
DFFARX1 I_41096 (I701570,I3035,I701423,I701415,);
not I_41097 (I701714,I191959);
nor I_41098 (I701731,I701714,I191932);
nor I_41099 (I701748,I701731,I701553);
DFFARX1 I_41100 (I701748,I3035,I701423,I701412,);
not I_41101 (I701779,I701731);
DFFARX1 I_41102 (I701779,I3035,I701423,I701805,);
not I_41103 (I701813,I701805);
nor I_41104 (I701409,I701813,I701731);
nor I_41105 (I701844,I701714,I191941);
and I_41106 (I701861,I701844,I191938);
or I_41107 (I701878,I701861,I191932);
DFFARX1 I_41108 (I701878,I3035,I701423,I701904,);
not I_41109 (I701912,I701904);
nand I_41110 (I701929,I701912,I701652);
not I_41111 (I701403,I701929);
nand I_41112 (I701397,I701929,I701669);
nand I_41113 (I701394,I701912,I701536);
not I_41114 (I702018,I3042);
DFFARX1 I_41115 (I215141,I3035,I702018,I702044,);
DFFARX1 I_41116 (I215135,I3035,I702018,I702061,);
not I_41117 (I702069,I702061);
nor I_41118 (I701986,I702044,I702069);
DFFARX1 I_41119 (I702069,I3035,I702018,I702001,);
nor I_41120 (I702114,I215123,I215144);
and I_41121 (I702131,I702114,I215138);
nor I_41122 (I702148,I702131,I215123);
not I_41123 (I702165,I215123);
and I_41124 (I702182,I702165,I215120);
nand I_41125 (I702199,I702182,I215132);
nor I_41126 (I702216,I702165,I702199);
DFFARX1 I_41127 (I702216,I3035,I702018,I701983,);
not I_41128 (I702247,I702199);
nand I_41129 (I702264,I702069,I702247);
nand I_41130 (I701995,I702131,I702247);
DFFARX1 I_41131 (I702165,I3035,I702018,I702010,);
not I_41132 (I702309,I215147);
nor I_41133 (I702326,I702309,I215120);
nor I_41134 (I702343,I702326,I702148);
DFFARX1 I_41135 (I702343,I3035,I702018,I702007,);
not I_41136 (I702374,I702326);
DFFARX1 I_41137 (I702374,I3035,I702018,I702400,);
not I_41138 (I702408,I702400);
nor I_41139 (I702004,I702408,I702326);
nor I_41140 (I702439,I702309,I215129);
and I_41141 (I702456,I702439,I215126);
or I_41142 (I702473,I702456,I215120);
DFFARX1 I_41143 (I702473,I3035,I702018,I702499,);
not I_41144 (I702507,I702499);
nand I_41145 (I702524,I702507,I702247);
not I_41146 (I701998,I702524);
nand I_41147 (I701992,I702524,I702264);
nand I_41148 (I701989,I702507,I702131);
not I_41149 (I702613,I3042);
DFFARX1 I_41150 (I603505,I3035,I702613,I702639,);
DFFARX1 I_41151 (I603517,I3035,I702613,I702656,);
not I_41152 (I702664,I702656);
nor I_41153 (I702581,I702639,I702664);
DFFARX1 I_41154 (I702664,I3035,I702613,I702596,);
nor I_41155 (I702709,I603514,I603508);
and I_41156 (I702726,I702709,I603502);
nor I_41157 (I702743,I702726,I603514);
not I_41158 (I702760,I603514);
and I_41159 (I702777,I702760,I603511);
nand I_41160 (I702794,I702777,I603502);
nor I_41161 (I702811,I702760,I702794);
DFFARX1 I_41162 (I702811,I3035,I702613,I702578,);
not I_41163 (I702842,I702794);
nand I_41164 (I702859,I702664,I702842);
nand I_41165 (I702590,I702726,I702842);
DFFARX1 I_41166 (I702760,I3035,I702613,I702605,);
not I_41167 (I702904,I603526);
nor I_41168 (I702921,I702904,I603511);
nor I_41169 (I702938,I702921,I702743);
DFFARX1 I_41170 (I702938,I3035,I702613,I702602,);
not I_41171 (I702969,I702921);
DFFARX1 I_41172 (I702969,I3035,I702613,I702995,);
not I_41173 (I703003,I702995);
nor I_41174 (I702599,I703003,I702921);
nor I_41175 (I703034,I702904,I603520);
and I_41176 (I703051,I703034,I603523);
or I_41177 (I703068,I703051,I603505);
DFFARX1 I_41178 (I703068,I3035,I702613,I703094,);
not I_41179 (I703102,I703094);
nand I_41180 (I703119,I703102,I702842);
not I_41181 (I702593,I703119);
nand I_41182 (I702587,I703119,I702859);
nand I_41183 (I702584,I703102,I702726);
not I_41184 (I703208,I3042);
DFFARX1 I_41185 (I588477,I3035,I703208,I703234,);
DFFARX1 I_41186 (I588489,I3035,I703208,I703251,);
not I_41187 (I703259,I703251);
nor I_41188 (I703176,I703234,I703259);
DFFARX1 I_41189 (I703259,I3035,I703208,I703191,);
nor I_41190 (I703304,I588486,I588480);
and I_41191 (I703321,I703304,I588474);
nor I_41192 (I703338,I703321,I588486);
not I_41193 (I703355,I588486);
and I_41194 (I703372,I703355,I588483);
nand I_41195 (I703389,I703372,I588474);
nor I_41196 (I703406,I703355,I703389);
DFFARX1 I_41197 (I703406,I3035,I703208,I703173,);
not I_41198 (I703437,I703389);
nand I_41199 (I703454,I703259,I703437);
nand I_41200 (I703185,I703321,I703437);
DFFARX1 I_41201 (I703355,I3035,I703208,I703200,);
not I_41202 (I703499,I588498);
nor I_41203 (I703516,I703499,I588483);
nor I_41204 (I703533,I703516,I703338);
DFFARX1 I_41205 (I703533,I3035,I703208,I703197,);
not I_41206 (I703564,I703516);
DFFARX1 I_41207 (I703564,I3035,I703208,I703590,);
not I_41208 (I703598,I703590);
nor I_41209 (I703194,I703598,I703516);
nor I_41210 (I703629,I703499,I588492);
and I_41211 (I703646,I703629,I588495);
or I_41212 (I703663,I703646,I588477);
DFFARX1 I_41213 (I703663,I3035,I703208,I703689,);
not I_41214 (I703697,I703689);
nand I_41215 (I703714,I703697,I703437);
not I_41216 (I703188,I703714);
nand I_41217 (I703182,I703714,I703454);
nand I_41218 (I703179,I703697,I703321);
not I_41219 (I703803,I3042);
DFFARX1 I_41220 (I507730,I3035,I703803,I703829,);
DFFARX1 I_41221 (I507748,I3035,I703803,I703846,);
not I_41222 (I703854,I703846);
nor I_41223 (I703771,I703829,I703854);
DFFARX1 I_41224 (I703854,I3035,I703803,I703786,);
nor I_41225 (I703899,I507727,I507739);
and I_41226 (I703916,I703899,I507724);
nor I_41227 (I703933,I703916,I507727);
not I_41228 (I703950,I507727);
and I_41229 (I703967,I703950,I507733);
nand I_41230 (I703984,I703967,I507745);
nor I_41231 (I704001,I703950,I703984);
DFFARX1 I_41232 (I704001,I3035,I703803,I703768,);
not I_41233 (I704032,I703984);
nand I_41234 (I704049,I703854,I704032);
nand I_41235 (I703780,I703916,I704032);
DFFARX1 I_41236 (I703950,I3035,I703803,I703795,);
not I_41237 (I704094,I507736);
nor I_41238 (I704111,I704094,I507733);
nor I_41239 (I704128,I704111,I703933);
DFFARX1 I_41240 (I704128,I3035,I703803,I703792,);
not I_41241 (I704159,I704111);
DFFARX1 I_41242 (I704159,I3035,I703803,I704185,);
not I_41243 (I704193,I704185);
nor I_41244 (I703789,I704193,I704111);
nor I_41245 (I704224,I704094,I507724);
and I_41246 (I704241,I704224,I507751);
or I_41247 (I704258,I704241,I507742);
DFFARX1 I_41248 (I704258,I3035,I703803,I704284,);
not I_41249 (I704292,I704284);
nand I_41250 (I704309,I704292,I704032);
not I_41251 (I703783,I704309);
nand I_41252 (I703777,I704309,I704049);
nand I_41253 (I703774,I704292,I703916);
not I_41254 (I704398,I3042);
DFFARX1 I_41255 (I659398,I3035,I704398,I704424,);
DFFARX1 I_41256 (I659401,I3035,I704398,I704441,);
not I_41257 (I704449,I704441);
nor I_41258 (I704366,I704424,I704449);
DFFARX1 I_41259 (I704449,I3035,I704398,I704381,);
nor I_41260 (I704494,I659401,I659416);
and I_41261 (I704511,I704494,I659410);
nor I_41262 (I704528,I704511,I659401);
not I_41263 (I704545,I659401);
and I_41264 (I704562,I704545,I659419);
nand I_41265 (I704579,I704562,I659407);
nor I_41266 (I704596,I704545,I704579);
DFFARX1 I_41267 (I704596,I3035,I704398,I704363,);
not I_41268 (I704627,I704579);
nand I_41269 (I704644,I704449,I704627);
nand I_41270 (I704375,I704511,I704627);
DFFARX1 I_41271 (I704545,I3035,I704398,I704390,);
not I_41272 (I704689,I659413);
nor I_41273 (I704706,I704689,I659419);
nor I_41274 (I704723,I704706,I704528);
DFFARX1 I_41275 (I704723,I3035,I704398,I704387,);
not I_41276 (I704754,I704706);
DFFARX1 I_41277 (I704754,I3035,I704398,I704780,);
not I_41278 (I704788,I704780);
nor I_41279 (I704384,I704788,I704706);
nor I_41280 (I704819,I704689,I659398);
and I_41281 (I704836,I704819,I659422);
or I_41282 (I704853,I704836,I659404);
DFFARX1 I_41283 (I704853,I3035,I704398,I704879,);
not I_41284 (I704887,I704879);
nand I_41285 (I704904,I704887,I704627);
not I_41286 (I704378,I704904);
nand I_41287 (I704372,I704904,I704644);
nand I_41288 (I704369,I704887,I704511);
not I_41289 (I704993,I3042);
DFFARX1 I_41290 (I2260,I3035,I704993,I705019,);
DFFARX1 I_41291 (I2452,I3035,I704993,I705036,);
not I_41292 (I705044,I705036);
nor I_41293 (I704961,I705019,I705044);
DFFARX1 I_41294 (I705044,I3035,I704993,I704976,);
nor I_41295 (I705089,I2460,I1412);
and I_41296 (I705106,I705089,I1444);
nor I_41297 (I705123,I705106,I2460);
not I_41298 (I705140,I2460);
and I_41299 (I705157,I705140,I2492);
nand I_41300 (I705174,I705157,I2628);
nor I_41301 (I705191,I705140,I705174);
DFFARX1 I_41302 (I705191,I3035,I704993,I704958,);
not I_41303 (I705222,I705174);
nand I_41304 (I705239,I705044,I705222);
nand I_41305 (I704970,I705106,I705222);
DFFARX1 I_41306 (I705140,I3035,I704993,I704985,);
not I_41307 (I705284,I1644);
nor I_41308 (I705301,I705284,I2492);
nor I_41309 (I705318,I705301,I705123);
DFFARX1 I_41310 (I705318,I3035,I704993,I704982,);
not I_41311 (I705349,I705301);
DFFARX1 I_41312 (I705349,I3035,I704993,I705375,);
not I_41313 (I705383,I705375);
nor I_41314 (I704979,I705383,I705301);
nor I_41315 (I705414,I705284,I2340);
and I_41316 (I705431,I705414,I2916);
or I_41317 (I705448,I705431,I2620);
DFFARX1 I_41318 (I705448,I3035,I704993,I705474,);
not I_41319 (I705482,I705474);
nand I_41320 (I705499,I705482,I705222);
not I_41321 (I704973,I705499);
nand I_41322 (I704967,I705499,I705239);
nand I_41323 (I704964,I705482,I705106);
not I_41324 (I705588,I3042);
DFFARX1 I_41325 (I600037,I3035,I705588,I705614,);
DFFARX1 I_41326 (I600049,I3035,I705588,I705631,);
not I_41327 (I705639,I705631);
nor I_41328 (I705556,I705614,I705639);
DFFARX1 I_41329 (I705639,I3035,I705588,I705571,);
nor I_41330 (I705684,I600046,I600040);
and I_41331 (I705701,I705684,I600034);
nor I_41332 (I705718,I705701,I600046);
not I_41333 (I705735,I600046);
and I_41334 (I705752,I705735,I600043);
nand I_41335 (I705769,I705752,I600034);
nor I_41336 (I705786,I705735,I705769);
DFFARX1 I_41337 (I705786,I3035,I705588,I705553,);
not I_41338 (I705817,I705769);
nand I_41339 (I705834,I705639,I705817);
nand I_41340 (I705565,I705701,I705817);
DFFARX1 I_41341 (I705735,I3035,I705588,I705580,);
not I_41342 (I705879,I600058);
nor I_41343 (I705896,I705879,I600043);
nor I_41344 (I705913,I705896,I705718);
DFFARX1 I_41345 (I705913,I3035,I705588,I705577,);
not I_41346 (I705944,I705896);
DFFARX1 I_41347 (I705944,I3035,I705588,I705970,);
not I_41348 (I705978,I705970);
nor I_41349 (I705574,I705978,I705896);
nor I_41350 (I706009,I705879,I600052);
and I_41351 (I706026,I706009,I600055);
or I_41352 (I706043,I706026,I600037);
DFFARX1 I_41353 (I706043,I3035,I705588,I706069,);
not I_41354 (I706077,I706069);
nand I_41355 (I706094,I706077,I705817);
not I_41356 (I705568,I706094);
nand I_41357 (I705562,I706094,I705834);
nand I_41358 (I705559,I706077,I705701);
not I_41359 (I706183,I3042);
DFFARX1 I_41360 (I460915,I3035,I706183,I706209,);
DFFARX1 I_41361 (I460912,I3035,I706183,I706226,);
not I_41362 (I706234,I706226);
nor I_41363 (I706151,I706209,I706234);
DFFARX1 I_41364 (I706234,I3035,I706183,I706166,);
nor I_41365 (I706279,I460927,I460909);
and I_41366 (I706296,I706279,I460906);
nor I_41367 (I706313,I706296,I460927);
not I_41368 (I706330,I460927);
and I_41369 (I706347,I706330,I460912);
nand I_41370 (I706364,I706347,I460924);
nor I_41371 (I706381,I706330,I706364);
DFFARX1 I_41372 (I706381,I3035,I706183,I706148,);
not I_41373 (I706412,I706364);
nand I_41374 (I706429,I706234,I706412);
nand I_41375 (I706160,I706296,I706412);
DFFARX1 I_41376 (I706330,I3035,I706183,I706175,);
not I_41377 (I706474,I460918);
nor I_41378 (I706491,I706474,I460912);
nor I_41379 (I706508,I706491,I706313);
DFFARX1 I_41380 (I706508,I3035,I706183,I706172,);
not I_41381 (I706539,I706491);
DFFARX1 I_41382 (I706539,I3035,I706183,I706565,);
not I_41383 (I706573,I706565);
nor I_41384 (I706169,I706573,I706491);
nor I_41385 (I706604,I706474,I460906);
and I_41386 (I706621,I706604,I460921);
or I_41387 (I706638,I706621,I460909);
DFFARX1 I_41388 (I706638,I3035,I706183,I706664,);
not I_41389 (I706672,I706664);
nand I_41390 (I706689,I706672,I706412);
not I_41391 (I706163,I706689);
nand I_41392 (I706157,I706689,I706429);
nand I_41393 (I706154,I706672,I706296);
not I_41394 (I706778,I3042);
DFFARX1 I_41395 (I357397,I3035,I706778,I706804,);
DFFARX1 I_41396 (I357379,I3035,I706778,I706821,);
not I_41397 (I706829,I706821);
nor I_41398 (I706746,I706804,I706829);
DFFARX1 I_41399 (I706829,I3035,I706778,I706761,);
nor I_41400 (I706874,I357385,I357388);
and I_41401 (I706891,I706874,I357376);
nor I_41402 (I706908,I706891,I357385);
not I_41403 (I706925,I357385);
and I_41404 (I706942,I706925,I357394);
nand I_41405 (I706959,I706942,I357382);
nor I_41406 (I706976,I706925,I706959);
DFFARX1 I_41407 (I706976,I3035,I706778,I706743,);
not I_41408 (I707007,I706959);
nand I_41409 (I707024,I706829,I707007);
nand I_41410 (I706755,I706891,I707007);
DFFARX1 I_41411 (I706925,I3035,I706778,I706770,);
not I_41412 (I707069,I357379);
nor I_41413 (I707086,I707069,I357394);
nor I_41414 (I707103,I707086,I706908);
DFFARX1 I_41415 (I707103,I3035,I706778,I706767,);
not I_41416 (I707134,I707086);
DFFARX1 I_41417 (I707134,I3035,I706778,I707160,);
not I_41418 (I707168,I707160);
nor I_41419 (I706764,I707168,I707086);
nor I_41420 (I707199,I707069,I357391);
and I_41421 (I707216,I707199,I357400);
or I_41422 (I707233,I707216,I357376);
DFFARX1 I_41423 (I707233,I3035,I706778,I707259,);
not I_41424 (I707267,I707259);
nand I_41425 (I707284,I707267,I707007);
not I_41426 (I706758,I707284);
nand I_41427 (I706752,I707284,I707024);
nand I_41428 (I706749,I707267,I706891);
not I_41429 (I707373,I3042);
DFFARX1 I_41430 (I27849,I3035,I707373,I707399,);
DFFARX1 I_41431 (I27831,I3035,I707373,I707416,);
not I_41432 (I707424,I707416);
nor I_41433 (I707341,I707399,I707424);
DFFARX1 I_41434 (I707424,I3035,I707373,I707356,);
nor I_41435 (I707469,I27831,I27846);
and I_41436 (I707486,I707469,I27840);
nor I_41437 (I707503,I707486,I27831);
not I_41438 (I707520,I27831);
and I_41439 (I707537,I707520,I27834);
nand I_41440 (I707554,I707537,I27837);
nor I_41441 (I707571,I707520,I707554);
DFFARX1 I_41442 (I707571,I3035,I707373,I707338,);
not I_41443 (I707602,I707554);
nand I_41444 (I707619,I707424,I707602);
nand I_41445 (I707350,I707486,I707602);
DFFARX1 I_41446 (I707520,I3035,I707373,I707365,);
not I_41447 (I707664,I27843);
nor I_41448 (I707681,I707664,I27834);
nor I_41449 (I707698,I707681,I707503);
DFFARX1 I_41450 (I707698,I3035,I707373,I707362,);
not I_41451 (I707729,I707681);
DFFARX1 I_41452 (I707729,I3035,I707373,I707755,);
not I_41453 (I707763,I707755);
nor I_41454 (I707359,I707763,I707681);
nor I_41455 (I707794,I707664,I27855);
and I_41456 (I707811,I707794,I27852);
or I_41457 (I707828,I707811,I27834);
DFFARX1 I_41458 (I707828,I3035,I707373,I707854,);
not I_41459 (I707862,I707854);
nand I_41460 (I707879,I707862,I707602);
not I_41461 (I707353,I707879);
nand I_41462 (I707347,I707879,I707619);
nand I_41463 (I707344,I707862,I707486);
not I_41464 (I707968,I3042);
DFFARX1 I_41465 (I192480,I3035,I707968,I707994,);
DFFARX1 I_41466 (I192474,I3035,I707968,I708011,);
not I_41467 (I708019,I708011);
nor I_41468 (I707936,I707994,I708019);
DFFARX1 I_41469 (I708019,I3035,I707968,I707951,);
nor I_41470 (I708064,I192462,I192483);
and I_41471 (I708081,I708064,I192477);
nor I_41472 (I708098,I708081,I192462);
not I_41473 (I708115,I192462);
and I_41474 (I708132,I708115,I192459);
nand I_41475 (I708149,I708132,I192471);
nor I_41476 (I708166,I708115,I708149);
DFFARX1 I_41477 (I708166,I3035,I707968,I707933,);
not I_41478 (I708197,I708149);
nand I_41479 (I708214,I708019,I708197);
nand I_41480 (I707945,I708081,I708197);
DFFARX1 I_41481 (I708115,I3035,I707968,I707960,);
not I_41482 (I708259,I192486);
nor I_41483 (I708276,I708259,I192459);
nor I_41484 (I708293,I708276,I708098);
DFFARX1 I_41485 (I708293,I3035,I707968,I707957,);
not I_41486 (I708324,I708276);
DFFARX1 I_41487 (I708324,I3035,I707968,I708350,);
not I_41488 (I708358,I708350);
nor I_41489 (I707954,I708358,I708276);
nor I_41490 (I708389,I708259,I192468);
and I_41491 (I708406,I708389,I192465);
or I_41492 (I708423,I708406,I192459);
DFFARX1 I_41493 (I708423,I3035,I707968,I708449,);
not I_41494 (I708457,I708449);
nand I_41495 (I708474,I708457,I708197);
not I_41496 (I707948,I708474);
nand I_41497 (I707942,I708474,I708214);
nand I_41498 (I707939,I708457,I708081);
not I_41499 (I708563,I3042);
DFFARX1 I_41500 (I68431,I3035,I708563,I708589,);
DFFARX1 I_41501 (I68419,I3035,I708563,I708606,);
not I_41502 (I708614,I708606);
nor I_41503 (I708531,I708589,I708614);
DFFARX1 I_41504 (I708614,I3035,I708563,I708546,);
nor I_41505 (I708659,I68410,I68434);
and I_41506 (I708676,I708659,I68413);
nor I_41507 (I708693,I708676,I68410);
not I_41508 (I708710,I68410);
and I_41509 (I708727,I708710,I68416);
nand I_41510 (I708744,I708727,I68428);
nor I_41511 (I708761,I708710,I708744);
DFFARX1 I_41512 (I708761,I3035,I708563,I708528,);
not I_41513 (I708792,I708744);
nand I_41514 (I708809,I708614,I708792);
nand I_41515 (I708540,I708676,I708792);
DFFARX1 I_41516 (I708710,I3035,I708563,I708555,);
not I_41517 (I708854,I68410);
nor I_41518 (I708871,I708854,I68416);
nor I_41519 (I708888,I708871,I708693);
DFFARX1 I_41520 (I708888,I3035,I708563,I708552,);
not I_41521 (I708919,I708871);
DFFARX1 I_41522 (I708919,I3035,I708563,I708945,);
not I_41523 (I708953,I708945);
nor I_41524 (I708549,I708953,I708871);
nor I_41525 (I708984,I708854,I68413);
and I_41526 (I709001,I708984,I68422);
or I_41527 (I709018,I709001,I68425);
DFFARX1 I_41528 (I709018,I3035,I708563,I709044,);
not I_41529 (I709052,I709044);
nand I_41530 (I709069,I709052,I708792);
not I_41531 (I708543,I709069);
nand I_41532 (I708537,I709069,I708809);
nand I_41533 (I708534,I709052,I708676);
not I_41534 (I709158,I3042);
DFFARX1 I_41535 (I655590,I3035,I709158,I709184,);
DFFARX1 I_41536 (I655593,I3035,I709158,I709201,);
not I_41537 (I709209,I709201);
nor I_41538 (I709126,I709184,I709209);
DFFARX1 I_41539 (I709209,I3035,I709158,I709141,);
nor I_41540 (I709254,I655593,I655608);
and I_41541 (I709271,I709254,I655602);
nor I_41542 (I709288,I709271,I655593);
not I_41543 (I709305,I655593);
and I_41544 (I709322,I709305,I655611);
nand I_41545 (I709339,I709322,I655599);
nor I_41546 (I709356,I709305,I709339);
DFFARX1 I_41547 (I709356,I3035,I709158,I709123,);
not I_41548 (I709387,I709339);
nand I_41549 (I709404,I709209,I709387);
nand I_41550 (I709135,I709271,I709387);
DFFARX1 I_41551 (I709305,I3035,I709158,I709150,);
not I_41552 (I709449,I655605);
nor I_41553 (I709466,I709449,I655611);
nor I_41554 (I709483,I709466,I709288);
DFFARX1 I_41555 (I709483,I3035,I709158,I709147,);
not I_41556 (I709514,I709466);
DFFARX1 I_41557 (I709514,I3035,I709158,I709540,);
not I_41558 (I709548,I709540);
nor I_41559 (I709144,I709548,I709466);
nor I_41560 (I709579,I709449,I655590);
and I_41561 (I709596,I709579,I655614);
or I_41562 (I709613,I709596,I655596);
DFFARX1 I_41563 (I709613,I3035,I709158,I709639,);
not I_41564 (I709647,I709639);
nand I_41565 (I709664,I709647,I709387);
not I_41566 (I709138,I709664);
nand I_41567 (I709132,I709664,I709404);
nand I_41568 (I709129,I709647,I709271);
not I_41569 (I709753,I3042);
DFFARX1 I_41570 (I352195,I3035,I709753,I709779,);
DFFARX1 I_41571 (I352177,I3035,I709753,I709796,);
not I_41572 (I709804,I709796);
nor I_41573 (I709721,I709779,I709804);
DFFARX1 I_41574 (I709804,I3035,I709753,I709736,);
nor I_41575 (I709849,I352183,I352186);
and I_41576 (I709866,I709849,I352174);
nor I_41577 (I709883,I709866,I352183);
not I_41578 (I709900,I352183);
and I_41579 (I709917,I709900,I352192);
nand I_41580 (I709934,I709917,I352180);
nor I_41581 (I709951,I709900,I709934);
DFFARX1 I_41582 (I709951,I3035,I709753,I709718,);
not I_41583 (I709982,I709934);
nand I_41584 (I709999,I709804,I709982);
nand I_41585 (I709730,I709866,I709982);
DFFARX1 I_41586 (I709900,I3035,I709753,I709745,);
not I_41587 (I710044,I352177);
nor I_41588 (I710061,I710044,I352192);
nor I_41589 (I710078,I710061,I709883);
DFFARX1 I_41590 (I710078,I3035,I709753,I709742,);
not I_41591 (I710109,I710061);
DFFARX1 I_41592 (I710109,I3035,I709753,I710135,);
not I_41593 (I710143,I710135);
nor I_41594 (I709739,I710143,I710061);
nor I_41595 (I710174,I710044,I352189);
and I_41596 (I710191,I710174,I352198);
or I_41597 (I710208,I710191,I352174);
DFFARX1 I_41598 (I710208,I3035,I709753,I710234,);
not I_41599 (I710242,I710234);
nand I_41600 (I710259,I710242,I709982);
not I_41601 (I709733,I710259);
nand I_41602 (I709727,I710259,I709999);
nand I_41603 (I709724,I710242,I709866);
not I_41604 (I710348,I3042);
DFFARX1 I_41605 (I393233,I3035,I710348,I710374,);
DFFARX1 I_41606 (I393215,I3035,I710348,I710391,);
not I_41607 (I710399,I710391);
nor I_41608 (I710316,I710374,I710399);
DFFARX1 I_41609 (I710399,I3035,I710348,I710331,);
nor I_41610 (I710444,I393221,I393224);
and I_41611 (I710461,I710444,I393212);
nor I_41612 (I710478,I710461,I393221);
not I_41613 (I710495,I393221);
and I_41614 (I710512,I710495,I393230);
nand I_41615 (I710529,I710512,I393218);
nor I_41616 (I710546,I710495,I710529);
DFFARX1 I_41617 (I710546,I3035,I710348,I710313,);
not I_41618 (I710577,I710529);
nand I_41619 (I710594,I710399,I710577);
nand I_41620 (I710325,I710461,I710577);
DFFARX1 I_41621 (I710495,I3035,I710348,I710340,);
not I_41622 (I710639,I393215);
nor I_41623 (I710656,I710639,I393230);
nor I_41624 (I710673,I710656,I710478);
DFFARX1 I_41625 (I710673,I3035,I710348,I710337,);
not I_41626 (I710704,I710656);
DFFARX1 I_41627 (I710704,I3035,I710348,I710730,);
not I_41628 (I710738,I710730);
nor I_41629 (I710334,I710738,I710656);
nor I_41630 (I710769,I710639,I393227);
and I_41631 (I710786,I710769,I393236);
or I_41632 (I710803,I710786,I393212);
DFFARX1 I_41633 (I710803,I3035,I710348,I710829,);
not I_41634 (I710837,I710829);
nand I_41635 (I710854,I710837,I710577);
not I_41636 (I710328,I710854);
nand I_41637 (I710322,I710854,I710594);
nand I_41638 (I710319,I710837,I710461);
not I_41639 (I710943,I3042);
DFFARX1 I_41640 (I521942,I3035,I710943,I710969,);
DFFARX1 I_41641 (I521960,I3035,I710943,I710986,);
not I_41642 (I710994,I710986);
nor I_41643 (I710911,I710969,I710994);
DFFARX1 I_41644 (I710994,I3035,I710943,I710926,);
nor I_41645 (I711039,I521939,I521951);
and I_41646 (I711056,I711039,I521936);
nor I_41647 (I711073,I711056,I521939);
not I_41648 (I711090,I521939);
and I_41649 (I711107,I711090,I521945);
nand I_41650 (I711124,I711107,I521957);
nor I_41651 (I711141,I711090,I711124);
DFFARX1 I_41652 (I711141,I3035,I710943,I710908,);
not I_41653 (I711172,I711124);
nand I_41654 (I711189,I710994,I711172);
nand I_41655 (I710920,I711056,I711172);
DFFARX1 I_41656 (I711090,I3035,I710943,I710935,);
not I_41657 (I711234,I521948);
nor I_41658 (I711251,I711234,I521945);
nor I_41659 (I711268,I711251,I711073);
DFFARX1 I_41660 (I711268,I3035,I710943,I710932,);
not I_41661 (I711299,I711251);
DFFARX1 I_41662 (I711299,I3035,I710943,I711325,);
not I_41663 (I711333,I711325);
nor I_41664 (I710929,I711333,I711251);
nor I_41665 (I711364,I711234,I521936);
and I_41666 (I711381,I711364,I521963);
or I_41667 (I711398,I711381,I521954);
DFFARX1 I_41668 (I711398,I3035,I710943,I711424,);
not I_41669 (I711432,I711424);
nand I_41670 (I711449,I711432,I711172);
not I_41671 (I710923,I711449);
nand I_41672 (I710917,I711449,I711189);
nand I_41673 (I710914,I711432,I711056);
not I_41674 (I711538,I3042);
DFFARX1 I_41675 (I126499,I3035,I711538,I711564,);
DFFARX1 I_41676 (I126502,I3035,I711538,I711581,);
not I_41677 (I711589,I711581);
nor I_41678 (I711506,I711564,I711589);
DFFARX1 I_41679 (I711589,I3035,I711538,I711521,);
nor I_41680 (I711634,I126508,I126502);
and I_41681 (I711651,I711634,I126505);
nor I_41682 (I711668,I711651,I126508);
not I_41683 (I711685,I126508);
and I_41684 (I711702,I711685,I126499);
nand I_41685 (I711719,I711702,I126517);
nor I_41686 (I711736,I711685,I711719);
DFFARX1 I_41687 (I711736,I3035,I711538,I711503,);
not I_41688 (I711767,I711719);
nand I_41689 (I711784,I711589,I711767);
nand I_41690 (I711515,I711651,I711767);
DFFARX1 I_41691 (I711685,I3035,I711538,I711530,);
not I_41692 (I711829,I126511);
nor I_41693 (I711846,I711829,I126499);
nor I_41694 (I711863,I711846,I711668);
DFFARX1 I_41695 (I711863,I3035,I711538,I711527,);
not I_41696 (I711894,I711846);
DFFARX1 I_41697 (I711894,I3035,I711538,I711920,);
not I_41698 (I711928,I711920);
nor I_41699 (I711524,I711928,I711846);
nor I_41700 (I711959,I711829,I126514);
and I_41701 (I711976,I711959,I126520);
or I_41702 (I711993,I711976,I126523);
DFFARX1 I_41703 (I711993,I3035,I711538,I712019,);
not I_41704 (I712027,I712019);
nand I_41705 (I712044,I712027,I711767);
not I_41706 (I711518,I712044);
nand I_41707 (I711512,I712044,I711784);
nand I_41708 (I711509,I712027,I711651);
not I_41709 (I712133,I3042);
DFFARX1 I_41710 (I144349,I3035,I712133,I712159,);
DFFARX1 I_41711 (I144352,I3035,I712133,I712176,);
not I_41712 (I712184,I712176);
nor I_41713 (I712101,I712159,I712184);
DFFARX1 I_41714 (I712184,I3035,I712133,I712116,);
nor I_41715 (I712229,I144358,I144352);
and I_41716 (I712246,I712229,I144355);
nor I_41717 (I712263,I712246,I144358);
not I_41718 (I712280,I144358);
and I_41719 (I712297,I712280,I144349);
nand I_41720 (I712314,I712297,I144367);
nor I_41721 (I712331,I712280,I712314);
DFFARX1 I_41722 (I712331,I3035,I712133,I712098,);
not I_41723 (I712362,I712314);
nand I_41724 (I712379,I712184,I712362);
nand I_41725 (I712110,I712246,I712362);
DFFARX1 I_41726 (I712280,I3035,I712133,I712125,);
not I_41727 (I712424,I144361);
nor I_41728 (I712441,I712424,I144349);
nor I_41729 (I712458,I712441,I712263);
DFFARX1 I_41730 (I712458,I3035,I712133,I712122,);
not I_41731 (I712489,I712441);
DFFARX1 I_41732 (I712489,I3035,I712133,I712515,);
not I_41733 (I712523,I712515);
nor I_41734 (I712119,I712523,I712441);
nor I_41735 (I712554,I712424,I144364);
and I_41736 (I712571,I712554,I144370);
or I_41737 (I712588,I712571,I144373);
DFFARX1 I_41738 (I712588,I3035,I712133,I712614,);
not I_41739 (I712622,I712614);
nand I_41740 (I712639,I712622,I712362);
not I_41741 (I712113,I712639);
nand I_41742 (I712107,I712639,I712379);
nand I_41743 (I712104,I712622,I712246);
not I_41744 (I712728,I3042);
DFFARX1 I_41745 (I498686,I3035,I712728,I712754,);
DFFARX1 I_41746 (I498704,I3035,I712728,I712771,);
not I_41747 (I712779,I712771);
nor I_41748 (I712696,I712754,I712779);
DFFARX1 I_41749 (I712779,I3035,I712728,I712711,);
nor I_41750 (I712824,I498683,I498695);
and I_41751 (I712841,I712824,I498680);
nor I_41752 (I712858,I712841,I498683);
not I_41753 (I712875,I498683);
and I_41754 (I712892,I712875,I498689);
nand I_41755 (I712909,I712892,I498701);
nor I_41756 (I712926,I712875,I712909);
DFFARX1 I_41757 (I712926,I3035,I712728,I712693,);
not I_41758 (I712957,I712909);
nand I_41759 (I712974,I712779,I712957);
nand I_41760 (I712705,I712841,I712957);
DFFARX1 I_41761 (I712875,I3035,I712728,I712720,);
not I_41762 (I713019,I498692);
nor I_41763 (I713036,I713019,I498689);
nor I_41764 (I713053,I713036,I712858);
DFFARX1 I_41765 (I713053,I3035,I712728,I712717,);
not I_41766 (I713084,I713036);
DFFARX1 I_41767 (I713084,I3035,I712728,I713110,);
not I_41768 (I713118,I713110);
nor I_41769 (I712714,I713118,I713036);
nor I_41770 (I713149,I713019,I498680);
and I_41771 (I713166,I713149,I498707);
or I_41772 (I713183,I713166,I498698);
DFFARX1 I_41773 (I713183,I3035,I712728,I713209,);
not I_41774 (I713217,I713209);
nand I_41775 (I713234,I713217,I712957);
not I_41776 (I712708,I713234);
nand I_41777 (I712702,I713234,I712974);
nand I_41778 (I712699,I713217,I712841);
not I_41779 (I713323,I3042);
DFFARX1 I_41780 (I578073,I3035,I713323,I713349,);
DFFARX1 I_41781 (I578085,I3035,I713323,I713366,);
not I_41782 (I713374,I713366);
nor I_41783 (I713291,I713349,I713374);
DFFARX1 I_41784 (I713374,I3035,I713323,I713306,);
nor I_41785 (I713419,I578082,I578076);
and I_41786 (I713436,I713419,I578070);
nor I_41787 (I713453,I713436,I578082);
not I_41788 (I713470,I578082);
and I_41789 (I713487,I713470,I578079);
nand I_41790 (I713504,I713487,I578070);
nor I_41791 (I713521,I713470,I713504);
DFFARX1 I_41792 (I713521,I3035,I713323,I713288,);
not I_41793 (I713552,I713504);
nand I_41794 (I713569,I713374,I713552);
nand I_41795 (I713300,I713436,I713552);
DFFARX1 I_41796 (I713470,I3035,I713323,I713315,);
not I_41797 (I713614,I578094);
nor I_41798 (I713631,I713614,I578079);
nor I_41799 (I713648,I713631,I713453);
DFFARX1 I_41800 (I713648,I3035,I713323,I713312,);
not I_41801 (I713679,I713631);
DFFARX1 I_41802 (I713679,I3035,I713323,I713705,);
not I_41803 (I713713,I713705);
nor I_41804 (I713309,I713713,I713631);
nor I_41805 (I713744,I713614,I578088);
and I_41806 (I713761,I713744,I578091);
or I_41807 (I713778,I713761,I578073);
DFFARX1 I_41808 (I713778,I3035,I713323,I713804,);
not I_41809 (I713812,I713804);
nand I_41810 (I713829,I713812,I713552);
not I_41811 (I713303,I713829);
nand I_41812 (I713297,I713829,I713569);
nand I_41813 (I713294,I713812,I713436);
not I_41814 (I713918,I3042);
DFFARX1 I_41815 (I395545,I3035,I713918,I713944,);
DFFARX1 I_41816 (I395527,I3035,I713918,I713961,);
not I_41817 (I713969,I713961);
nor I_41818 (I713886,I713944,I713969);
DFFARX1 I_41819 (I713969,I3035,I713918,I713901,);
nor I_41820 (I714014,I395533,I395536);
and I_41821 (I714031,I714014,I395524);
nor I_41822 (I714048,I714031,I395533);
not I_41823 (I714065,I395533);
and I_41824 (I714082,I714065,I395542);
nand I_41825 (I714099,I714082,I395530);
nor I_41826 (I714116,I714065,I714099);
DFFARX1 I_41827 (I714116,I3035,I713918,I713883,);
not I_41828 (I714147,I714099);
nand I_41829 (I714164,I713969,I714147);
nand I_41830 (I713895,I714031,I714147);
DFFARX1 I_41831 (I714065,I3035,I713918,I713910,);
not I_41832 (I714209,I395527);
nor I_41833 (I714226,I714209,I395542);
nor I_41834 (I714243,I714226,I714048);
DFFARX1 I_41835 (I714243,I3035,I713918,I713907,);
not I_41836 (I714274,I714226);
DFFARX1 I_41837 (I714274,I3035,I713918,I714300,);
not I_41838 (I714308,I714300);
nor I_41839 (I713904,I714308,I714226);
nor I_41840 (I714339,I714209,I395539);
and I_41841 (I714356,I714339,I395548);
or I_41842 (I714373,I714356,I395524);
DFFARX1 I_41843 (I714373,I3035,I713918,I714399,);
not I_41844 (I714407,I714399);
nand I_41845 (I714424,I714407,I714147);
not I_41846 (I713898,I714424);
nand I_41847 (I713892,I714424,I714164);
nand I_41848 (I713889,I714407,I714031);
not I_41849 (I714513,I3042);
DFFARX1 I_41850 (I248933,I3035,I714513,I714539,);
DFFARX1 I_41851 (I248939,I3035,I714513,I714556,);
not I_41852 (I714564,I714556);
nor I_41853 (I714481,I714539,I714564);
DFFARX1 I_41854 (I714564,I3035,I714513,I714496,);
nor I_41855 (I714609,I248948,I248933);
and I_41856 (I714626,I714609,I248960);
nor I_41857 (I714643,I714626,I248948);
not I_41858 (I714660,I248948);
and I_41859 (I714677,I714660,I248936);
nand I_41860 (I714694,I714677,I248957);
nor I_41861 (I714711,I714660,I714694);
DFFARX1 I_41862 (I714711,I3035,I714513,I714478,);
not I_41863 (I714742,I714694);
nand I_41864 (I714759,I714564,I714742);
nand I_41865 (I714490,I714626,I714742);
DFFARX1 I_41866 (I714660,I3035,I714513,I714505,);
not I_41867 (I714804,I248945);
nor I_41868 (I714821,I714804,I248936);
nor I_41869 (I714838,I714821,I714643);
DFFARX1 I_41870 (I714838,I3035,I714513,I714502,);
not I_41871 (I714869,I714821);
DFFARX1 I_41872 (I714869,I3035,I714513,I714895,);
not I_41873 (I714903,I714895);
nor I_41874 (I714499,I714903,I714821);
nor I_41875 (I714934,I714804,I248942);
and I_41876 (I714951,I714934,I248954);
or I_41877 (I714968,I714951,I248951);
DFFARX1 I_41878 (I714968,I3035,I714513,I714994,);
not I_41879 (I715002,I714994);
nand I_41880 (I715019,I715002,I714742);
not I_41881 (I714493,I715019);
nand I_41882 (I714487,I715019,I714759);
nand I_41883 (I714484,I715002,I714626);
not I_41884 (I715108,I3042);
DFFARX1 I_41885 (I503854,I3035,I715108,I715134,);
DFFARX1 I_41886 (I503872,I3035,I715108,I715151,);
not I_41887 (I715159,I715151);
nor I_41888 (I715076,I715134,I715159);
DFFARX1 I_41889 (I715159,I3035,I715108,I715091,);
nor I_41890 (I715204,I503851,I503863);
and I_41891 (I715221,I715204,I503848);
nor I_41892 (I715238,I715221,I503851);
not I_41893 (I715255,I503851);
and I_41894 (I715272,I715255,I503857);
nand I_41895 (I715289,I715272,I503869);
nor I_41896 (I715306,I715255,I715289);
DFFARX1 I_41897 (I715306,I3035,I715108,I715073,);
not I_41898 (I715337,I715289);
nand I_41899 (I715354,I715159,I715337);
nand I_41900 (I715085,I715221,I715337);
DFFARX1 I_41901 (I715255,I3035,I715108,I715100,);
not I_41902 (I715399,I503860);
nor I_41903 (I715416,I715399,I503857);
nor I_41904 (I715433,I715416,I715238);
DFFARX1 I_41905 (I715433,I3035,I715108,I715097,);
not I_41906 (I715464,I715416);
DFFARX1 I_41907 (I715464,I3035,I715108,I715490,);
not I_41908 (I715498,I715490);
nor I_41909 (I715094,I715498,I715416);
nor I_41910 (I715529,I715399,I503848);
and I_41911 (I715546,I715529,I503875);
or I_41912 (I715563,I715546,I503866);
DFFARX1 I_41913 (I715563,I3035,I715108,I715589,);
not I_41914 (I715597,I715589);
nand I_41915 (I715614,I715597,I715337);
not I_41916 (I715088,I715614);
nand I_41917 (I715082,I715614,I715354);
nand I_41918 (I715079,I715597,I715221);
not I_41919 (I715703,I3042);
DFFARX1 I_41920 (I581541,I3035,I715703,I715729,);
DFFARX1 I_41921 (I581553,I3035,I715703,I715746,);
not I_41922 (I715754,I715746);
nor I_41923 (I715671,I715729,I715754);
DFFARX1 I_41924 (I715754,I3035,I715703,I715686,);
nor I_41925 (I715799,I581550,I581544);
and I_41926 (I715816,I715799,I581538);
nor I_41927 (I715833,I715816,I581550);
not I_41928 (I715850,I581550);
and I_41929 (I715867,I715850,I581547);
nand I_41930 (I715884,I715867,I581538);
nor I_41931 (I715901,I715850,I715884);
DFFARX1 I_41932 (I715901,I3035,I715703,I715668,);
not I_41933 (I715932,I715884);
nand I_41934 (I715949,I715754,I715932);
nand I_41935 (I715680,I715816,I715932);
DFFARX1 I_41936 (I715850,I3035,I715703,I715695,);
not I_41937 (I715994,I581562);
nor I_41938 (I716011,I715994,I581547);
nor I_41939 (I716028,I716011,I715833);
DFFARX1 I_41940 (I716028,I3035,I715703,I715692,);
not I_41941 (I716059,I716011);
DFFARX1 I_41942 (I716059,I3035,I715703,I716085,);
not I_41943 (I716093,I716085);
nor I_41944 (I715689,I716093,I716011);
nor I_41945 (I716124,I715994,I581556);
and I_41946 (I716141,I716124,I581559);
or I_41947 (I716158,I716141,I581541);
DFFARX1 I_41948 (I716158,I3035,I715703,I716184,);
not I_41949 (I716192,I716184);
nand I_41950 (I716209,I716192,I715932);
not I_41951 (I715683,I716209);
nand I_41952 (I715677,I716209,I715949);
nand I_41953 (I715674,I716192,I715816);
not I_41954 (I716298,I3042);
DFFARX1 I_41955 (I136614,I3035,I716298,I716324,);
DFFARX1 I_41956 (I136617,I3035,I716298,I716341,);
not I_41957 (I716349,I716341);
nor I_41958 (I716266,I716324,I716349);
DFFARX1 I_41959 (I716349,I3035,I716298,I716281,);
nor I_41960 (I716394,I136623,I136617);
and I_41961 (I716411,I716394,I136620);
nor I_41962 (I716428,I716411,I136623);
not I_41963 (I716445,I136623);
and I_41964 (I716462,I716445,I136614);
nand I_41965 (I716479,I716462,I136632);
nor I_41966 (I716496,I716445,I716479);
DFFARX1 I_41967 (I716496,I3035,I716298,I716263,);
not I_41968 (I716527,I716479);
nand I_41969 (I716544,I716349,I716527);
nand I_41970 (I716275,I716411,I716527);
DFFARX1 I_41971 (I716445,I3035,I716298,I716290,);
not I_41972 (I716589,I136626);
nor I_41973 (I716606,I716589,I136614);
nor I_41974 (I716623,I716606,I716428);
DFFARX1 I_41975 (I716623,I3035,I716298,I716287,);
not I_41976 (I716654,I716606);
DFFARX1 I_41977 (I716654,I3035,I716298,I716680,);
not I_41978 (I716688,I716680);
nor I_41979 (I716284,I716688,I716606);
nor I_41980 (I716719,I716589,I136629);
and I_41981 (I716736,I716719,I136635);
or I_41982 (I716753,I716736,I136638);
DFFARX1 I_41983 (I716753,I3035,I716298,I716779,);
not I_41984 (I716787,I716779);
nand I_41985 (I716804,I716787,I716527);
not I_41986 (I716278,I716804);
nand I_41987 (I716272,I716804,I716544);
nand I_41988 (I716269,I716787,I716411);
not I_41989 (I716893,I3042);
DFFARX1 I_41990 (I364333,I3035,I716893,I716919,);
DFFARX1 I_41991 (I364315,I3035,I716893,I716936,);
not I_41992 (I716944,I716936);
nor I_41993 (I716861,I716919,I716944);
DFFARX1 I_41994 (I716944,I3035,I716893,I716876,);
nor I_41995 (I716989,I364321,I364324);
and I_41996 (I717006,I716989,I364312);
nor I_41997 (I717023,I717006,I364321);
not I_41998 (I717040,I364321);
and I_41999 (I717057,I717040,I364330);
nand I_42000 (I717074,I717057,I364318);
nor I_42001 (I717091,I717040,I717074);
DFFARX1 I_42002 (I717091,I3035,I716893,I716858,);
not I_42003 (I717122,I717074);
nand I_42004 (I717139,I716944,I717122);
nand I_42005 (I716870,I717006,I717122);
DFFARX1 I_42006 (I717040,I3035,I716893,I716885,);
not I_42007 (I717184,I364315);
nor I_42008 (I717201,I717184,I364330);
nor I_42009 (I717218,I717201,I717023);
DFFARX1 I_42010 (I717218,I3035,I716893,I716882,);
not I_42011 (I717249,I717201);
DFFARX1 I_42012 (I717249,I3035,I716893,I717275,);
not I_42013 (I717283,I717275);
nor I_42014 (I716879,I717283,I717201);
nor I_42015 (I717314,I717184,I364327);
and I_42016 (I717331,I717314,I364336);
or I_42017 (I717348,I717331,I364312);
DFFARX1 I_42018 (I717348,I3035,I716893,I717374,);
not I_42019 (I717382,I717374);
nand I_42020 (I717399,I717382,I717122);
not I_42021 (I716873,I717399);
nand I_42022 (I716867,I717399,I717139);
nand I_42023 (I716864,I717382,I717006);
not I_42024 (I717488,I3042);
DFFARX1 I_42025 (I152955,I3035,I717488,I717514,);
DFFARX1 I_42026 (I152949,I3035,I717488,I717531,);
not I_42027 (I717539,I717531);
nor I_42028 (I717456,I717514,I717539);
DFFARX1 I_42029 (I717539,I3035,I717488,I717471,);
nor I_42030 (I717584,I152937,I152958);
and I_42031 (I717601,I717584,I152952);
nor I_42032 (I717618,I717601,I152937);
not I_42033 (I717635,I152937);
and I_42034 (I717652,I717635,I152934);
nand I_42035 (I717669,I717652,I152946);
nor I_42036 (I717686,I717635,I717669);
DFFARX1 I_42037 (I717686,I3035,I717488,I717453,);
not I_42038 (I717717,I717669);
nand I_42039 (I717734,I717539,I717717);
nand I_42040 (I717465,I717601,I717717);
DFFARX1 I_42041 (I717635,I3035,I717488,I717480,);
not I_42042 (I717779,I152961);
nor I_42043 (I717796,I717779,I152934);
nor I_42044 (I717813,I717796,I717618);
DFFARX1 I_42045 (I717813,I3035,I717488,I717477,);
not I_42046 (I717844,I717796);
DFFARX1 I_42047 (I717844,I3035,I717488,I717870,);
not I_42048 (I717878,I717870);
nor I_42049 (I717474,I717878,I717796);
nor I_42050 (I717909,I717779,I152943);
and I_42051 (I717926,I717909,I152940);
or I_42052 (I717943,I717926,I152934);
DFFARX1 I_42053 (I717943,I3035,I717488,I717969,);
not I_42054 (I717977,I717969);
nand I_42055 (I717994,I717977,I717717);
not I_42056 (I717468,I717994);
nand I_42057 (I717462,I717994,I717734);
nand I_42058 (I717459,I717977,I717601);
not I_42059 (I718083,I3042);
DFFARX1 I_42060 (I140779,I3035,I718083,I718109,);
DFFARX1 I_42061 (I140782,I3035,I718083,I718126,);
not I_42062 (I718134,I718126);
nor I_42063 (I718051,I718109,I718134);
DFFARX1 I_42064 (I718134,I3035,I718083,I718066,);
nor I_42065 (I718179,I140788,I140782);
and I_42066 (I718196,I718179,I140785);
nor I_42067 (I718213,I718196,I140788);
not I_42068 (I718230,I140788);
and I_42069 (I718247,I718230,I140779);
nand I_42070 (I718264,I718247,I140797);
nor I_42071 (I718281,I718230,I718264);
DFFARX1 I_42072 (I718281,I3035,I718083,I718048,);
not I_42073 (I718312,I718264);
nand I_42074 (I718329,I718134,I718312);
nand I_42075 (I718060,I718196,I718312);
DFFARX1 I_42076 (I718230,I3035,I718083,I718075,);
not I_42077 (I718374,I140791);
nor I_42078 (I718391,I718374,I140779);
nor I_42079 (I718408,I718391,I718213);
DFFARX1 I_42080 (I718408,I3035,I718083,I718072,);
not I_42081 (I718439,I718391);
DFFARX1 I_42082 (I718439,I3035,I718083,I718465,);
not I_42083 (I718473,I718465);
nor I_42084 (I718069,I718473,I718391);
nor I_42085 (I718504,I718374,I140794);
and I_42086 (I718521,I718504,I140800);
or I_42087 (I718538,I718521,I140803);
DFFARX1 I_42088 (I718538,I3035,I718083,I718564,);
not I_42089 (I718572,I718564);
nand I_42090 (I718589,I718572,I718312);
not I_42091 (I718063,I718589);
nand I_42092 (I718057,I718589,I718329);
nand I_42093 (I718054,I718572,I718196);
not I_42094 (I718678,I3042);
DFFARX1 I_42095 (I523234,I3035,I718678,I718704,);
DFFARX1 I_42096 (I523252,I3035,I718678,I718721,);
not I_42097 (I718729,I718721);
nor I_42098 (I718646,I718704,I718729);
DFFARX1 I_42099 (I718729,I3035,I718678,I718661,);
nor I_42100 (I718774,I523231,I523243);
and I_42101 (I718791,I718774,I523228);
nor I_42102 (I718808,I718791,I523231);
not I_42103 (I718825,I523231);
and I_42104 (I718842,I718825,I523237);
nand I_42105 (I718859,I718842,I523249);
nor I_42106 (I718876,I718825,I718859);
DFFARX1 I_42107 (I718876,I3035,I718678,I718643,);
not I_42108 (I718907,I718859);
nand I_42109 (I718924,I718729,I718907);
nand I_42110 (I718655,I718791,I718907);
DFFARX1 I_42111 (I718825,I3035,I718678,I718670,);
not I_42112 (I718969,I523240);
nor I_42113 (I718986,I718969,I523237);
nor I_42114 (I719003,I718986,I718808);
DFFARX1 I_42115 (I719003,I3035,I718678,I718667,);
not I_42116 (I719034,I718986);
DFFARX1 I_42117 (I719034,I3035,I718678,I719060,);
not I_42118 (I719068,I719060);
nor I_42119 (I718664,I719068,I718986);
nor I_42120 (I719099,I718969,I523228);
and I_42121 (I719116,I719099,I523255);
or I_42122 (I719133,I719116,I523246);
DFFARX1 I_42123 (I719133,I3035,I718678,I719159,);
not I_42124 (I719167,I719159);
nand I_42125 (I719184,I719167,I718907);
not I_42126 (I718658,I719184);
nand I_42127 (I718652,I719184,I718924);
nand I_42128 (I718649,I719167,I718791);
not I_42129 (I719273,I3042);
DFFARX1 I_42130 (I37865,I3035,I719273,I719299,);
DFFARX1 I_42131 (I37853,I3035,I719273,I719316,);
not I_42132 (I719324,I719316);
nor I_42133 (I719241,I719299,I719324);
DFFARX1 I_42134 (I719324,I3035,I719273,I719256,);
nor I_42135 (I719369,I37844,I37868);
and I_42136 (I719386,I719369,I37847);
nor I_42137 (I719403,I719386,I37844);
not I_42138 (I719420,I37844);
and I_42139 (I719437,I719420,I37850);
nand I_42140 (I719454,I719437,I37862);
nor I_42141 (I719471,I719420,I719454);
DFFARX1 I_42142 (I719471,I3035,I719273,I719238,);
not I_42143 (I719502,I719454);
nand I_42144 (I719519,I719324,I719502);
nand I_42145 (I719250,I719386,I719502);
DFFARX1 I_42146 (I719420,I3035,I719273,I719265,);
not I_42147 (I719564,I37844);
nor I_42148 (I719581,I719564,I37850);
nor I_42149 (I719598,I719581,I719403);
DFFARX1 I_42150 (I719598,I3035,I719273,I719262,);
not I_42151 (I719629,I719581);
DFFARX1 I_42152 (I719629,I3035,I719273,I719655,);
not I_42153 (I719663,I719655);
nor I_42154 (I719259,I719663,I719581);
nor I_42155 (I719694,I719564,I37847);
and I_42156 (I719711,I719694,I37856);
or I_42157 (I719728,I719711,I37859);
DFFARX1 I_42158 (I719728,I3035,I719273,I719754,);
not I_42159 (I719762,I719754);
nand I_42160 (I719779,I719762,I719502);
not I_42161 (I719253,I719779);
nand I_42162 (I719247,I719779,I719519);
nand I_42163 (I719244,I719762,I719386);
not I_42164 (I719868,I3042);
DFFARX1 I_42165 (I492872,I3035,I719868,I719894,);
DFFARX1 I_42166 (I492890,I3035,I719868,I719911,);
not I_42167 (I719919,I719911);
nor I_42168 (I719836,I719894,I719919);
DFFARX1 I_42169 (I719919,I3035,I719868,I719851,);
nor I_42170 (I719964,I492869,I492881);
and I_42171 (I719981,I719964,I492866);
nor I_42172 (I719998,I719981,I492869);
not I_42173 (I720015,I492869);
and I_42174 (I720032,I720015,I492875);
nand I_42175 (I720049,I720032,I492887);
nor I_42176 (I720066,I720015,I720049);
DFFARX1 I_42177 (I720066,I3035,I719868,I719833,);
not I_42178 (I720097,I720049);
nand I_42179 (I720114,I719919,I720097);
nand I_42180 (I719845,I719981,I720097);
DFFARX1 I_42181 (I720015,I3035,I719868,I719860,);
not I_42182 (I720159,I492878);
nor I_42183 (I720176,I720159,I492875);
nor I_42184 (I720193,I720176,I719998);
DFFARX1 I_42185 (I720193,I3035,I719868,I719857,);
not I_42186 (I720224,I720176);
DFFARX1 I_42187 (I720224,I3035,I719868,I720250,);
not I_42188 (I720258,I720250);
nor I_42189 (I719854,I720258,I720176);
nor I_42190 (I720289,I720159,I492866);
and I_42191 (I720306,I720289,I492893);
or I_42192 (I720323,I720306,I492884);
DFFARX1 I_42193 (I720323,I3035,I719868,I720349,);
not I_42194 (I720357,I720349);
nand I_42195 (I720374,I720357,I720097);
not I_42196 (I719848,I720374);
nand I_42197 (I719842,I720374,I720114);
nand I_42198 (I719839,I720357,I719981);
not I_42199 (I720463,I3042);
DFFARX1 I_42200 (I388609,I3035,I720463,I720489,);
DFFARX1 I_42201 (I388591,I3035,I720463,I720506,);
not I_42202 (I720514,I720506);
nor I_42203 (I720431,I720489,I720514);
DFFARX1 I_42204 (I720514,I3035,I720463,I720446,);
nor I_42205 (I720559,I388597,I388600);
and I_42206 (I720576,I720559,I388588);
nor I_42207 (I720593,I720576,I388597);
not I_42208 (I720610,I388597);
and I_42209 (I720627,I720610,I388606);
nand I_42210 (I720644,I720627,I388594);
nor I_42211 (I720661,I720610,I720644);
DFFARX1 I_42212 (I720661,I3035,I720463,I720428,);
not I_42213 (I720692,I720644);
nand I_42214 (I720709,I720514,I720692);
nand I_42215 (I720440,I720576,I720692);
DFFARX1 I_42216 (I720610,I3035,I720463,I720455,);
not I_42217 (I720754,I388591);
nor I_42218 (I720771,I720754,I388606);
nor I_42219 (I720788,I720771,I720593);
DFFARX1 I_42220 (I720788,I3035,I720463,I720452,);
not I_42221 (I720819,I720771);
DFFARX1 I_42222 (I720819,I3035,I720463,I720845,);
not I_42223 (I720853,I720845);
nor I_42224 (I720449,I720853,I720771);
nor I_42225 (I720884,I720754,I388603);
and I_42226 (I720901,I720884,I388612);
or I_42227 (I720918,I720901,I388588);
DFFARX1 I_42228 (I720918,I3035,I720463,I720944,);
not I_42229 (I720952,I720944);
nand I_42230 (I720969,I720952,I720692);
not I_42231 (I720443,I720969);
nand I_42232 (I720437,I720969,I720709);
nand I_42233 (I720434,I720952,I720576);
not I_42234 (I721058,I3042);
DFFARX1 I_42235 (I99724,I3035,I721058,I721084,);
DFFARX1 I_42236 (I99727,I3035,I721058,I721101,);
not I_42237 (I721109,I721101);
nor I_42238 (I721026,I721084,I721109);
DFFARX1 I_42239 (I721109,I3035,I721058,I721041,);
nor I_42240 (I721154,I99733,I99727);
and I_42241 (I721171,I721154,I99730);
nor I_42242 (I721188,I721171,I99733);
not I_42243 (I721205,I99733);
and I_42244 (I721222,I721205,I99724);
nand I_42245 (I721239,I721222,I99742);
nor I_42246 (I721256,I721205,I721239);
DFFARX1 I_42247 (I721256,I3035,I721058,I721023,);
not I_42248 (I721287,I721239);
nand I_42249 (I721304,I721109,I721287);
nand I_42250 (I721035,I721171,I721287);
DFFARX1 I_42251 (I721205,I3035,I721058,I721050,);
not I_42252 (I721349,I99736);
nor I_42253 (I721366,I721349,I99724);
nor I_42254 (I721383,I721366,I721188);
DFFARX1 I_42255 (I721383,I3035,I721058,I721047,);
not I_42256 (I721414,I721366);
DFFARX1 I_42257 (I721414,I3035,I721058,I721440,);
not I_42258 (I721448,I721440);
nor I_42259 (I721044,I721448,I721366);
nor I_42260 (I721479,I721349,I99739);
and I_42261 (I721496,I721479,I99745);
or I_42262 (I721513,I721496,I99748);
DFFARX1 I_42263 (I721513,I3035,I721058,I721539,);
not I_42264 (I721547,I721539);
nand I_42265 (I721564,I721547,I721287);
not I_42266 (I721038,I721564);
nand I_42267 (I721032,I721564,I721304);
nand I_42268 (I721029,I721547,I721171);
not I_42269 (I721653,I3042);
DFFARX1 I_42270 (I166657,I3035,I721653,I721679,);
DFFARX1 I_42271 (I166651,I3035,I721653,I721696,);
not I_42272 (I721704,I721696);
nor I_42273 (I721621,I721679,I721704);
DFFARX1 I_42274 (I721704,I3035,I721653,I721636,);
nor I_42275 (I721749,I166639,I166660);
and I_42276 (I721766,I721749,I166654);
nor I_42277 (I721783,I721766,I166639);
not I_42278 (I721800,I166639);
and I_42279 (I721817,I721800,I166636);
nand I_42280 (I721834,I721817,I166648);
nor I_42281 (I721851,I721800,I721834);
DFFARX1 I_42282 (I721851,I3035,I721653,I721618,);
not I_42283 (I721882,I721834);
nand I_42284 (I721899,I721704,I721882);
nand I_42285 (I721630,I721766,I721882);
DFFARX1 I_42286 (I721800,I3035,I721653,I721645,);
not I_42287 (I721944,I166663);
nor I_42288 (I721961,I721944,I166636);
nor I_42289 (I721978,I721961,I721783);
DFFARX1 I_42290 (I721978,I3035,I721653,I721642,);
not I_42291 (I722009,I721961);
DFFARX1 I_42292 (I722009,I3035,I721653,I722035,);
not I_42293 (I722043,I722035);
nor I_42294 (I721639,I722043,I721961);
nor I_42295 (I722074,I721944,I166645);
and I_42296 (I722091,I722074,I166642);
or I_42297 (I722108,I722091,I166636);
DFFARX1 I_42298 (I722108,I3035,I721653,I722134,);
not I_42299 (I722142,I722134);
nand I_42300 (I722159,I722142,I721882);
not I_42301 (I721633,I722159);
nand I_42302 (I721627,I722159,I721899);
nand I_42303 (I721624,I722142,I721766);
not I_42304 (I722248,I3042);
DFFARX1 I_42305 (I487058,I3035,I722248,I722274,);
DFFARX1 I_42306 (I487076,I3035,I722248,I722291,);
not I_42307 (I722299,I722291);
nor I_42308 (I722216,I722274,I722299);
DFFARX1 I_42309 (I722299,I3035,I722248,I722231,);
nor I_42310 (I722344,I487055,I487067);
and I_42311 (I722361,I722344,I487052);
nor I_42312 (I722378,I722361,I487055);
not I_42313 (I722395,I487055);
and I_42314 (I722412,I722395,I487061);
nand I_42315 (I722429,I722412,I487073);
nor I_42316 (I722446,I722395,I722429);
DFFARX1 I_42317 (I722446,I3035,I722248,I722213,);
not I_42318 (I722477,I722429);
nand I_42319 (I722494,I722299,I722477);
nand I_42320 (I722225,I722361,I722477);
DFFARX1 I_42321 (I722395,I3035,I722248,I722240,);
not I_42322 (I722539,I487064);
nor I_42323 (I722556,I722539,I487061);
nor I_42324 (I722573,I722556,I722378);
DFFARX1 I_42325 (I722573,I3035,I722248,I722237,);
not I_42326 (I722604,I722556);
DFFARX1 I_42327 (I722604,I3035,I722248,I722630,);
not I_42328 (I722638,I722630);
nor I_42329 (I722234,I722638,I722556);
nor I_42330 (I722669,I722539,I487052);
and I_42331 (I722686,I722669,I487079);
or I_42332 (I722703,I722686,I487070);
DFFARX1 I_42333 (I722703,I3035,I722248,I722729,);
not I_42334 (I722737,I722729);
nand I_42335 (I722754,I722737,I722477);
not I_42336 (I722228,I722754);
nand I_42337 (I722222,I722754,I722494);
nand I_42338 (I722219,I722737,I722361);
not I_42339 (I722843,I3042);
DFFARX1 I_42340 (I462496,I3035,I722843,I722869,);
DFFARX1 I_42341 (I462493,I3035,I722843,I722886,);
not I_42342 (I722894,I722886);
nor I_42343 (I722811,I722869,I722894);
DFFARX1 I_42344 (I722894,I3035,I722843,I722826,);
nor I_42345 (I722939,I462508,I462490);
and I_42346 (I722956,I722939,I462487);
nor I_42347 (I722973,I722956,I462508);
not I_42348 (I722990,I462508);
and I_42349 (I723007,I722990,I462493);
nand I_42350 (I723024,I723007,I462505);
nor I_42351 (I723041,I722990,I723024);
DFFARX1 I_42352 (I723041,I3035,I722843,I722808,);
not I_42353 (I723072,I723024);
nand I_42354 (I723089,I722894,I723072);
nand I_42355 (I722820,I722956,I723072);
DFFARX1 I_42356 (I722990,I3035,I722843,I722835,);
not I_42357 (I723134,I462499);
nor I_42358 (I723151,I723134,I462493);
nor I_42359 (I723168,I723151,I722973);
DFFARX1 I_42360 (I723168,I3035,I722843,I722832,);
not I_42361 (I723199,I723151);
DFFARX1 I_42362 (I723199,I3035,I722843,I723225,);
not I_42363 (I723233,I723225);
nor I_42364 (I722829,I723233,I723151);
nor I_42365 (I723264,I723134,I462487);
and I_42366 (I723281,I723264,I462502);
or I_42367 (I723298,I723281,I462490);
DFFARX1 I_42368 (I723298,I3035,I722843,I723324,);
not I_42369 (I723332,I723324);
nand I_42370 (I723349,I723332,I723072);
not I_42371 (I722823,I723349);
nand I_42372 (I722817,I723349,I723089);
nand I_42373 (I722814,I723332,I722956);
not I_42374 (I723438,I3042);
DFFARX1 I_42375 (I389187,I3035,I723438,I723464,);
DFFARX1 I_42376 (I389169,I3035,I723438,I723481,);
not I_42377 (I723489,I723481);
nor I_42378 (I723406,I723464,I723489);
DFFARX1 I_42379 (I723489,I3035,I723438,I723421,);
nor I_42380 (I723534,I389175,I389178);
and I_42381 (I723551,I723534,I389166);
nor I_42382 (I723568,I723551,I389175);
not I_42383 (I723585,I389175);
and I_42384 (I723602,I723585,I389184);
nand I_42385 (I723619,I723602,I389172);
nor I_42386 (I723636,I723585,I723619);
DFFARX1 I_42387 (I723636,I3035,I723438,I723403,);
not I_42388 (I723667,I723619);
nand I_42389 (I723684,I723489,I723667);
nand I_42390 (I723415,I723551,I723667);
DFFARX1 I_42391 (I723585,I3035,I723438,I723430,);
not I_42392 (I723729,I389169);
nor I_42393 (I723746,I723729,I389184);
nor I_42394 (I723763,I723746,I723568);
DFFARX1 I_42395 (I723763,I3035,I723438,I723427,);
not I_42396 (I723794,I723746);
DFFARX1 I_42397 (I723794,I3035,I723438,I723820,);
not I_42398 (I723828,I723820);
nor I_42399 (I723424,I723828,I723746);
nor I_42400 (I723859,I723729,I389181);
and I_42401 (I723876,I723859,I389190);
or I_42402 (I723893,I723876,I389166);
DFFARX1 I_42403 (I723893,I3035,I723438,I723919,);
not I_42404 (I723927,I723919);
nand I_42405 (I723944,I723927,I723667);
not I_42406 (I723418,I723944);
nand I_42407 (I723412,I723944,I723684);
nand I_42408 (I723409,I723927,I723551);
not I_42409 (I724033,I3042);
DFFARX1 I_42410 (I461442,I3035,I724033,I724059,);
DFFARX1 I_42411 (I461439,I3035,I724033,I724076,);
not I_42412 (I724084,I724076);
nor I_42413 (I724001,I724059,I724084);
DFFARX1 I_42414 (I724084,I3035,I724033,I724016,);
nor I_42415 (I724129,I461454,I461436);
and I_42416 (I724146,I724129,I461433);
nor I_42417 (I724163,I724146,I461454);
not I_42418 (I724180,I461454);
and I_42419 (I724197,I724180,I461439);
nand I_42420 (I724214,I724197,I461451);
nor I_42421 (I724231,I724180,I724214);
DFFARX1 I_42422 (I724231,I3035,I724033,I723998,);
not I_42423 (I724262,I724214);
nand I_42424 (I724279,I724084,I724262);
nand I_42425 (I724010,I724146,I724262);
DFFARX1 I_42426 (I724180,I3035,I724033,I724025,);
not I_42427 (I724324,I461445);
nor I_42428 (I724341,I724324,I461439);
nor I_42429 (I724358,I724341,I724163);
DFFARX1 I_42430 (I724358,I3035,I724033,I724022,);
not I_42431 (I724389,I724341);
DFFARX1 I_42432 (I724389,I3035,I724033,I724415,);
not I_42433 (I724423,I724415);
nor I_42434 (I724019,I724423,I724341);
nor I_42435 (I724454,I724324,I461433);
and I_42436 (I724471,I724454,I461448);
or I_42437 (I724488,I724471,I461436);
DFFARX1 I_42438 (I724488,I3035,I724033,I724514,);
not I_42439 (I724522,I724514);
nand I_42440 (I724539,I724522,I724262);
not I_42441 (I724013,I724539);
nand I_42442 (I724007,I724539,I724279);
nand I_42443 (I724004,I724522,I724146);
not I_42444 (I724628,I3042);
DFFARX1 I_42445 (I658310,I3035,I724628,I724654,);
DFFARX1 I_42446 (I658313,I3035,I724628,I724671,);
not I_42447 (I724679,I724671);
nor I_42448 (I724596,I724654,I724679);
DFFARX1 I_42449 (I724679,I3035,I724628,I724611,);
nor I_42450 (I724724,I658313,I658328);
and I_42451 (I724741,I724724,I658322);
nor I_42452 (I724758,I724741,I658313);
not I_42453 (I724775,I658313);
and I_42454 (I724792,I724775,I658331);
nand I_42455 (I724809,I724792,I658319);
nor I_42456 (I724826,I724775,I724809);
DFFARX1 I_42457 (I724826,I3035,I724628,I724593,);
not I_42458 (I724857,I724809);
nand I_42459 (I724874,I724679,I724857);
nand I_42460 (I724605,I724741,I724857);
DFFARX1 I_42461 (I724775,I3035,I724628,I724620,);
not I_42462 (I724919,I658325);
nor I_42463 (I724936,I724919,I658331);
nor I_42464 (I724953,I724936,I724758);
DFFARX1 I_42465 (I724953,I3035,I724628,I724617,);
not I_42466 (I724984,I724936);
DFFARX1 I_42467 (I724984,I3035,I724628,I725010,);
not I_42468 (I725018,I725010);
nor I_42469 (I724614,I725018,I724936);
nor I_42470 (I725049,I724919,I658310);
and I_42471 (I725066,I725049,I658334);
or I_42472 (I725083,I725066,I658316);
DFFARX1 I_42473 (I725083,I3035,I724628,I725109,);
not I_42474 (I725117,I725109);
nand I_42475 (I725134,I725117,I724857);
not I_42476 (I724608,I725134);
nand I_42477 (I724602,I725134,I724874);
nand I_42478 (I724599,I725117,I724741);
not I_42479 (I725223,I3042);
DFFARX1 I_42480 (I641653,I3035,I725223,I725249,);
DFFARX1 I_42481 (I641665,I3035,I725223,I725266,);
not I_42482 (I725274,I725266);
nor I_42483 (I725191,I725249,I725274);
DFFARX1 I_42484 (I725274,I3035,I725223,I725206,);
nor I_42485 (I725319,I641662,I641656);
and I_42486 (I725336,I725319,I641650);
nor I_42487 (I725353,I725336,I641662);
not I_42488 (I725370,I641662);
and I_42489 (I725387,I725370,I641659);
nand I_42490 (I725404,I725387,I641650);
nor I_42491 (I725421,I725370,I725404);
DFFARX1 I_42492 (I725421,I3035,I725223,I725188,);
not I_42493 (I725452,I725404);
nand I_42494 (I725469,I725274,I725452);
nand I_42495 (I725200,I725336,I725452);
DFFARX1 I_42496 (I725370,I3035,I725223,I725215,);
not I_42497 (I725514,I641674);
nor I_42498 (I725531,I725514,I641659);
nor I_42499 (I725548,I725531,I725353);
DFFARX1 I_42500 (I725548,I3035,I725223,I725212,);
not I_42501 (I725579,I725531);
DFFARX1 I_42502 (I725579,I3035,I725223,I725605,);
not I_42503 (I725613,I725605);
nor I_42504 (I725209,I725613,I725531);
nor I_42505 (I725644,I725514,I641668);
and I_42506 (I725661,I725644,I641671);
or I_42507 (I725678,I725661,I641653);
DFFARX1 I_42508 (I725678,I3035,I725223,I725704,);
not I_42509 (I725712,I725704);
nand I_42510 (I725729,I725712,I725452);
not I_42511 (I725203,I725729);
nand I_42512 (I725197,I725729,I725469);
nand I_42513 (I725194,I725712,I725336);
not I_42514 (I725818,I3042);
DFFARX1 I_42515 (I55783,I3035,I725818,I725844,);
DFFARX1 I_42516 (I55771,I3035,I725818,I725861,);
not I_42517 (I725869,I725861);
nor I_42518 (I725786,I725844,I725869);
DFFARX1 I_42519 (I725869,I3035,I725818,I725801,);
nor I_42520 (I725914,I55762,I55786);
and I_42521 (I725931,I725914,I55765);
nor I_42522 (I725948,I725931,I55762);
not I_42523 (I725965,I55762);
and I_42524 (I725982,I725965,I55768);
nand I_42525 (I725999,I725982,I55780);
nor I_42526 (I726016,I725965,I725999);
DFFARX1 I_42527 (I726016,I3035,I725818,I725783,);
not I_42528 (I726047,I725999);
nand I_42529 (I726064,I725869,I726047);
nand I_42530 (I725795,I725931,I726047);
DFFARX1 I_42531 (I725965,I3035,I725818,I725810,);
not I_42532 (I726109,I55762);
nor I_42533 (I726126,I726109,I55768);
nor I_42534 (I726143,I726126,I725948);
DFFARX1 I_42535 (I726143,I3035,I725818,I725807,);
not I_42536 (I726174,I726126);
DFFARX1 I_42537 (I726174,I3035,I725818,I726200,);
not I_42538 (I726208,I726200);
nor I_42539 (I725804,I726208,I726126);
nor I_42540 (I726239,I726109,I55765);
and I_42541 (I726256,I726239,I55774);
or I_42542 (I726273,I726256,I55777);
DFFARX1 I_42543 (I726273,I3035,I725818,I726299,);
not I_42544 (I726307,I726299);
nand I_42545 (I726324,I726307,I726047);
not I_42546 (I725798,I726324);
nand I_42547 (I725792,I726324,I726064);
nand I_42548 (I725789,I726307,I725931);
not I_42549 (I726413,I3042);
DFFARX1 I_42550 (I217249,I3035,I726413,I726439,);
DFFARX1 I_42551 (I217243,I3035,I726413,I726456,);
not I_42552 (I726464,I726456);
nor I_42553 (I726381,I726439,I726464);
DFFARX1 I_42554 (I726464,I3035,I726413,I726396,);
nor I_42555 (I726509,I217231,I217252);
and I_42556 (I726526,I726509,I217246);
nor I_42557 (I726543,I726526,I217231);
not I_42558 (I726560,I217231);
and I_42559 (I726577,I726560,I217228);
nand I_42560 (I726594,I726577,I217240);
nor I_42561 (I726611,I726560,I726594);
DFFARX1 I_42562 (I726611,I3035,I726413,I726378,);
not I_42563 (I726642,I726594);
nand I_42564 (I726659,I726464,I726642);
nand I_42565 (I726390,I726526,I726642);
DFFARX1 I_42566 (I726560,I3035,I726413,I726405,);
not I_42567 (I726704,I217255);
nor I_42568 (I726721,I726704,I217228);
nor I_42569 (I726738,I726721,I726543);
DFFARX1 I_42570 (I726738,I3035,I726413,I726402,);
not I_42571 (I726769,I726721);
DFFARX1 I_42572 (I726769,I3035,I726413,I726795,);
not I_42573 (I726803,I726795);
nor I_42574 (I726399,I726803,I726721);
nor I_42575 (I726834,I726704,I217237);
and I_42576 (I726851,I726834,I217234);
or I_42577 (I726868,I726851,I217228);
DFFARX1 I_42578 (I726868,I3035,I726413,I726894,);
not I_42579 (I726902,I726894);
nand I_42580 (I726919,I726902,I726642);
not I_42581 (I726393,I726919);
nand I_42582 (I726387,I726919,I726659);
nand I_42583 (I726384,I726902,I726526);
not I_42584 (I727008,I3042);
DFFARX1 I_42585 (I352773,I3035,I727008,I727034,);
DFFARX1 I_42586 (I352755,I3035,I727008,I727051,);
not I_42587 (I727059,I727051);
nor I_42588 (I726976,I727034,I727059);
DFFARX1 I_42589 (I727059,I3035,I727008,I726991,);
nor I_42590 (I727104,I352761,I352764);
and I_42591 (I727121,I727104,I352752);
nor I_42592 (I727138,I727121,I352761);
not I_42593 (I727155,I352761);
and I_42594 (I727172,I727155,I352770);
nand I_42595 (I727189,I727172,I352758);
nor I_42596 (I727206,I727155,I727189);
DFFARX1 I_42597 (I727206,I3035,I727008,I726973,);
not I_42598 (I727237,I727189);
nand I_42599 (I727254,I727059,I727237);
nand I_42600 (I726985,I727121,I727237);
DFFARX1 I_42601 (I727155,I3035,I727008,I727000,);
not I_42602 (I727299,I352755);
nor I_42603 (I727316,I727299,I352770);
nor I_42604 (I727333,I727316,I727138);
DFFARX1 I_42605 (I727333,I3035,I727008,I726997,);
not I_42606 (I727364,I727316);
DFFARX1 I_42607 (I727364,I3035,I727008,I727390,);
not I_42608 (I727398,I727390);
nor I_42609 (I726994,I727398,I727316);
nor I_42610 (I727429,I727299,I352767);
and I_42611 (I727446,I727429,I352776);
or I_42612 (I727463,I727446,I352752);
DFFARX1 I_42613 (I727463,I3035,I727008,I727489,);
not I_42614 (I727497,I727489);
nand I_42615 (I727514,I727497,I727237);
not I_42616 (I726988,I727514);
nand I_42617 (I726982,I727514,I727254);
nand I_42618 (I726979,I727497,I727121);
not I_42619 (I727603,I3042);
DFFARX1 I_42620 (I545198,I3035,I727603,I727629,);
DFFARX1 I_42621 (I545216,I3035,I727603,I727646,);
not I_42622 (I727654,I727646);
nor I_42623 (I727571,I727629,I727654);
DFFARX1 I_42624 (I727654,I3035,I727603,I727586,);
nor I_42625 (I727699,I545195,I545207);
and I_42626 (I727716,I727699,I545192);
nor I_42627 (I727733,I727716,I545195);
not I_42628 (I727750,I545195);
and I_42629 (I727767,I727750,I545201);
nand I_42630 (I727784,I727767,I545213);
nor I_42631 (I727801,I727750,I727784);
DFFARX1 I_42632 (I727801,I3035,I727603,I727568,);
not I_42633 (I727832,I727784);
nand I_42634 (I727849,I727654,I727832);
nand I_42635 (I727580,I727716,I727832);
DFFARX1 I_42636 (I727750,I3035,I727603,I727595,);
not I_42637 (I727894,I545204);
nor I_42638 (I727911,I727894,I545201);
nor I_42639 (I727928,I727911,I727733);
DFFARX1 I_42640 (I727928,I3035,I727603,I727592,);
not I_42641 (I727959,I727911);
DFFARX1 I_42642 (I727959,I3035,I727603,I727985,);
not I_42643 (I727993,I727985);
nor I_42644 (I727589,I727993,I727911);
nor I_42645 (I728024,I727894,I545192);
and I_42646 (I728041,I728024,I545219);
or I_42647 (I728058,I728041,I545210);
DFFARX1 I_42648 (I728058,I3035,I727603,I728084,);
not I_42649 (I728092,I728084);
nand I_42650 (I728109,I728092,I727832);
not I_42651 (I727583,I728109);
nand I_42652 (I727577,I728109,I727849);
nand I_42653 (I727574,I728092,I727716);
not I_42654 (I728198,I3042);
DFFARX1 I_42655 (I100914,I3035,I728198,I728224,);
DFFARX1 I_42656 (I100917,I3035,I728198,I728241,);
not I_42657 (I728249,I728241);
nor I_42658 (I728166,I728224,I728249);
DFFARX1 I_42659 (I728249,I3035,I728198,I728181,);
nor I_42660 (I728294,I100923,I100917);
and I_42661 (I728311,I728294,I100920);
nor I_42662 (I728328,I728311,I100923);
not I_42663 (I728345,I100923);
and I_42664 (I728362,I728345,I100914);
nand I_42665 (I728379,I728362,I100932);
nor I_42666 (I728396,I728345,I728379);
DFFARX1 I_42667 (I728396,I3035,I728198,I728163,);
not I_42668 (I728427,I728379);
nand I_42669 (I728444,I728249,I728427);
nand I_42670 (I728175,I728311,I728427);
DFFARX1 I_42671 (I728345,I3035,I728198,I728190,);
not I_42672 (I728489,I100926);
nor I_42673 (I728506,I728489,I100914);
nor I_42674 (I728523,I728506,I728328);
DFFARX1 I_42675 (I728523,I3035,I728198,I728187,);
not I_42676 (I728554,I728506);
DFFARX1 I_42677 (I728554,I3035,I728198,I728580,);
not I_42678 (I728588,I728580);
nor I_42679 (I728184,I728588,I728506);
nor I_42680 (I728619,I728489,I100929);
and I_42681 (I728636,I728619,I100935);
or I_42682 (I728653,I728636,I100938);
DFFARX1 I_42683 (I728653,I3035,I728198,I728679,);
not I_42684 (I728687,I728679);
nand I_42685 (I728704,I728687,I728427);
not I_42686 (I728178,I728704);
nand I_42687 (I728172,I728704,I728444);
nand I_42688 (I728169,I728687,I728311);
not I_42689 (I728793,I3042);
DFFARX1 I_42690 (I527110,I3035,I728793,I728819,);
DFFARX1 I_42691 (I527128,I3035,I728793,I728836,);
not I_42692 (I728844,I728836);
nor I_42693 (I728761,I728819,I728844);
DFFARX1 I_42694 (I728844,I3035,I728793,I728776,);
nor I_42695 (I728889,I527107,I527119);
and I_42696 (I728906,I728889,I527104);
nor I_42697 (I728923,I728906,I527107);
not I_42698 (I728940,I527107);
and I_42699 (I728957,I728940,I527113);
nand I_42700 (I728974,I728957,I527125);
nor I_42701 (I728991,I728940,I728974);
DFFARX1 I_42702 (I728991,I3035,I728793,I728758,);
not I_42703 (I729022,I728974);
nand I_42704 (I729039,I728844,I729022);
nand I_42705 (I728770,I728906,I729022);
DFFARX1 I_42706 (I728940,I3035,I728793,I728785,);
not I_42707 (I729084,I527116);
nor I_42708 (I729101,I729084,I527113);
nor I_42709 (I729118,I729101,I728923);
DFFARX1 I_42710 (I729118,I3035,I728793,I728782,);
not I_42711 (I729149,I729101);
DFFARX1 I_42712 (I729149,I3035,I728793,I729175,);
not I_42713 (I729183,I729175);
nor I_42714 (I728779,I729183,I729101);
nor I_42715 (I729214,I729084,I527104);
and I_42716 (I729231,I729214,I527131);
or I_42717 (I729248,I729231,I527122);
DFFARX1 I_42718 (I729248,I3035,I728793,I729274,);
not I_42719 (I729282,I729274);
nand I_42720 (I729299,I729282,I729022);
not I_42721 (I728773,I729299);
nand I_42722 (I728767,I729299,I729039);
nand I_42723 (I728764,I729282,I728906);
not I_42724 (I729388,I3042);
DFFARX1 I_42725 (I553228,I3035,I729388,I729414,);
DFFARX1 I_42726 (I553219,I3035,I729388,I729431,);
not I_42727 (I729439,I729431);
nor I_42728 (I729356,I729414,I729439);
DFFARX1 I_42729 (I729439,I3035,I729388,I729371,);
nor I_42730 (I729484,I553225,I553234);
and I_42731 (I729501,I729484,I553237);
nor I_42732 (I729518,I729501,I553225);
not I_42733 (I729535,I553225);
and I_42734 (I729552,I729535,I553216);
nand I_42735 (I729569,I729552,I553222);
nor I_42736 (I729586,I729535,I729569);
DFFARX1 I_42737 (I729586,I3035,I729388,I729353,);
not I_42738 (I729617,I729569);
nand I_42739 (I729634,I729439,I729617);
nand I_42740 (I729365,I729501,I729617);
DFFARX1 I_42741 (I729535,I3035,I729388,I729380,);
not I_42742 (I729679,I553231);
nor I_42743 (I729696,I729679,I553216);
nor I_42744 (I729713,I729696,I729518);
DFFARX1 I_42745 (I729713,I3035,I729388,I729377,);
not I_42746 (I729744,I729696);
DFFARX1 I_42747 (I729744,I3035,I729388,I729770,);
not I_42748 (I729778,I729770);
nor I_42749 (I729374,I729778,I729696);
nor I_42750 (I729809,I729679,I553216);
and I_42751 (I729826,I729809,I553219);
or I_42752 (I729843,I729826,I553222);
DFFARX1 I_42753 (I729843,I3035,I729388,I729869,);
not I_42754 (I729877,I729869);
nand I_42755 (I729894,I729877,I729617);
not I_42756 (I729368,I729894);
nand I_42757 (I729362,I729894,I729634);
nand I_42758 (I729359,I729877,I729501);
not I_42759 (I729983,I3042);
DFFARX1 I_42760 (I23106,I3035,I729983,I730009,);
DFFARX1 I_42761 (I23088,I3035,I729983,I730026,);
not I_42762 (I730034,I730026);
nor I_42763 (I729951,I730009,I730034);
DFFARX1 I_42764 (I730034,I3035,I729983,I729966,);
nor I_42765 (I730079,I23088,I23103);
and I_42766 (I730096,I730079,I23097);
nor I_42767 (I730113,I730096,I23088);
not I_42768 (I730130,I23088);
and I_42769 (I730147,I730130,I23091);
nand I_42770 (I730164,I730147,I23094);
nor I_42771 (I730181,I730130,I730164);
DFFARX1 I_42772 (I730181,I3035,I729983,I729948,);
not I_42773 (I730212,I730164);
nand I_42774 (I730229,I730034,I730212);
nand I_42775 (I729960,I730096,I730212);
DFFARX1 I_42776 (I730130,I3035,I729983,I729975,);
not I_42777 (I730274,I23100);
nor I_42778 (I730291,I730274,I23091);
nor I_42779 (I730308,I730291,I730113);
DFFARX1 I_42780 (I730308,I3035,I729983,I729972,);
not I_42781 (I730339,I730291);
DFFARX1 I_42782 (I730339,I3035,I729983,I730365,);
not I_42783 (I730373,I730365);
nor I_42784 (I729969,I730373,I730291);
nor I_42785 (I730404,I730274,I23112);
and I_42786 (I730421,I730404,I23109);
or I_42787 (I730438,I730421,I23091);
DFFARX1 I_42788 (I730438,I3035,I729983,I730464,);
not I_42789 (I730472,I730464);
nand I_42790 (I730489,I730472,I730212);
not I_42791 (I729963,I730489);
nand I_42792 (I729957,I730489,I730229);
nand I_42793 (I729954,I730472,I730096);
not I_42794 (I730578,I3042);
DFFARX1 I_42795 (I454064,I3035,I730578,I730604,);
DFFARX1 I_42796 (I454061,I3035,I730578,I730621,);
not I_42797 (I730629,I730621);
nor I_42798 (I730546,I730604,I730629);
DFFARX1 I_42799 (I730629,I3035,I730578,I730561,);
nor I_42800 (I730674,I454076,I454058);
and I_42801 (I730691,I730674,I454055);
nor I_42802 (I730708,I730691,I454076);
not I_42803 (I730725,I454076);
and I_42804 (I730742,I730725,I454061);
nand I_42805 (I730759,I730742,I454073);
nor I_42806 (I730776,I730725,I730759);
DFFARX1 I_42807 (I730776,I3035,I730578,I730543,);
not I_42808 (I730807,I730759);
nand I_42809 (I730824,I730629,I730807);
nand I_42810 (I730555,I730691,I730807);
DFFARX1 I_42811 (I730725,I3035,I730578,I730570,);
not I_42812 (I730869,I454067);
nor I_42813 (I730886,I730869,I454061);
nor I_42814 (I730903,I730886,I730708);
DFFARX1 I_42815 (I730903,I3035,I730578,I730567,);
not I_42816 (I730934,I730886);
DFFARX1 I_42817 (I730934,I3035,I730578,I730960,);
not I_42818 (I730968,I730960);
nor I_42819 (I730564,I730968,I730886);
nor I_42820 (I730999,I730869,I454055);
and I_42821 (I731016,I730999,I454070);
or I_42822 (I731033,I731016,I454058);
DFFARX1 I_42823 (I731033,I3035,I730578,I731059,);
not I_42824 (I731067,I731059);
nand I_42825 (I731084,I731067,I730807);
not I_42826 (I730558,I731084);
nand I_42827 (I730552,I731084,I730824);
nand I_42828 (I730549,I731067,I730691);
not I_42829 (I731173,I3042);
DFFARX1 I_42830 (I235333,I3035,I731173,I731199,);
DFFARX1 I_42831 (I235339,I3035,I731173,I731216,);
not I_42832 (I731224,I731216);
nor I_42833 (I731141,I731199,I731224);
DFFARX1 I_42834 (I731224,I3035,I731173,I731156,);
nor I_42835 (I731269,I235348,I235333);
and I_42836 (I731286,I731269,I235360);
nor I_42837 (I731303,I731286,I235348);
not I_42838 (I731320,I235348);
and I_42839 (I731337,I731320,I235336);
nand I_42840 (I731354,I731337,I235357);
nor I_42841 (I731371,I731320,I731354);
DFFARX1 I_42842 (I731371,I3035,I731173,I731138,);
not I_42843 (I731402,I731354);
nand I_42844 (I731419,I731224,I731402);
nand I_42845 (I731150,I731286,I731402);
DFFARX1 I_42846 (I731320,I3035,I731173,I731165,);
not I_42847 (I731464,I235345);
nor I_42848 (I731481,I731464,I235336);
nor I_42849 (I731498,I731481,I731303);
DFFARX1 I_42850 (I731498,I3035,I731173,I731162,);
not I_42851 (I731529,I731481);
DFFARX1 I_42852 (I731529,I3035,I731173,I731555,);
not I_42853 (I731563,I731555);
nor I_42854 (I731159,I731563,I731481);
nor I_42855 (I731594,I731464,I235342);
and I_42856 (I731611,I731594,I235354);
or I_42857 (I731628,I731611,I235351);
DFFARX1 I_42858 (I731628,I3035,I731173,I731654,);
not I_42859 (I731662,I731654);
nand I_42860 (I731679,I731662,I731402);
not I_42861 (I731153,I731679);
nand I_42862 (I731147,I731679,I731419);
nand I_42863 (I731144,I731662,I731286);
not I_42864 (I731768,I3042);
DFFARX1 I_42865 (I288866,I3035,I731768,I731794,);
DFFARX1 I_42866 (I288869,I3035,I731768,I731811,);
not I_42867 (I731819,I731811);
nor I_42868 (I731736,I731794,I731819);
DFFARX1 I_42869 (I731819,I3035,I731768,I731751,);
nor I_42870 (I731864,I288872,I288890);
and I_42871 (I731881,I731864,I288875);
nor I_42872 (I731898,I731881,I288872);
not I_42873 (I731915,I288872);
and I_42874 (I731932,I731915,I288884);
nand I_42875 (I731949,I731932,I288887);
nor I_42876 (I731966,I731915,I731949);
DFFARX1 I_42877 (I731966,I3035,I731768,I731733,);
not I_42878 (I731997,I731949);
nand I_42879 (I732014,I731819,I731997);
nand I_42880 (I731745,I731881,I731997);
DFFARX1 I_42881 (I731915,I3035,I731768,I731760,);
not I_42882 (I732059,I288878);
nor I_42883 (I732076,I732059,I288884);
nor I_42884 (I732093,I732076,I731898);
DFFARX1 I_42885 (I732093,I3035,I731768,I731757,);
not I_42886 (I732124,I732076);
DFFARX1 I_42887 (I732124,I3035,I731768,I732150,);
not I_42888 (I732158,I732150);
nor I_42889 (I731754,I732158,I732076);
nor I_42890 (I732189,I732059,I288866);
and I_42891 (I732206,I732189,I288881);
or I_42892 (I732223,I732206,I288869);
DFFARX1 I_42893 (I732223,I3035,I731768,I732249,);
not I_42894 (I732257,I732249);
nand I_42895 (I732274,I732257,I731997);
not I_42896 (I731748,I732274);
nand I_42897 (I731742,I732274,I732014);
nand I_42898 (I731739,I732257,I731881);
not I_42899 (I732363,I3042);
DFFARX1 I_42900 (I220938,I3035,I732363,I732389,);
DFFARX1 I_42901 (I220932,I3035,I732363,I732406,);
not I_42902 (I732414,I732406);
nor I_42903 (I732331,I732389,I732414);
DFFARX1 I_42904 (I732414,I3035,I732363,I732346,);
nor I_42905 (I732459,I220920,I220941);
and I_42906 (I732476,I732459,I220935);
nor I_42907 (I732493,I732476,I220920);
not I_42908 (I732510,I220920);
and I_42909 (I732527,I732510,I220917);
nand I_42910 (I732544,I732527,I220929);
nor I_42911 (I732561,I732510,I732544);
DFFARX1 I_42912 (I732561,I3035,I732363,I732328,);
not I_42913 (I732592,I732544);
nand I_42914 (I732609,I732414,I732592);
nand I_42915 (I732340,I732476,I732592);
DFFARX1 I_42916 (I732510,I3035,I732363,I732355,);
not I_42917 (I732654,I220944);
nor I_42918 (I732671,I732654,I220917);
nor I_42919 (I732688,I732671,I732493);
DFFARX1 I_42920 (I732688,I3035,I732363,I732352,);
not I_42921 (I732719,I732671);
DFFARX1 I_42922 (I732719,I3035,I732363,I732745,);
not I_42923 (I732753,I732745);
nor I_42924 (I732349,I732753,I732671);
nor I_42925 (I732784,I732654,I220926);
and I_42926 (I732801,I732784,I220923);
or I_42927 (I732818,I732801,I220917);
DFFARX1 I_42928 (I732818,I3035,I732363,I732844,);
not I_42929 (I732852,I732844);
nand I_42930 (I732869,I732852,I732592);
not I_42931 (I732343,I732869);
nand I_42932 (I732337,I732869,I732609);
nand I_42933 (I732334,I732852,I732476);
not I_42934 (I732958,I3042);
DFFARX1 I_42935 (I558277,I3035,I732958,I732984,);
DFFARX1 I_42936 (I558268,I3035,I732958,I733001,);
not I_42937 (I733009,I733001);
nor I_42938 (I732926,I732984,I733009);
DFFARX1 I_42939 (I733009,I3035,I732958,I732941,);
nor I_42940 (I733054,I558274,I558283);
and I_42941 (I733071,I733054,I558286);
nor I_42942 (I733088,I733071,I558274);
not I_42943 (I733105,I558274);
and I_42944 (I733122,I733105,I558265);
nand I_42945 (I733139,I733122,I558271);
nor I_42946 (I733156,I733105,I733139);
DFFARX1 I_42947 (I733156,I3035,I732958,I732923,);
not I_42948 (I733187,I733139);
nand I_42949 (I733204,I733009,I733187);
nand I_42950 (I732935,I733071,I733187);
DFFARX1 I_42951 (I733105,I3035,I732958,I732950,);
not I_42952 (I733249,I558280);
nor I_42953 (I733266,I733249,I558265);
nor I_42954 (I733283,I733266,I733088);
DFFARX1 I_42955 (I733283,I3035,I732958,I732947,);
not I_42956 (I733314,I733266);
DFFARX1 I_42957 (I733314,I3035,I732958,I733340,);
not I_42958 (I733348,I733340);
nor I_42959 (I732944,I733348,I733266);
nor I_42960 (I733379,I733249,I558265);
and I_42961 (I733396,I733379,I558268);
or I_42962 (I733413,I733396,I558271);
DFFARX1 I_42963 (I733413,I3035,I732958,I733439,);
not I_42964 (I733447,I733439);
nand I_42965 (I733464,I733447,I733187);
not I_42966 (I732938,I733464);
nand I_42967 (I732932,I733464,I733204);
nand I_42968 (I732929,I733447,I733071);
not I_42969 (I733553,I3042);
DFFARX1 I_42970 (I549301,I3035,I733553,I733579,);
DFFARX1 I_42971 (I549292,I3035,I733553,I733596,);
not I_42972 (I733604,I733596);
nor I_42973 (I733521,I733579,I733604);
DFFARX1 I_42974 (I733604,I3035,I733553,I733536,);
nor I_42975 (I733649,I549298,I549307);
and I_42976 (I733666,I733649,I549310);
nor I_42977 (I733683,I733666,I549298);
not I_42978 (I733700,I549298);
and I_42979 (I733717,I733700,I549289);
nand I_42980 (I733734,I733717,I549295);
nor I_42981 (I733751,I733700,I733734);
DFFARX1 I_42982 (I733751,I3035,I733553,I733518,);
not I_42983 (I733782,I733734);
nand I_42984 (I733799,I733604,I733782);
nand I_42985 (I733530,I733666,I733782);
DFFARX1 I_42986 (I733700,I3035,I733553,I733545,);
not I_42987 (I733844,I549304);
nor I_42988 (I733861,I733844,I549289);
nor I_42989 (I733878,I733861,I733683);
DFFARX1 I_42990 (I733878,I3035,I733553,I733542,);
not I_42991 (I733909,I733861);
DFFARX1 I_42992 (I733909,I3035,I733553,I733935,);
not I_42993 (I733943,I733935);
nor I_42994 (I733539,I733943,I733861);
nor I_42995 (I733974,I733844,I549289);
and I_42996 (I733991,I733974,I549292);
or I_42997 (I734008,I733991,I549295);
DFFARX1 I_42998 (I734008,I3035,I733553,I734034,);
not I_42999 (I734042,I734034);
nand I_43000 (I734059,I734042,I733782);
not I_43001 (I733533,I734059);
nand I_43002 (I733527,I734059,I733799);
nand I_43003 (I733524,I734042,I733666);
not I_43004 (I734148,I3042);
DFFARX1 I_43005 (I1668,I3035,I734148,I734174,);
DFFARX1 I_43006 (I2604,I3035,I734148,I734191,);
not I_43007 (I734199,I734191);
nor I_43008 (I734116,I734174,I734199);
DFFARX1 I_43009 (I734199,I3035,I734148,I734131,);
nor I_43010 (I734244,I2868,I2652);
and I_43011 (I734261,I734244,I1764);
nor I_43012 (I734278,I734261,I2868);
not I_43013 (I734295,I2868);
and I_43014 (I734312,I734295,I2332);
nand I_43015 (I734329,I734312,I2164);
nor I_43016 (I734346,I734295,I734329);
DFFARX1 I_43017 (I734346,I3035,I734148,I734113,);
not I_43018 (I734377,I734329);
nand I_43019 (I734394,I734199,I734377);
nand I_43020 (I734125,I734261,I734377);
DFFARX1 I_43021 (I734295,I3035,I734148,I734140,);
not I_43022 (I734439,I2724);
nor I_43023 (I734456,I734439,I2332);
nor I_43024 (I734473,I734456,I734278);
DFFARX1 I_43025 (I734473,I3035,I734148,I734137,);
not I_43026 (I734504,I734456);
DFFARX1 I_43027 (I734504,I3035,I734148,I734530,);
not I_43028 (I734538,I734530);
nor I_43029 (I734134,I734538,I734456);
nor I_43030 (I734569,I734439,I1884);
and I_43031 (I734586,I734569,I2548);
or I_43032 (I734603,I734586,I1652);
DFFARX1 I_43033 (I734603,I3035,I734148,I734629,);
not I_43034 (I734637,I734629);
nand I_43035 (I734654,I734637,I734377);
not I_43036 (I734128,I734654);
nand I_43037 (I734122,I734654,I734394);
nand I_43038 (I734119,I734637,I734261);
not I_43039 (I734743,I3042);
DFFARX1 I_43040 (I604661,I3035,I734743,I734769,);
DFFARX1 I_43041 (I604673,I3035,I734743,I734786,);
not I_43042 (I734794,I734786);
nor I_43043 (I734711,I734769,I734794);
DFFARX1 I_43044 (I734794,I3035,I734743,I734726,);
nor I_43045 (I734839,I604670,I604664);
and I_43046 (I734856,I734839,I604658);
nor I_43047 (I734873,I734856,I604670);
not I_43048 (I734890,I604670);
and I_43049 (I734907,I734890,I604667);
nand I_43050 (I734924,I734907,I604658);
nor I_43051 (I734941,I734890,I734924);
DFFARX1 I_43052 (I734941,I3035,I734743,I734708,);
not I_43053 (I734972,I734924);
nand I_43054 (I734989,I734794,I734972);
nand I_43055 (I734720,I734856,I734972);
DFFARX1 I_43056 (I734890,I3035,I734743,I734735,);
not I_43057 (I735034,I604682);
nor I_43058 (I735051,I735034,I604667);
nor I_43059 (I735068,I735051,I734873);
DFFARX1 I_43060 (I735068,I3035,I734743,I734732,);
not I_43061 (I735099,I735051);
DFFARX1 I_43062 (I735099,I3035,I734743,I735125,);
not I_43063 (I735133,I735125);
nor I_43064 (I734729,I735133,I735051);
nor I_43065 (I735164,I735034,I604676);
and I_43066 (I735181,I735164,I604679);
or I_43067 (I735198,I735181,I604661);
DFFARX1 I_43068 (I735198,I3035,I734743,I735224,);
not I_43069 (I735232,I735224);
nand I_43070 (I735249,I735232,I734972);
not I_43071 (I734723,I735249);
nand I_43072 (I734717,I735249,I734989);
nand I_43073 (I734714,I735232,I734856);
not I_43074 (I735338,I3042);
DFFARX1 I_43075 (I379361,I3035,I735338,I735364,);
DFFARX1 I_43076 (I379343,I3035,I735338,I735381,);
not I_43077 (I735389,I735381);
nor I_43078 (I735306,I735364,I735389);
DFFARX1 I_43079 (I735389,I3035,I735338,I735321,);
nor I_43080 (I735434,I379349,I379352);
and I_43081 (I735451,I735434,I379340);
nor I_43082 (I735468,I735451,I379349);
not I_43083 (I735485,I379349);
and I_43084 (I735502,I735485,I379358);
nand I_43085 (I735519,I735502,I379346);
nor I_43086 (I735536,I735485,I735519);
DFFARX1 I_43087 (I735536,I3035,I735338,I735303,);
not I_43088 (I735567,I735519);
nand I_43089 (I735584,I735389,I735567);
nand I_43090 (I735315,I735451,I735567);
DFFARX1 I_43091 (I735485,I3035,I735338,I735330,);
not I_43092 (I735629,I379343);
nor I_43093 (I735646,I735629,I379358);
nor I_43094 (I735663,I735646,I735468);
DFFARX1 I_43095 (I735663,I3035,I735338,I735327,);
not I_43096 (I735694,I735646);
DFFARX1 I_43097 (I735694,I3035,I735338,I735720,);
not I_43098 (I735728,I735720);
nor I_43099 (I735324,I735728,I735646);
nor I_43100 (I735759,I735629,I379355);
and I_43101 (I735776,I735759,I379364);
or I_43102 (I735793,I735776,I379340);
DFFARX1 I_43103 (I735793,I3035,I735338,I735819,);
not I_43104 (I735827,I735819);
nand I_43105 (I735844,I735827,I735567);
not I_43106 (I735318,I735844);
nand I_43107 (I735312,I735844,I735584);
nand I_43108 (I735309,I735827,I735451);
not I_43109 (I735933,I3042);
DFFARX1 I_43110 (I620267,I3035,I735933,I735959,);
DFFARX1 I_43111 (I620279,I3035,I735933,I735976,);
not I_43112 (I735984,I735976);
nor I_43113 (I735901,I735959,I735984);
DFFARX1 I_43114 (I735984,I3035,I735933,I735916,);
nor I_43115 (I736029,I620276,I620270);
and I_43116 (I736046,I736029,I620264);
nor I_43117 (I736063,I736046,I620276);
not I_43118 (I736080,I620276);
and I_43119 (I736097,I736080,I620273);
nand I_43120 (I736114,I736097,I620264);
nor I_43121 (I736131,I736080,I736114);
DFFARX1 I_43122 (I736131,I3035,I735933,I735898,);
not I_43123 (I736162,I736114);
nand I_43124 (I736179,I735984,I736162);
nand I_43125 (I735910,I736046,I736162);
DFFARX1 I_43126 (I736080,I3035,I735933,I735925,);
not I_43127 (I736224,I620288);
nor I_43128 (I736241,I736224,I620273);
nor I_43129 (I736258,I736241,I736063);
DFFARX1 I_43130 (I736258,I3035,I735933,I735922,);
not I_43131 (I736289,I736241);
DFFARX1 I_43132 (I736289,I3035,I735933,I736315,);
not I_43133 (I736323,I736315);
nor I_43134 (I735919,I736323,I736241);
nor I_43135 (I736354,I736224,I620282);
and I_43136 (I736371,I736354,I620285);
or I_43137 (I736388,I736371,I620267);
DFFARX1 I_43138 (I736388,I3035,I735933,I736414,);
not I_43139 (I736422,I736414);
nand I_43140 (I736439,I736422,I736162);
not I_43141 (I735913,I736439);
nand I_43142 (I735907,I736439,I736179);
nand I_43143 (I735904,I736422,I736046);
not I_43144 (I736528,I3042);
DFFARX1 I_43145 (I179832,I3035,I736528,I736554,);
DFFARX1 I_43146 (I179826,I3035,I736528,I736571,);
not I_43147 (I736579,I736571);
nor I_43148 (I736496,I736554,I736579);
DFFARX1 I_43149 (I736579,I3035,I736528,I736511,);
nor I_43150 (I736624,I179814,I179835);
and I_43151 (I736641,I736624,I179829);
nor I_43152 (I736658,I736641,I179814);
not I_43153 (I736675,I179814);
and I_43154 (I736692,I736675,I179811);
nand I_43155 (I736709,I736692,I179823);
nor I_43156 (I736726,I736675,I736709);
DFFARX1 I_43157 (I736726,I3035,I736528,I736493,);
not I_43158 (I736757,I736709);
nand I_43159 (I736774,I736579,I736757);
nand I_43160 (I736505,I736641,I736757);
DFFARX1 I_43161 (I736675,I3035,I736528,I736520,);
not I_43162 (I736819,I179838);
nor I_43163 (I736836,I736819,I179811);
nor I_43164 (I736853,I736836,I736658);
DFFARX1 I_43165 (I736853,I3035,I736528,I736517,);
not I_43166 (I736884,I736836);
DFFARX1 I_43167 (I736884,I3035,I736528,I736910,);
not I_43168 (I736918,I736910);
nor I_43169 (I736514,I736918,I736836);
nor I_43170 (I736949,I736819,I179820);
and I_43171 (I736966,I736949,I179817);
or I_43172 (I736983,I736966,I179811);
DFFARX1 I_43173 (I736983,I3035,I736528,I737009,);
not I_43174 (I737017,I737009);
nand I_43175 (I737034,I737017,I736757);
not I_43176 (I736508,I737034);
nand I_43177 (I736502,I737034,I736774);
nand I_43178 (I736499,I737017,I736641);
not I_43179 (I737123,I3042);
DFFARX1 I_43180 (I86039,I3035,I737123,I737149,);
DFFARX1 I_43181 (I86042,I3035,I737123,I737166,);
not I_43182 (I737174,I737166);
nor I_43183 (I737091,I737149,I737174);
DFFARX1 I_43184 (I737174,I3035,I737123,I737106,);
nor I_43185 (I737219,I86048,I86042);
and I_43186 (I737236,I737219,I86045);
nor I_43187 (I737253,I737236,I86048);
not I_43188 (I737270,I86048);
and I_43189 (I737287,I737270,I86039);
nand I_43190 (I737304,I737287,I86057);
nor I_43191 (I737321,I737270,I737304);
DFFARX1 I_43192 (I737321,I3035,I737123,I737088,);
not I_43193 (I737352,I737304);
nand I_43194 (I737369,I737174,I737352);
nand I_43195 (I737100,I737236,I737352);
DFFARX1 I_43196 (I737270,I3035,I737123,I737115,);
not I_43197 (I737414,I86051);
nor I_43198 (I737431,I737414,I86039);
nor I_43199 (I737448,I737431,I737253);
DFFARX1 I_43200 (I737448,I3035,I737123,I737112,);
not I_43201 (I737479,I737431);
DFFARX1 I_43202 (I737479,I3035,I737123,I737505,);
not I_43203 (I737513,I737505);
nor I_43204 (I737109,I737513,I737431);
nor I_43205 (I737544,I737414,I86054);
and I_43206 (I737561,I737544,I86060);
or I_43207 (I737578,I737561,I86063);
DFFARX1 I_43208 (I737578,I3035,I737123,I737604,);
not I_43209 (I737612,I737604);
nand I_43210 (I737629,I737612,I737352);
not I_43211 (I737103,I737629);
nand I_43212 (I737097,I737629,I737369);
nand I_43213 (I737094,I737612,I737236);
not I_43214 (I737718,I3042);
DFFARX1 I_43215 (I129474,I3035,I737718,I737744,);
DFFARX1 I_43216 (I129477,I3035,I737718,I737761,);
not I_43217 (I737769,I737761);
nor I_43218 (I737686,I737744,I737769);
DFFARX1 I_43219 (I737769,I3035,I737718,I737701,);
nor I_43220 (I737814,I129483,I129477);
and I_43221 (I737831,I737814,I129480);
nor I_43222 (I737848,I737831,I129483);
not I_43223 (I737865,I129483);
and I_43224 (I737882,I737865,I129474);
nand I_43225 (I737899,I737882,I129492);
nor I_43226 (I737916,I737865,I737899);
DFFARX1 I_43227 (I737916,I3035,I737718,I737683,);
not I_43228 (I737947,I737899);
nand I_43229 (I737964,I737769,I737947);
nand I_43230 (I737695,I737831,I737947);
DFFARX1 I_43231 (I737865,I3035,I737718,I737710,);
not I_43232 (I738009,I129486);
nor I_43233 (I738026,I738009,I129474);
nor I_43234 (I738043,I738026,I737848);
DFFARX1 I_43235 (I738043,I3035,I737718,I737707,);
not I_43236 (I738074,I738026);
DFFARX1 I_43237 (I738074,I3035,I737718,I738100,);
not I_43238 (I738108,I738100);
nor I_43239 (I737704,I738108,I738026);
nor I_43240 (I738139,I738009,I129489);
and I_43241 (I738156,I738139,I129495);
or I_43242 (I738173,I738156,I129498);
DFFARX1 I_43243 (I738173,I3035,I737718,I738199,);
not I_43244 (I738207,I738199);
nand I_43245 (I738224,I738207,I737947);
not I_43246 (I737698,I738224);
nand I_43247 (I737692,I738224,I737964);
nand I_43248 (I737689,I738207,I737831);
not I_43249 (I738313,I3042);
DFFARX1 I_43250 (I70539,I3035,I738313,I738339,);
DFFARX1 I_43251 (I70527,I3035,I738313,I738356,);
not I_43252 (I738364,I738356);
nor I_43253 (I738281,I738339,I738364);
DFFARX1 I_43254 (I738364,I3035,I738313,I738296,);
nor I_43255 (I738409,I70518,I70542);
and I_43256 (I738426,I738409,I70521);
nor I_43257 (I738443,I738426,I70518);
not I_43258 (I738460,I70518);
and I_43259 (I738477,I738460,I70524);
nand I_43260 (I738494,I738477,I70536);
nor I_43261 (I738511,I738460,I738494);
DFFARX1 I_43262 (I738511,I3035,I738313,I738278,);
not I_43263 (I738542,I738494);
nand I_43264 (I738559,I738364,I738542);
nand I_43265 (I738290,I738426,I738542);
DFFARX1 I_43266 (I738460,I3035,I738313,I738305,);
not I_43267 (I738604,I70518);
nor I_43268 (I738621,I738604,I70524);
nor I_43269 (I738638,I738621,I738443);
DFFARX1 I_43270 (I738638,I3035,I738313,I738302,);
not I_43271 (I738669,I738621);
DFFARX1 I_43272 (I738669,I3035,I738313,I738695,);
not I_43273 (I738703,I738695);
nor I_43274 (I738299,I738703,I738621);
nor I_43275 (I738734,I738604,I70521);
and I_43276 (I738751,I738734,I70530);
or I_43277 (I738768,I738751,I70533);
DFFARX1 I_43278 (I738768,I3035,I738313,I738794,);
not I_43279 (I738802,I738794);
nand I_43280 (I738819,I738802,I738542);
not I_43281 (I738293,I738819);
nand I_43282 (I738287,I738819,I738559);
nand I_43283 (I738284,I738802,I738426);
not I_43284 (I738908,I3042);
DFFARX1 I_43285 (I580963,I3035,I738908,I738934,);
DFFARX1 I_43286 (I580975,I3035,I738908,I738951,);
not I_43287 (I738959,I738951);
nor I_43288 (I738876,I738934,I738959);
DFFARX1 I_43289 (I738959,I3035,I738908,I738891,);
nor I_43290 (I739004,I580972,I580966);
and I_43291 (I739021,I739004,I580960);
nor I_43292 (I739038,I739021,I580972);
not I_43293 (I739055,I580972);
and I_43294 (I739072,I739055,I580969);
nand I_43295 (I739089,I739072,I580960);
nor I_43296 (I739106,I739055,I739089);
DFFARX1 I_43297 (I739106,I3035,I738908,I738873,);
not I_43298 (I739137,I739089);
nand I_43299 (I739154,I738959,I739137);
nand I_43300 (I738885,I739021,I739137);
DFFARX1 I_43301 (I739055,I3035,I738908,I738900,);
not I_43302 (I739199,I580984);
nor I_43303 (I739216,I739199,I580969);
nor I_43304 (I739233,I739216,I739038);
DFFARX1 I_43305 (I739233,I3035,I738908,I738897,);
not I_43306 (I739264,I739216);
DFFARX1 I_43307 (I739264,I3035,I738908,I739290,);
not I_43308 (I739298,I739290);
nor I_43309 (I738894,I739298,I739216);
nor I_43310 (I739329,I739199,I580978);
and I_43311 (I739346,I739329,I580981);
or I_43312 (I739363,I739346,I580963);
DFFARX1 I_43313 (I739363,I3035,I738908,I739389,);
not I_43314 (I739397,I739389);
nand I_43315 (I739414,I739397,I739137);
not I_43316 (I738888,I739414);
nand I_43317 (I738882,I739414,I739154);
nand I_43318 (I738879,I739397,I739021);
not I_43319 (I739503,I3042);
DFFARX1 I_43320 (I289461,I3035,I739503,I739529,);
DFFARX1 I_43321 (I289464,I3035,I739503,I739546,);
not I_43322 (I739554,I739546);
nor I_43323 (I739471,I739529,I739554);
DFFARX1 I_43324 (I739554,I3035,I739503,I739486,);
nor I_43325 (I739599,I289467,I289485);
and I_43326 (I739616,I739599,I289470);
nor I_43327 (I739633,I739616,I289467);
not I_43328 (I739650,I289467);
and I_43329 (I739667,I739650,I289479);
nand I_43330 (I739684,I739667,I289482);
nor I_43331 (I739701,I739650,I739684);
DFFARX1 I_43332 (I739701,I3035,I739503,I739468,);
not I_43333 (I739732,I739684);
nand I_43334 (I739749,I739554,I739732);
nand I_43335 (I739480,I739616,I739732);
DFFARX1 I_43336 (I739650,I3035,I739503,I739495,);
not I_43337 (I739794,I289473);
nor I_43338 (I739811,I739794,I289479);
nor I_43339 (I739828,I739811,I739633);
DFFARX1 I_43340 (I739828,I3035,I739503,I739492,);
not I_43341 (I739859,I739811);
DFFARX1 I_43342 (I739859,I3035,I739503,I739885,);
not I_43343 (I739893,I739885);
nor I_43344 (I739489,I739893,I739811);
nor I_43345 (I739924,I739794,I289461);
and I_43346 (I739941,I739924,I289476);
or I_43347 (I739958,I739941,I289464);
DFFARX1 I_43348 (I739958,I3035,I739503,I739984,);
not I_43349 (I739992,I739984);
nand I_43350 (I740009,I739992,I739732);
not I_43351 (I739483,I740009);
nand I_43352 (I739477,I740009,I739749);
nand I_43353 (I739474,I739992,I739616);
not I_43354 (I740098,I3042);
DFFARX1 I_43355 (I86634,I3035,I740098,I740124,);
DFFARX1 I_43356 (I86637,I3035,I740098,I740141,);
not I_43357 (I740149,I740141);
nor I_43358 (I740066,I740124,I740149);
DFFARX1 I_43359 (I740149,I3035,I740098,I740081,);
nor I_43360 (I740194,I86643,I86637);
and I_43361 (I740211,I740194,I86640);
nor I_43362 (I740228,I740211,I86643);
not I_43363 (I740245,I86643);
and I_43364 (I740262,I740245,I86634);
nand I_43365 (I740279,I740262,I86652);
nor I_43366 (I740296,I740245,I740279);
DFFARX1 I_43367 (I740296,I3035,I740098,I740063,);
not I_43368 (I740327,I740279);
nand I_43369 (I740344,I740149,I740327);
nand I_43370 (I740075,I740211,I740327);
DFFARX1 I_43371 (I740245,I3035,I740098,I740090,);
not I_43372 (I740389,I86646);
nor I_43373 (I740406,I740389,I86634);
nor I_43374 (I740423,I740406,I740228);
DFFARX1 I_43375 (I740423,I3035,I740098,I740087,);
not I_43376 (I740454,I740406);
DFFARX1 I_43377 (I740454,I3035,I740098,I740480,);
not I_43378 (I740488,I740480);
nor I_43379 (I740084,I740488,I740406);
nor I_43380 (I740519,I740389,I86649);
and I_43381 (I740536,I740519,I86655);
or I_43382 (I740553,I740536,I86658);
DFFARX1 I_43383 (I740553,I3035,I740098,I740579,);
not I_43384 (I740587,I740579);
nand I_43385 (I740604,I740587,I740327);
not I_43386 (I740078,I740604);
nand I_43387 (I740072,I740604,I740344);
nand I_43388 (I740069,I740587,I740211);
not I_43389 (I740693,I3042);
DFFARX1 I_43390 (I400747,I3035,I740693,I740719,);
DFFARX1 I_43391 (I400729,I3035,I740693,I740736,);
not I_43392 (I740744,I740736);
nor I_43393 (I740661,I740719,I740744);
DFFARX1 I_43394 (I740744,I3035,I740693,I740676,);
nor I_43395 (I740789,I400735,I400738);
and I_43396 (I740806,I740789,I400726);
nor I_43397 (I740823,I740806,I400735);
not I_43398 (I740840,I400735);
and I_43399 (I740857,I740840,I400744);
nand I_43400 (I740874,I740857,I400732);
nor I_43401 (I740891,I740840,I740874);
DFFARX1 I_43402 (I740891,I3035,I740693,I740658,);
not I_43403 (I740922,I740874);
nand I_43404 (I740939,I740744,I740922);
nand I_43405 (I740670,I740806,I740922);
DFFARX1 I_43406 (I740840,I3035,I740693,I740685,);
not I_43407 (I740984,I400729);
nor I_43408 (I741001,I740984,I400744);
nor I_43409 (I741018,I741001,I740823);
DFFARX1 I_43410 (I741018,I3035,I740693,I740682,);
not I_43411 (I741049,I741001);
DFFARX1 I_43412 (I741049,I3035,I740693,I741075,);
not I_43413 (I741083,I741075);
nor I_43414 (I740679,I741083,I741001);
nor I_43415 (I741114,I740984,I400741);
and I_43416 (I741131,I741114,I400750);
or I_43417 (I741148,I741131,I400726);
DFFARX1 I_43418 (I741148,I3035,I740693,I741174,);
not I_43419 (I741182,I741174);
nand I_43420 (I741199,I741182,I740922);
not I_43421 (I740673,I741199);
nand I_43422 (I740667,I741199,I740939);
nand I_43423 (I740664,I741182,I740806);
not I_43424 (I741288,I3042);
DFFARX1 I_43425 (I337167,I3035,I741288,I741314,);
DFFARX1 I_43426 (I337161,I3035,I741288,I741331,);
not I_43427 (I741339,I741331);
nor I_43428 (I741256,I741314,I741339);
DFFARX1 I_43429 (I741339,I3035,I741288,I741271,);
nor I_43430 (I741384,I337158,I337149);
and I_43431 (I741401,I741384,I337146);
nor I_43432 (I741418,I741401,I337158);
not I_43433 (I741435,I337158);
and I_43434 (I741452,I741435,I337152);
nand I_43435 (I741469,I741452,I337164);
nor I_43436 (I741486,I741435,I741469);
DFFARX1 I_43437 (I741486,I3035,I741288,I741253,);
not I_43438 (I741517,I741469);
nand I_43439 (I741534,I741339,I741517);
nand I_43440 (I741265,I741401,I741517);
DFFARX1 I_43441 (I741435,I3035,I741288,I741280,);
not I_43442 (I741579,I337170);
nor I_43443 (I741596,I741579,I337152);
nor I_43444 (I741613,I741596,I741418);
DFFARX1 I_43445 (I741613,I3035,I741288,I741277,);
not I_43446 (I741644,I741596);
DFFARX1 I_43447 (I741644,I3035,I741288,I741670,);
not I_43448 (I741678,I741670);
nor I_43449 (I741274,I741678,I741596);
nor I_43450 (I741709,I741579,I337149);
and I_43451 (I741726,I741709,I337155);
or I_43452 (I741743,I741726,I337146);
DFFARX1 I_43453 (I741743,I3035,I741288,I741769,);
not I_43454 (I741777,I741769);
nand I_43455 (I741794,I741777,I741517);
not I_43456 (I741268,I741794);
nand I_43457 (I741262,I741794,I741534);
nand I_43458 (I741259,I741777,I741401);
not I_43459 (I741883,I3042);
DFFARX1 I_43460 (I33122,I3035,I741883,I741909,);
DFFARX1 I_43461 (I33110,I3035,I741883,I741926,);
not I_43462 (I741934,I741926);
nor I_43463 (I741851,I741909,I741934);
DFFARX1 I_43464 (I741934,I3035,I741883,I741866,);
nor I_43465 (I741979,I33101,I33125);
and I_43466 (I741996,I741979,I33104);
nor I_43467 (I742013,I741996,I33101);
not I_43468 (I742030,I33101);
and I_43469 (I742047,I742030,I33107);
nand I_43470 (I742064,I742047,I33119);
nor I_43471 (I742081,I742030,I742064);
DFFARX1 I_43472 (I742081,I3035,I741883,I741848,);
not I_43473 (I742112,I742064);
nand I_43474 (I742129,I741934,I742112);
nand I_43475 (I741860,I741996,I742112);
DFFARX1 I_43476 (I742030,I3035,I741883,I741875,);
not I_43477 (I742174,I33101);
nor I_43478 (I742191,I742174,I33107);
nor I_43479 (I742208,I742191,I742013);
DFFARX1 I_43480 (I742208,I3035,I741883,I741872,);
not I_43481 (I742239,I742191);
DFFARX1 I_43482 (I742239,I3035,I741883,I742265,);
not I_43483 (I742273,I742265);
nor I_43484 (I741869,I742273,I742191);
nor I_43485 (I742304,I742174,I33104);
and I_43486 (I742321,I742304,I33113);
or I_43487 (I742338,I742321,I33116);
DFFARX1 I_43488 (I742338,I3035,I741883,I742364,);
not I_43489 (I742372,I742364);
nand I_43490 (I742389,I742372,I742112);
not I_43491 (I741863,I742389);
nand I_43492 (I741857,I742389,I742129);
nand I_43493 (I741854,I742372,I741996);
not I_43494 (I742478,I3042);
DFFARX1 I_43495 (I598881,I3035,I742478,I742504,);
DFFARX1 I_43496 (I598893,I3035,I742478,I742521,);
not I_43497 (I742529,I742521);
nor I_43498 (I742446,I742504,I742529);
DFFARX1 I_43499 (I742529,I3035,I742478,I742461,);
nor I_43500 (I742574,I598890,I598884);
and I_43501 (I742591,I742574,I598878);
nor I_43502 (I742608,I742591,I598890);
not I_43503 (I742625,I598890);
and I_43504 (I742642,I742625,I598887);
nand I_43505 (I742659,I742642,I598878);
nor I_43506 (I742676,I742625,I742659);
DFFARX1 I_43507 (I742676,I3035,I742478,I742443,);
not I_43508 (I742707,I742659);
nand I_43509 (I742724,I742529,I742707);
nand I_43510 (I742455,I742591,I742707);
DFFARX1 I_43511 (I742625,I3035,I742478,I742470,);
not I_43512 (I742769,I598902);
nor I_43513 (I742786,I742769,I598887);
nor I_43514 (I742803,I742786,I742608);
DFFARX1 I_43515 (I742803,I3035,I742478,I742467,);
not I_43516 (I742834,I742786);
DFFARX1 I_43517 (I742834,I3035,I742478,I742860,);
not I_43518 (I742868,I742860);
nor I_43519 (I742464,I742868,I742786);
nor I_43520 (I742899,I742769,I598896);
and I_43521 (I742916,I742899,I598899);
or I_43522 (I742933,I742916,I598881);
DFFARX1 I_43523 (I742933,I3035,I742478,I742959,);
not I_43524 (I742967,I742959);
nand I_43525 (I742984,I742967,I742707);
not I_43526 (I742458,I742984);
nand I_43527 (I742452,I742984,I742724);
nand I_43528 (I742449,I742967,I742591);
not I_43529 (I743073,I3042);
DFFARX1 I_43530 (I116979,I3035,I743073,I743099,);
DFFARX1 I_43531 (I116982,I3035,I743073,I743116,);
not I_43532 (I743124,I743116);
nor I_43533 (I743041,I743099,I743124);
DFFARX1 I_43534 (I743124,I3035,I743073,I743056,);
nor I_43535 (I743169,I116988,I116982);
and I_43536 (I743186,I743169,I116985);
nor I_43537 (I743203,I743186,I116988);
not I_43538 (I743220,I116988);
and I_43539 (I743237,I743220,I116979);
nand I_43540 (I743254,I743237,I116997);
nor I_43541 (I743271,I743220,I743254);
DFFARX1 I_43542 (I743271,I3035,I743073,I743038,);
not I_43543 (I743302,I743254);
nand I_43544 (I743319,I743124,I743302);
nand I_43545 (I743050,I743186,I743302);
DFFARX1 I_43546 (I743220,I3035,I743073,I743065,);
not I_43547 (I743364,I116991);
nor I_43548 (I743381,I743364,I116979);
nor I_43549 (I743398,I743381,I743203);
DFFARX1 I_43550 (I743398,I3035,I743073,I743062,);
not I_43551 (I743429,I743381);
DFFARX1 I_43552 (I743429,I3035,I743073,I743455,);
not I_43553 (I743463,I743455);
nor I_43554 (I743059,I743463,I743381);
nor I_43555 (I743494,I743364,I116994);
and I_43556 (I743511,I743494,I117000);
or I_43557 (I743528,I743511,I117003);
DFFARX1 I_43558 (I743528,I3035,I743073,I743554,);
not I_43559 (I743562,I743554);
nand I_43560 (I743579,I743562,I743302);
not I_43561 (I743053,I743579);
nand I_43562 (I743047,I743579,I743319);
nand I_43563 (I743044,I743562,I743186);
not I_43564 (I743668,I3042);
DFFARX1 I_43565 (I64742,I3035,I743668,I743694,);
DFFARX1 I_43566 (I64730,I3035,I743668,I743711,);
not I_43567 (I743719,I743711);
nor I_43568 (I743636,I743694,I743719);
DFFARX1 I_43569 (I743719,I3035,I743668,I743651,);
nor I_43570 (I743764,I64721,I64745);
and I_43571 (I743781,I743764,I64724);
nor I_43572 (I743798,I743781,I64721);
not I_43573 (I743815,I64721);
and I_43574 (I743832,I743815,I64727);
nand I_43575 (I743849,I743832,I64739);
nor I_43576 (I743866,I743815,I743849);
DFFARX1 I_43577 (I743866,I3035,I743668,I743633,);
not I_43578 (I743897,I743849);
nand I_43579 (I743914,I743719,I743897);
nand I_43580 (I743645,I743781,I743897);
DFFARX1 I_43581 (I743815,I3035,I743668,I743660,);
not I_43582 (I743959,I64721);
nor I_43583 (I743976,I743959,I64727);
nor I_43584 (I743993,I743976,I743798);
DFFARX1 I_43585 (I743993,I3035,I743668,I743657,);
not I_43586 (I744024,I743976);
DFFARX1 I_43587 (I744024,I3035,I743668,I744050,);
not I_43588 (I744058,I744050);
nor I_43589 (I743654,I744058,I743976);
nor I_43590 (I744089,I743959,I64724);
and I_43591 (I744106,I744089,I64733);
or I_43592 (I744123,I744106,I64736);
DFFARX1 I_43593 (I744123,I3035,I743668,I744149,);
not I_43594 (I744157,I744149);
nand I_43595 (I744174,I744157,I743897);
not I_43596 (I743648,I744174);
nand I_43597 (I743642,I744174,I743914);
nand I_43598 (I743639,I744157,I743781);
not I_43599 (I744263,I3042);
DFFARX1 I_43600 (I34703,I3035,I744263,I744289,);
DFFARX1 I_43601 (I34691,I3035,I744263,I744306,);
not I_43602 (I744314,I744306);
nor I_43603 (I744231,I744289,I744314);
DFFARX1 I_43604 (I744314,I3035,I744263,I744246,);
nor I_43605 (I744359,I34682,I34706);
and I_43606 (I744376,I744359,I34685);
nor I_43607 (I744393,I744376,I34682);
not I_43608 (I744410,I34682);
and I_43609 (I744427,I744410,I34688);
nand I_43610 (I744444,I744427,I34700);
nor I_43611 (I744461,I744410,I744444);
DFFARX1 I_43612 (I744461,I3035,I744263,I744228,);
not I_43613 (I744492,I744444);
nand I_43614 (I744509,I744314,I744492);
nand I_43615 (I744240,I744376,I744492);
DFFARX1 I_43616 (I744410,I3035,I744263,I744255,);
not I_43617 (I744554,I34682);
nor I_43618 (I744571,I744554,I34688);
nor I_43619 (I744588,I744571,I744393);
DFFARX1 I_43620 (I744588,I3035,I744263,I744252,);
not I_43621 (I744619,I744571);
DFFARX1 I_43622 (I744619,I3035,I744263,I744645,);
not I_43623 (I744653,I744645);
nor I_43624 (I744249,I744653,I744571);
nor I_43625 (I744684,I744554,I34685);
and I_43626 (I744701,I744684,I34694);
or I_43627 (I744718,I744701,I34697);
DFFARX1 I_43628 (I744718,I3035,I744263,I744744,);
not I_43629 (I744752,I744744);
nand I_43630 (I744769,I744752,I744492);
not I_43631 (I744243,I744769);
nand I_43632 (I744237,I744769,I744509);
nand I_43633 (I744234,I744752,I744376);
not I_43634 (I744858,I3042);
DFFARX1 I_43635 (I18890,I3035,I744858,I744884,);
DFFARX1 I_43636 (I18872,I3035,I744858,I744901,);
not I_43637 (I744909,I744901);
nor I_43638 (I744826,I744884,I744909);
DFFARX1 I_43639 (I744909,I3035,I744858,I744841,);
nor I_43640 (I744954,I18872,I18887);
and I_43641 (I744971,I744954,I18881);
nor I_43642 (I744988,I744971,I18872);
not I_43643 (I745005,I18872);
and I_43644 (I745022,I745005,I18875);
nand I_43645 (I745039,I745022,I18878);
nor I_43646 (I745056,I745005,I745039);
DFFARX1 I_43647 (I745056,I3035,I744858,I744823,);
not I_43648 (I745087,I745039);
nand I_43649 (I745104,I744909,I745087);
nand I_43650 (I744835,I744971,I745087);
DFFARX1 I_43651 (I745005,I3035,I744858,I744850,);
not I_43652 (I745149,I18884);
nor I_43653 (I745166,I745149,I18875);
nor I_43654 (I745183,I745166,I744988);
DFFARX1 I_43655 (I745183,I3035,I744858,I744847,);
not I_43656 (I745214,I745166);
DFFARX1 I_43657 (I745214,I3035,I744858,I745240,);
not I_43658 (I745248,I745240);
nor I_43659 (I744844,I745248,I745166);
nor I_43660 (I745279,I745149,I18896);
and I_43661 (I745296,I745279,I18893);
or I_43662 (I745313,I745296,I18875);
DFFARX1 I_43663 (I745313,I3035,I744858,I745339,);
not I_43664 (I745347,I745339);
nand I_43665 (I745364,I745347,I745087);
not I_43666 (I744838,I745364);
nand I_43667 (I744832,I745364,I745104);
nand I_43668 (I744829,I745347,I744971);
not I_43669 (I745453,I3042);
DFFARX1 I_43670 (I369535,I3035,I745453,I745479,);
DFFARX1 I_43671 (I369517,I3035,I745453,I745496,);
not I_43672 (I745504,I745496);
nor I_43673 (I745421,I745479,I745504);
DFFARX1 I_43674 (I745504,I3035,I745453,I745436,);
nor I_43675 (I745549,I369523,I369526);
and I_43676 (I745566,I745549,I369514);
nor I_43677 (I745583,I745566,I369523);
not I_43678 (I745600,I369523);
and I_43679 (I745617,I745600,I369532);
nand I_43680 (I745634,I745617,I369520);
nor I_43681 (I745651,I745600,I745634);
DFFARX1 I_43682 (I745651,I3035,I745453,I745418,);
not I_43683 (I745682,I745634);
nand I_43684 (I745699,I745504,I745682);
nand I_43685 (I745430,I745566,I745682);
DFFARX1 I_43686 (I745600,I3035,I745453,I745445,);
not I_43687 (I745744,I369517);
nor I_43688 (I745761,I745744,I369532);
nor I_43689 (I745778,I745761,I745583);
DFFARX1 I_43690 (I745778,I3035,I745453,I745442,);
not I_43691 (I745809,I745761);
DFFARX1 I_43692 (I745809,I3035,I745453,I745835,);
not I_43693 (I745843,I745835);
nor I_43694 (I745439,I745843,I745761);
nor I_43695 (I745874,I745744,I369529);
and I_43696 (I745891,I745874,I369538);
or I_43697 (I745908,I745891,I369514);
DFFARX1 I_43698 (I745908,I3035,I745453,I745934,);
not I_43699 (I745942,I745934);
nand I_43700 (I745959,I745942,I745682);
not I_43701 (I745433,I745959);
nand I_43702 (I745427,I745959,I745699);
nand I_43703 (I745424,I745942,I745566);
not I_43704 (I746048,I3042);
DFFARX1 I_43705 (I529048,I3035,I746048,I746074,);
DFFARX1 I_43706 (I529066,I3035,I746048,I746091,);
not I_43707 (I746099,I746091);
nor I_43708 (I746016,I746074,I746099);
DFFARX1 I_43709 (I746099,I3035,I746048,I746031,);
nor I_43710 (I746144,I529045,I529057);
and I_43711 (I746161,I746144,I529042);
nor I_43712 (I746178,I746161,I529045);
not I_43713 (I746195,I529045);
and I_43714 (I746212,I746195,I529051);
nand I_43715 (I746229,I746212,I529063);
nor I_43716 (I746246,I746195,I746229);
DFFARX1 I_43717 (I746246,I3035,I746048,I746013,);
not I_43718 (I746277,I746229);
nand I_43719 (I746294,I746099,I746277);
nand I_43720 (I746025,I746161,I746277);
DFFARX1 I_43721 (I746195,I3035,I746048,I746040,);
not I_43722 (I746339,I529054);
nor I_43723 (I746356,I746339,I529051);
nor I_43724 (I746373,I746356,I746178);
DFFARX1 I_43725 (I746373,I3035,I746048,I746037,);
not I_43726 (I746404,I746356);
DFFARX1 I_43727 (I746404,I3035,I746048,I746430,);
not I_43728 (I746438,I746430);
nor I_43729 (I746034,I746438,I746356);
nor I_43730 (I746469,I746339,I529042);
and I_43731 (I746486,I746469,I529069);
or I_43732 (I746503,I746486,I529060);
DFFARX1 I_43733 (I746503,I3035,I746048,I746529,);
not I_43734 (I746537,I746529);
nand I_43735 (I746554,I746537,I746277);
not I_43736 (I746028,I746554);
nand I_43737 (I746022,I746554,I746294);
nand I_43738 (I746019,I746537,I746161);
not I_43739 (I746643,I3042);
DFFARX1 I_43740 (I692736,I3035,I746643,I746669,);
DFFARX1 I_43741 (I692727,I3035,I746643,I746686,);
not I_43742 (I746694,I746686);
nor I_43743 (I746611,I746669,I746694);
DFFARX1 I_43744 (I746694,I3035,I746643,I746626,);
nor I_43745 (I746739,I692718,I692733);
and I_43746 (I746756,I746739,I692721);
nor I_43747 (I746773,I746756,I692718);
not I_43748 (I746790,I692718);
and I_43749 (I746807,I746790,I692724);
nand I_43750 (I746824,I746807,I692742);
nor I_43751 (I746841,I746790,I746824);
DFFARX1 I_43752 (I746841,I3035,I746643,I746608,);
not I_43753 (I746872,I746824);
nand I_43754 (I746889,I746694,I746872);
nand I_43755 (I746620,I746756,I746872);
DFFARX1 I_43756 (I746790,I3035,I746643,I746635,);
not I_43757 (I746934,I692718);
nor I_43758 (I746951,I746934,I692724);
nor I_43759 (I746968,I746951,I746773);
DFFARX1 I_43760 (I746968,I3035,I746643,I746632,);
not I_43761 (I746999,I746951);
DFFARX1 I_43762 (I746999,I3035,I746643,I747025,);
not I_43763 (I747033,I747025);
nor I_43764 (I746629,I747033,I746951);
nor I_43765 (I747064,I746934,I692721);
and I_43766 (I747081,I747064,I692730);
or I_43767 (I747098,I747081,I692739);
DFFARX1 I_43768 (I747098,I3035,I746643,I747124,);
not I_43769 (I747132,I747124);
nand I_43770 (I747149,I747132,I746872);
not I_43771 (I746623,I747149);
nand I_43772 (I746617,I747149,I746889);
nand I_43773 (I746614,I747132,I746756);
endmodule


