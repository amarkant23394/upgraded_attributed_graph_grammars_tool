module test_I2733(I1351,I1447,I1431,I1477,I1470,I1359,I2776,I2733);
input I1351,I1447,I1431,I1477,I1470,I1359,I2776;
output I2733;
wire I3217,I2759,I3107,I3200,I3076,I2844,I2827;
nand I_0(I2733,I3217,I3107);
not I_1(I3217,I3200);
not I_2(I2759,I1477);
nor I_3(I3107,I3076,I2844);
DFFARX1 I_4(I1431,I1470,I2759,,,I3200,);
DFFARX1 I_5(I1447,I1470,I2759,,,I3076,);
nand I_6(I2844,I2827,I1359);
nor I_7(I2827,I2776,I1351);
endmodule


