module test_I15423(I14982,I1477,I1470,I15423);
input I14982,I1477,I1470;
output I15423;
wire I12619,I12602,I12670,I12913,I12584,I12930,I15047,I15064,I15389,I15406,I12587,I14965,I15372,I10609;
not I_0(I12619,I1477);
not I_1(I12602,I12930);
DFFARX1 I_2(I1470,I12619,,,I12670,);
DFFARX1 I_3(I1470,I12619,,,I12913,);
and I_4(I12584,I12670);
and I_5(I12930,I12913,I10609);
nor I_6(I15047,I14982,I12584);
nand I_7(I15064,I15047,I12587);
not I_8(I15389,I15372);
nor I_9(I15406,I15064,I15389);
DFFARX1 I_10(I12670,I1470,I12619,,,I12587,);
not I_11(I14965,I1477);
DFFARX1 I_12(I12602,I1470,I14965,,,I15372,);
and I_13(I15423,I15372,I15406);
DFFARX1 I_14(I1470,,,I10609,);
endmodule


