module test_I7652(I3966,I6589,I1477,I6442,I1470,I7652);
input I3966,I6589,I1477,I6442,I1470;
output I7652;
wire I6606,I6781,I6297,I6826,I7587,I6329,I6843,I6493,I6300;
DFFARX1 I_0(I6589,I1470,I6329,,,I6606,);
DFFARX1 I_1(I1470,I6329,,,I6781,);
DFFARX1 I_2(I6843,I1470,I6329,,,I6297,);
nor I_3(I7652,I7587,I6297);
nand I_4(I6826,I6781,I6442);
not I_5(I7587,I6300);
not I_6(I6329,I1477);
and I_7(I6843,I6493,I6826);
DFFARX1 I_8(I3966,I1470,I6329,,,I6493,);
DFFARX1 I_9(I6606,I1470,I6329,,,I6300,);
endmodule


