module test_I2440(I1223,I1294,I1207,I1239,I1301,I2440);
input I1223,I1294,I1207,I1239,I1301;
output I2440;
wire I1410,I1328,I1622,I2313,I1310,I1937,I2087,I2423,I1331,I2070,I2389,I1639,I2406;
nor I_0(I1410,I1223,I1239);
nand I_1(I1328,I1639);
DFFARX1 I_2(I1294,,,I1622,);
and I_3(I2440,I2313,I2423);
DFFARX1 I_4(I1331,I1294,I1937,,,I2313,);
DFFARX1 I_5(I1294,,,I1310,);
not I_6(I1937,I1301);
not I_7(I2087,I2070);
nor I_8(I2423,I2406,I2087);
nor I_9(I1331,I1639,I1410);
not I_10(I2070,I1310);
DFFARX1 I_11(I1328,I1294,I1937,,,I2389,);
and I_12(I1639,I1622,I1207);
not I_13(I2406,I2389);
endmodule


