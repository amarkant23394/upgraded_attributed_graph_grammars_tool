module test_final(IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_4_2_l_6,IN_5_2_l_6,IN_1_6_l_6,IN_2_6_l_6,IN_3_6_l_6,IN_4_6_l_6,IN_5_6_l_6,IN_1_9_l_6,IN_2_9_l_6,IN_3_9_l_6,IN_4_9_l_6,IN_5_9_l_6,blif_clk_net_8_r_10,blif_reset_net_8_r_10,N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10);
input IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_4_2_l_6,IN_5_2_l_6,IN_1_6_l_6,IN_2_6_l_6,IN_3_6_l_6,IN_4_6_l_6,IN_5_6_l_6,IN_1_9_l_6,IN_2_9_l_6,IN_3_9_l_6,IN_4_9_l_6,IN_5_9_l_6,blif_clk_net_8_r_10,blif_reset_net_8_r_10;
output N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10;
wire N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,I_BUFF_1_9_r_6,N1372_10_r_6,N1508_10_r_6,N3_8_r_6,n30_6,n31_6,n32_6,n33_6,n34_6,n35_6,n36_6,n37_6,n38_6,n39_6,n40_6,n41_6,n42_6,n43_6,n44_6,n45_6,n46_6,n47_6,n48_6,n49_6,n50_6,n51_6,n52_6,n53_6,n54_6,N1372_4_r_10,I_BUFF_1_9_r_10,N3_8_r_10,n11_10,n35_10,n36_10,n37_10,n38_10,n39_10,n40_10,n41_10,n42_10,n43_10,n44_10,n45_10,n46_10,n47_10,n48_10,n49_10,n50_10,n51_10,n52_10,n53_10,n54_10,n55_10,n56_10,n57_10,n58_10,n59_10,n60_10,n61_10,n62_10,n63_10,n64_10;
nor I_0(N1371_0_r_6,n30_6,n33_6);
nor I_1(N1508_0_r_6,n33_6,n44_6);
not I_2(N1372_1_r_6,n41_6);
nor I_3(N1508_1_r_6,n40_6,n41_6);
nor I_4(N1507_6_r_6,n39_6,n45_6);
nor I_5(N1508_6_r_6,n37_6,n38_6);
nor I_6(n_42_8_r_6,n30_6,n31_6);
DFFARX1 I_7(N3_8_r_6,blif_clk_net_8_r_10,n11_10,G199_8_r_6,);
nor I_8(N6147_9_r_6,n32_6,n33_6);
nor I_9(N6134_9_r_6,I_BUFF_1_9_r_6,n35_6);
not I_10(I_BUFF_1_9_r_6,n37_6);
not I_11(N1372_10_r_6,n43_6);
nor I_12(N1508_10_r_6,n42_6,n43_6);
nor I_13(N3_8_r_6,IN_1_9_l_6,n36_6);
nor I_14(n30_6,IN_5_9_l_6,n53_6);
not I_15(n31_6,n36_6);
nor I_16(n32_6,I_BUFF_1_9_r_6,n34_6);
not I_17(n33_6,IN_1_9_l_6);
not I_18(n34_6,n35_6);
nand I_19(n35_6,IN_2_6_l_6,n49_6);
nand I_20(n36_6,IN_5_6_l_6,n51_6);
nand I_21(n37_6,IN_2_9_l_6,n54_6);
or I_22(n38_6,n35_6,n39_6);
nor I_23(n39_6,n40_6,n45_6);
and I_24(n40_6,n46_6,n47_6);
nand I_25(n41_6,n30_6,n31_6);
nor I_26(n42_6,n34_6,n40_6);
nand I_27(n43_6,IN_1_9_l_6,n30_6);
nor I_28(n44_6,n31_6,n40_6);
nor I_29(n45_6,n35_6,n36_6);
nor I_30(n46_6,IN_1_2_l_6,IN_2_2_l_6);
or I_31(n47_6,IN_5_2_l_6,n48_6);
nor I_32(n48_6,IN_3_2_l_6,IN_4_2_l_6);
and I_33(n49_6,IN_1_6_l_6,n50_6);
nand I_34(n50_6,n51_6,n52_6);
nand I_35(n51_6,IN_3_6_l_6,IN_4_6_l_6);
not I_36(n52_6,IN_5_6_l_6);
nor I_37(n53_6,IN_3_9_l_6,IN_4_9_l_6);
or I_38(n54_6,IN_3_9_l_6,IN_4_9_l_6);
nor I_39(N1371_0_r_10,n37_10,n38_10);
nor I_40(N1508_0_r_10,n37_10,n58_10);
nand I_41(N6147_2_r_10,n39_10,n40_10);
not I_42(N6147_3_r_10,n39_10);
nor I_43(N1372_4_r_10,n46_10,n49_10);
nor I_44(N1508_4_r_10,n51_10,n52_10);
nor I_45(N1507_6_r_10,n49_10,n60_10);
nor I_46(N1508_6_r_10,n49_10,n50_10);
nor I_47(n_42_8_r_10,I_BUFF_1_9_r_10,n35_10);
DFFARX1 I_48(N3_8_r_10,blif_clk_net_8_r_10,n11_10,G199_8_r_10,);
nor I_49(N6147_9_r_10,n36_10,n37_10);
nor I_50(N6134_9_r_10,I_BUFF_1_9_r_10,n46_10);
not I_51(I_BUFF_1_9_r_10,n48_10);
nor I_52(N3_8_r_10,n44_10,n47_10);
not I_53(n11_10,blif_reset_net_8_r_10);
not I_54(n35_10,n49_10);
nor I_55(n36_10,I_BUFF_1_9_r_10,n38_10);
not I_56(n37_10,N1371_0_r_6);
not I_57(n38_10,n46_10);
nand I_58(n39_10,n43_10,n44_10);
nand I_59(n40_10,I_BUFF_1_9_r_10,n41_10);
nor I_60(n41_10,n42_10,N1371_0_r_6);
not I_61(n42_10,n44_10);
nor I_62(n43_10,n45_10,N1371_0_r_6);
nand I_63(n44_10,n54_10,N1372_1_r_6);
nor I_64(n45_10,n59_10,N1507_6_r_6);
nand I_65(n46_10,n61_10,N1508_6_r_6);
nor I_66(n47_10,n46_10,n48_10);
nand I_67(n48_10,n62_10,n63_10);
nand I_68(n49_10,n56_10,N6147_9_r_6);
not I_69(n50_10,n45_10);
nor I_70(n51_10,n42_10,n53_10);
not I_71(n52_10,N1372_4_r_10);
nor I_72(n53_10,n48_10,n50_10);
and I_73(n54_10,n55_10,N1372_10_r_6);
nand I_74(n55_10,n56_10,n57_10);
nand I_75(n56_10,N1508_0_r_6,N1508_1_r_6);
not I_76(n57_10,N6147_9_r_6);
nor I_77(n58_10,n35_10,n45_10);
nor I_78(n59_10,N1372_1_r_6,G199_8_r_6);
nor I_79(n60_10,n37_10,n46_10);
or I_80(n61_10,N1372_1_r_6,G199_8_r_6);
nor I_81(n62_10,N1371_0_r_6,N6134_9_r_6);
or I_82(n63_10,n64_10,N1508_0_r_6);
nor I_83(n64_10,n_42_8_r_6,N1508_10_r_6);
endmodule


