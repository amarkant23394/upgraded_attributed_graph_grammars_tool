module test_I5450(I1477,I3521,I1470,I5317,I3685,I3572,I5450);
input I1477,I3521,I1470,I5317,I3685,I3572;
output I5450;
wire I5416,I3388,I5351,I3362,I3350,I5334,I5122,I5433,I3589,I3356,I5105;
nand I_0(I5416,I5122,I3356);
and I_1(I5450,I5416,I5433);
not I_2(I3388,I1477);
DFFARX1 I_3(I5334,I1470,I5105,,,I5351,);
DFFARX1 I_4(I1470,I3388,,,I3362,);
DFFARX1 I_5(I3685,I1470,I3388,,,I3350,);
or I_6(I5334,I5317,I3362);
not I_7(I5122,I3350);
nand I_8(I5433,I5416,I5351);
and I_9(I3589,I3521,I3572);
DFFARX1 I_10(I3589,I1470,I3388,,,I3356,);
not I_11(I5105,I1477);
endmodule


