module test_I5091(I1477,I3521,I3405,I5317,I3798,I1470,I5091);
input I1477,I3521,I3405,I5317,I3798,I1470;
output I5091;
wire I5266,I5385,I3815,I5249,I3747,I5156,I3388,I3846,I3362,I5334,I3371,I3380,I5139,I5105,I3359,I5351;
not I_0(I5266,I5249);
nor I_1(I5385,I5351,I5266);
or I_2(I3815,I3405,I3798);
not I_3(I5249,I3380);
DFFARX1 I_4(I1470,I3388,,,I3747,);
nand I_5(I5156,I5139,I3371);
not I_6(I3388,I1477);
nand I_7(I5091,I5156,I5385);
nor I_8(I3846,I3747);
DFFARX1 I_9(I1470,I3388,,,I3362,);
or I_10(I5334,I5317,I3362);
DFFARX1 I_11(I3815,I1470,I3388,,,I3371,);
nand I_12(I3380,I3521,I3846);
nor I_13(I5139,I3380,I3359);
not I_14(I5105,I1477);
DFFARX1 I_15(I3747,I1470,I3388,,,I3359,);
DFFARX1 I_16(I5334,I1470,I5105,,,I5351,);
endmodule


