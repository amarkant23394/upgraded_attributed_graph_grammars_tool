module test_final(IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_6_2_l_6,IN_1_3_l_6,IN_2_3_l_6,IN_4_3_l_6,IN_1_4_l_6,IN_2_4_l_6,IN_3_4_l_6,IN_6_4_l_6,blif_clk_net_1_r_10,blif_reset_net_1_r_10,G42_1_r_10,n_572_1_r_10,n_573_1_r_10,n_549_1_r_10,n_42_2_r_10,G199_2_r_10,ACVQN2_3_r_10,n_266_and_0_3_r_10);
input IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_6_2_l_6,IN_1_3_l_6,IN_2_3_l_6,IN_4_3_l_6,IN_1_4_l_6,IN_2_4_l_6,IN_3_4_l_6,IN_6_4_l_6,blif_clk_net_1_r_10,blif_reset_net_1_r_10;
output G42_1_r_10,n_572_1_r_10,n_573_1_r_10,n_549_1_r_10,n_42_2_r_10,G199_2_r_10,ACVQN2_3_r_10,n_266_and_0_3_r_10;
wire G42_1_r_6,n_572_1_r_6,n_573_1_r_6,n_549_1_r_6,n_569_1_r_6,n_452_1_r_6,G199_4_r_6,G214_4_r_6,ACVQN1_5_r_6,P6_5_r_6,N3_2_l_6,n27_6,n17_6,n28_6,n26_6,N1_4_l_6,n29_6,n18_6,G214_4_l_6,n12_6,n4_1_r_6,N1_4_r_6,n_42_2_l_6,P6_5_r_internal_6,n19_6,n20_6,n21_6,n22_6,n23_6,n24_6,n25_6,n_452_1_r_10,N3_2_l_10,n4_10,n25_10,n16_10,n26_10,ACVQN1_3_l_10,N1_4_l_10,G199_4_l_10,n27_10,n17_10,n4_1_r_10,N3_2_r_10,n3_10,n13_internal_10,n13_10,n18_10,n19_10,n20_10,n21_10,n22_10,n23_10,n24_10;
DFFARX1 I_0(n4_1_r_6,blif_clk_net_1_r_10,n4_10,G42_1_r_6,);
nor I_1(n_572_1_r_6,n27_6,n28_6);
nand I_2(n_573_1_r_6,n18_6,n19_6);
nor I_3(n_549_1_r_6,n_42_2_l_6,n21_6);
nand I_4(n_569_1_r_6,n19_6,n20_6);
nor I_5(n_452_1_r_6,n28_6,n29_6);
DFFARX1 I_6(N1_4_r_6,blif_clk_net_1_r_10,n4_10,G199_4_r_6,);
DFFARX1 I_7(n_42_2_l_6,blif_clk_net_1_r_10,n4_10,G214_4_r_6,);
DFFARX1 I_8(n_42_2_l_6,blif_clk_net_1_r_10,n4_10,ACVQN1_5_r_6,);
not I_9(P6_5_r_6,P6_5_r_internal_6);
and I_10(N3_2_l_6,IN_6_2_l_6,n23_6);
DFFARX1 I_11(N3_2_l_6,blif_clk_net_1_r_10,n4_10,n27_6,);
not I_12(n17_6,n27_6);
DFFARX1 I_13(IN_1_3_l_6,blif_clk_net_1_r_10,n4_10,n28_6,);
DFFARX1 I_14(IN_2_3_l_6,blif_clk_net_1_r_10,n4_10,n26_6,);
and I_15(N1_4_l_6,IN_6_4_l_6,n25_6);
DFFARX1 I_16(N1_4_l_6,blif_clk_net_1_r_10,n4_10,n29_6,);
not I_17(n18_6,n29_6);
DFFARX1 I_18(IN_3_4_l_6,blif_clk_net_1_r_10,n4_10,G214_4_l_6,);
not I_19(n12_6,G214_4_l_6);
nor I_20(n4_1_r_6,n28_6,n22_6);
nor I_21(N1_4_r_6,n12_6,n24_6);
nor I_22(n_42_2_l_6,IN_1_2_l_6,IN_3_2_l_6);
DFFARX1 I_23(G214_4_l_6,blif_clk_net_1_r_10,n4_10,P6_5_r_internal_6,);
nand I_24(n19_6,IN_4_3_l_6,n26_6);
not I_25(n20_6,n_42_2_l_6);
nor I_26(n21_6,n17_6,n28_6);
and I_27(n22_6,IN_4_3_l_6,n26_6);
nand I_28(n23_6,IN_2_2_l_6,IN_3_2_l_6);
nor I_29(n24_6,n17_6,n18_6);
nand I_30(n25_6,IN_1_4_l_6,IN_2_4_l_6);
DFFARX1 I_31(n4_1_r_10,blif_clk_net_1_r_10,n4_10,G42_1_r_10,);
nor I_32(n_572_1_r_10,n26_10,n3_10);
nand I_33(n_573_1_r_10,n16_10,n18_10);
nand I_34(n_549_1_r_10,n19_10,n20_10);
nor I_35(n_452_1_r_10,n25_10,n21_10);
nor I_36(n_42_2_r_10,n26_10,G199_4_l_10);
DFFARX1 I_37(N3_2_r_10,blif_clk_net_1_r_10,n4_10,G199_2_r_10,);
DFFARX1 I_38(G199_4_l_10,blif_clk_net_1_r_10,n4_10,ACVQN2_3_r_10,);
nor I_39(n_266_and_0_3_r_10,n17_10,n13_10);
and I_40(N3_2_l_10,n23_10,G42_1_r_6);
not I_41(n4_10,blif_reset_net_1_r_10);
DFFARX1 I_42(N3_2_l_10,blif_clk_net_1_r_10,n4_10,n25_10,);
not I_43(n16_10,n25_10);
DFFARX1 I_44(n_569_1_r_6,blif_clk_net_1_r_10,n4_10,n26_10,);
DFFARX1 I_45(n_549_1_r_6,blif_clk_net_1_r_10,n4_10,ACVQN1_3_l_10,);
and I_46(N1_4_l_10,n24_10,n_452_1_r_6);
DFFARX1 I_47(N1_4_l_10,blif_clk_net_1_r_10,n4_10,G199_4_l_10,);
DFFARX1 I_48(G42_1_r_6,blif_clk_net_1_r_10,n4_10,n27_10,);
not I_49(n17_10,n27_10);
nor I_50(n4_1_r_10,n27_10,n21_10);
nor I_51(N3_2_r_10,n16_10,n22_10);
not I_52(n3_10,n18_10);
DFFARX1 I_53(n3_10,blif_clk_net_1_r_10,n4_10,n13_internal_10,);
not I_54(n13_10,n13_internal_10);
nand I_55(n18_10,ACVQN1_3_l_10,ACVQN1_5_r_6);
not I_56(n19_10,n_452_1_r_10);
nand I_57(n20_10,n16_10,n26_10);
nor I_58(n21_10,n_572_1_r_6,G199_4_r_6);
and I_59(n22_10,n26_10,n21_10);
nand I_60(n23_10,n_572_1_r_6,G214_4_r_6);
nand I_61(n24_10,n_573_1_r_6,P6_5_r_6);
endmodule


