module test_I4869(I1477,I2294,I1470,I1375,I4869);
input I1477,I2294,I1470,I1375;
output I4869;
wire I2181,I4544,I2149,I2678,I2345,I2633,I2695;
not I_0(I2181,I1477);
not I_1(I4544,I1477);
DFFARX1 I_2(I2149,I1470,I4544,,,I4869,);
DFFARX1 I_3(I2695,I1470,I2181,,,I2149,);
nand I_4(I2678,I2633,I2294);
DFFARX1 I_5(I1375,I1470,I2181,,,I2345,);
DFFARX1 I_6(I1470,I2181,,,I2633,);
and I_7(I2695,I2345,I2678);
endmodule


