module test_I10630(I1477,I1470,I10630);
input I1477,I1470;
output I10630;
wire I10647,I9491,I9816,I9468,I11009,I9621,I9864;
not I_0(I10647,I1477);
not I_1(I9491,I1477);
DFFARX1 I_2(I1470,I9491,,,I9816,);
DFFARX1 I_3(I9864,I1470,I9491,,,I9468,);
not I_4(I10630,I11009);
DFFARX1 I_5(I9468,I1470,I10647,,,I11009,);
DFFARX1 I_6(I1470,I9491,,,I9621,);
nor I_7(I9864,I9816,I9621);
endmodule


