module Benchmark_testing100(I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1294,I1301,I1316,I1310,I1307,I1319,I1304,I1325,I1334,I1328,I1331,I1322,I1313);
input I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1294,I1301;
output I1316,I1310,I1307,I1319,I1304,I1325,I1334,I1328,I1331,I1322,I1313;
wire I1207,I1215,I1223,I1231,I1239,I1247,I1255,I1263,I1271,I1279,I1287,I1294,I1301,I1342,I1359,I1899,I1914,I1376,I1902,I1407,I1905,I1920,I1424,I1441,I1458,I1908,I1475,I1492,I1911,I1929,I1509,I1526,I1543,I1574,I1591,I1622,I1926,I1639,I1917,I1656,I1701,I1923,I1718,I1735,I1752,I1769,I1800,I1831,I1937,I1954,I3237,I1971,I3234,I3252,I1988,I3255,I2005,I2022,I3240,I2039,I2056,I2087,I2118,I3249,I2135,I3231,I2152,I3225,I2169,I3243,I2186,I2203,I2220,I2251,I2268,I2299,I3228,I2316,I2347,I2378,I2395,I2440,I3246,I2457,I2474,I2491,I2522,I2600,I2617,I2634,I2651,I2668,I2685,I2702,I2719,I2589,I2750,I2574,I2781,I2798,I2815,I2832,I2849,I2866,I2883,I2571,I2914,I2931,I2568,I2962,I2979,I2586,I3010,I2583,I3041,I3058,I2562,I2565,I3103,I3120,I3137,I3154,I2592,I3185,I2577,I2580,I3263,I3280,I3297,I3314,I3331,I3348,I3365,I3396,I3413,I3430,I3447,I3464,I3481,I3498,I3529,I3560,I3577,I3594,I3639,I3670,I3715,I3732,I3749,I3766,I3783,I3814,I3831;
not I_0 (I1342,I1301);
or I_1 (I1359,I1899,I1914);
or I_2 (I1376,I1902,I1899);
DFFARX1 I_3  ( .D(I1376), .CLK(I1294), .RSTB(I1342), .Q(I1316) );
nor I_4 (I1407,I1905,I1920);
not I_5 (I1424,I1407);
not I_6 (I1441,I1905);
and I_7 (I1458,I1441,I1908);
nor I_8 (I1475,I1458,I1914);
nor I_9 (I1492,I1911,I1929);
DFFARX1 I_10  ( .D(I1492), .CLK(I1294), .RSTB(I1342), .Q(I1509) );
nand I_11 (I1526,I1509,I1359);
and I_12 (I1543,I1475,I1526);
DFFARX1 I_13  ( .D(I1543), .CLK(I1294), .RSTB(I1342), .Q(I1310) );
nor I_14 (I1574,I1911,I1902);
DFFARX1 I_15  ( .D(I1574), .CLK(I1294), .RSTB(I1342), .Q(I1591) );
and I_16 (I1307,I1407,I1591);
DFFARX1 I_17  ( .D(I1926), .CLK(I1294), .RSTB(I1342), .Q(I1622) );
and I_18 (I1639,I1622,I1917);
DFFARX1 I_19  ( .D(I1639), .CLK(I1294), .RSTB(I1342), .Q(I1656) );
not I_20 (I1319,I1656);
DFFARX1 I_21  ( .D(I1639), .CLK(I1294), .RSTB(I1342), .Q(I1304) );
DFFARX1 I_22  ( .D(I1923), .CLK(I1294), .RSTB(I1342), .Q(I1701) );
not I_23 (I1718,I1701);
nor I_24 (I1735,I1376,I1718);
and I_25 (I1752,I1639,I1735);
or I_26 (I1769,I1359,I1752);
DFFARX1 I_27  ( .D(I1769), .CLK(I1294), .RSTB(I1342), .Q(I1325) );
nor I_28 (I1800,I1701,I1509);
nand I_29 (I1334,I1475,I1800);
nor I_30 (I1831,I1701,I1424);
nand I_31 (I1328,I1574,I1831);
not I_32 (I1331,I1701);
nand I_33 (I1322,I1701,I1424);
DFFARX1 I_34  ( .D(I1701), .CLK(I1294), .RSTB(I1342), .Q(I1313) );
not I_35 (I1937,I1301);
not I_36 (I1954,I3237);
nor I_37 (I1971,I3234,I3252);
nand I_38 (I1988,I1971,I3255);
nor I_39 (I2005,I1954,I3234);
nand I_40 (I2022,I2005,I3240);
not I_41 (I2039,I2022);
not I_42 (I2056,I3234);
nor I_43 (I1926,I2022,I2056);
not I_44 (I2087,I2056);
nand I_45 (I1911,I2022,I2087);
not I_46 (I2118,I3249);
nor I_47 (I2135,I2118,I3231);
and I_48 (I2152,I2135,I3225);
or I_49 (I2169,I2152,I3243);
DFFARX1 I_50  ( .D(I2169), .CLK(I1294), .RSTB(I1937), .Q(I2186) );
nor I_51 (I2203,I2186,I2039);
DFFARX1 I_52  ( .D(I2186), .CLK(I1294), .RSTB(I1937), .Q(I2220) );
not I_53 (I1908,I2220);
nand I_54 (I2251,I1954,I3249);
and I_55 (I2268,I2251,I2203);
DFFARX1 I_56  ( .D(I2251), .CLK(I1294), .RSTB(I1937), .Q(I1905) );
DFFARX1 I_57  ( .D(I3228), .CLK(I1294), .RSTB(I1937), .Q(I2299) );
nor I_58 (I2316,I2299,I2022);
nand I_59 (I1923,I2186,I2316);
nor I_60 (I2347,I2299,I2087);
not I_61 (I1920,I2299);
nand I_62 (I2378,I2299,I1988);
and I_63 (I2395,I2056,I2378);
DFFARX1 I_64  ( .D(I2395), .CLK(I1294), .RSTB(I1937), .Q(I1899) );
DFFARX1 I_65  ( .D(I2299), .CLK(I1294), .RSTB(I1937), .Q(I1902) );
DFFARX1 I_66  ( .D(I3246), .CLK(I1294), .RSTB(I1937), .Q(I2440) );
not I_67 (I2457,I2440);
nand I_68 (I2474,I2457,I2022);
and I_69 (I2491,I2251,I2474);
DFFARX1 I_70  ( .D(I2491), .CLK(I1294), .RSTB(I1937), .Q(I1929) );
or I_71 (I2522,I2457,I2268);
DFFARX1 I_72  ( .D(I2522), .CLK(I1294), .RSTB(I1937), .Q(I1914) );
nand I_73 (I1917,I2457,I2347);
not I_74 (I2600,I1301);
not I_75 (I2617,I1287);
nor I_76 (I2634,I1271,I1231);
nand I_77 (I2651,I2634,I1215);
nor I_78 (I2668,I2617,I1271);
nand I_79 (I2685,I2668,I1255);
not I_80 (I2702,I2685);
not I_81 (I2719,I1271);
nor I_82 (I2589,I2685,I2719);
not I_83 (I2750,I2719);
nand I_84 (I2574,I2685,I2750);
not I_85 (I2781,I1279);
nor I_86 (I2798,I2781,I1239);
and I_87 (I2815,I2798,I1207);
or I_88 (I2832,I2815,I1263);
DFFARX1 I_89  ( .D(I2832), .CLK(I1294), .RSTB(I2600), .Q(I2849) );
nor I_90 (I2866,I2849,I2702);
DFFARX1 I_91  ( .D(I2849), .CLK(I1294), .RSTB(I2600), .Q(I2883) );
not I_92 (I2571,I2883);
nand I_93 (I2914,I2617,I1279);
and I_94 (I2931,I2914,I2866);
DFFARX1 I_95  ( .D(I2914), .CLK(I1294), .RSTB(I2600), .Q(I2568) );
DFFARX1 I_96  ( .D(I1223), .CLK(I1294), .RSTB(I2600), .Q(I2962) );
nor I_97 (I2979,I2962,I2685);
nand I_98 (I2586,I2849,I2979);
nor I_99 (I3010,I2962,I2750);
not I_100 (I2583,I2962);
nand I_101 (I3041,I2962,I2651);
and I_102 (I3058,I2719,I3041);
DFFARX1 I_103  ( .D(I3058), .CLK(I1294), .RSTB(I2600), .Q(I2562) );
DFFARX1 I_104  ( .D(I2962), .CLK(I1294), .RSTB(I2600), .Q(I2565) );
DFFARX1 I_105  ( .D(I1247), .CLK(I1294), .RSTB(I2600), .Q(I3103) );
not I_106 (I3120,I3103);
nand I_107 (I3137,I3120,I2685);
and I_108 (I3154,I2914,I3137);
DFFARX1 I_109  ( .D(I3154), .CLK(I1294), .RSTB(I2600), .Q(I2592) );
or I_110 (I3185,I3120,I2931);
DFFARX1 I_111  ( .D(I3185), .CLK(I1294), .RSTB(I2600), .Q(I2577) );
nand I_112 (I2580,I3120,I3010);
not I_113 (I3263,I1301);
not I_114 (I3280,I2586);
nor I_115 (I3297,I2565,I2577);
nand I_116 (I3314,I3297,I2580);
nor I_117 (I3331,I3280,I2565);
nand I_118 (I3348,I3331,I2562);
DFFARX1 I_119  ( .D(I3348), .CLK(I1294), .RSTB(I3263), .Q(I3365) );
not I_120 (I3234,I3365);
not I_121 (I3396,I2565);
not I_122 (I3413,I3396);
not I_123 (I3430,I2583);
nor I_124 (I3447,I3430,I2574);
and I_125 (I3464,I3447,I2568);
or I_126 (I3481,I3464,I2592);
DFFARX1 I_127  ( .D(I3481), .CLK(I1294), .RSTB(I3263), .Q(I3498) );
DFFARX1 I_128  ( .D(I3498), .CLK(I1294), .RSTB(I3263), .Q(I3231) );
DFFARX1 I_129  ( .D(I3498), .CLK(I1294), .RSTB(I3263), .Q(I3529) );
DFFARX1 I_130  ( .D(I3498), .CLK(I1294), .RSTB(I3263), .Q(I3225) );
nand I_131 (I3560,I3280,I2583);
nand I_132 (I3577,I3560,I3314);
and I_133 (I3594,I3396,I3577);
DFFARX1 I_134  ( .D(I3594), .CLK(I1294), .RSTB(I3263), .Q(I3255) );
and I_135 (I3228,I3560,I3529);
DFFARX1 I_136  ( .D(I2589), .CLK(I1294), .RSTB(I3263), .Q(I3639) );
nor I_137 (I3252,I3639,I3560);
nor I_138 (I3670,I3639,I3314);
nand I_139 (I3249,I3348,I3670);
not I_140 (I3246,I3639);
DFFARX1 I_141  ( .D(I2571), .CLK(I1294), .RSTB(I3263), .Q(I3715) );
not I_142 (I3732,I3715);
nor I_143 (I3749,I3732,I3413);
and I_144 (I3766,I3639,I3749);
or I_145 (I3783,I3560,I3766);
DFFARX1 I_146  ( .D(I3783), .CLK(I1294), .RSTB(I3263), .Q(I3240) );
not I_147 (I3814,I3732);
nor I_148 (I3831,I3639,I3814);
nand I_149 (I3243,I3732,I3831);
nand I_150 (I3237,I3396,I3814);
endmodule


