module test_I10397(I8107,I6321,I7714,I1477,I1470,I10397);
input I8107,I6321,I7714,I1477,I1470;
output I10397;
wire I10349,I7550,I7570,I7977,I7731,I10052,I7532,I10332;
and I_0(I10349,I10332,I7550);
nand I_1(I7550,I7977,I7731);
not I_2(I7570,I1477);
not I_3(I10397,I10349);
DFFARX1 I_4(I6321,I1470,I7570,,,I7977,);
not I_5(I7731,I7714);
not I_6(I10052,I1477);
DFFARX1 I_7(I8107,I1470,I7570,,,I7532,);
DFFARX1 I_8(I7532,I1470,I10052,,,I10332,);
endmodule


