module test_final(IN_1_1_l_9,IN_2_1_l_9,IN_3_1_l_9,G18_7_l_9,G15_7_l_9,IN_1_7_l_9,IN_4_7_l_9,IN_5_7_l_9,IN_7_7_l_9,IN_9_7_l_9,IN_10_7_l_9,IN_1_8_l_9,IN_2_8_l_9,IN_3_8_l_9,IN_6_8_l_9,blif_clk_net_8_r_8,blif_reset_net_8_r_8,N1371_0_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,N1508_10_r_8);
input IN_1_1_l_9,IN_2_1_l_9,IN_3_1_l_9,G18_7_l_9,G15_7_l_9,IN_1_7_l_9,IN_4_7_l_9,IN_5_7_l_9,IN_7_7_l_9,IN_9_7_l_9,IN_10_7_l_9,IN_1_8_l_9,IN_2_8_l_9,IN_3_8_l_9,IN_6_8_l_9,blif_clk_net_8_r_8,blif_reset_net_8_r_8;
output N1371_0_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,N1508_10_r_8;
wire N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,n_429_or_0_5_r_9,G78_5_r_9,n_576_5_r_9,n_102_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9,I_BUFF_1_9_r_9,n4_7_l_9,n62_9,N3_8_l_9,n63_9,n38_9,n_431_5_r_9,N3_8_r_9,n39_9,n40_9,n41_9,n42_9,n43_9,n44_9,n45_9,n46_9,n47_9,n48_9,n49_9,n50_9,n51_9,n52_9,n53_9,n54_9,n55_9,n56_9,n57_9,n58_9,n59_9,n60_9,n61_9,N1508_0_r_8,N1372_1_r_8,I_BUFF_1_9_r_8,N1372_10_r_8,N3_8_l_8,n8_8,n53_8,n29_8,N3_8_r_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8,n38_8,n39_8,n40_8,n41_8,n42_8,n43_8,n44_8,n45_8,n46_8,n47_8,n48_8,n49_8,n50_8,n51_8,n52_8;
nor I_0(N6147_2_r_9,n62_9,n46_9);
not I_1(N1372_4_r_9,n59_9);
nor I_2(N1508_4_r_9,n58_9,n59_9);
nand I_3(n_429_or_0_5_r_9,n_431_5_r_9,n42_9);
DFFARX1 I_4(n_431_5_r_9,blif_clk_net_8_r_8,n8_8,G78_5_r_9,);
nand I_5(n_576_5_r_9,n39_9,n40_9);
not I_6(n_102_5_r_9,I_BUFF_1_9_r_9);
nand I_7(n_547_5_r_9,IN_3_1_l_9,n43_9);
and I_8(n_42_8_r_9,G18_7_l_9,n44_9);
DFFARX1 I_9(N3_8_r_9,blif_clk_net_8_r_8,n8_8,G199_8_r_9,);
nor I_10(N6147_9_r_9,n41_9,n45_9);
nor I_11(N6134_9_r_9,n45_9,n51_9);
nor I_12(I_BUFF_1_9_r_9,IN_3_1_l_9,n41_9);
nor I_13(n4_7_l_9,G18_7_l_9,IN_1_7_l_9);
DFFARX1 I_14(n4_7_l_9,blif_clk_net_8_r_8,n8_8,n62_9,);
and I_15(N3_8_l_9,IN_6_8_l_9,n57_9);
DFFARX1 I_16(N3_8_l_9,blif_clk_net_8_r_8,n8_8,n63_9,);
not I_17(n38_9,n63_9);
nor I_18(n_431_5_r_9,G15_7_l_9,IN_7_7_l_9);
nor I_19(N3_8_r_9,n_102_5_r_9,n53_9);
nor I_20(n39_9,I_BUFF_1_9_r_9,n42_9);
not I_21(n40_9,n41_9);
nand I_22(n41_9,IN_1_1_l_9,IN_2_1_l_9);
nor I_23(n42_9,IN_9_7_l_9,IN_10_7_l_9);
nor I_24(n43_9,n63_9,n41_9);
nor I_25(n44_9,IN_5_7_l_9,IN_9_7_l_9);
and I_26(n45_9,IN_4_7_l_9,n52_9);
nor I_27(n46_9,n47_9,n48_9);
nor I_28(n47_9,n49_9,n50_9);
not I_29(n48_9,n_429_or_0_5_r_9);
not I_30(n49_9,n42_9);
or I_31(n50_9,n63_9,n51_9);
nor I_32(n51_9,IN_1_8_l_9,IN_3_8_l_9);
nor I_33(n52_9,G15_7_l_9,n49_9);
nor I_34(n53_9,n54_9,n55_9);
nor I_35(n54_9,G15_7_l_9,n56_9);
or I_36(n55_9,IN_10_7_l_9,n44_9);
not I_37(n56_9,IN_4_7_l_9);
nand I_38(n57_9,IN_2_8_l_9,IN_3_8_l_9);
nor I_39(n58_9,n62_9,n60_9);
nand I_40(n59_9,n51_9,n61_9);
nor I_41(n60_9,n38_9,n44_9);
nor I_42(n61_9,G18_7_l_9,IN_5_7_l_9);
nor I_43(N1371_0_r_8,n46_8,n51_8);
not I_44(N1508_0_r_8,n46_8);
nor I_45(N1372_1_r_8,n37_8,n49_8);
and I_46(N1508_1_r_8,N1372_1_r_8,n29_8);
nor I_47(N1507_6_r_8,n47_8,n48_8);
nor I_48(N1508_6_r_8,n37_8,n38_8);
nor I_49(n_42_8_r_8,I_BUFF_1_9_r_8,n53_8);
DFFARX1 I_50(N3_8_r_8,blif_clk_net_8_r_8,n8_8,G199_8_r_8,);
nor I_51(N6147_9_r_8,n29_8,n30_8);
nor I_52(N6134_9_r_8,n30_8,n31_8);
not I_53(I_BUFF_1_9_r_8,n35_8);
nor I_54(N1372_10_r_8,n46_8,n49_8);
nor I_55(N1508_10_r_8,n40_8,n41_8);
and I_56(N3_8_l_8,n36_8,n_576_5_r_9);
not I_57(n8_8,blif_reset_net_8_r_8);
DFFARX1 I_58(N3_8_l_8,blif_clk_net_8_r_8,n8_8,n53_8,);
not I_59(n29_8,n53_8);
nor I_60(N3_8_r_8,n33_8,n34_8);
and I_61(n30_8,n32_8,n33_8);
nor I_62(n31_8,n_42_8_r_9,N6147_2_r_9);
nand I_63(n32_8,n42_8,N1372_4_r_9);
or I_64(n33_8,n46_8,N1508_4_r_9);
nor I_65(n34_8,n32_8,n35_8);
nand I_66(n35_8,n44_8,n_547_5_r_9);
nand I_67(n36_8,N6134_9_r_9,N6147_2_r_9);
not I_68(n37_8,n31_8);
nand I_69(n38_8,N1508_0_r_8,n39_8);
nand I_70(n39_8,n33_8,n50_8);
and I_71(n40_8,n32_8,n35_8);
not I_72(n41_8,N1372_10_r_8);
and I_73(n42_8,n43_8,N6147_9_r_9);
nand I_74(n43_8,n44_8,n45_8);
nand I_75(n44_8,G78_5_r_9,n_576_5_r_9);
not I_76(n45_8,n_547_5_r_9);
nand I_77(n46_8,N1372_4_r_9,G78_5_r_9);
not I_78(n47_8,n39_8);
nor I_79(n48_8,n35_8,n49_8);
not I_80(n49_8,n51_8);
nand I_81(n50_8,I_BUFF_1_9_r_8,n51_8);
nor I_82(n51_8,n52_8,N1508_4_r_9);
or I_83(n52_8,N6147_2_r_9,G199_8_r_9);
endmodule


