module test_I13361(I8836,I1477,I1470,I13361);
input I8836,I1477,I1470;
output I13361;
wire I13313,I11672,I13197,I11293,I11310;
DFFARX1 I_0(I13313,I1470,I13197,,,I13361,);
DFFARX1 I_1(I11293,I1470,I13197,,,I13313,);
DFFARX1 I_2(I8836,I1470,I11310,,,I11672,);
not I_3(I13197,I1477);
not I_4(I11293,I11672);
not I_5(I11310,I1477);
endmodule


