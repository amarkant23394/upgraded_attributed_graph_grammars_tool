module test_I8827(I6893,I6992,I1477,I7026,I9114,I1470,I8827);
input I6893,I6992,I1477,I7026,I9114,I1470;
output I8827;
wire I9148,I9131,I9066,I9179,I8862,I9258,I8964,I6896;
and I_0(I9148,I8964,I9131);
nor I_1(I9131,I9066,I9114);
DFFARX1 I_2(I9258,I1470,I8862,,,I8827,);
DFFARX1 I_3(I1470,I8862,,,I9066,);
DFFARX1 I_4(I6896,I1470,I8862,,,I9179,);
not I_5(I8862,I1477);
or I_6(I9258,I9179,I9148);
not I_7(I8964,I6893);
nor I_8(I6896,I6992,I7026);
endmodule


