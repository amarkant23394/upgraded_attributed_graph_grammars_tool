module test_final(IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_6_2_l_10,IN_1_3_l_10,IN_2_3_l_10,IN_4_3_l_10,IN_1_4_l_10,IN_2_4_l_10,IN_3_4_l_10,IN_6_4_l_10,blif_clk_net_1_r_1,blif_reset_net_1_r_1,G42_1_r_1,n_572_1_r_1,n_573_1_r_1,n_549_1_r_1,n_452_1_r_1,ACVQN2_3_r_1,n_266_and_0_3_r_1,G199_4_r_1,G214_4_r_1);
input IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_6_2_l_10,IN_1_3_l_10,IN_2_3_l_10,IN_4_3_l_10,IN_1_4_l_10,IN_2_4_l_10,IN_3_4_l_10,IN_6_4_l_10,blif_clk_net_1_r_1,blif_reset_net_1_r_1;
output G42_1_r_1,n_572_1_r_1,n_573_1_r_1,n_549_1_r_1,n_452_1_r_1,ACVQN2_3_r_1,n_266_and_0_3_r_1,G199_4_r_1,G214_4_r_1;
wire G42_1_r_10,n_572_1_r_10,n_573_1_r_10,n_549_1_r_10,n_452_1_r_10,n_42_2_r_10,G199_2_r_10,ACVQN2_3_r_10,n_266_and_0_3_r_10,N3_2_l_10,n25_10,n16_10,n26_10,ACVQN1_3_l_10,N1_4_l_10,G199_4_l_10,n27_10,n17_10,n4_1_r_10,N3_2_r_10,n3_10,n13_internal_10,n13_10,n18_10,n19_10,n20_10,n21_10,n22_10,n23_10,n24_10,N3_2_l_1,n5_1,n26_1,n17_1,n16_internal_1,n16_1,ACVQN1_3_l_1,N1_4_l_1,G199_4_l_1,G214_4_l_1,n4_1_r_1,n14_internal_1,n14_1,N1_4_r_1,n18_1,n19_1,n20_1,n21_1,n22_1,n23_1,n24_1,n25_1;
DFFARX1 I_0(n4_1_r_10,blif_clk_net_1_r_1,n5_1,G42_1_r_10,);
nor I_1(n_572_1_r_10,n26_10,n3_10);
nand I_2(n_573_1_r_10,n16_10,n18_10);
nand I_3(n_549_1_r_10,n19_10,n20_10);
nor I_4(n_452_1_r_10,n25_10,n21_10);
nor I_5(n_42_2_r_10,n26_10,G199_4_l_10);
DFFARX1 I_6(N3_2_r_10,blif_clk_net_1_r_1,n5_1,G199_2_r_10,);
DFFARX1 I_7(G199_4_l_10,blif_clk_net_1_r_1,n5_1,ACVQN2_3_r_10,);
nor I_8(n_266_and_0_3_r_10,n17_10,n13_10);
and I_9(N3_2_l_10,IN_6_2_l_10,n23_10);
DFFARX1 I_10(N3_2_l_10,blif_clk_net_1_r_1,n5_1,n25_10,);
not I_11(n16_10,n25_10);
DFFARX1 I_12(IN_1_3_l_10,blif_clk_net_1_r_1,n5_1,n26_10,);
DFFARX1 I_13(IN_2_3_l_10,blif_clk_net_1_r_1,n5_1,ACVQN1_3_l_10,);
and I_14(N1_4_l_10,IN_6_4_l_10,n24_10);
DFFARX1 I_15(N1_4_l_10,blif_clk_net_1_r_1,n5_1,G199_4_l_10,);
DFFARX1 I_16(IN_3_4_l_10,blif_clk_net_1_r_1,n5_1,n27_10,);
not I_17(n17_10,n27_10);
nor I_18(n4_1_r_10,n27_10,n21_10);
nor I_19(N3_2_r_10,n16_10,n22_10);
not I_20(n3_10,n18_10);
DFFARX1 I_21(n3_10,blif_clk_net_1_r_1,n5_1,n13_internal_10,);
not I_22(n13_10,n13_internal_10);
nand I_23(n18_10,IN_4_3_l_10,ACVQN1_3_l_10);
not I_24(n19_10,n_452_1_r_10);
nand I_25(n20_10,n16_10,n26_10);
nor I_26(n21_10,IN_1_2_l_10,IN_3_2_l_10);
and I_27(n22_10,n26_10,n21_10);
nand I_28(n23_10,IN_2_2_l_10,IN_3_2_l_10);
nand I_29(n24_10,IN_1_4_l_10,IN_2_4_l_10);
DFFARX1 I_30(n4_1_r_1,blif_clk_net_1_r_1,n5_1,G42_1_r_1,);
nor I_31(n_572_1_r_1,n26_1,n19_1);
nand I_32(n_573_1_r_1,n16_1,n18_1);
nor I_33(n_549_1_r_1,n20_1,n21_1);
nor I_34(n_452_1_r_1,G214_4_l_1,n20_1);
DFFARX1 I_35(G199_4_l_1,blif_clk_net_1_r_1,n5_1,ACVQN2_3_r_1,);
nor I_36(n_266_and_0_3_r_1,n16_1,n14_1);
DFFARX1 I_37(N1_4_r_1,blif_clk_net_1_r_1,n5_1,G199_4_r_1,);
DFFARX1 I_38(G199_4_l_1,blif_clk_net_1_r_1,n5_1,G214_4_r_1,);
and I_39(N3_2_l_1,n23_1,n_266_and_0_3_r_10);
not I_40(n5_1,blif_reset_net_1_r_1);
DFFARX1 I_41(N3_2_l_1,blif_clk_net_1_r_1,n5_1,n26_1,);
not I_42(n17_1,n26_1);
DFFARX1 I_43(n_549_1_r_10,blif_clk_net_1_r_1,n5_1,n16_internal_1,);
not I_44(n16_1,n16_internal_1);
DFFARX1 I_45(n_573_1_r_10,blif_clk_net_1_r_1,n5_1,ACVQN1_3_l_1,);
and I_46(N1_4_l_1,n25_1,n_572_1_r_10);
DFFARX1 I_47(N1_4_l_1,blif_clk_net_1_r_1,n5_1,G199_4_l_1,);
DFFARX1 I_48(n_573_1_r_10,blif_clk_net_1_r_1,n5_1,G214_4_l_1,);
nor I_49(n4_1_r_1,n26_1,G214_4_l_1);
DFFARX1 I_50(G214_4_l_1,blif_clk_net_1_r_1,n5_1,n14_internal_1,);
not I_51(n14_1,n14_internal_1);
nor I_52(N1_4_r_1,n17_1,n24_1);
nand I_53(n18_1,ACVQN1_3_l_1,n_42_2_r_10);
nor I_54(n19_1,n_572_1_r_10,G199_2_r_10);
not I_55(n20_1,n18_1);
nor I_56(n21_1,n26_1,n22_1);
not I_57(n22_1,n19_1);
nand I_58(n23_1,n_572_1_r_10,G42_1_r_10);
nor I_59(n24_1,n18_1,n22_1);
nand I_60(n25_1,G42_1_r_10,ACVQN2_3_r_10);
endmodule


