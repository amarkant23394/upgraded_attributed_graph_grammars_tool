module test_final(IN_1_2_l_3,IN_2_2_l_3,IN_3_2_l_3,IN_4_2_l_3,IN_5_2_l_3,IN_1_6_l_3,IN_2_6_l_3,IN_3_6_l_3,IN_4_6_l_3,IN_5_6_l_3,IN_1_9_l_3,IN_2_9_l_3,IN_3_9_l_3,IN_4_9_l_3,IN_5_9_l_3,blif_clk_net_5_r_13,blif_reset_net_5_r_13,N1371_0_r_13,N1508_0_r_13,n_429_or_0_5_r_13,G78_5_r_13,n_576_5_r_13,n_547_5_r_13,G42_7_r_13,n_572_7_r_13,n_573_7_r_13,n_549_7_r_13,n_569_7_r_13,n_452_7_r_13);
input IN_1_2_l_3,IN_2_2_l_3,IN_3_2_l_3,IN_4_2_l_3,IN_5_2_l_3,IN_1_6_l_3,IN_2_6_l_3,IN_3_6_l_3,IN_4_6_l_3,IN_5_6_l_3,IN_1_9_l_3,IN_2_9_l_3,IN_3_9_l_3,IN_4_9_l_3,IN_5_9_l_3,blif_clk_net_5_r_13,blif_reset_net_5_r_13;
output N1371_0_r_13,N1508_0_r_13,n_429_or_0_5_r_13,G78_5_r_13,n_576_5_r_13,n_547_5_r_13,G42_7_r_13,n_572_7_r_13,n_573_7_r_13,n_549_7_r_13,n_569_7_r_13,n_452_7_r_13;
wire N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_572_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6147_9_r_3,N6134_9_r_3,I_BUFF_1_9_r_3,n4_7_r_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3,n40_3,n41_3,n42_3,n43_3,n44_3,n45_3,n46_3,n47_3,n48_3,n49_3,n50_3,n51_3,n_102_5_r_13,n4_7_l_13,n9_13,n62_13,n33_13,n_431_5_r_13,n1_13,n34_13,n35_13,n36_13,n37_13,n38_13,n39_13,n40_13,n41_13,n42_13,n43_13,n44_13,n45_13,n46_13,n47_13,n48_13,n49_13,n50_13,n51_13,n52_13,n53_13,n54_13,n55_13,n56_13,n57_13,n58_13,n59_13,n60_13,n61_13;
not I_0(N1372_1_r_3,n40_3);
nor I_1(N1508_1_r_3,N6147_9_r_3,n40_3);
nor I_2(N1507_6_r_3,n31_3,n42_3);
nor I_3(N1508_6_r_3,n30_3,n38_3);
DFFARX1 I_4(n4_7_r_3,blif_clk_net_5_r_13,n9_13,G42_7_r_3,);
nor I_5(n_572_7_r_3,I_BUFF_1_9_r_3,n35_3);
nand I_6(n_573_7_r_3,n30_3,n31_3);
nor I_7(n_549_7_r_3,N6147_9_r_3,n33_3);
nand I_8(n_569_7_r_3,n30_3,n32_3);
nor I_9(n_452_7_r_3,IN_1_9_l_3,n35_3);
not I_10(N6147_9_r_3,n32_3);
nor I_11(N6134_9_r_3,n36_3,n37_3);
not I_12(I_BUFF_1_9_r_3,n45_3);
nor I_13(n4_7_r_3,IN_1_9_l_3,I_BUFF_1_9_r_3);
not I_14(n30_3,n39_3);
not I_15(n31_3,n35_3);
nand I_16(n32_3,IN_5_6_l_3,n41_3);
nor I_17(n33_3,I_BUFF_1_9_r_3,n34_3);
nand I_18(n34_3,IN_2_6_l_3,n46_3);
nor I_19(n35_3,n43_3,n44_3);
not I_20(n36_3,n34_3);
nor I_21(n37_3,IN_1_9_l_3,N6147_9_r_3);
or I_22(n38_3,n_572_7_r_3,n34_3);
nor I_23(n39_3,IN_5_9_l_3,n44_3);
nand I_24(n40_3,IN_1_9_l_3,n39_3);
nand I_25(n41_3,IN_3_6_l_3,IN_4_6_l_3);
nor I_26(n42_3,n34_3,n45_3);
not I_27(n43_3,IN_2_9_l_3);
nor I_28(n44_3,IN_3_9_l_3,IN_4_9_l_3);
nand I_29(n45_3,n49_3,n50_3);
and I_30(n46_3,IN_1_6_l_3,n47_3);
nand I_31(n47_3,n41_3,n48_3);
not I_32(n48_3,IN_5_6_l_3);
nor I_33(n49_3,IN_1_2_l_3,IN_2_2_l_3);
or I_34(n50_3,IN_5_2_l_3,n51_3);
nor I_35(n51_3,IN_3_2_l_3,IN_4_2_l_3);
nor I_36(N1371_0_r_13,n59_13,n61_13);
nor I_37(N1508_0_r_13,n59_13,n60_13);
not I_38(n_429_or_0_5_r_13,n46_13);
DFFARX1 I_39(n_431_5_r_13,blif_clk_net_5_r_13,n9_13,G78_5_r_13,);
nand I_40(n_576_5_r_13,n_102_5_r_13,n34_13);
nor I_41(n_102_5_r_13,N1508_1_r_3,N1508_6_r_3);
nand I_42(n_547_5_r_13,n48_13,n49_13);
DFFARX1 I_43(n1_13,blif_clk_net_5_r_13,n9_13,G42_7_r_13,);
nor I_44(n_572_7_r_13,n40_13,n41_13);
nand I_45(n_573_7_r_13,n37_13,n38_13);
nor I_46(n_549_7_r_13,n46_13,n47_13);
nand I_47(n_569_7_r_13,n37_13,n43_13);
nand I_48(n_452_7_r_13,n52_13,n53_13);
nor I_49(n4_7_l_13,N1508_1_r_3,N1507_6_r_3);
not I_50(n9_13,blif_reset_net_5_r_13);
DFFARX1 I_51(n4_7_l_13,blif_clk_net_5_r_13,n9_13,n62_13,);
not I_52(n33_13,n62_13);
nand I_53(n_431_5_r_13,n54_13,n55_13);
not I_54(n1_13,n52_13);
nor I_55(n34_13,n35_13,n36_13);
nor I_56(n35_13,n42_13,G42_7_r_3);
nand I_57(n36_13,n50_13,n58_13);
nand I_58(n37_13,n44_13,n45_13);
or I_59(n38_13,n39_13,n_452_7_r_3);
nand I_60(n39_13,n_573_7_r_3,G42_7_r_3);
not I_61(n40_13,n36_13);
nor I_62(n41_13,n35_13,N1508_6_r_3);
not I_63(n42_13,n_569_7_r_3);
or I_64(n43_13,n_549_7_r_3,N1507_6_r_3);
not I_65(n44_13,G42_7_r_3);
not I_66(n45_13,N1372_1_r_3);
nor I_67(n46_13,n39_13,n40_13);
nor I_68(n47_13,n_549_7_r_3,N1507_6_r_3);
nor I_69(n48_13,n50_13,n51_13);
nor I_70(n49_13,G42_7_r_3,N1372_1_r_3);
not I_71(n50_13,n59_13);
not I_72(n51_13,n_102_5_r_13);
nand I_73(n52_13,n33_13,n39_13);
nand I_74(n53_13,n33_13,n_452_7_r_3);
nor I_75(n54_13,N1508_1_r_3,n_549_7_r_3);
nand I_76(n55_13,n62_13,n56_13);
nor I_77(n56_13,n39_13,n57_13);
not I_78(n57_13,N1507_6_r_3);
or I_79(n58_13,N1507_6_r_3,N1508_6_r_3);
nand I_80(n59_13,N1372_1_r_3,N6134_9_r_3);
nor I_81(n60_13,n51_13,n_549_7_r_3);
nor I_82(n61_13,n39_13,n_452_7_r_3);
endmodule


