module test_final(IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_4_2_l_10,IN_5_2_l_10,IN_1_6_l_10,IN_2_6_l_10,IN_3_6_l_10,IN_4_6_l_10,IN_5_6_l_10,IN_1_9_l_10,IN_2_9_l_10,IN_3_9_l_10,IN_4_9_l_10,IN_5_9_l_10,blif_clk_net_7_r_16,blif_reset_net_7_r_16,N1371_0_r_16,N1508_0_r_16,N1372_1_r_16,N1508_1_r_16,N6147_2_r_16,N1507_6_r_16,N1508_6_r_16,G42_7_r_16,n_572_7_r_16,n_573_7_r_16,n_569_7_r_16,n_452_7_r_16);
input IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_4_2_l_10,IN_5_2_l_10,IN_1_6_l_10,IN_2_6_l_10,IN_3_6_l_10,IN_4_6_l_10,IN_5_6_l_10,IN_1_9_l_10,IN_2_9_l_10,IN_3_9_l_10,IN_4_9_l_10,IN_5_9_l_10,blif_clk_net_7_r_16,blif_reset_net_7_r_16;
output N1371_0_r_16,N1508_0_r_16,N1372_1_r_16,N1508_1_r_16,N6147_2_r_16,N1507_6_r_16,N1508_6_r_16,G42_7_r_16,n_572_7_r_16,n_573_7_r_16,n_569_7_r_16,n_452_7_r_16;
wire N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1372_4_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10,I_BUFF_1_9_r_10,N3_8_r_10,n35_10,n36_10,n37_10,n38_10,n39_10,n40_10,n41_10,n42_10,n43_10,n44_10,n45_10,n46_10,n47_10,n48_10,n49_10,n50_10,n51_10,n52_10,n53_10,n54_10,n55_10,n56_10,n57_10,n58_10,n59_10,n60_10,n61_10,n62_10,n63_10,n64_10,n_549_7_r_16,N3_8_l_16,n8_16,n53_16,n29_16,n4_7_r_16,n30_16,n31_16,n32_16,n33_16,n34_16,n35_16,n36_16,n37_16,n38_16,n39_16,n40_16,n41_16,n42_16,n43_16,n44_16,n45_16,n46_16,n47_16,n48_16,n49_16,n50_16,n51_16,n52_16;
nor I_0(N1371_0_r_10,n37_10,n38_10);
nor I_1(N1508_0_r_10,n37_10,n58_10);
nand I_2(N6147_2_r_10,n39_10,n40_10);
not I_3(N6147_3_r_10,n39_10);
nor I_4(N1372_4_r_10,n46_10,n49_10);
nor I_5(N1508_4_r_10,n51_10,n52_10);
nor I_6(N1507_6_r_10,n49_10,n60_10);
nor I_7(N1508_6_r_10,n49_10,n50_10);
nor I_8(n_42_8_r_10,I_BUFF_1_9_r_10,n35_10);
DFFARX1 I_9(N3_8_r_10,blif_clk_net_7_r_16,n8_16,G199_8_r_10,);
nor I_10(N6147_9_r_10,n36_10,n37_10);
nor I_11(N6134_9_r_10,I_BUFF_1_9_r_10,n46_10);
not I_12(I_BUFF_1_9_r_10,n48_10);
nor I_13(N3_8_r_10,n44_10,n47_10);
not I_14(n35_10,n49_10);
nor I_15(n36_10,I_BUFF_1_9_r_10,n38_10);
not I_16(n37_10,IN_1_9_l_10);
not I_17(n38_10,n46_10);
nand I_18(n39_10,n43_10,n44_10);
nand I_19(n40_10,I_BUFF_1_9_r_10,n41_10);
nor I_20(n41_10,IN_1_9_l_10,n42_10);
not I_21(n42_10,n44_10);
nor I_22(n43_10,IN_1_9_l_10,n45_10);
nand I_23(n44_10,IN_2_6_l_10,n54_10);
nor I_24(n45_10,IN_5_9_l_10,n59_10);
nand I_25(n46_10,IN_2_9_l_10,n61_10);
nor I_26(n47_10,n46_10,n48_10);
nand I_27(n48_10,n62_10,n63_10);
nand I_28(n49_10,IN_5_6_l_10,n56_10);
not I_29(n50_10,n45_10);
nor I_30(n51_10,n42_10,n53_10);
not I_31(n52_10,N1372_4_r_10);
nor I_32(n53_10,n48_10,n50_10);
and I_33(n54_10,IN_1_6_l_10,n55_10);
nand I_34(n55_10,n56_10,n57_10);
nand I_35(n56_10,IN_3_6_l_10,IN_4_6_l_10);
not I_36(n57_10,IN_5_6_l_10);
nor I_37(n58_10,n35_10,n45_10);
nor I_38(n59_10,IN_3_9_l_10,IN_4_9_l_10);
nor I_39(n60_10,n37_10,n46_10);
or I_40(n61_10,IN_3_9_l_10,IN_4_9_l_10);
nor I_41(n62_10,IN_1_2_l_10,IN_2_2_l_10);
or I_42(n63_10,IN_5_2_l_10,n64_10);
nor I_43(n64_10,IN_3_2_l_10,IN_4_2_l_10);
nor I_44(N1371_0_r_16,n35_16,n39_16);
nor I_45(N1508_0_r_16,n39_16,n46_16);
not I_46(N1372_1_r_16,n45_16);
nor I_47(N1508_1_r_16,n53_16,n45_16);
nor I_48(N6147_2_r_16,n37_16,n38_16);
nor I_49(N1507_6_r_16,n44_16,n49_16);
nor I_50(N1508_6_r_16,n29_16,n42_16);
DFFARX1 I_51(n4_7_r_16,blif_clk_net_7_r_16,n8_16,G42_7_r_16,);
nor I_52(n_572_7_r_16,n32_16,n33_16);
nand I_53(n_573_7_r_16,n30_16,n31_16);
nand I_54(n_549_7_r_16,n47_16,N6147_3_r_10);
nand I_55(n_569_7_r_16,n_549_7_r_16,n30_16);
nor I_56(n_452_7_r_16,n34_16,n35_16);
and I_57(N3_8_l_16,n41_16,N1508_4_r_10);
not I_58(n8_16,blif_reset_net_7_r_16);
DFFARX1 I_59(N3_8_l_16,blif_clk_net_7_r_16,n8_16,n53_16,);
not I_60(n29_16,n53_16);
nor I_61(n4_7_r_16,n35_16,n36_16);
nand I_62(n30_16,N1508_0_r_10,N6147_2_r_10);
not I_63(n31_16,n34_16);
nor I_64(n32_16,n30_16,G199_8_r_10);
not I_65(n33_16,n_549_7_r_16);
nor I_66(n34_16,n48_16,N6147_3_r_10);
and I_67(n35_16,n50_16,N1507_6_r_10);
not I_68(n36_16,n30_16);
nor I_69(n37_16,n31_16,n40_16);
nand I_70(n38_16,n29_16,n39_16);
not I_71(n39_16,n32_16);
nor I_72(n40_16,N1508_6_r_10,N1508_0_r_10);
nand I_73(n41_16,N1371_0_r_10,N1508_0_r_10);
nand I_74(n42_16,n35_16,n43_16);
not I_75(n43_16,n44_16);
nor I_76(n44_16,n32_16,n49_16);
nand I_77(n45_16,n36_16,n40_16);
nor I_78(n46_16,n33_16,n34_16);
nand I_79(n47_16,N6134_9_r_10,N6147_2_r_10);
or I_80(n48_16,n_42_8_r_10,N6147_9_r_10);
and I_81(n49_16,n35_16,n36_16);
and I_82(n50_16,n51_16,N1371_0_r_10);
nand I_83(n51_16,n47_16,n52_16);
not I_84(n52_16,N6147_3_r_10);
endmodule


