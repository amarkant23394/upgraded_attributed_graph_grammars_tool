module test_I8428(I5864,I6045,I1477,I4518,I4533,I1470,I8428);
input I5864,I6045,I1477,I4518,I4533,I1470;
output I8428;
wire I8394,I6062,I5751,I5713,I6203,I8411,I5725,I6127,I6110,I5734,I6144;
not I_0(I8394,I5713);
and I_1(I8428,I8411,I5734);
and I_2(I6062,I5864,I6045);
not I_3(I5751,I1477);
DFFARX1 I_4(I6127,I1470,I5751,,,I5713,);
DFFARX1 I_5(I4518,I1470,I5751,,,I6203,);
nor I_6(I8411,I8394,I5725);
DFFARX1 I_7(I6203,I1470,I5751,,,I5725,);
and I_8(I6127,I6110,I4533);
DFFARX1 I_9(I1470,I5751,,,I6110,);
DFFARX1 I_10(I6144,I1470,I5751,,,I5734,);
or I_11(I6144,I6127,I6062);
endmodule


