module test_I16786(I12602,I15109,I1477,I1470,I16786);
input I12602,I15109,I1477,I1470;
output I16786;
wire I16934,I14945,I16818,I15126,I14965,I15372;
DFFARX1 I_0(I14945,I1470,I16818,,,I16934,);
nand I_1(I14945,I15372,I15126);
not I_2(I16818,I1477);
not I_3(I15126,I15109);
not I_4(I14965,I1477);
DFFARX1 I_5(I12602,I1470,I14965,,,I15372,);
DFFARX1 I_6(I16934,I1470,I16818,,,I16786,);
endmodule


