module test_final(IN_1_0_l_1,IN_2_0_l_1,IN_3_0_l_1,IN_4_0_l_1,IN_1_1_l_1,IN_2_1_l_1,IN_3_1_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_3_3_l_1,IN_1_6_l_1,IN_2_6_l_1,IN_3_6_l_1,IN_4_6_l_1,IN_5_6_l_1,blif_clk_net_5_r_15,blif_reset_net_5_r_15,N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15);
input IN_1_0_l_1,IN_2_0_l_1,IN_3_0_l_1,IN_4_0_l_1,IN_1_1_l_1,IN_2_1_l_1,IN_3_1_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_3_3_l_1,IN_1_6_l_1,IN_2_6_l_1,IN_3_6_l_1,IN_4_6_l_1,IN_5_6_l_1,blif_clk_net_5_r_15,blif_reset_net_5_r_15;
output N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15;
wire N1371_0_r_1,N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,n_452_7_r_1,N6147_9_r_1,N6134_9_r_1,I_BUFF_1_9_r_1,n4_7_r_1,n29_1,n30_1,n31_1,n32_1,n33_1,n34_1,n35_1,n36_1,n37_1,n38_1,n39_1,n40_1,n41_1,n42_1,n43_1,n44_1,n45_1,n46_1,n47_1,n48_1,n49_1,n50_1,n51_1,n52_1,n53_1,n54_1,n55_1,N1371_0_r_15,N1508_0_r_15,N1372_1_r_15,n_102_5_r_15,n_431_5_r_15,n9_15,n31_15,n32_15,n33_15,n34_15,n35_15,n36_15,n37_15,n38_15,n39_15,n40_15,n41_15,n42_15,n43_15,n44_15,n45_15,n46_15,n47_15,n48_15,n49_15,n50_15,n51_15,n52_15,n53_15,n54_15,n55_15;
and I_0(N1371_0_r_1,I_BUFF_1_9_r_1,n55_1);
nor I_1(N1508_0_r_1,n40_1,n44_1);
nor I_2(N1507_6_r_1,n43_1,n49_1);
nor I_3(N1508_6_r_1,n41_1,n42_1);
DFFARX1 I_4(n4_7_r_1,blif_clk_net_5_r_15,n9_15,G42_7_r_1,);
nor I_5(n_572_7_r_1,n29_1,n30_1);
not I_6(n_573_7_r_1,n_452_7_r_1);
nor I_7(n_549_7_r_1,N1371_0_r_1,n31_1);
or I_8(n_569_7_r_1,n30_1,n31_1);
nor I_9(n_452_7_r_1,n30_1,n32_1);
nor I_10(N6147_9_r_1,n35_1,n36_1);
nand I_11(N6134_9_r_1,n38_1,n39_1);
not I_12(I_BUFF_1_9_r_1,n40_1);
nor I_13(n4_7_r_1,I_BUFF_1_9_r_1,n30_1);
nor I_14(n29_1,IN_2_0_l_1,n34_1);
nor I_15(n30_1,n33_1,n34_1);
nor I_16(n31_1,IN_1_3_l_1,n54_1);
not I_17(n32_1,n48_1);
nor I_18(n33_1,IN_3_0_l_1,IN_4_0_l_1);
not I_19(n34_1,IN_1_0_l_1);
nor I_20(n35_1,I_BUFF_1_9_r_1,n37_1);
not I_21(n36_1,n29_1);
not I_22(n37_1,n41_1);
nand I_23(n38_1,IN_3_1_l_1,I_BUFF_1_9_r_1);
nand I_24(n39_1,n37_1,n40_1);
nand I_25(n40_1,IN_1_1_l_1,IN_2_1_l_1);
nand I_26(n41_1,IN_5_6_l_1,n52_1);
or I_27(n42_1,n36_1,n43_1);
nor I_28(n43_1,n32_1,n49_1);
nand I_29(n44_1,n45_1,n46_1);
nand I_30(n45_1,n47_1,n48_1);
not I_31(n46_1,IN_3_1_l_1);
not I_32(n47_1,n31_1);
nand I_33(n48_1,IN_2_6_l_1,n50_1);
nor I_34(n49_1,n41_1,n47_1);
and I_35(n50_1,IN_1_6_l_1,n51_1);
nand I_36(n51_1,n52_1,n53_1);
nand I_37(n52_1,IN_3_6_l_1,IN_4_6_l_1);
not I_38(n53_1,IN_5_6_l_1);
or I_39(n54_1,IN_2_3_l_1,IN_3_3_l_1);
nor I_40(n55_1,IN_3_1_l_1,n29_1);
and I_41(N1371_0_r_15,N1508_0_r_15,n_102_5_r_15);
nor I_42(N1508_0_r_15,n55_15,n_573_7_r_1);
nor I_43(N1372_1_r_15,n_102_5_r_15,n46_15);
nor I_44(N1508_1_r_15,N1508_0_r_15,n45_15);
not I_45(N1372_4_r_15,n39_15);
nor I_46(N1508_4_r_15,n39_15,n43_15);
nand I_47(n_429_or_0_5_r_15,n36_15,n38_15);
DFFARX1 I_48(n_431_5_r_15,blif_clk_net_5_r_15,n9_15,G78_5_r_15,);
nand I_49(n_576_5_r_15,n31_15,n32_15);
not I_50(n_102_5_r_15,n33_15);
nand I_51(n_547_5_r_15,N1371_0_r_15,n35_15);
nor I_52(N1507_6_r_15,n42_15,n46_15);
nand I_53(N1508_6_r_15,n39_15,n40_15);
nand I_54(n_431_5_r_15,n36_15,n37_15);
not I_55(n9_15,blif_reset_net_5_r_15);
nor I_56(n31_15,n33_15,n34_15);
nor I_57(n32_15,n44_15,n_569_7_r_1);
nor I_58(n33_15,n54_15,n55_15);
nand I_59(n34_15,n49_15,n_572_7_r_1);
nand I_60(n35_15,G42_7_r_1,n_549_7_r_1);
not I_61(n36_15,n32_15);
nand I_62(n37_15,n34_15,n38_15);
not I_63(n38_15,n46_15);
nand I_64(n39_15,n38_15,n41_15);
nand I_65(n40_15,n41_15,n42_15);
and I_66(n41_15,n51_15,N1508_0_r_1);
and I_67(n42_15,n47_15,G42_7_r_1);
and I_68(n43_15,n34_15,n36_15);
or I_69(n44_15,N1508_6_r_1,G42_7_r_1);
not I_70(n45_15,N1372_1_r_15);
nand I_71(n46_15,n53_15,G42_7_r_1);
nor I_72(n47_15,n34_15,n48_15);
not I_73(n48_15,n_549_7_r_1);
and I_74(n49_15,n50_15,N1507_6_r_1);
nand I_75(n50_15,n51_15,n52_15);
nand I_76(n51_15,N6134_9_r_1,n_573_7_r_1);
not I_77(n52_15,N1508_0_r_1);
nor I_78(n53_15,n48_15,N1508_0_r_1);
nor I_79(n54_15,N1507_6_r_1,n_572_7_r_1);
not I_80(n55_15,N6147_9_r_1);
endmodule


