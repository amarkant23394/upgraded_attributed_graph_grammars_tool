module test_final(G1_0_l_7,G2_0_l_7,IN_2_0_l_7,IN_4_0_l_7,IN_5_0_l_7,IN_7_0_l_7,IN_8_0_l_7,IN_10_0_l_7,IN_11_0_l_7,IN_1_5_l_7,IN_2_5_l_7,blif_clk_net_1_r_2,blif_reset_net_1_r_2,G42_1_r_2,n_572_1_r_2,n_549_1_r_2,n_569_1_r_2,n_452_1_r_2,n_42_2_r_2,G199_2_r_2,ACVQN1_5_r_2,P6_5_r_2);
input G1_0_l_7,G2_0_l_7,IN_2_0_l_7,IN_4_0_l_7,IN_5_0_l_7,IN_7_0_l_7,IN_8_0_l_7,IN_10_0_l_7,IN_11_0_l_7,IN_1_5_l_7,IN_2_5_l_7,blif_clk_net_1_r_2,blif_reset_net_1_r_2;
output G42_1_r_2,n_572_1_r_2,n_549_1_r_2,n_569_1_r_2,n_452_1_r_2,n_42_2_r_2,G199_2_r_2,ACVQN1_5_r_2,P6_5_r_2;
wire G42_1_r_7,n_572_1_r_7,n_573_1_r_7,n_549_1_r_7,n_569_1_r_7,G199_4_r_7,G214_4_r_7,ACVQN1_5_r_7,P6_5_r_7,n_431_0_l_7,n43_7,n27_7,ACVQN1_5_l_7,n44_7,n4_1_r_7,N1_4_r_7,n26_7,n5_7,P6_5_r_internal_7,n28_7,n29_7,n30_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7,n_573_1_r_2,N3_2_l_2,n5_2,G199_2_l_2,n13_2,ACVQN2_3_l_2,n16_2,N1_4_l_2,n26_2,n17_internal_2,n17_2,n4_1_r_2,N3_2_r_2,P6_5_r_internal_2,n18_2,n19_2,n20_2,n21_2,n22_2,n23_2,n24_2,n25_2;
DFFARX1 I_0(n4_1_r_7,blif_clk_net_1_r_2,n5_2,G42_1_r_7,);
nor I_1(n_572_1_r_7,n30_7,n31_7);
nand I_2(n_573_1_r_7,IN_7_0_l_7,n28_7);
nor I_3(n_549_1_r_7,ACVQN1_5_l_7,n35_7);
nand I_4(n_569_1_r_7,n32_7,n33_7);
DFFARX1 I_5(N1_4_r_7,blif_clk_net_1_r_2,n5_2,G199_4_r_7,);
DFFARX1 I_6(n26_7,blif_clk_net_1_r_2,n5_2,G214_4_r_7,);
DFFARX1 I_7(n5_7,blif_clk_net_1_r_2,n5_2,ACVQN1_5_r_7,);
not I_8(P6_5_r_7,P6_5_r_internal_7);
or I_9(n_431_0_l_7,IN_8_0_l_7,n36_7);
DFFARX1 I_10(n_431_0_l_7,blif_clk_net_1_r_2,n5_2,n43_7,);
not I_11(n27_7,n43_7);
DFFARX1 I_12(IN_2_5_l_7,blif_clk_net_1_r_2,n5_2,ACVQN1_5_l_7,);
DFFARX1 I_13(IN_1_5_l_7,blif_clk_net_1_r_2,n5_2,n44_7,);
nor I_14(n4_1_r_7,n30_7,n38_7);
nor I_15(N1_4_r_7,n27_7,n40_7);
nand I_16(n26_7,IN_11_0_l_7,n39_7);
not I_17(n5_7,G2_0_l_7);
DFFARX1 I_18(ACVQN1_5_l_7,blif_clk_net_1_r_2,n5_2,P6_5_r_internal_7,);
nor I_19(n28_7,n26_7,n29_7);
not I_20(n29_7,IN_5_0_l_7);
not I_21(n30_7,G1_0_l_7);
nand I_22(n31_7,n27_7,n29_7);
nor I_23(n32_7,ACVQN1_5_l_7,n34_7);
nor I_24(n33_7,G2_0_l_7,n29_7);
not I_25(n34_7,IN_7_0_l_7);
nor I_26(n35_7,n43_7,n44_7);
and I_27(n36_7,IN_2_0_l_7,n37_7);
nor I_28(n37_7,IN_4_0_l_7,n30_7);
nand I_29(n38_7,G2_0_l_7,n29_7);
nor I_30(n39_7,G2_0_l_7,IN_10_0_l_7);
nor I_31(n40_7,n44_7,n41_7);
nor I_32(n41_7,n34_7,n42_7);
nand I_33(n42_7,IN_5_0_l_7,n5_7);
DFFARX1 I_34(n4_1_r_2,blif_clk_net_1_r_2,n5_2,G42_1_r_2,);
nor I_35(n_572_1_r_2,n26_2,n18_2);
nand I_36(n_573_1_r_2,n17_2,n19_2);
nor I_37(n_549_1_r_2,G199_2_l_2,n20_2);
nand I_38(n_569_1_r_2,n13_2,n19_2);
not I_39(n_452_1_r_2,n_573_1_r_2);
nor I_40(n_42_2_r_2,ACVQN2_3_l_2,n18_2);
DFFARX1 I_41(N3_2_r_2,blif_clk_net_1_r_2,n5_2,G199_2_r_2,);
DFFARX1 I_42(ACVQN2_3_l_2,blif_clk_net_1_r_2,n5_2,ACVQN1_5_r_2,);
not I_43(P6_5_r_2,P6_5_r_internal_2);
and I_44(N3_2_l_2,n24_2,G214_4_r_7);
not I_45(n5_2,blif_reset_net_1_r_2);
DFFARX1 I_46(N3_2_l_2,blif_clk_net_1_r_2,n5_2,G199_2_l_2,);
not I_47(n13_2,G199_2_l_2);
DFFARX1 I_48(G42_1_r_7,blif_clk_net_1_r_2,n5_2,ACVQN2_3_l_2,);
DFFARX1 I_49(G199_4_r_7,blif_clk_net_1_r_2,n5_2,n16_2,);
and I_50(N1_4_l_2,n25_2,n_549_1_r_7);
DFFARX1 I_51(N1_4_l_2,blif_clk_net_1_r_2,n5_2,n26_2,);
DFFARX1 I_52(ACVQN1_5_r_7,blif_clk_net_1_r_2,n5_2,n17_internal_2,);
not I_53(n17_2,n17_internal_2);
nor I_54(n4_1_r_2,n26_2,n22_2);
nor I_55(N3_2_r_2,n17_2,n23_2);
DFFARX1 I_56(G199_2_l_2,blif_clk_net_1_r_2,n5_2,P6_5_r_internal_2,);
nor I_57(n18_2,n_572_1_r_7,n_569_1_r_7);
nand I_58(n19_2,n16_2,n_572_1_r_7);
nor I_59(n20_2,n26_2,n21_2);
not I_60(n21_2,n18_2);
and I_61(n22_2,n16_2,n_572_1_r_7);
nor I_62(n23_2,n13_2,n21_2);
nand I_63(n24_2,n_572_1_r_7,n_573_1_r_7);
nand I_64(n25_2,G42_1_r_7,P6_5_r_7);
endmodule


