module test_final(IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_6_2_l_6,IN_1_3_l_6,IN_2_3_l_6,IN_4_3_l_6,IN_1_4_l_6,IN_2_4_l_6,IN_3_4_l_6,IN_6_4_l_6,blif_clk_net_1_r_3,blif_reset_net_1_r_3,G42_1_r_3,n_572_1_r_3,n_573_1_r_3,n_549_1_r_3,n_569_1_r_3,n_452_1_r_3,n_42_2_r_3,G199_2_r_3,ACVQN2_3_r_3,n_266_and_0_3_r_3);
input IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_6_2_l_6,IN_1_3_l_6,IN_2_3_l_6,IN_4_3_l_6,IN_1_4_l_6,IN_2_4_l_6,IN_3_4_l_6,IN_6_4_l_6,blif_clk_net_1_r_3,blif_reset_net_1_r_3;
output G42_1_r_3,n_572_1_r_3,n_573_1_r_3,n_549_1_r_3,n_569_1_r_3,n_452_1_r_3,n_42_2_r_3,G199_2_r_3,ACVQN2_3_r_3,n_266_and_0_3_r_3;
wire G42_1_r_6,n_572_1_r_6,n_573_1_r_6,n_549_1_r_6,n_569_1_r_6,n_452_1_r_6,G199_4_r_6,G214_4_r_6,ACVQN1_5_r_6,P6_5_r_6,N3_2_l_6,n27_6,n17_6,n28_6,n26_6,N1_4_l_6,n29_6,n18_6,G214_4_l_6,n12_6,n4_1_r_6,N1_4_r_6,n_42_2_l_6,P6_5_r_internal_6,n19_6,n20_6,n21_6,n22_6,n23_6,n24_6,n25_6,n4_1_l_3,n9_3,G42_1_l_3,n22_3,n40_3,n25_internal_3,n25_3,n4_1_r_3,N3_2_r_3,n_572_1_l_3,ACVQN1_3_r_3,n26_3,n27_3,n28_3,n29_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3;
DFFARX1 I_0(n4_1_r_6,blif_clk_net_1_r_3,n9_3,G42_1_r_6,);
nor I_1(n_572_1_r_6,n27_6,n28_6);
nand I_2(n_573_1_r_6,n18_6,n19_6);
nor I_3(n_549_1_r_6,n_42_2_l_6,n21_6);
nand I_4(n_569_1_r_6,n19_6,n20_6);
nor I_5(n_452_1_r_6,n28_6,n29_6);
DFFARX1 I_6(N1_4_r_6,blif_clk_net_1_r_3,n9_3,G199_4_r_6,);
DFFARX1 I_7(n_42_2_l_6,blif_clk_net_1_r_3,n9_3,G214_4_r_6,);
DFFARX1 I_8(n_42_2_l_6,blif_clk_net_1_r_3,n9_3,ACVQN1_5_r_6,);
not I_9(P6_5_r_6,P6_5_r_internal_6);
and I_10(N3_2_l_6,IN_6_2_l_6,n23_6);
DFFARX1 I_11(N3_2_l_6,blif_clk_net_1_r_3,n9_3,n27_6,);
not I_12(n17_6,n27_6);
DFFARX1 I_13(IN_1_3_l_6,blif_clk_net_1_r_3,n9_3,n28_6,);
DFFARX1 I_14(IN_2_3_l_6,blif_clk_net_1_r_3,n9_3,n26_6,);
and I_15(N1_4_l_6,IN_6_4_l_6,n25_6);
DFFARX1 I_16(N1_4_l_6,blif_clk_net_1_r_3,n9_3,n29_6,);
not I_17(n18_6,n29_6);
DFFARX1 I_18(IN_3_4_l_6,blif_clk_net_1_r_3,n9_3,G214_4_l_6,);
not I_19(n12_6,G214_4_l_6);
nor I_20(n4_1_r_6,n28_6,n22_6);
nor I_21(N1_4_r_6,n12_6,n24_6);
nor I_22(n_42_2_l_6,IN_1_2_l_6,IN_3_2_l_6);
DFFARX1 I_23(G214_4_l_6,blif_clk_net_1_r_3,n9_3,P6_5_r_internal_6,);
nand I_24(n19_6,IN_4_3_l_6,n26_6);
not I_25(n20_6,n_42_2_l_6);
nor I_26(n21_6,n17_6,n28_6);
and I_27(n22_6,IN_4_3_l_6,n26_6);
nand I_28(n23_6,IN_2_2_l_6,IN_3_2_l_6);
nor I_29(n24_6,n17_6,n18_6);
nand I_30(n25_6,IN_1_4_l_6,IN_2_4_l_6);
DFFARX1 I_31(n4_1_r_3,blif_clk_net_1_r_3,n9_3,G42_1_r_3,);
nor I_32(n_572_1_r_3,G42_1_l_3,n28_3);
nand I_33(n_573_1_r_3,n26_3,n27_3);
nor I_34(n_549_1_r_3,n40_3,n32_3);
nand I_35(n_569_1_r_3,n27_3,n31_3);
and I_36(n_452_1_r_3,n26_3,P6_5_r_6);
nor I_37(n_42_2_r_3,n_572_1_l_3,n34_3);
DFFARX1 I_38(N3_2_r_3,blif_clk_net_1_r_3,n9_3,G199_2_r_3,);
DFFARX1 I_39(n_572_1_l_3,blif_clk_net_1_r_3,n9_3,ACVQN2_3_r_3,);
nor I_40(n_266_and_0_3_r_3,n25_3,n35_3);
nor I_41(n4_1_l_3,n_573_1_r_6,P6_5_r_6);
not I_42(n9_3,blif_reset_net_1_r_3);
DFFARX1 I_43(n4_1_l_3,blif_clk_net_1_r_3,n9_3,G42_1_l_3,);
not I_44(n22_3,G42_1_l_3);
DFFARX1 I_45(G42_1_r_6,blif_clk_net_1_r_3,n9_3,n40_3,);
DFFARX1 I_46(G42_1_r_6,blif_clk_net_1_r_3,n9_3,n25_internal_3,);
not I_47(n25_3,n25_internal_3);
nor I_48(n4_1_r_3,n40_3,n36_3);
nor I_49(N3_2_r_3,n26_3,n37_3);
nor I_50(n_572_1_l_3,n_569_1_r_6,G214_4_r_6);
DFFARX1 I_51(G42_1_l_3,blif_clk_net_1_r_3,n9_3,ACVQN1_3_r_3,);
nor I_52(n26_3,n_572_1_r_6,n_452_1_r_6);
not I_53(n27_3,n_549_1_r_6);
nor I_54(n28_3,n29_3,n_549_1_r_6);
nor I_55(n29_3,n30_3,G214_4_r_6);
not I_56(n30_3,ACVQN1_5_r_6);
nor I_57(n31_3,n40_3,n_572_1_r_6);
nor I_58(n32_3,n25_3,n33_3);
nand I_59(n33_3,n22_3,G199_4_r_6);
or I_60(n34_3,n_572_1_r_6,n_549_1_r_6);
nand I_61(n35_3,ACVQN1_3_r_3,G199_4_r_6);
nor I_62(n36_3,n_452_1_r_6,P6_5_r_6);
nor I_63(n37_3,n38_3,n39_3);
not I_64(n38_3,n_572_1_l_3);
nand I_65(n39_3,n27_3,n30_3);
endmodule


