module test_I6265(I2167,I1477,I2173,I1470,I4578,I6265);
input I2167,I1477,I2173,I1470,I4578;
output I6265;
wire I4629,I6248,I5864,I5751,I6203,I4595,I4518,I4527,I4536,I4515,I4544,I4869,I5915,I4691;
nor I_0(I4629,I2167,I2173);
and I_1(I6265,I5915,I6248);
nand I_2(I6248,I6203,I5864);
nor I_3(I5864,I4536,I4515);
not I_4(I5751,I1477);
DFFARX1 I_5(I4518,I1470,I5751,,,I6203,);
DFFARX1 I_6(I4578,I1470,I4544,,,I4595,);
nand I_7(I4518,I4869,I4691);
or I_8(I4527,I4629,I4595);
nor I_9(I4536,I4869,I4595);
not I_10(I4515,I4629);
not I_11(I4544,I1477);
DFFARX1 I_12(I1470,I4544,,,I4869,);
DFFARX1 I_13(I4527,I1470,I5751,,,I5915,);
nor I_14(I4691,I4629);
endmodule


