module test_final(G1_0_l_17,G2_0_l_17,IN_2_0_l_17,IN_4_0_l_17,IN_5_0_l_17,IN_7_0_l_17,IN_8_0_l_17,IN_10_0_l_17,IN_11_0_l_17,IN_1_5_l_17,IN_2_5_l_17,blif_clk_net_1_r_4,blif_reset_net_1_r_4,G42_1_r_4,n_572_1_r_4,n_573_1_r_4,n_549_1_r_4,n_569_1_r_4,ACVQN2_3_r_4,n_266_and_0_3_r_4,ACVQN1_5_r_4,P6_5_r_4);
input G1_0_l_17,G2_0_l_17,IN_2_0_l_17,IN_4_0_l_17,IN_5_0_l_17,IN_7_0_l_17,IN_8_0_l_17,IN_10_0_l_17,IN_11_0_l_17,IN_1_5_l_17,IN_2_5_l_17,blif_clk_net_1_r_4,blif_reset_net_1_r_4;
output G42_1_r_4,n_572_1_r_4,n_573_1_r_4,n_549_1_r_4,n_569_1_r_4,ACVQN2_3_r_4,n_266_and_0_3_r_4,ACVQN1_5_r_4,P6_5_r_4;
wire G42_1_r_17,n_572_1_r_17,n_573_1_r_17,n_549_1_r_17,n_569_1_r_17,n_452_1_r_17,ACVQN2_3_r_17,n_266_and_0_3_r_17,G199_4_r_17,G214_4_r_17,n_431_0_l_17,n20_internal_17,n20_17,ACVQN1_5_l_17,n19_internal_17,n19_17,n4_1_r_17,n2_17,n17_internal_17,n17_17,N1_4_r_17,n5_17,n21_17,n22_17,n23_17,n24_17,n25_17,n26_17,n27_17,n28_17,n29_17,n30_17,n31_17,n32_17,n_431_0_l_4,n6_4,G78_0_l_4,ACVQN1_5_l_4,n16_4,n17_internal_4,n17_4,n4_1_r_4,n19_4,n15_internal_4,n15_4,P6_5_r_internal_4,n20_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4;
DFFARX1 I_0(n4_1_r_17,blif_clk_net_1_r_4,n6_4,G42_1_r_17,);
nor I_1(n_572_1_r_17,ACVQN1_5_l_17,n19_17);
nand I_2(n_573_1_r_17,n20_17,n21_17);
nand I_3(n_549_1_r_17,n23_17,n24_17);
nand I_4(n_569_1_r_17,n21_17,n22_17);
not I_5(n_452_1_r_17,n23_17);
DFFARX1 I_6(n19_17,blif_clk_net_1_r_4,n6_4,ACVQN2_3_r_17,);
nor I_7(n_266_and_0_3_r_17,n17_17,n29_17);
DFFARX1 I_8(N1_4_r_17,blif_clk_net_1_r_4,n6_4,G199_4_r_17,);
DFFARX1 I_9(n5_17,blif_clk_net_1_r_4,n6_4,G214_4_r_17,);
or I_10(n_431_0_l_17,IN_8_0_l_17,n26_17);
DFFARX1 I_11(n_431_0_l_17,blif_clk_net_1_r_4,n6_4,n20_internal_17,);
not I_12(n20_17,n20_internal_17);
DFFARX1 I_13(IN_2_5_l_17,blif_clk_net_1_r_4,n6_4,ACVQN1_5_l_17,);
DFFARX1 I_14(IN_1_5_l_17,blif_clk_net_1_r_4,n6_4,n19_internal_17,);
not I_15(n19_17,n19_internal_17);
nor I_16(n4_1_r_17,n5_17,n25_17);
not I_17(n2_17,n29_17);
DFFARX1 I_18(n2_17,blif_clk_net_1_r_4,n6_4,n17_internal_17,);
not I_19(n17_17,n17_internal_17);
nor I_20(N1_4_r_17,n29_17,n31_17);
not I_21(n5_17,G2_0_l_17);
and I_22(n21_17,IN_11_0_l_17,n32_17);
not I_23(n22_17,n25_17);
nand I_24(n23_17,n20_17,n22_17);
nand I_25(n24_17,n19_17,n22_17);
nand I_26(n25_17,IN_7_0_l_17,n30_17);
and I_27(n26_17,IN_2_0_l_17,n27_17);
nor I_28(n27_17,IN_4_0_l_17,n28_17);
not I_29(n28_17,G1_0_l_17);
nor I_30(n29_17,IN_5_0_l_17,n28_17);
and I_31(n30_17,IN_5_0_l_17,n5_17);
nor I_32(n31_17,G2_0_l_17,n21_17);
nor I_33(n32_17,G2_0_l_17,IN_10_0_l_17);
DFFARX1 I_34(n4_1_r_4,blif_clk_net_1_r_4,n6_4,G42_1_r_4,);
nor I_35(n_572_1_r_4,G78_0_l_4,n17_4);
nand I_36(n_573_1_r_4,n16_4,ACVQN2_3_r_17);
nor I_37(n_549_1_r_4,n22_4,n23_4);
nand I_38(n_569_1_r_4,n20_4,n21_4);
DFFARX1 I_39(n19_4,blif_clk_net_1_r_4,n6_4,ACVQN2_3_r_4,);
nor I_40(n_266_and_0_3_r_4,n15_4,n29_4);
DFFARX1 I_41(n19_4,blif_clk_net_1_r_4,n6_4,ACVQN1_5_r_4,);
not I_42(P6_5_r_4,P6_5_r_internal_4);
or I_43(n_431_0_l_4,n26_4,n_266_and_0_3_r_17);
not I_44(n6_4,blif_reset_net_1_r_4);
DFFARX1 I_45(n_431_0_l_4,blif_clk_net_1_r_4,n6_4,G78_0_l_4,);
DFFARX1 I_46(n_572_1_r_17,blif_clk_net_1_r_4,n6_4,ACVQN1_5_l_4,);
not I_47(n16_4,ACVQN1_5_l_4);
DFFARX1 I_48(n_573_1_r_17,blif_clk_net_1_r_4,n6_4,n17_internal_4,);
not I_49(n17_4,n17_internal_4);
nor I_50(n4_1_r_4,n30_4,n31_4);
nand I_51(n19_4,n33_4,G199_4_r_17);
DFFARX1 I_52(G78_0_l_4,blif_clk_net_1_r_4,n6_4,n15_internal_4,);
not I_53(n15_4,n15_internal_4);
DFFARX1 I_54(ACVQN1_5_l_4,blif_clk_net_1_r_4,n6_4,P6_5_r_internal_4,);
and I_55(n20_4,n16_4,n_452_1_r_17);
nor I_56(n21_4,ACVQN2_3_r_17,G214_4_r_17);
nand I_57(n22_4,G78_0_l_4,n25_4);
nand I_58(n23_4,n24_4,n_452_1_r_17);
not I_59(n24_4,ACVQN2_3_r_17);
not I_60(n25_4,G214_4_r_17);
and I_61(n26_4,n27_4,n_549_1_r_17);
nor I_62(n27_4,n28_4,n_569_1_r_17);
not I_63(n28_4,G199_4_r_17);
not I_64(n29_4,n30_4);
nand I_65(n30_4,n32_4,G42_1_r_17);
nand I_66(n31_4,n25_4,n_452_1_r_17);
nor I_67(n32_4,n33_4,ACVQN2_3_r_17);
not I_68(n33_4,G42_1_r_17);
endmodule


