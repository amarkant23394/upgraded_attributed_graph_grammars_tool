module test_I14957(I12947,I1477,I14982,I15177,I1470,I14957);
input I12947,I1477,I14982,I15177,I1470;
output I14957;
wire I12670,I15064,I14965,I15485,I13023,I12608,I15194,I12587,I12619,I12605,I15047,I15211,I15228,I12584,I15502;
DFFARX1 I_0(I1470,I12619,,,I12670,);
nand I_1(I15064,I15047,I12587);
not I_2(I14965,I1477);
DFFARX1 I_3(I12605,I1470,I14965,,,I15485,);
DFFARX1 I_4(I1470,I12619,,,I13023,);
nor I_5(I12608,I13023);
or I_6(I15194,I15177,I12608);
DFFARX1 I_7(I12670,I1470,I12619,,,I12587,);
nand I_8(I14957,I15502,I15228);
not I_9(I12619,I1477);
nand I_10(I12605,I13023,I12947);
nor I_11(I15047,I14982,I12584);
DFFARX1 I_12(I15194,I1470,I14965,,,I15211,);
nor I_13(I15228,I15211,I15064);
and I_14(I12584,I12670);
not I_15(I15502,I15485);
endmodule


