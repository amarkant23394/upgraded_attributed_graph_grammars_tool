module test_I11624(I9131,I8896,I1477,I8964,I1470,I6878,I6896,I11624);
input I9131,I8896,I1477,I8964,I1470,I6878,I6896;
output I11624;
wire I9148,I8830,I8827,I8913,I8981,I8862,I9227,I9179,I9258,I11327;
and I_0(I9148,I8964,I9131);
nand I_1(I8830,I8913,I9227);
DFFARX1 I_2(I9258,I1470,I8862,,,I8827,);
nand I_3(I8913,I8896,I6878);
not I_4(I8981,I8964);
not I_5(I8862,I1477);
nor I_6(I9227,I9179,I8981);
DFFARX1 I_7(I6896,I1470,I8862,,,I9179,);
or I_8(I9258,I9179,I9148);
not I_9(I11327,I8830);
nand I_10(I11624,I11327,I8827);
endmodule


