module test_I17413_rst(I1477_rst,I17413_rst);
,I17413_rst);
input I1477_rst;
output I17413_rst;
wire ;
not I_0(I17413_rst,I1477_rst);
endmodule


