module test_final(IN_1_2_l_3,IN_2_2_l_3,IN_3_2_l_3,IN_4_2_l_3,IN_5_2_l_3,IN_1_6_l_3,IN_2_6_l_3,IN_3_6_l_3,IN_4_6_l_3,IN_5_6_l_3,IN_1_9_l_3,IN_2_9_l_3,IN_3_9_l_3,IN_4_9_l_3,IN_5_9_l_3,blif_clk_net_5_r_15,blif_reset_net_5_r_15,N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15);
input IN_1_2_l_3,IN_2_2_l_3,IN_3_2_l_3,IN_4_2_l_3,IN_5_2_l_3,IN_1_6_l_3,IN_2_6_l_3,IN_3_6_l_3,IN_4_6_l_3,IN_5_6_l_3,IN_1_9_l_3,IN_2_9_l_3,IN_3_9_l_3,IN_4_9_l_3,IN_5_9_l_3,blif_clk_net_5_r_15,blif_reset_net_5_r_15;
output N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15;
wire N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_572_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6147_9_r_3,N6134_9_r_3,I_BUFF_1_9_r_3,n4_7_r_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3,n40_3,n41_3,n42_3,n43_3,n44_3,n45_3,n46_3,n47_3,n48_3,n49_3,n50_3,n51_3,N1371_0_r_15,N1508_0_r_15,N1372_1_r_15,n_102_5_r_15,n_431_5_r_15,n9_15,n31_15,n32_15,n33_15,n34_15,n35_15,n36_15,n37_15,n38_15,n39_15,n40_15,n41_15,n42_15,n43_15,n44_15,n45_15,n46_15,n47_15,n48_15,n49_15,n50_15,n51_15,n52_15,n53_15,n54_15,n55_15;
not I_0(N1372_1_r_3,n40_3);
nor I_1(N1508_1_r_3,N6147_9_r_3,n40_3);
nor I_2(N1507_6_r_3,n31_3,n42_3);
nor I_3(N1508_6_r_3,n30_3,n38_3);
DFFARX1 I_4(n4_7_r_3,blif_clk_net_5_r_15,n9_15,G42_7_r_3,);
nor I_5(n_572_7_r_3,I_BUFF_1_9_r_3,n35_3);
nand I_6(n_573_7_r_3,n30_3,n31_3);
nor I_7(n_549_7_r_3,N6147_9_r_3,n33_3);
nand I_8(n_569_7_r_3,n30_3,n32_3);
nor I_9(n_452_7_r_3,IN_1_9_l_3,n35_3);
not I_10(N6147_9_r_3,n32_3);
nor I_11(N6134_9_r_3,n36_3,n37_3);
not I_12(I_BUFF_1_9_r_3,n45_3);
nor I_13(n4_7_r_3,IN_1_9_l_3,I_BUFF_1_9_r_3);
not I_14(n30_3,n39_3);
not I_15(n31_3,n35_3);
nand I_16(n32_3,IN_5_6_l_3,n41_3);
nor I_17(n33_3,I_BUFF_1_9_r_3,n34_3);
nand I_18(n34_3,IN_2_6_l_3,n46_3);
nor I_19(n35_3,n43_3,n44_3);
not I_20(n36_3,n34_3);
nor I_21(n37_3,IN_1_9_l_3,N6147_9_r_3);
or I_22(n38_3,n_572_7_r_3,n34_3);
nor I_23(n39_3,IN_5_9_l_3,n44_3);
nand I_24(n40_3,IN_1_9_l_3,n39_3);
nand I_25(n41_3,IN_3_6_l_3,IN_4_6_l_3);
nor I_26(n42_3,n34_3,n45_3);
not I_27(n43_3,IN_2_9_l_3);
nor I_28(n44_3,IN_3_9_l_3,IN_4_9_l_3);
nand I_29(n45_3,n49_3,n50_3);
and I_30(n46_3,IN_1_6_l_3,n47_3);
nand I_31(n47_3,n41_3,n48_3);
not I_32(n48_3,IN_5_6_l_3);
nor I_33(n49_3,IN_1_2_l_3,IN_2_2_l_3);
or I_34(n50_3,IN_5_2_l_3,n51_3);
nor I_35(n51_3,IN_3_2_l_3,IN_4_2_l_3);
and I_36(N1371_0_r_15,N1508_0_r_15,n_102_5_r_15);
nor I_37(N1508_0_r_15,n55_15,N1508_6_r_3);
nor I_38(N1372_1_r_15,n_102_5_r_15,n46_15);
nor I_39(N1508_1_r_15,N1508_0_r_15,n45_15);
not I_40(N1372_4_r_15,n39_15);
nor I_41(N1508_4_r_15,n39_15,n43_15);
nand I_42(n_429_or_0_5_r_15,n36_15,n38_15);
DFFARX1 I_43(n_431_5_r_15,blif_clk_net_5_r_15,n9_15,G78_5_r_15,);
nand I_44(n_576_5_r_15,n31_15,n32_15);
not I_45(n_102_5_r_15,n33_15);
nand I_46(n_547_5_r_15,N1371_0_r_15,n35_15);
nor I_47(N1507_6_r_15,n42_15,n46_15);
nand I_48(N1508_6_r_15,n39_15,n40_15);
nand I_49(n_431_5_r_15,n36_15,n37_15);
not I_50(n9_15,blif_reset_net_5_r_15);
nor I_51(n31_15,n33_15,n34_15);
nor I_52(n32_15,n44_15,n_573_7_r_3);
nor I_53(n33_15,n54_15,n55_15);
nand I_54(n34_15,n49_15,N6134_9_r_3);
nand I_55(n35_15,N1507_6_r_3,n_573_7_r_3);
not I_56(n36_15,n32_15);
nand I_57(n37_15,n34_15,n38_15);
not I_58(n38_15,n46_15);
nand I_59(n39_15,n38_15,n41_15);
nand I_60(n40_15,n41_15,n42_15);
and I_61(n41_15,n51_15,N1372_1_r_3);
and I_62(n42_15,n47_15,N1507_6_r_3);
and I_63(n43_15,n34_15,n36_15);
or I_64(n44_15,G42_7_r_3,n_452_7_r_3);
not I_65(n45_15,N1372_1_r_15);
nand I_66(n46_15,n53_15,N1507_6_r_3);
nor I_67(n47_15,n34_15,n48_15);
not I_68(n48_15,n_573_7_r_3);
and I_69(n49_15,n50_15,N1508_6_r_3);
nand I_70(n50_15,n51_15,n52_15);
nand I_71(n51_15,N1508_1_r_3,N1507_6_r_3);
not I_72(n52_15,N1372_1_r_3);
nor I_73(n53_15,n48_15,n_549_7_r_3);
nor I_74(n54_15,N1372_1_r_3,G42_7_r_3);
not I_75(n55_15,n_569_7_r_3);
endmodule


