module test_I2328(I1231,I1343,I1477,I1470,I1271,I1287,I2328);
input I1231,I1343,I1477,I1470,I1271,I1287;
output I2328;
wire I2181,I2232,I2294,I2311,I2198,I2215;
not I_0(I2181,I1477);
nor I_1(I2328,I2232,I2311);
DFFARX1 I_2(I2215,I1470,I2181,,,I2232,);
nor I_3(I2294,I1287,I1231);
not I_4(I2311,I2294);
nand I_5(I2198,I1343,I1231);
and I_6(I2215,I2198,I1271);
endmodule


