module test_I16469(I14667,I1477,I1470,I14438,I14732,I16469);
input I14667,I1477,I1470,I14438,I14732;
output I16469;
wire I14362,I14350,I16452,I14684,I14455,I16240,I16435,I14808,I14825,I14359,I14370;
DFFARX1 I_0(I14825,I1470,I14370,,,I14362,);
nand I_1(I14350,I14455,I14732);
and I_2(I16452,I16435,I14362);
nand I_3(I14684,I14667);
DFFARX1 I_4(I16452,I1470,I16240,,,I16469,);
DFFARX1 I_5(I1470,I14370,,,I14455,);
not I_6(I16240,I1477);
nand I_7(I16435,I14359,I14350);
DFFARX1 I_8(I1470,I14370,,,I14808,);
and I_9(I14825,I14808,I14684);
nor I_10(I14359,I14667,I14438);
not I_11(I14370,I1477);
endmodule


