module test_I5642(I1504,I1477,I1470,I5642);
input I1504,I1477,I1470;
output I5642;
wire I3388,I5625,I3377,I3747,I5105;
not I_0(I3388,I1477);
DFFARX1 I_1(I3377,I1470,I5105,,,I5625,);
not I_2(I3377,I3747);
DFFARX1 I_3(I1504,I1470,I3388,,,I3747,);
not I_4(I5105,I1477);
not I_5(I5642,I5625);
endmodule


