module test_I16069(I1477,I1470,I14261,I14066,I16069);
input I1477,I1470,I14261,I14066;
output I16069;
wire I13752,I16052,I13775,I15611,I14278;
DFFARX1 I_0(I14278,I1470,I13775,,,I13752,);
DFFARX1 I_1(I13752,I1470,I15611,,,I16052,);
not I_2(I13775,I1477);
not I_3(I15611,I1477);
or I_4(I14278,I14066,I14261);
not I_5(I16069,I16052);
endmodule


