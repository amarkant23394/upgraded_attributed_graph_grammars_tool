module test_final(IN_1_1_l_7,IN_2_1_l_7,IN_3_1_l_7,G18_7_l_7,G15_7_l_7,IN_1_7_l_7,IN_4_7_l_7,IN_5_7_l_7,IN_7_7_l_7,IN_9_7_l_7,IN_10_7_l_7,IN_1_8_l_7,IN_2_8_l_7,IN_3_8_l_7,IN_6_8_l_7,blif_clk_net_7_r_2,blif_reset_net_7_r_2,N1371_0_r_2,N1508_0_r_2,N1372_1_r_2,N1508_1_r_2,N6147_2_r_2,N1507_6_r_2,N1508_6_r_2,G42_7_r_2,n_572_7_r_2,n_573_7_r_2,n_549_7_r_2,n_569_7_r_2,n_452_7_r_2);
input IN_1_1_l_7,IN_2_1_l_7,IN_3_1_l_7,G18_7_l_7,G15_7_l_7,IN_1_7_l_7,IN_4_7_l_7,IN_5_7_l_7,IN_7_7_l_7,IN_9_7_l_7,IN_10_7_l_7,IN_1_8_l_7,IN_2_8_l_7,IN_3_8_l_7,IN_6_8_l_7,blif_clk_net_7_r_2,blif_reset_net_7_r_2;
output N1371_0_r_2,N1508_0_r_2,N1372_1_r_2,N1508_1_r_2,N6147_2_r_2,N1507_6_r_2,N1508_6_r_2,G42_7_r_2,n_572_7_r_2,n_573_7_r_2,n_549_7_r_2,n_569_7_r_2,n_452_7_r_2;
wire N1371_0_r_7,N1508_0_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_102_5_r_7,n_547_5_r_7,G42_7_r_7,n_572_7_r_7,n_573_7_r_7,n_549_7_r_7,n_569_7_r_7,n_452_7_r_7,n4_7_l_7,n53_7,n30_7,N3_8_l_7,n54_7,n_431_5_r_7,n4_7_r_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7,n43_7,n44_7,n45_7,n46_7,n47_7,n48_7,n49_7,n50_7,n51_7,n52_7,n4_7_l_2,n10_2,n59_2,n33_2,N3_8_l_2,n32_internal_2,n32_2,n4_7_r_2,n34_2,n35_2,n36_2,n37_2,n38_2,n39_2,n40_2,n41_2,n42_2,n43_2,n44_2,n45_2,n46_2,n47_2,n48_2,n49_2,n50_2,n51_2,n52_2,n53_2,n54_2,n55_2,n56_2,n57_2,n58_2;
nor I_0(N1371_0_r_7,n53_7,n52_7);
nor I_1(N1508_0_r_7,n51_7,n52_7);
nand I_2(n_429_or_0_5_r_7,n43_7,n48_7);
DFFARX1 I_3(n_431_5_r_7,blif_clk_net_7_r_2,n10_2,G78_5_r_7,);
nand I_4(n_576_5_r_7,n31_7,n32_7);
nor I_5(n_102_5_r_7,IN_5_7_l_7,IN_9_7_l_7);
nand I_6(n_547_5_r_7,n31_7,n38_7);
DFFARX1 I_7(n4_7_r_7,blif_clk_net_7_r_2,n10_2,G42_7_r_7,);
nor I_8(n_572_7_r_7,n54_7,n33_7);
nand I_9(n_573_7_r_7,n_102_5_r_7,n_452_7_r_7);
nor I_10(n_549_7_r_7,n53_7,n36_7);
nand I_11(n_569_7_r_7,n_102_5_r_7,n30_7);
nand I_12(n_452_7_r_7,IN_1_1_l_7,IN_2_1_l_7);
nor I_13(n4_7_l_7,G18_7_l_7,IN_1_7_l_7);
DFFARX1 I_14(n4_7_l_7,blif_clk_net_7_r_2,n10_2,n53_7,);
not I_15(n30_7,n53_7);
and I_16(N3_8_l_7,IN_6_8_l_7,n50_7);
DFFARX1 I_17(N3_8_l_7,blif_clk_net_7_r_2,n10_2,n54_7,);
nand I_18(n_431_5_r_7,n40_7,n41_7);
nor I_19(n4_7_r_7,n54_7,n49_7);
and I_20(n31_7,n_102_5_r_7,n39_7);
not I_21(n32_7,G18_7_l_7);
nor I_22(n33_7,IN_10_7_l_7,n34_7);
and I_23(n34_7,IN_4_7_l_7,n35_7);
not I_24(n35_7,G15_7_l_7);
nor I_25(n36_7,G18_7_l_7,n37_7);
or I_26(n37_7,IN_5_7_l_7,n54_7);
or I_27(n38_7,IN_1_8_l_7,IN_3_8_l_7);
nor I_28(n39_7,IN_3_1_l_7,n_452_7_r_7);
nand I_29(n40_7,n46_7,n47_7);
nand I_30(n41_7,n42_7,n43_7);
nor I_31(n42_7,n44_7,n45_7);
nor I_32(n43_7,IN_1_8_l_7,IN_3_8_l_7);
nor I_33(n44_7,G15_7_l_7,IN_7_7_l_7);
nor I_34(n45_7,IN_9_7_l_7,IN_10_7_l_7);
nand I_35(n46_7,IN_4_7_l_7,n35_7);
not I_36(n47_7,IN_10_7_l_7);
or I_37(n48_7,IN_3_1_l_7,n_452_7_r_7);
not I_38(n49_7,n_452_7_r_7);
nand I_39(n50_7,IN_2_8_l_7,IN_3_8_l_7);
and I_40(n51_7,n_452_7_r_7,n45_7);
not I_41(n52_7,n44_7);
nor I_42(N1371_0_r_2,n32_2,n35_2);
nor I_43(N1508_0_r_2,n32_2,n55_2);
not I_44(N1372_1_r_2,n54_2);
nor I_45(N1508_1_r_2,n59_2,n54_2);
nor I_46(N6147_2_r_2,n42_2,n43_2);
nor I_47(N1507_6_r_2,n40_2,n53_2);
nor I_48(N1508_6_r_2,n33_2,n50_2);
DFFARX1 I_49(n4_7_r_2,blif_clk_net_7_r_2,n10_2,G42_7_r_2,);
nor I_50(n_572_7_r_2,n36_2,n37_2);
or I_51(n_573_7_r_2,n34_2,n35_2);
nor I_52(n_549_7_r_2,n40_2,n41_2);
nand I_53(n_569_7_r_2,n38_2,n39_2);
nor I_54(n_452_7_r_2,n59_2,n35_2);
nor I_55(n4_7_l_2,N1508_0_r_7,n_429_or_0_5_r_7);
not I_56(n10_2,blif_reset_net_7_r_2);
DFFARX1 I_57(n4_7_l_2,blif_clk_net_7_r_2,n10_2,n59_2,);
not I_58(n33_2,n59_2);
and I_59(N3_8_l_2,n49_2,N1371_0_r_7);
DFFARX1 I_60(N3_8_l_2,blif_clk_net_7_r_2,n10_2,n32_internal_2,);
not I_61(n32_2,n32_internal_2);
nor I_62(n4_7_r_2,n59_2,n36_2);
not I_63(n34_2,n39_2);
nor I_64(n35_2,n_429_or_0_5_r_7,N1371_0_r_7);
nor I_65(n36_2,N1508_0_r_7,n_576_5_r_7);
or I_66(n37_2,n_573_7_r_7,n_549_7_r_7);
not I_67(n38_2,n40_2);
nand I_68(n39_2,n45_2,n57_2);
nor I_69(n40_2,n47_2,G78_5_r_7);
nor I_70(n41_2,n32_2,n36_2);
not I_71(n42_2,n53_2);
nand I_72(n43_2,n44_2,n45_2);
nand I_73(n44_2,n38_2,n46_2);
not I_74(n45_2,n_573_7_r_7);
nand I_75(n46_2,n47_2,n48_2);
nand I_76(n47_2,G42_7_r_7,n_572_7_r_7);
or I_77(n48_2,n_569_7_r_7,G78_5_r_7);
nand I_78(n49_2,n_547_5_r_7,N1371_0_r_7);
nand I_79(n50_2,n51_2,n52_2);
not I_80(n51_2,n47_2);
nand I_81(n52_2,n38_2,n53_2);
nor I_82(n53_2,n_576_5_r_7,n_549_7_r_7);
nand I_83(n54_2,n42_2,n56_2);
nor I_84(n55_2,n34_2,n56_2);
nor I_85(n56_2,n_569_7_r_7,G78_5_r_7);
nand I_86(n57_2,n58_2,n_576_5_r_7);
not I_87(n58_2,G78_5_r_7);
endmodule


