module test_I10414(I7621,I1477,I7559,I7535,I1470,I7731,I10414);
input I7621,I1477,I7559,I7535,I1470,I7731;
output I10414;
wire I10349,I10086,I7550,I7570,I7532,I10397,I7977,I7544,I10052,I10103,I10332,I10069;
and I_0(I10349,I10332,I7550);
and I_1(I10086,I10069,I7544);
nand I_2(I7550,I7977,I7731);
not I_3(I7570,I1477);
nor I_4(I10414,I10103,I10397);
DFFARX1 I_5(I1470,I7570,,,I7532,);
not I_6(I10397,I10349);
DFFARX1 I_7(I1470,I7570,,,I7977,);
DFFARX1 I_8(I7621,I1470,I7570,,,I7544,);
not I_9(I10052,I1477);
DFFARX1 I_10(I10086,I1470,I10052,,,I10103,);
DFFARX1 I_11(I7532,I1470,I10052,,,I10332,);
nand I_12(I10069,I7559,I7535);
endmodule


