module test_I10349(I1477,I1470,I6705,I6657,I10349);
input I1477,I1470,I6705,I6657;
output I10349;
wire I8107,I7550,I6321,I6297,I7714,I8090,I7570,I7977,I7731,I10052,I7532,I10332;
and I_0(I10349,I10332,I7550);
not I_1(I8107,I8090);
nand I_2(I7550,I7977,I7731);
nand I_3(I6321,I6705,I6657);
DFFARX1 I_4(I1470,,,I6297,);
not I_5(I7714,I6297);
DFFARX1 I_6(I1470,I7570,,,I8090,);
not I_7(I7570,I1477);
DFFARX1 I_8(I6321,I1470,I7570,,,I7977,);
not I_9(I7731,I7714);
not I_10(I10052,I1477);
DFFARX1 I_11(I8107,I1470,I7570,,,I7532,);
DFFARX1 I_12(I7532,I1470,I10052,,,I10332,);
endmodule


