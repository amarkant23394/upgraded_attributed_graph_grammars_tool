module test_I8394(I4629,I1477,I1470,I4824,I8394);
input I4629,I1477,I1470,I4824;
output I8394;
wire I5751,I5713,I6110,I6127,I4533,I4509;
not I_0(I8394,I5713);
not I_1(I5751,I1477);
DFFARX1 I_2(I6127,I1470,I5751,,,I5713,);
DFFARX1 I_3(I4509,I1470,I5751,,,I6110,);
and I_4(I6127,I6110,I4533);
or I_5(I4533,I4824,I4629);
DFFARX1 I_6(I1470,,,I4509,);
endmodule


