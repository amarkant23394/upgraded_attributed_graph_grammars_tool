module test_I1359(I1239,I1287,I1359);
input I1239,I1287;
output I1359;
wire ;
nand I_0(I1359,I1287,I1239);
endmodule


