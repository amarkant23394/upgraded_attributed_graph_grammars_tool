module test_final(IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_4_2_l_10,IN_5_2_l_10,IN_1_6_l_10,IN_2_6_l_10,IN_3_6_l_10,IN_4_6_l_10,IN_5_6_l_10,IN_1_9_l_10,IN_2_9_l_10,IN_3_9_l_10,IN_4_9_l_10,IN_5_9_l_10,blif_clk_net_7_r_1,blif_reset_net_7_r_1,N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,N6147_9_r_1,N6134_9_r_1);
input IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_4_2_l_10,IN_5_2_l_10,IN_1_6_l_10,IN_2_6_l_10,IN_3_6_l_10,IN_4_6_l_10,IN_5_6_l_10,IN_1_9_l_10,IN_2_9_l_10,IN_3_9_l_10,IN_4_9_l_10,IN_5_9_l_10,blif_clk_net_7_r_1,blif_reset_net_7_r_1;
output N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,N6147_9_r_1,N6134_9_r_1;
wire N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1372_4_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10,I_BUFF_1_9_r_10,N3_8_r_10,n35_10,n36_10,n37_10,n38_10,n39_10,n40_10,n41_10,n42_10,n43_10,n44_10,n45_10,n46_10,n47_10,n48_10,n49_10,n50_10,n51_10,n52_10,n53_10,n54_10,n55_10,n56_10,n57_10,n58_10,n59_10,n60_10,n61_10,n62_10,n63_10,n64_10,N1371_0_r_1,n_452_7_r_1,I_BUFF_1_9_r_1,n4_7_r_1,n9_1,n29_1,n30_1,n31_1,n32_1,n33_1,n34_1,n35_1,n36_1,n37_1,n38_1,n39_1,n40_1,n41_1,n42_1,n43_1,n44_1,n45_1,n46_1,n47_1,n48_1,n49_1,n50_1,n51_1,n52_1,n53_1,n54_1,n55_1;
nor I_0(N1371_0_r_10,n37_10,n38_10);
nor I_1(N1508_0_r_10,n37_10,n58_10);
nand I_2(N6147_2_r_10,n39_10,n40_10);
not I_3(N6147_3_r_10,n39_10);
nor I_4(N1372_4_r_10,n46_10,n49_10);
nor I_5(N1508_4_r_10,n51_10,n52_10);
nor I_6(N1507_6_r_10,n49_10,n60_10);
nor I_7(N1508_6_r_10,n49_10,n50_10);
nor I_8(n_42_8_r_10,I_BUFF_1_9_r_10,n35_10);
DFFARX1 I_9(N3_8_r_10,blif_clk_net_7_r_1,n9_1,G199_8_r_10,);
nor I_10(N6147_9_r_10,n36_10,n37_10);
nor I_11(N6134_9_r_10,I_BUFF_1_9_r_10,n46_10);
not I_12(I_BUFF_1_9_r_10,n48_10);
nor I_13(N3_8_r_10,n44_10,n47_10);
not I_14(n35_10,n49_10);
nor I_15(n36_10,I_BUFF_1_9_r_10,n38_10);
not I_16(n37_10,IN_1_9_l_10);
not I_17(n38_10,n46_10);
nand I_18(n39_10,n43_10,n44_10);
nand I_19(n40_10,I_BUFF_1_9_r_10,n41_10);
nor I_20(n41_10,IN_1_9_l_10,n42_10);
not I_21(n42_10,n44_10);
nor I_22(n43_10,IN_1_9_l_10,n45_10);
nand I_23(n44_10,IN_2_6_l_10,n54_10);
nor I_24(n45_10,IN_5_9_l_10,n59_10);
nand I_25(n46_10,IN_2_9_l_10,n61_10);
nor I_26(n47_10,n46_10,n48_10);
nand I_27(n48_10,n62_10,n63_10);
nand I_28(n49_10,IN_5_6_l_10,n56_10);
not I_29(n50_10,n45_10);
nor I_30(n51_10,n42_10,n53_10);
not I_31(n52_10,N1372_4_r_10);
nor I_32(n53_10,n48_10,n50_10);
and I_33(n54_10,IN_1_6_l_10,n55_10);
nand I_34(n55_10,n56_10,n57_10);
nand I_35(n56_10,IN_3_6_l_10,IN_4_6_l_10);
not I_36(n57_10,IN_5_6_l_10);
nor I_37(n58_10,n35_10,n45_10);
nor I_38(n59_10,IN_3_9_l_10,IN_4_9_l_10);
nor I_39(n60_10,n37_10,n46_10);
or I_40(n61_10,IN_3_9_l_10,IN_4_9_l_10);
nor I_41(n62_10,IN_1_2_l_10,IN_2_2_l_10);
or I_42(n63_10,IN_5_2_l_10,n64_10);
nor I_43(n64_10,IN_3_2_l_10,IN_4_2_l_10);
and I_44(N1371_0_r_1,I_BUFF_1_9_r_1,n55_1);
nor I_45(N1508_0_r_1,n40_1,n44_1);
nor I_46(N1507_6_r_1,n43_1,n49_1);
nor I_47(N1508_6_r_1,n41_1,n42_1);
DFFARX1 I_48(n4_7_r_1,blif_clk_net_7_r_1,n9_1,G42_7_r_1,);
nor I_49(n_572_7_r_1,n29_1,n30_1);
not I_50(n_573_7_r_1,n_452_7_r_1);
nor I_51(n_549_7_r_1,N1371_0_r_1,n31_1);
or I_52(n_569_7_r_1,n30_1,n31_1);
nor I_53(n_452_7_r_1,n30_1,n32_1);
nor I_54(N6147_9_r_1,n35_1,n36_1);
nand I_55(N6134_9_r_1,n38_1,n39_1);
not I_56(I_BUFF_1_9_r_1,n40_1);
nor I_57(n4_7_r_1,I_BUFF_1_9_r_1,n30_1);
not I_58(n9_1,blif_reset_net_7_r_1);
nor I_59(n29_1,n34_1,N6147_3_r_10);
nor I_60(n30_1,n33_1,n34_1);
nor I_61(n31_1,n54_1,N6147_2_r_10);
not I_62(n32_1,n48_1);
nor I_63(n33_1,N6147_2_r_10,N1508_6_r_10);
not I_64(n34_1,G199_8_r_10);
nor I_65(n35_1,I_BUFF_1_9_r_1,n37_1);
not I_66(n36_1,n29_1);
not I_67(n37_1,n41_1);
nand I_68(n38_1,I_BUFF_1_9_r_1,N6134_9_r_10);
nand I_69(n39_1,n37_1,n40_1);
nand I_70(n40_1,N1371_0_r_10,N1508_0_r_10);
nand I_71(n41_1,n52_1,N1507_6_r_10);
or I_72(n42_1,n36_1,n43_1);
nor I_73(n43_1,n32_1,n49_1);
nand I_74(n44_1,n45_1,n46_1);
nand I_75(n45_1,n47_1,n48_1);
not I_76(n46_1,N6134_9_r_10);
not I_77(n47_1,n31_1);
nand I_78(n48_1,n50_1,N1508_0_r_10);
nor I_79(n49_1,n41_1,n47_1);
and I_80(n50_1,n51_1,N6147_9_r_10);
nand I_81(n51_1,n52_1,n53_1);
nand I_82(n52_1,n_42_8_r_10,N6147_3_r_10);
not I_83(n53_1,N1507_6_r_10);
or I_84(n54_1,N1508_4_r_10,N1371_0_r_10);
nor I_85(n55_1,n29_1,N6134_9_r_10);
endmodule


