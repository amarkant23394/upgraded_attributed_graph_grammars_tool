module test_I2152(I1327,I1223,I1255,I1477,I1470,I2152);
input I1327,I1223,I1255,I1477,I1470;
output I2152;
wire I2441,I2181,I2458,I2424;
and I_0(I2441,I2424,I1327);
not I_1(I2181,I1477);
DFFARX1 I_2(I2441,I1470,I2181,,,I2458,);
DFFARX1 I_3(I2458,I1470,I2181,,,I2152,);
nand I_4(I2424,I1223,I1255);
endmodule


