module test_I14049(I10349,I10120,I10032,I1477,I1470,I14049);
input I10349,I10120,I10032,I1477,I1470;
output I14049;
wire I12270,I10219,I10014,I12349,I10041,I13775,I11973,I11990,I10052,I11962;
nand I_0(I12270,I11990,I10014);
DFFARX1 I_1(I1470,I10052,,,I10219,);
DFFARX1 I_2(I10219,I1470,I10052,,,I10014,);
DFFARX1 I_3(I10041,I1470,I11973,,,I12349,);
nor I_4(I10041,I10349,I10120);
DFFARX1 I_5(I11962,I1470,I13775,,,I14049,);
not I_6(I13775,I1477);
not I_7(I11973,I1477);
not I_8(I11990,I10032);
not I_9(I10052,I1477);
nor I_10(I11962,I12349,I12270);
endmodule


