module test_final(IN_1_1_l_2,IN_2_1_l_2,IN_3_1_l_2,G18_7_l_2,G15_7_l_2,IN_1_7_l_2,IN_4_7_l_2,IN_5_7_l_2,IN_7_7_l_2,IN_9_7_l_2,IN_10_7_l_2,IN_1_8_l_2,IN_2_8_l_2,IN_3_8_l_2,IN_6_8_l_2,blif_clk_net_7_r_1,blif_reset_net_7_r_1,N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,N6147_9_r_1,N6134_9_r_1);
input IN_1_1_l_2,IN_2_1_l_2,IN_3_1_l_2,G18_7_l_2,G15_7_l_2,IN_1_7_l_2,IN_4_7_l_2,IN_5_7_l_2,IN_7_7_l_2,IN_9_7_l_2,IN_10_7_l_2,IN_1_8_l_2,IN_2_8_l_2,IN_3_8_l_2,IN_6_8_l_2,blif_clk_net_7_r_1,blif_reset_net_7_r_1;
output N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,N6147_9_r_1,N6134_9_r_1;
wire N1371_0_r_2,N1508_0_r_2,N1372_1_r_2,N1508_1_r_2,N6147_2_r_2,N1507_6_r_2,N1508_6_r_2,G42_7_r_2,n_572_7_r_2,n_573_7_r_2,n_549_7_r_2,n_569_7_r_2,n_452_7_r_2,n4_7_l_2,n59_2,n33_2,N3_8_l_2,n32_internal_2,n32_2,n4_7_r_2,n34_2,n35_2,n36_2,n37_2,n38_2,n39_2,n40_2,n41_2,n42_2,n43_2,n44_2,n45_2,n46_2,n47_2,n48_2,n49_2,n50_2,n51_2,n52_2,n53_2,n54_2,n55_2,n56_2,n57_2,n58_2,N1371_0_r_1,n_452_7_r_1,I_BUFF_1_9_r_1,n4_7_r_1,n9_1,n29_1,n30_1,n31_1,n32_1,n33_1,n34_1,n35_1,n36_1,n37_1,n38_1,n39_1,n40_1,n41_1,n42_1,n43_1,n44_1,n45_1,n46_1,n47_1,n48_1,n49_1,n50_1,n51_1,n52_1,n53_1,n54_1,n55_1;
nor I_0(N1371_0_r_2,n32_2,n35_2);
nor I_1(N1508_0_r_2,n32_2,n55_2);
not I_2(N1372_1_r_2,n54_2);
nor I_3(N1508_1_r_2,n59_2,n54_2);
nor I_4(N6147_2_r_2,n42_2,n43_2);
nor I_5(N1507_6_r_2,n40_2,n53_2);
nor I_6(N1508_6_r_2,n33_2,n50_2);
DFFARX1 I_7(n4_7_r_2,blif_clk_net_7_r_1,n9_1,G42_7_r_2,);
nor I_8(n_572_7_r_2,n36_2,n37_2);
or I_9(n_573_7_r_2,n34_2,n35_2);
nor I_10(n_549_7_r_2,n40_2,n41_2);
nand I_11(n_569_7_r_2,n38_2,n39_2);
nor I_12(n_452_7_r_2,n59_2,n35_2);
nor I_13(n4_7_l_2,G18_7_l_2,IN_1_7_l_2);
DFFARX1 I_14(n4_7_l_2,blif_clk_net_7_r_1,n9_1,n59_2,);
not I_15(n33_2,n59_2);
and I_16(N3_8_l_2,IN_6_8_l_2,n49_2);
DFFARX1 I_17(N3_8_l_2,blif_clk_net_7_r_1,n9_1,n32_internal_2,);
not I_18(n32_2,n32_internal_2);
nor I_19(n4_7_r_2,n59_2,n36_2);
not I_20(n34_2,n39_2);
nor I_21(n35_2,IN_1_8_l_2,IN_3_8_l_2);
nor I_22(n36_2,G18_7_l_2,IN_5_7_l_2);
or I_23(n37_2,IN_9_7_l_2,IN_10_7_l_2);
not I_24(n38_2,n40_2);
nand I_25(n39_2,n45_2,n57_2);
nor I_26(n40_2,IN_3_1_l_2,n47_2);
nor I_27(n41_2,n32_2,n36_2);
not I_28(n42_2,n53_2);
nand I_29(n43_2,n44_2,n45_2);
nand I_30(n44_2,n38_2,n46_2);
not I_31(n45_2,IN_10_7_l_2);
nand I_32(n46_2,n47_2,n48_2);
nand I_33(n47_2,IN_1_1_l_2,IN_2_1_l_2);
or I_34(n48_2,G15_7_l_2,IN_7_7_l_2);
nand I_35(n49_2,IN_2_8_l_2,IN_3_8_l_2);
nand I_36(n50_2,n51_2,n52_2);
not I_37(n51_2,n47_2);
nand I_38(n52_2,n38_2,n53_2);
nor I_39(n53_2,IN_5_7_l_2,IN_9_7_l_2);
nand I_40(n54_2,n42_2,n56_2);
nor I_41(n55_2,n34_2,n56_2);
nor I_42(n56_2,G15_7_l_2,IN_7_7_l_2);
nand I_43(n57_2,IN_4_7_l_2,n58_2);
not I_44(n58_2,G15_7_l_2);
and I_45(N1371_0_r_1,I_BUFF_1_9_r_1,n55_1);
nor I_46(N1508_0_r_1,n40_1,n44_1);
nor I_47(N1507_6_r_1,n43_1,n49_1);
nor I_48(N1508_6_r_1,n41_1,n42_1);
DFFARX1 I_49(n4_7_r_1,blif_clk_net_7_r_1,n9_1,G42_7_r_1,);
nor I_50(n_572_7_r_1,n29_1,n30_1);
not I_51(n_573_7_r_1,n_452_7_r_1);
nor I_52(n_549_7_r_1,N1371_0_r_1,n31_1);
or I_53(n_569_7_r_1,n30_1,n31_1);
nor I_54(n_452_7_r_1,n30_1,n32_1);
nor I_55(N6147_9_r_1,n35_1,n36_1);
nand I_56(N6134_9_r_1,n38_1,n39_1);
not I_57(I_BUFF_1_9_r_1,n40_1);
nor I_58(n4_7_r_1,I_BUFF_1_9_r_1,n30_1);
not I_59(n9_1,blif_reset_net_7_r_1);
nor I_60(n29_1,n34_1,n_452_7_r_2);
nor I_61(n30_1,n33_1,n34_1);
nor I_62(n31_1,n54_1,N6147_2_r_2);
not I_63(n32_1,n48_1);
nor I_64(n33_1,N1508_1_r_2,N1508_0_r_2);
not I_65(n34_1,n_569_7_r_2);
nor I_66(n35_1,I_BUFF_1_9_r_1,n37_1);
not I_67(n36_1,n29_1);
not I_68(n37_1,n41_1);
nand I_69(n38_1,I_BUFF_1_9_r_1,n_572_7_r_2);
nand I_70(n39_1,n37_1,n40_1);
nand I_71(n40_1,N1372_1_r_2,n_549_7_r_2);
nand I_72(n41_1,n52_1,N1371_0_r_2);
or I_73(n42_1,n36_1,n43_1);
nor I_74(n43_1,n32_1,n49_1);
nand I_75(n44_1,n45_1,n46_1);
nand I_76(n45_1,n47_1,n48_1);
not I_77(n46_1,n_572_7_r_2);
not I_78(n47_1,n31_1);
nand I_79(n48_1,n50_1,n_573_7_r_2);
nor I_80(n49_1,n41_1,n47_1);
and I_81(n50_1,n51_1,N1507_6_r_2);
nand I_82(n51_1,n52_1,n53_1);
nand I_83(n52_1,G42_7_r_2,N1371_0_r_2);
not I_84(n53_1,N1371_0_r_2);
or I_85(n54_1,N1508_0_r_2,N1508_6_r_2);
nor I_86(n55_1,n29_1,n_572_7_r_2);
endmodule


