module test_I12590(I1477,I1470,I12590);
input I1477,I1470;
output I12590;
wire I12619,I12752,I12735,I10630,I11009;
not I_0(I12619,I1477);
not I_1(I12590,I12752);
DFFARX1 I_2(I12735,I1470,I12619,,,I12752,);
DFFARX1 I_3(I10630,I1470,I12619,,,I12735,);
not I_4(I10630,I11009);
DFFARX1 I_5(I1470,,,I11009,);
endmodule


