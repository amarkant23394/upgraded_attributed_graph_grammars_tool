module test_I2294(I1287,I1231,I2294);
input I1287,I1231;
output I2294;
wire ;
nor I_0(I2294,I1287,I1231);
endmodule


