module test_final(IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_6_2_l_10,IN_1_3_l_10,IN_2_3_l_10,IN_4_3_l_10,IN_1_4_l_10,IN_2_4_l_10,IN_3_4_l_10,IN_6_4_l_10,blif_clk_net_1_r_5,blif_reset_net_1_r_5,G42_1_r_5,n_572_1_r_5,n_573_1_r_5,n_549_1_r_5,n_569_1_r_5,n_452_1_r_5,ACVQN2_3_r_5,n_266_and_0_3_r_5,ACVQN1_5_r_5,P6_5_r_5);
input IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_6_2_l_10,IN_1_3_l_10,IN_2_3_l_10,IN_4_3_l_10,IN_1_4_l_10,IN_2_4_l_10,IN_3_4_l_10,IN_6_4_l_10,blif_clk_net_1_r_5,blif_reset_net_1_r_5;
output G42_1_r_5,n_572_1_r_5,n_573_1_r_5,n_549_1_r_5,n_569_1_r_5,n_452_1_r_5,ACVQN2_3_r_5,n_266_and_0_3_r_5,ACVQN1_5_r_5,P6_5_r_5;
wire G42_1_r_10,n_572_1_r_10,n_573_1_r_10,n_549_1_r_10,n_452_1_r_10,n_42_2_r_10,G199_2_r_10,ACVQN2_3_r_10,n_266_and_0_3_r_10,N3_2_l_10,n25_10,n16_10,n26_10,ACVQN1_3_l_10,N1_4_l_10,G199_4_l_10,n27_10,n17_10,n4_1_r_10,N3_2_r_10,n3_10,n13_internal_10,n13_10,n18_10,n19_10,n20_10,n21_10,n22_10,n23_10,n24_10,N3_2_l_5,n5_5,G199_2_l_5,ACVQN2_3_l_5,n13_5,ACVQN1_3_l_5,N1_4_l_5,n21_5,n15_5,n22_5,n4_1_r_5,n11_internal_5,n11_5,n_42_2_l_5,n1_5,P6_5_r_internal_5,n16_5,n17_5,n18_5,n19_5,n20_5;
DFFARX1 I_0(n4_1_r_10,blif_clk_net_1_r_5,n5_5,G42_1_r_10,);
nor I_1(n_572_1_r_10,n26_10,n3_10);
nand I_2(n_573_1_r_10,n16_10,n18_10);
nand I_3(n_549_1_r_10,n19_10,n20_10);
nor I_4(n_452_1_r_10,n25_10,n21_10);
nor I_5(n_42_2_r_10,n26_10,G199_4_l_10);
DFFARX1 I_6(N3_2_r_10,blif_clk_net_1_r_5,n5_5,G199_2_r_10,);
DFFARX1 I_7(G199_4_l_10,blif_clk_net_1_r_5,n5_5,ACVQN2_3_r_10,);
nor I_8(n_266_and_0_3_r_10,n17_10,n13_10);
and I_9(N3_2_l_10,IN_6_2_l_10,n23_10);
DFFARX1 I_10(N3_2_l_10,blif_clk_net_1_r_5,n5_5,n25_10,);
not I_11(n16_10,n25_10);
DFFARX1 I_12(IN_1_3_l_10,blif_clk_net_1_r_5,n5_5,n26_10,);
DFFARX1 I_13(IN_2_3_l_10,blif_clk_net_1_r_5,n5_5,ACVQN1_3_l_10,);
and I_14(N1_4_l_10,IN_6_4_l_10,n24_10);
DFFARX1 I_15(N1_4_l_10,blif_clk_net_1_r_5,n5_5,G199_4_l_10,);
DFFARX1 I_16(IN_3_4_l_10,blif_clk_net_1_r_5,n5_5,n27_10,);
not I_17(n17_10,n27_10);
nor I_18(n4_1_r_10,n27_10,n21_10);
nor I_19(N3_2_r_10,n16_10,n22_10);
not I_20(n3_10,n18_10);
DFFARX1 I_21(n3_10,blif_clk_net_1_r_5,n5_5,n13_internal_10,);
not I_22(n13_10,n13_internal_10);
nand I_23(n18_10,IN_4_3_l_10,ACVQN1_3_l_10);
not I_24(n19_10,n_452_1_r_10);
nand I_25(n20_10,n16_10,n26_10);
nor I_26(n21_10,IN_1_2_l_10,IN_3_2_l_10);
and I_27(n22_10,n26_10,n21_10);
nand I_28(n23_10,IN_2_2_l_10,IN_3_2_l_10);
nand I_29(n24_10,IN_1_4_l_10,IN_2_4_l_10);
DFFARX1 I_30(n4_1_r_5,blif_clk_net_1_r_5,n5_5,G42_1_r_5,);
nor I_31(n_572_1_r_5,n21_5,n22_5);
nand I_32(n_573_1_r_5,n13_5,n16_5);
nor I_33(n_549_1_r_5,n21_5,n17_5);
nand I_34(n_569_1_r_5,n13_5,n15_5);
nor I_35(n_452_1_r_5,n22_5,n_42_2_l_5);
DFFARX1 I_36(G199_2_l_5,blif_clk_net_1_r_5,n5_5,ACVQN2_3_r_5,);
nor I_37(n_266_and_0_3_r_5,n11_5,n16_5);
DFFARX1 I_38(n_42_2_l_5,blif_clk_net_1_r_5,n5_5,ACVQN1_5_r_5,);
not I_39(P6_5_r_5,P6_5_r_internal_5);
and I_40(N3_2_l_5,n19_5,n_572_1_r_10);
not I_41(n5_5,blif_reset_net_1_r_5);
DFFARX1 I_42(N3_2_l_5,blif_clk_net_1_r_5,n5_5,G199_2_l_5,);
DFFARX1 I_43(ACVQN2_3_r_10,blif_clk_net_1_r_5,n5_5,ACVQN2_3_l_5,);
not I_44(n13_5,ACVQN2_3_l_5);
DFFARX1 I_45(G199_2_r_10,blif_clk_net_1_r_5,n5_5,ACVQN1_3_l_5,);
and I_46(N1_4_l_5,n20_5,n_42_2_r_10);
DFFARX1 I_47(N1_4_l_5,blif_clk_net_1_r_5,n5_5,n21_5,);
not I_48(n15_5,n21_5);
DFFARX1 I_49(n_572_1_r_10,blif_clk_net_1_r_5,n5_5,n22_5,);
nor I_50(n4_1_r_5,G199_2_l_5,n22_5);
DFFARX1 I_51(ACVQN2_3_l_5,blif_clk_net_1_r_5,n5_5,n11_internal_5,);
not I_52(n11_5,n11_internal_5);
nor I_53(n_42_2_l_5,n_549_1_r_10,n_266_and_0_3_r_10);
not I_54(n1_5,n18_5);
DFFARX1 I_55(n1_5,blif_clk_net_1_r_5,n5_5,P6_5_r_internal_5,);
not I_56(n16_5,n_42_2_l_5);
nor I_57(n17_5,n22_5,n18_5);
nand I_58(n18_5,ACVQN1_3_l_5,n_573_1_r_10);
nand I_59(n19_5,G42_1_r_10,n_549_1_r_10);
nand I_60(n20_5,G42_1_r_10,n_573_1_r_10);
endmodule


