module test_I1749(I1223,I1255,I1376,I1294,I1239,I1207,I1301,I1749);
input I1223,I1255,I1376,I1294,I1239,I1207,I1301;
output I1749;
wire I1410,I1560,I1622,I1543,I1526,I1342,I1393,I1509,I1639;
nor I_0(I1410,I1223,I1239);
and I_1(I1560,I1410,I1543);
DFFARX1 I_2(I1255,I1294,I1342,,,I1622,);
or I_3(I1749,I1639,I1560);
nor I_4(I1543,I1393,I1526);
not I_5(I1526,I1509);
not I_6(I1342,I1301);
DFFARX1 I_7(I1376,I1294,I1342,,,I1393,);
DFFARX1 I_8(I1294,I1342,,,I1509,);
and I_9(I1639,I1622,I1207);
endmodule


