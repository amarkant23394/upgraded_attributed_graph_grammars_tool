module test_I2055(I1215,I1423,I1295,I1470,I1477,I1455,I2055);
input I1215,I1423,I1295,I1470,I1477,I1455;
output I2055;
wire I1518,I2038,I2021,I1586,I1603,I1535;
not I_0(I1518,I1477);
not I_1(I2038,I2021);
DFFARX1 I_2(I1295,I1470,I1518,,,I2021,);
nor I_3(I1586,I1535,I1215);
nand I_4(I1603,I1586,I1423);
not I_5(I1535,I1455);
nand I_6(I2055,I2038,I1603);
endmodule


