module test_final(G1_0_l_12,G2_0_l_12,IN_2_0_l_12,IN_4_0_l_12,IN_5_0_l_12,IN_7_0_l_12,IN_8_0_l_12,IN_10_0_l_12,IN_11_0_l_12,IN_1_5_l_12,IN_2_5_l_12,blif_clk_net_1_r_15,blif_reset_net_1_r_15,G42_1_r_15,n_572_1_r_15,n_573_1_r_15,n_549_1_r_15,n_569_1_r_15,ACVQN2_3_r_15,n_266_and_0_3_r_15,G199_4_r_15,G214_4_r_15);
input G1_0_l_12,G2_0_l_12,IN_2_0_l_12,IN_4_0_l_12,IN_5_0_l_12,IN_7_0_l_12,IN_8_0_l_12,IN_10_0_l_12,IN_11_0_l_12,IN_1_5_l_12,IN_2_5_l_12,blif_clk_net_1_r_15,blif_reset_net_1_r_15;
output G42_1_r_15,n_572_1_r_15,n_573_1_r_15,n_549_1_r_15,n_569_1_r_15,ACVQN2_3_r_15,n_266_and_0_3_r_15,G199_4_r_15,G214_4_r_15;
wire G42_1_r_12,n_572_1_r_12,n_573_1_r_12,n_549_1_r_12,n_42_2_r_12,G199_2_r_12,ACVQN1_5_r_12,P6_5_r_12,n_431_0_l_12,n41_12,ACVQN1_5_l_12,n22_12,n42_12,n4_1_r_12,N3_2_r_12,n3_12,P6_5_r_internal_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12,n_452_1_r_15,n4_1_l_15,n4_15,G42_1_l_15,n15_15,n17_internal_15,n17_15,n30_15,n_572_1_l_15,n14_internal_15,n14_15,N1_4_r_15,n_573_1_l_15,n18_15,n19_15,n20_15,n21_15,n22_15,n23_15,n24_15,n25_15,n26_15,n27_15,n28_15,n29_15;
DFFARX1 I_0(n4_1_r_12,blif_clk_net_1_r_15,n4_15,G42_1_r_12,);
nor I_1(n_572_1_r_12,n29_12,n30_12);
nand I_2(n_573_1_r_12,n26_12,n27_12);
nor I_3(n_549_1_r_12,n33_12,n34_12);
and I_4(n_42_2_r_12,n42_12,n39_12);
DFFARX1 I_5(N3_2_r_12,blif_clk_net_1_r_15,n4_15,G199_2_r_12,);
DFFARX1 I_6(n3_12,blif_clk_net_1_r_15,n4_15,ACVQN1_5_r_12,);
not I_7(P6_5_r_12,P6_5_r_internal_12);
or I_8(n_431_0_l_12,IN_8_0_l_12,n36_12);
DFFARX1 I_9(n_431_0_l_12,blif_clk_net_1_r_15,n4_15,n41_12,);
DFFARX1 I_10(IN_2_5_l_12,blif_clk_net_1_r_15,n4_15,ACVQN1_5_l_12,);
not I_11(n22_12,ACVQN1_5_l_12);
DFFARX1 I_12(IN_1_5_l_12,blif_clk_net_1_r_15,n4_15,n42_12,);
nor I_13(n4_1_r_12,n41_12,n31_12);
nor I_14(N3_2_r_12,n22_12,n40_12);
not I_15(n3_12,n39_12);
DFFARX1 I_16(ACVQN1_5_l_12,blif_clk_net_1_r_15,n4_15,P6_5_r_internal_12,);
and I_17(n26_12,IN_5_0_l_12,IN_7_0_l_12);
nor I_18(n27_12,n28_12,n29_12);
not I_19(n28_12,IN_11_0_l_12);
nand I_20(n29_12,n31_12,n32_12);
nand I_21(n30_12,IN_11_0_l_12,n42_12);
not I_22(n31_12,G2_0_l_12);
not I_23(n32_12,IN_10_0_l_12);
nand I_24(n33_12,n31_12,n35_12);
nand I_25(n34_12,IN_5_0_l_12,IN_7_0_l_12);
nand I_26(n35_12,n41_12,n42_12);
and I_27(n36_12,IN_2_0_l_12,n37_12);
nor I_28(n37_12,IN_4_0_l_12,n38_12);
not I_29(n38_12,G1_0_l_12);
nor I_30(n39_12,IN_5_0_l_12,n38_12);
nor I_31(n40_12,G2_0_l_12,n39_12);
DFFARX1 I_32(n_452_1_r_15,blif_clk_net_1_r_15,n4_15,G42_1_r_15,);
and I_33(n_572_1_r_15,n17_15,n19_15);
nand I_34(n_573_1_r_15,n15_15,n18_15);
nor I_35(n_549_1_r_15,n21_15,n22_15);
nand I_36(n_569_1_r_15,n15_15,n20_15);
nor I_37(n_452_1_r_15,n23_15,n24_15);
DFFARX1 I_38(G42_1_l_15,blif_clk_net_1_r_15,n4_15,ACVQN2_3_r_15,);
nor I_39(n_266_and_0_3_r_15,n17_15,n14_15);
DFFARX1 I_40(N1_4_r_15,blif_clk_net_1_r_15,n4_15,G199_4_r_15,);
DFFARX1 I_41(n_573_1_l_15,blif_clk_net_1_r_15,n4_15,G214_4_r_15,);
nor I_42(n4_1_l_15,G42_1_r_12,P6_5_r_12);
not I_43(n4_15,blif_reset_net_1_r_15);
DFFARX1 I_44(n4_1_l_15,blif_clk_net_1_r_15,n4_15,G42_1_l_15,);
not I_45(n15_15,G42_1_l_15);
DFFARX1 I_46(n_573_1_r_12,blif_clk_net_1_r_15,n4_15,n17_internal_15,);
not I_47(n17_15,n17_internal_15);
DFFARX1 I_48(n_549_1_r_12,blif_clk_net_1_r_15,n4_15,n30_15,);
nor I_49(n_572_1_l_15,ACVQN1_5_r_12,n_572_1_r_12);
DFFARX1 I_50(n_572_1_l_15,blif_clk_net_1_r_15,n4_15,n14_internal_15,);
not I_51(n14_15,n14_internal_15);
nand I_52(N1_4_r_15,n25_15,n26_15);
or I_53(n_573_1_l_15,n_42_2_r_12,G199_2_r_12);
nor I_54(n18_15,n_572_1_r_12,n_42_2_r_12);
nand I_55(n19_15,n27_15,n28_15);
nand I_56(n20_15,n30_15,n_573_1_r_12);
not I_57(n21_15,n20_15);
and I_58(n22_15,n17_15,n_572_1_l_15);
nor I_59(n23_15,G199_2_r_12,P6_5_r_12);
or I_60(n24_15,n_572_1_r_12,n_42_2_r_12);
or I_61(n25_15,n_573_1_l_15,P6_5_r_12);
nand I_62(n26_15,n19_15,n23_15);
not I_63(n27_15,n_572_1_r_12);
nand I_64(n28_15,n29_15,G42_1_r_12);
not I_65(n29_15,n_572_1_r_12);
endmodule


