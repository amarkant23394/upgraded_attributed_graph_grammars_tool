module test_final(G18_1_l_16,G15_1_l_16,IN_1_1_l_16,IN_4_1_l_16,IN_5_1_l_16,IN_7_1_l_16,IN_9_1_l_16,IN_10_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_4_3_l_16,blif_clk_net_1_r_6,blif_reset_net_1_r_6,G42_1_r_6,n_572_1_r_6,n_573_1_r_6,n_549_1_r_6,n_569_1_r_6,n_452_1_r_6,G199_4_r_6,G214_4_r_6,ACVQN1_5_r_6,P6_5_r_6);
input G18_1_l_16,G15_1_l_16,IN_1_1_l_16,IN_4_1_l_16,IN_5_1_l_16,IN_7_1_l_16,IN_9_1_l_16,IN_10_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_4_3_l_16,blif_clk_net_1_r_6,blif_reset_net_1_r_6;
output G42_1_r_6,n_572_1_r_6,n_573_1_r_6,n_549_1_r_6,n_569_1_r_6,n_452_1_r_6,G199_4_r_6,G214_4_r_6,ACVQN1_5_r_6,P6_5_r_6;
wire G42_1_r_16,n_572_1_r_16,n_573_1_r_16,n_549_1_r_16,n_569_1_r_16,n_452_1_r_16,G199_4_r_16,G214_4_r_16,ACVQN1_5_r_16,P6_5_r_16,n4_1_l_16,n29_16,n16_internal_16,n16_16,ACVQN1_3_l_16,n4_1_r_16,N1_4_r_16,n6_16,n_573_1_l_16,n_452_1_l_16,P6_5_r_internal_16,n18_16,n19_16,n20_16,n21_16,n22_16,n23_16,n24_16,n25_16,n26_16,n27_16,n28_16,N3_2_l_6,n4_6,n27_6,n17_6,n28_6,n26_6,N1_4_l_6,n29_6,n18_6,G214_4_l_6,n12_6,n4_1_r_6,N1_4_r_6,n_42_2_l_6,P6_5_r_internal_6,n19_6,n20_6,n21_6,n22_6,n23_6,n24_6,n25_6;
DFFARX1 I_0(n4_1_r_16,blif_clk_net_1_r_6,n4_6,G42_1_r_16,);
nor I_1(n_572_1_r_16,n20_16,n21_16);
nand I_2(n_573_1_r_16,n18_16,n19_16);
nor I_3(n_549_1_r_16,n23_16,n24_16);
nand I_4(n_569_1_r_16,n18_16,n22_16);
nor I_5(n_452_1_r_16,n29_16,n6_16);
DFFARX1 I_6(N1_4_r_16,blif_clk_net_1_r_6,n4_6,G199_4_r_16,);
DFFARX1 I_7(n6_16,blif_clk_net_1_r_6,n4_6,G214_4_r_16,);
DFFARX1 I_8(n_573_1_l_16,blif_clk_net_1_r_6,n4_6,ACVQN1_5_r_16,);
not I_9(P6_5_r_16,P6_5_r_internal_16);
nor I_10(n4_1_l_16,G18_1_l_16,IN_1_1_l_16);
DFFARX1 I_11(n4_1_l_16,blif_clk_net_1_r_6,n4_6,n29_16,);
DFFARX1 I_12(IN_1_3_l_16,blif_clk_net_1_r_6,n4_6,n16_internal_16,);
not I_13(n16_16,n16_internal_16);
DFFARX1 I_14(IN_2_3_l_16,blif_clk_net_1_r_6,n4_6,ACVQN1_3_l_16,);
nor I_15(n4_1_r_16,n29_16,n21_16);
nor I_16(N1_4_r_16,n27_16,n28_16);
not I_17(n6_16,n19_16);
or I_18(n_573_1_l_16,IN_5_1_l_16,IN_9_1_l_16);
nor I_19(n_452_1_l_16,G18_1_l_16,IN_5_1_l_16);
DFFARX1 I_20(n_452_1_l_16,blif_clk_net_1_r_6,n4_6,P6_5_r_internal_16,);
not I_21(n18_16,n20_16);
nor I_22(n19_16,IN_9_1_l_16,IN_10_1_l_16);
nor I_23(n20_16,G15_1_l_16,IN_7_1_l_16);
nor I_24(n21_16,IN_10_1_l_16,n25_16);
nand I_25(n22_16,IN_4_3_l_16,ACVQN1_3_l_16);
not I_26(n23_16,n22_16);
nor I_27(n24_16,n16_16,n20_16);
nor I_28(n25_16,G15_1_l_16,n26_16);
not I_29(n26_16,IN_4_1_l_16);
and I_30(n27_16,IN_9_1_l_16,n29_16);
not I_31(n28_16,n_452_1_l_16);
DFFARX1 I_32(n4_1_r_6,blif_clk_net_1_r_6,n4_6,G42_1_r_6,);
nor I_33(n_572_1_r_6,n27_6,n28_6);
nand I_34(n_573_1_r_6,n18_6,n19_6);
nor I_35(n_549_1_r_6,n_42_2_l_6,n21_6);
nand I_36(n_569_1_r_6,n19_6,n20_6);
nor I_37(n_452_1_r_6,n28_6,n29_6);
DFFARX1 I_38(N1_4_r_6,blif_clk_net_1_r_6,n4_6,G199_4_r_6,);
DFFARX1 I_39(n_42_2_l_6,blif_clk_net_1_r_6,n4_6,G214_4_r_6,);
DFFARX1 I_40(n_42_2_l_6,blif_clk_net_1_r_6,n4_6,ACVQN1_5_r_6,);
not I_41(P6_5_r_6,P6_5_r_internal_6);
and I_42(N3_2_l_6,n23_6,G199_4_r_16);
not I_43(n4_6,blif_reset_net_1_r_6);
DFFARX1 I_44(N3_2_l_6,blif_clk_net_1_r_6,n4_6,n27_6,);
not I_45(n17_6,n27_6);
DFFARX1 I_46(n_573_1_r_16,blif_clk_net_1_r_6,n4_6,n28_6,);
DFFARX1 I_47(P6_5_r_16,blif_clk_net_1_r_6,n4_6,n26_6,);
and I_48(N1_4_l_6,n25_6,G42_1_r_16);
DFFARX1 I_49(N1_4_l_6,blif_clk_net_1_r_6,n4_6,n29_6,);
not I_50(n18_6,n29_6);
DFFARX1 I_51(n_452_1_r_16,blif_clk_net_1_r_6,n4_6,G214_4_l_6,);
not I_52(n12_6,G214_4_l_6);
nor I_53(n4_1_r_6,n28_6,n22_6);
nor I_54(N1_4_r_6,n12_6,n24_6);
nor I_55(n_42_2_l_6,n_569_1_r_16,G42_1_r_16);
DFFARX1 I_56(G214_4_l_6,blif_clk_net_1_r_6,n4_6,P6_5_r_internal_6,);
nand I_57(n19_6,n26_6,n_549_1_r_16);
not I_58(n20_6,n_42_2_l_6);
nor I_59(n21_6,n17_6,n28_6);
and I_60(n22_6,n26_6,n_549_1_r_16);
nand I_61(n23_6,n_572_1_r_16,n_569_1_r_16);
nor I_62(n24_6,n17_6,n18_6);
nand I_63(n25_6,G214_4_r_16,ACVQN1_5_r_16);
endmodule


