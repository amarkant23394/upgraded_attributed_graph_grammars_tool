module test_I10797(I9754,I9816,I9559,I8178,I10797);
input I9754,I9816,I9559,I8178;
output I10797;
wire I9477,I10766,I9771,I9833;
nor I_0(I9477,I9771,I9833);
not I_1(I10797,I10766);
not I_2(I10766,I9477);
and I_3(I9771,I9754,I8178);
and I_4(I9833,I9816,I9559);
endmodule


