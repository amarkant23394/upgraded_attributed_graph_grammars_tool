module test_I6062(I2167,I1477,I5994,I4578,I2173,I1470,I6062);
input I2167,I1477,I5994,I4578,I2173,I1470;
output I6062;
wire I4629,I6045,I6028,I4595,I4544,I4869,I2149,I4527,I5932,I4536,I6011,I5751,I4521,I5915,I5864,I4515;
nor I_0(I4629,I2167,I2173);
nor I_1(I6045,I6028,I5932);
DFFARX1 I_2(I6011,I1470,I5751,,,I6028,);
DFFARX1 I_3(I4578,I1470,I4544,,,I4595,);
not I_4(I4544,I1477);
DFFARX1 I_5(I2149,I1470,I4544,,,I4869,);
DFFARX1 I_6(I1470,,,I2149,);
or I_7(I4527,I4629,I4595);
not I_8(I5932,I5915);
and I_9(I6062,I5864,I6045);
nor I_10(I4536,I4869,I4595);
and I_11(I6011,I5994,I4521);
not I_12(I5751,I1477);
DFFARX1 I_13(I1470,I4544,,,I4521,);
DFFARX1 I_14(I4527,I1470,I5751,,,I5915,);
nor I_15(I5864,I4536,I4515);
not I_16(I4515,I4629);
endmodule


