// Verilog
// c880
// Ninputs 60
// Noutputs 26
// NtotalGates 383

module c880(G1,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G2,G20,G21,G22,G23,G24,G25,G26,G27,G28,G29,G3,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,G4,G40,G41,G42,G43,G44,G45,G46,G47,G48,G49,G5,G50,G51,G52,G53,G54,G55,G56,G57,G58,G59,G6,G60,G7,G8,G855,G856,G857,G858,G859,G860,G861,G862,G863,G864,G865,G866,G867,G868,G869,G870,G871,G872,G873,G874,G875,G876,G877,G878,G879,G880,G9);
input G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,G40,G41,G42,G43,G44,G45,G46,G47,G48,G49,G50,G51,G52,G53,G54,G55,G56,G57,G58,G59,G60;
output G855,G856,G857,G858,G859,G860,G861,G862,G863,G864,G865,G866,G867,G868,G869,G870,G871,G872,G873,G874,G875,G876,G877,G878,G879,G880;

wire G269,G270,G273,G276,G279,G280,G284,G285,G286,G287,G290,G291,G292,G293,G294,G295,G296,G297,G298,G301,G302,G303,G304,G305,G306,G307,G308,G309,G310,G316,G317,G318,G319,G322,G323,G324,G325,G326,G327,G328,G329,G330,G331,G332,G333,G334,G335,G336,G337,G338,G339,G340,G341,G342,G343,G344,G345,G346,G347,G348,G349,G350,G351,G352,G353,G354,G355,G356,G357,G360,G363,G366,G369,G375,G376,G379,G382,G385,G388,G389,G395,G396,G397,G398,G399,G400,G401,G402,G403,G404,G405,G406,G407,G408,G409,G410,G411,G412,G413,G414,G415,G416,G417,G422,G427,G432,G433,G434,G435,G436,G445,G448,G451,G460,G461,G462,G463,G464,G465,G466,G467,G468,G473,G474,G475,G476,G477,G480,G483,G484,G485,G486,G487,G488,G489,G490,G491,G492,G493,G494,G495,G496,G497,G498,G499,G500,G501,G502,G503,G504,G505,G506,G507,G508,G509,G510,G511,G512,G513,G514,G515,G518,G521,G522,G523,G524,G525,G526,G527,G528,G529,G532,G535,G536,G537,G538,G542,G546,G550,G554,G558,G562,G566,G570,G571,G572,G573,G574,G575,G578,G581,G582,G585,G590,G591,G594,G600,G601,G604,G609,G610,G613,G616,G617,G620,G625,G626,G629,G635,G636,G639,G644,G645,G646,G647,G650,G654,G655,G658,G662,G663,G667,G671,G672,G677,G681,G682,G685,G689,G690,G693,G697,G698,G702,G706,G707,G712,G716,G717,G718,G719,G720,G721,G722,G723,G724,G725,G726,G727,G728,G729,G730,G731,G732,G733,G734,G735,G736,G737,G738,G739,G740,G741,G742,G743,G744,G745,G746,G747,G748,G749,G750,G751,G752,G753,G754,G755,G756,G760,G761,G764,G765,G768,G769,G770,G771,G772,G773,G774,G775,G776,G777,G778,G779,G785,G786,G787,G788,G789,G790,G791,G792,G793,G794,G795,G796,G797,G798,G802,G805,G808,G809,G810,G811,G812,G813,G814,G815,G816,G817,G818,G819,G820,G821,G822,G823,G824,G825,G826,G827,G828,G829,G830,G831,G832,G833,G834,G835,G836,G837,G838,G839,G840,G841,G842,G843,G844,G845,G846,G847,G848,G849,G850,G851,G852,G853,G854;

nand NAND4_0(G269,G1,G2,G3,G4);
nand NAND4_1(G270,G1,G5,G3,G4);
and AND3_0(G273,G6,G7,G8);
and AND3_1(G276,G1,G5,G9);
nand NAND4_2(G279,G1,G2,G9,G4);
nand NAND4_3(G280,G1,G2,G3,G10);
nand NAND4_4(G284,G11,G8,G12,G13);
nand NAND2_0(G285,G6,G12);
nand NAND3_0(G286,G11,G12,G15);
and AND3_2(G287,G6,G16,G17);
and AND3_3(G290,G6,G16,G8);
and AND3_4(G291,G6,G7,G17);
and AND3_5(G292,G6,G7,G8);
and AND3_6(G293,G11,G16,G17);
and AND3_7(G294,G11,G16,G8);
and AND3_8(G295,G11,G7,G17);
and AND3_9(G296,G11,G7,G8);
and AND2_0(G297,G18,G19);
or OR2_0(G298,G20,G21);
nand NAND2_1(G301,G24,G25);
or OR2_1(G302,G24,G25);
nand NAND2_2(G303,G26,G27);
or OR2_2(G304,G26,G27);
nand NAND2_3(G305,G28,G29);
or OR2_3(G306,G28,G29);
nand NAND2_4(G307,G30,G31);
or OR2_4(G308,G30,G31);
and AND2_1(G309,G2,G34);
not NOT_0(G310,G60);
and AND2_2(G316,G9,G34);
and AND2_3(G317,G4,G34);
and AND2_4(G318,G38,G34);
nand NAND2_5(G319,G11,G40);
nor NOR2_0(G322,G4,G8);
and AND2_5(G323,G4,G8);
nand NAND2_6(G324,G41,G42);
or OR2_5(G325,G41,G42);
nand NAND2_7(G326,G43,G44);
or OR2_6(G327,G43,G44);
nand NAND2_8(G328,G45,G46);
or OR2_7(G329,G45,G46);
nand NAND2_9(G330,G47,G48);
or OR2_8(G331,G47,G48);
and AND2_6(G332,G50,G24);
and AND2_7(G333,G50,G25);
and AND2_8(G334,G50,G26);
and AND2_9(G335,G50,G27);
and AND2_10(G336,G50,G28);
and AND2_11(G337,G55,G56);
and AND2_12(G338,G50,G29);
and AND2_13(G339,G55,G57);
and AND2_14(G340,G50,G30);
and AND2_15(G341,G55,G59);
not NOT_1(G342,G269);
not NOT_2(G343,G273);
or OR2_9(G344,G270,G273);
not NOT_3(G345,G276);
not NOT_4(G346,G276);
not NOT_5(G347,G279);
nor NOR2_1(G348,G280,G284);
or OR2_10(G349,G280,G285);
or OR2_11(G350,G280,G286);
not NOT_6(G351,G293);
not NOT_7(G352,G294);
not NOT_8(G353,G295);
not NOT_9(G354,G296);
nand NAND2_10(G355,G22,G298);
and AND2_16(G356,G23,G298);
nand NAND2_11(G357,G301,G302);
nand NAND2_12(G360,G303,G304);
nand NAND2_13(G363,G305,G306);
nand NAND2_14(G366,G307,G308);
not NOT_10(G369,G310);
nor NOR2_2(G375,G322,G323);
nand NAND2_15(G376,G324,G325);
nand NAND2_16(G379,G326,G327);
nand NAND2_17(G382,G328,G329);
nand NAND2_18(G385,G330,G331);
or OR2_12(G388,G270,G343);
not NOT_11(G389,G345);
not NOT_12(G395,G346);
and AND2_17(G396,G348,G14);
not NOT_13(G397,G349);
not NOT_14(G398,G350);
not NOT_15(G399,G355);
not NOT_16(G400,G357);
not NOT_17(G401,G360);
and AND2_18(G402,G357,G360);
not NOT_18(G403,G363);
not NOT_19(G404,G366);
and AND2_19(G405,G363,G366);
nand NAND2_19(G406,G347,G352);
not NOT_20(G407,G376);
not NOT_21(G408,G379);
and AND2_20(G409,G376,G379);
not NOT_22(G410,G382);
not NOT_23(G411,G385);
and AND2_21(G412,G382,G385);
and AND2_22(G413,G50,G369);
not NOT_24(G414,G396);
and AND2_23(G415,G400,G401);
and AND2_24(G416,G403,G404);
and AND3_10(G417,G319,G389,G10);
and AND3_11(G422,G389,G4,G287);
nand NAND3_1(G427,G389,G287,G10);
nand NAND4_5(G432,G375,G11,G40,G389);
nand NAND3_2(G433,G389,G319,G4);
and AND2_25(G434,G407,G408);
and AND2_26(G435,G410,G411);
not NOT_25(G436,G414);
nor NOR2_3(G445,G402,G415);
nor NOR2_4(G448,G405,G416);
nand NAND2_20(G451,G432,G406);
and AND2_27(G460,G35,G417);
and AND2_28(G461,G310,G422);
and AND2_29(G462,G36,G417);
and AND2_30(G463,G310,G422);
and AND2_31(G464,G37,G417);
and AND2_32(G465,G310,G422);
and AND2_33(G466,G39,G417);
and AND2_34(G467,G310,G422);
nand NAND2_21(G468,G433,G1);
or OR2_13(G473,G369,G427);
or OR2_14(G474,G369,G427);
or OR2_15(G475,G369,G427);
or OR2_16(G476,G369,G427);
nor NOR2_5(G477,G409,G434);
nor NOR2_6(G480,G412,G435);
nand NAND2_22(G483,G32,G445);
or OR2_17(G484,G32,G445);
nand NAND2_23(G485,G448,G33);
or OR2_18(G486,G448,G33);
and AND2_35(G487,G24,G451);
nor NOR2_7(G488,G460,G461);
and AND2_36(G489,G25,G451);
nor NOR2_8(G490,G462,G463);
and AND2_37(G491,G26,G451);
nor NOR2_9(G492,G464,G465);
and AND2_38(G493,G27,G451);
nor NOR2_10(G494,G466,G467);
and AND2_39(G495,G35,G468);
and AND2_40(G496,G28,G451);
and AND2_41(G497,G36,G468);
and AND2_42(G498,G29,G451);
and AND2_43(G499,G37,G468);
and AND2_44(G500,G30,G451);
and AND2_45(G501,G39,G468);
and AND2_46(G502,G31,G451);
nand NAND2_24(G503,G32,G477);
or OR2_19(G504,G32,G477);
nand NAND2_25(G505,G480,G49);
or OR2_20(G506,G480,G49);
and AND2_47(G507,G436,G41);
and AND2_48(G508,G436,G42);
and AND2_49(G509,G436,G43);
and AND2_50(G510,G436,G44);
and AND2_51(G511,G436,G45);
nand NAND2_26(G512,G436,G46);
nand NAND2_27(G513,G436,G47);
nand NAND2_28(G514,G436,G48);
nand NAND2_29(G515,G483,G484);
nand NAND2_30(G518,G485,G486);
nor NOR2_11(G521,G309,G487);
nor NOR2_12(G522,G316,G489);
nor NOR2_13(G523,G317,G491);
nor NOR2_14(G524,G318,G493);
nor NOR2_15(G525,G495,G496);
nor NOR2_16(G526,G497,G498);
nor NOR2_17(G527,G499,G500);
nor NOR2_18(G528,G501,G502);
nand NAND2_31(G529,G503,G504);
nand NAND2_32(G532,G505,G506);
not NOT_26(G535,G515);
not NOT_27(G536,G518);
and AND2_52(G537,G515,G518);
nand NAND2_33(G538,G521,G488);
nand NAND2_34(G542,G522,G490);
nand NAND2_35(G546,G523,G492);
nand NAND2_36(G550,G524,G494);
nand NAND2_37(G554,G473,G525);
nand NAND2_38(G558,G474,G526);
nand NAND2_39(G562,G475,G527);
nand NAND2_40(G566,G476,G528);
not NOT_28(G570,G529);
not NOT_29(G571,G532);
and AND2_53(G572,G529,G532);
and AND2_54(G573,G535,G536);
and AND2_55(G574,G570,G571);
nand NAND2_41(G575,G538,G41);
or OR2_21(G578,G538,G41);
and AND2_56(G581,G54,G538);
nand NAND2_42(G582,G542,G42);
or OR2_22(G585,G542,G42);
and AND2_57(G590,G54,G542);
nand NAND2_43(G591,G546,G43);
or OR2_23(G594,G546,G43);
and AND2_58(G600,G54,G546);
nand NAND2_44(G601,G550,G44);
or OR2_24(G604,G550,G44);
and AND2_59(G609,G54,G550);
nand NAND2_45(G610,G554,G45);
or OR2_25(G613,G554,G45);
and AND2_60(G616,G54,G554);
nand NAND2_46(G617,G558,G46);
or OR2_26(G620,G558,G46);
and AND2_61(G625,G54,G558);
nand NAND2_47(G626,G562,G47);
or OR2_27(G629,G562,G47);
and AND2_62(G635,G54,G562);
nand NAND2_48(G636,G566,G48);
or OR2_28(G639,G566,G48);
and AND2_63(G644,G54,G566);
nor NOR2_19(G645,G537,G573);
nor NOR2_20(G646,G572,G574);
not NOT_30(G647,G575);
and AND2_64(G650,G578,G575);
nor NOR2_21(G654,G581,G507);
not NOT_31(G655,G582);
and AND2_65(G658,G585,G582);
nor NOR2_22(G662,G590,G508);
not NOT_32(G663,G591);
and AND2_66(G667,G594,G591);
nor NOR2_23(G671,G600,G509);
not NOT_33(G672,G601);
and AND2_67(G677,G604,G601);
nor NOR2_24(G681,G609,G510);
not NOT_34(G682,G610);
and AND2_68(G685,G613,G610);
nor NOR2_25(G689,G616,G511);
not NOT_35(G690,G617);
and AND2_69(G693,G620,G617);
nor NOR2_26(G697,G337,G625);
not NOT_36(G698,G626);
and AND2_70(G702,G629,G626);
nor NOR2_27(G706,G339,G635);
not NOT_37(G707,G636);
and AND2_71(G712,G639,G636);
nor NOR2_28(G716,G341,G644);
nand NAND2_49(G717,G639,G58);
nand NAND3_3(G718,G629,G639,G58);
nand NAND4_6(G719,G620,G629,G639,G58);
not NOT_38(G720,G647);
and AND2_72(G721,G52,G650);
and AND2_73(G722,G53,G647);
not NOT_39(G723,G655);
and AND2_74(G724,G52,G658);
and AND2_75(G725,G53,G655);
not NOT_40(G726,G663);
and AND2_76(G727,G52,G667);
and AND2_77(G728,G53,G663);
not NOT_41(G729,G672);
and AND2_78(G730,G52,G677);
and AND2_79(G731,G53,G672);
not NOT_42(G732,G682);
and AND2_80(G733,G52,G685);
and AND2_81(G734,G53,G682);
not NOT_43(G735,G690);
and AND2_82(G736,G52,G693);
and AND2_83(G737,G53,G690);
not NOT_44(G738,G698);
and AND2_84(G739,G52,G702);
and AND2_85(G740,G53,G698);
not NOT_45(G741,G707);
nor NOR2_29(G742,G712,G58);
and AND2_86(G743,G712,G58);
and AND2_87(G744,G52,G712);
and AND2_88(G745,G53,G707);
nand NAND2_50(G746,G629,G707);
nand NAND2_51(G747,G620,G698);
nand NAND3_4(G748,G620,G629,G707);
nand NAND2_52(G749,G594,G672);
nand NAND2_53(G750,G585,G663);
nand NAND3_5(G751,G585,G594,G672);
nor NOR2_30(G752,G721,G722);
nor NOR2_31(G753,G724,G725);
nor NOR2_32(G754,G727,G728);
nor NOR2_33(G755,G730,G731);
nand NAND4_7(G756,G735,G747,G748,G719);
nor NOR2_34(G760,G733,G734);
nand NAND3_6(G761,G738,G746,G718);
nor NOR2_35(G764,G736,G737);
nand NAND2_54(G765,G741,G717);
nor NOR2_36(G768,G739,G740);
nor NOR2_37(G769,G742,G743);
nor NOR2_38(G770,G744,G745);
nor NOR2_39(G771,G685,G756);
and AND2_89(G772,G685,G756);
nor NOR2_40(G773,G693,G761);
and AND2_90(G774,G693,G761);
nor NOR2_41(G775,G702,G765);
and AND2_91(G776,G702,G765);
and AND2_92(G777,G51,G769);
nand NAND2_55(G778,G613,G756);
nand NAND2_56(G779,G778,G732);
nor NOR2_42(G785,G771,G772);
nor NOR2_43(G786,G773,G774);
nor NOR2_44(G787,G775,G776);
nor NOR2_45(G788,G340,G777);
nor NOR2_46(G789,G677,G779);
and AND2_93(G790,G677,G779);
and AND2_94(G791,G51,G785);
and AND2_95(G792,G51,G786);
and AND2_96(G793,G51,G787);
nand NAND4_8(G794,G788,G770,G716,G514);
nand NAND2_57(G795,G604,G779);
nand NAND3_7(G796,G594,G604,G779);
nand NAND4_9(G797,G585,G594,G604,G779);
nand NAND4_10(G798,G723,G750,G751,G797);
nand NAND3_8(G802,G726,G749,G796);
nand NAND2_58(G805,G729,G795);
nor NOR2_47(G808,G789,G790);
nor NOR2_48(G809,G335,G791);
nor NOR2_49(G810,G336,G792);
nor NOR2_50(G811,G338,G793);
not NOT_46(G812,G794);
nor NOR2_51(G813,G650,G798);
and AND2_97(G814,G650,G798);
nor NOR2_52(G815,G658,G802);
and AND2_98(G816,G658,G802);
nor NOR2_53(G817,G667,G805);
and AND2_99(G818,G667,G805);
and AND2_100(G819,G51,G808);
nand NAND3_9(G820,G809,G760,G689);
nand NAND4_11(G821,G810,G764,G697,G512);
nand NAND4_12(G822,G811,G768,G706,G513);
not NOT_47(G823,G812);
nand NAND2_59(G824,G798,G578);
nor NOR2_54(G825,G813,G814);
nor NOR2_55(G826,G815,G816);
nor NOR2_56(G827,G817,G818);
nor NOR2_57(G828,G334,G819);
not NOT_48(G829,G820);
not NOT_49(G830,G821);
not NOT_50(G831,G822);
and AND2_101(G832,G720,G824);
and AND2_102(G833,G51,G825);
and AND2_103(G834,G51,G826);
and AND2_104(G835,G51,G827);
nand NAND3_10(G836,G828,G755,G681);
not NOT_51(G837,G829);
not NOT_52(G838,G830);
not NOT_53(G839,G831);
not NOT_54(G840,G832);
nor NOR2_58(G841,G413,G833);
nor NOR2_59(G842,G332,G834);
nor NOR2_60(G843,G333,G835);
not NOT_55(G844,G836);
nand NAND3_11(G845,G841,G752,G654);
nand NAND3_12(G846,G842,G753,G662);
nand NAND3_13(G847,G843,G754,G671);
not NOT_56(G848,G844);
not NOT_57(G849,G845);
not NOT_58(G850,G846);
not NOT_59(G851,G847);
not NOT_60(G852,G849);
not NOT_61(G853,G850);
not NOT_62(G854,G851);
not NOT_63(G855,G290);
not NOT_64(G856,G291);
not NOT_65(G857,G292);
not NOT_66(G858,G297);
not NOT_67(G859,G342);
not NOT_68(G860,G344);
not NOT_69(G861,G351);
not NOT_70(G862,G353);
not NOT_71(G863,G354);
not NOT_72(G864,G356);
not NOT_73(G865,G388);
not NOT_74(G866,G395);
not NOT_75(G867,G397);
not NOT_76(G868,G398);
not NOT_77(G869,G399);
not NOT_78(G870,G645);
not NOT_79(G871,G646);
not NOT_80(G872,G823);
not NOT_81(G873,G837);
not NOT_82(G874,G838);
not NOT_83(G875,G839);
not NOT_84(G876,G840);
not NOT_85(G877,G848);
not NOT_86(G878,G852);
not NOT_87(G879,G853);
not NOT_88(G880,G854);

endmodule