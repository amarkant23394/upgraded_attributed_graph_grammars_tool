module test_I13826(I12442,I1477,I1470,I13826);
input I12442,I1477,I1470;
output I13826;
wire I11947,I12541,I12304,I11953,I13792,I10020,I13809,I13775,I12106,I11965,I12524,I11973;
DFFARX1 I_0(I13809,I1470,I13775,,,I13826,);
nand I_1(I11947,I12106,I12524);
nor I_2(I12541,I12524);
and I_3(I12304,I12106);
nand I_4(I11953,I12442,I12541);
nand I_5(I13792,I11953,I11965);
DFFARX1 I_6(I1470,,,I10020,);
and I_7(I13809,I13792,I11947);
not I_8(I13775,I1477);
not I_9(I12106,I10020);
DFFARX1 I_10(I12304,I1470,I11973,,,I11965,);
not I_11(I12524,I12442);
not I_12(I11973,I1477);
endmodule


