module test_I8298(I5864,I6011,I1477,I4527,I1470,I8298);
input I5864,I6011,I1477,I4527,I1470;
output I8298;
wire I8233,I6265,I6248,I5751,I6028,I6203,I5915,I5719,I5722;
not I_0(I8233,I5722);
and I_1(I6265,I5915,I6248);
nand I_2(I6248,I6203,I5864);
not I_3(I5751,I1477);
DFFARX1 I_4(I6011,I1470,I5751,,,I6028,);
DFFARX1 I_5(I1470,I5751,,,I6203,);
DFFARX1 I_6(I4527,I1470,I5751,,,I5915,);
nor I_7(I8298,I8233,I5719);
DFFARX1 I_8(I6265,I1470,I5751,,,I5719,);
DFFARX1 I_9(I6028,I1470,I5751,,,I5722,);
endmodule


