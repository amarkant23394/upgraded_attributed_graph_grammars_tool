module test_final(IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_6_2_l_10,IN_1_3_l_10,IN_2_3_l_10,IN_4_3_l_10,IN_1_4_l_10,IN_2_4_l_10,IN_3_4_l_10,IN_6_4_l_10,blif_clk_net_1_r_13,blif_reset_net_1_r_13,G42_1_r_13,n_572_1_r_13,n_573_1_r_13,n_549_1_r_13,n_452_1_r_13,ACVQN2_3_r_13,n_266_and_0_3_r_13,ACVQN1_5_r_13,P6_5_r_13);
input IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_6_2_l_10,IN_1_3_l_10,IN_2_3_l_10,IN_4_3_l_10,IN_1_4_l_10,IN_2_4_l_10,IN_3_4_l_10,IN_6_4_l_10,blif_clk_net_1_r_13,blif_reset_net_1_r_13;
output G42_1_r_13,n_572_1_r_13,n_573_1_r_13,n_549_1_r_13,n_452_1_r_13,ACVQN2_3_r_13,n_266_and_0_3_r_13,ACVQN1_5_r_13,P6_5_r_13;
wire G42_1_r_10,n_572_1_r_10,n_573_1_r_10,n_549_1_r_10,n_452_1_r_10,n_42_2_r_10,G199_2_r_10,ACVQN2_3_r_10,n_266_and_0_3_r_10,N3_2_l_10,n25_10,n16_10,n26_10,ACVQN1_3_l_10,N1_4_l_10,G199_4_l_10,n27_10,n17_10,n4_1_r_10,N3_2_r_10,n3_10,n13_internal_10,n13_10,n18_10,n19_10,n20_10,n21_10,n22_10,n23_10,n24_10,n_569_1_r_13,n4_1_l_13,n7_13,n17_internal_13,n17_13,n28_13,ACVQN1_3_l_13,n4_1_r_13,n_266_and_0_3_l_13,n_573_1_l_13,n14_internal_13,n14_13,n_549_1_l_13,n_569_1_l_13,P6_5_r_internal_13,n18_13,n19_13,n20_13,n21_13,n22_13,n23_13,n24_13,n25_13,n26_13,n27_13;
DFFARX1 I_0(n4_1_r_10,blif_clk_net_1_r_13,n7_13,G42_1_r_10,);
nor I_1(n_572_1_r_10,n26_10,n3_10);
nand I_2(n_573_1_r_10,n16_10,n18_10);
nand I_3(n_549_1_r_10,n19_10,n20_10);
nor I_4(n_452_1_r_10,n25_10,n21_10);
nor I_5(n_42_2_r_10,n26_10,G199_4_l_10);
DFFARX1 I_6(N3_2_r_10,blif_clk_net_1_r_13,n7_13,G199_2_r_10,);
DFFARX1 I_7(G199_4_l_10,blif_clk_net_1_r_13,n7_13,ACVQN2_3_r_10,);
nor I_8(n_266_and_0_3_r_10,n17_10,n13_10);
and I_9(N3_2_l_10,IN_6_2_l_10,n23_10);
DFFARX1 I_10(N3_2_l_10,blif_clk_net_1_r_13,n7_13,n25_10,);
not I_11(n16_10,n25_10);
DFFARX1 I_12(IN_1_3_l_10,blif_clk_net_1_r_13,n7_13,n26_10,);
DFFARX1 I_13(IN_2_3_l_10,blif_clk_net_1_r_13,n7_13,ACVQN1_3_l_10,);
and I_14(N1_4_l_10,IN_6_4_l_10,n24_10);
DFFARX1 I_15(N1_4_l_10,blif_clk_net_1_r_13,n7_13,G199_4_l_10,);
DFFARX1 I_16(IN_3_4_l_10,blif_clk_net_1_r_13,n7_13,n27_10,);
not I_17(n17_10,n27_10);
nor I_18(n4_1_r_10,n27_10,n21_10);
nor I_19(N3_2_r_10,n16_10,n22_10);
not I_20(n3_10,n18_10);
DFFARX1 I_21(n3_10,blif_clk_net_1_r_13,n7_13,n13_internal_10,);
not I_22(n13_10,n13_internal_10);
nand I_23(n18_10,IN_4_3_l_10,ACVQN1_3_l_10);
not I_24(n19_10,n_452_1_r_10);
nand I_25(n20_10,n16_10,n26_10);
nor I_26(n21_10,IN_1_2_l_10,IN_3_2_l_10);
and I_27(n22_10,n26_10,n21_10);
nand I_28(n23_10,IN_2_2_l_10,IN_3_2_l_10);
nand I_29(n24_10,IN_1_4_l_10,IN_2_4_l_10);
DFFARX1 I_30(n4_1_r_13,blif_clk_net_1_r_13,n7_13,G42_1_r_13,);
nor I_31(n_572_1_r_13,n28_13,n_569_1_l_13);
nand I_32(n_573_1_r_13,n18_13,n19_13);
nand I_33(n_549_1_r_13,n_569_1_r_13,n22_13);
nand I_34(n_569_1_r_13,n17_13,n18_13);
nor I_35(n_452_1_r_13,n_573_1_l_13,n25_13);
DFFARX1 I_36(n_266_and_0_3_l_13,blif_clk_net_1_r_13,n7_13,ACVQN2_3_r_13,);
nor I_37(n_266_and_0_3_r_13,n17_13,n14_13);
DFFARX1 I_38(n_549_1_l_13,blif_clk_net_1_r_13,n7_13,ACVQN1_5_r_13,);
not I_39(P6_5_r_13,P6_5_r_internal_13);
nor I_40(n4_1_l_13,n_573_1_r_10,n_549_1_r_10);
not I_41(n7_13,blif_reset_net_1_r_13);
DFFARX1 I_42(n4_1_l_13,blif_clk_net_1_r_13,n7_13,n17_internal_13,);
not I_43(n17_13,n17_internal_13);
DFFARX1 I_44(G199_2_r_10,blif_clk_net_1_r_13,n7_13,n28_13,);
DFFARX1 I_45(n_572_1_r_10,blif_clk_net_1_r_13,n7_13,ACVQN1_3_l_13,);
nor I_46(n4_1_r_13,n_573_1_l_13,n_549_1_l_13);
and I_47(n_266_and_0_3_l_13,ACVQN1_3_l_13,n_549_1_r_10);
nand I_48(n_573_1_l_13,n20_13,n24_13);
DFFARX1 I_49(n_573_1_l_13,blif_clk_net_1_r_13,n7_13,n14_internal_13,);
not I_50(n14_13,n14_internal_13);
and I_51(n_549_1_l_13,n21_13,n26_13);
nand I_52(n_569_1_l_13,n20_13,n21_13);
DFFARX1 I_53(n_569_1_l_13,blif_clk_net_1_r_13,n7_13,P6_5_r_internal_13,);
nand I_54(n18_13,n23_13,n24_13);
or I_55(n19_13,n_42_2_r_10,n_266_and_0_3_r_10);
not I_56(n20_13,G42_1_r_10);
not I_57(n21_13,G42_1_r_10);
nand I_58(n22_13,n17_13,n28_13);
not I_59(n23_13,n_573_1_r_10);
not I_60(n24_13,ACVQN2_3_r_10);
nor I_61(n25_13,n_42_2_r_10,n_266_and_0_3_r_10);
nand I_62(n26_13,n27_13,n_572_1_r_10);
not I_63(n27_13,n_42_2_r_10);
endmodule


