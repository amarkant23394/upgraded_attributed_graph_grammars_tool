module test_final(IN_1_2_l_0,IN_2_2_l_0,IN_3_2_l_0,IN_4_2_l_0,IN_5_2_l_0,IN_1_4_l_0,IN_2_4_l_0,IN_3_4_l_0,IN_4_4_l_0,IN_5_4_l_0,IN_1_9_l_0,IN_2_9_l_0,IN_3_9_l_0,IN_4_9_l_0,IN_5_9_l_0,blif_clk_net_7_r_2,blif_reset_net_7_r_2,N1371_0_r_2,N1508_0_r_2,N1372_1_r_2,N1508_1_r_2,N6147_2_r_2,N1507_6_r_2,N1508_6_r_2,G42_7_r_2,n_572_7_r_2,n_573_7_r_2,n_549_7_r_2,n_569_7_r_2,n_452_7_r_2);
input IN_1_2_l_0,IN_2_2_l_0,IN_3_2_l_0,IN_4_2_l_0,IN_5_2_l_0,IN_1_4_l_0,IN_2_4_l_0,IN_3_4_l_0,IN_4_4_l_0,IN_5_4_l_0,IN_1_9_l_0,IN_2_9_l_0,IN_3_9_l_0,IN_4_9_l_0,IN_5_9_l_0,blif_clk_net_7_r_2,blif_reset_net_7_r_2;
output N1371_0_r_2,N1508_0_r_2,N1372_1_r_2,N1508_1_r_2,N6147_2_r_2,N1507_6_r_2,N1508_6_r_2,G42_7_r_2,n_572_7_r_2,n_573_7_r_2,n_549_7_r_2,n_569_7_r_2,n_452_7_r_2;
wire N1371_0_r_0,N1508_0_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_102_5_r_0,n_547_5_r_0,G42_7_r_0,n_572_7_r_0,n_573_7_r_0,n_549_7_r_0,n_569_7_r_0,n_452_7_r_0,n_431_5_r_0,n4_7_r_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0,n37_0,n38_0,n39_0,n40_0,n41_0,n42_0,n43_0,n44_0,n45_0,n4_7_l_2,n10_2,n59_2,n33_2,N3_8_l_2,n32_internal_2,n32_2,n4_7_r_2,n34_2,n35_2,n36_2,n37_2,n38_2,n39_2,n40_2,n41_2,n42_2,n43_2,n44_2,n45_2,n46_2,n47_2,n48_2,n49_2,n50_2,n51_2,n52_2,n53_2,n54_2,n55_2,n56_2,n57_2,n58_2;
nor I_0(N1371_0_r_0,n_102_5_r_0,n29_0);
nor I_1(N1508_0_r_0,n_102_5_r_0,n_452_7_r_0);
or I_2(n_429_or_0_5_r_0,IN_1_9_l_0,n38_0);
DFFARX1 I_3(n_431_5_r_0,blif_clk_net_7_r_2,n10_2,G78_5_r_0,);
nand I_4(n_576_5_r_0,IN_1_9_l_0,n26_0);
not I_5(n_102_5_r_0,n27_0);
nand I_6(n_547_5_r_0,n30_0,n34_0);
DFFARX1 I_7(n4_7_r_0,blif_clk_net_7_r_2,n10_2,G42_7_r_0,);
nor I_8(n_572_7_r_0,IN_1_9_l_0,n31_0);
or I_9(n_573_7_r_0,n29_0,n30_0);
nor I_10(n_549_7_r_0,n29_0,n33_0);
nand I_11(n_569_7_r_0,n28_0,n32_0);
nor I_12(n_452_7_r_0,n30_0,n31_0);
nand I_13(n_431_5_r_0,n_102_5_r_0,n35_0);
nor I_14(n4_7_r_0,n31_0,n37_0);
nor I_15(n26_0,n27_0,n28_0);
nor I_16(n27_0,n28_0,n44_0);
nand I_17(n28_0,IN_1_4_l_0,IN_2_4_l_0);
not I_18(n29_0,n32_0);
nor I_19(n30_0,IN_5_9_l_0,n39_0);
not I_20(n31_0,n38_0);
nand I_21(n32_0,n41_0,n42_0);
nor I_22(n33_0,IN_1_9_l_0,n_102_5_r_0);
nor I_23(n34_0,IN_1_9_l_0,n27_0);
nand I_24(n35_0,n29_0,n36_0);
nor I_25(n36_0,n37_0,n38_0);
not I_26(n37_0,n28_0);
nand I_27(n38_0,IN_2_9_l_0,n40_0);
nor I_28(n39_0,IN_3_9_l_0,IN_4_9_l_0);
or I_29(n40_0,IN_3_9_l_0,IN_4_9_l_0);
nor I_30(n41_0,IN_1_2_l_0,IN_2_2_l_0);
or I_31(n42_0,IN_5_2_l_0,n43_0);
nor I_32(n43_0,IN_3_2_l_0,IN_4_2_l_0);
nor I_33(n44_0,IN_5_4_l_0,n45_0);
and I_34(n45_0,IN_3_4_l_0,IN_4_4_l_0);
nor I_35(N1371_0_r_2,n32_2,n35_2);
nor I_36(N1508_0_r_2,n32_2,n55_2);
not I_37(N1372_1_r_2,n54_2);
nor I_38(N1508_1_r_2,n59_2,n54_2);
nor I_39(N6147_2_r_2,n42_2,n43_2);
nor I_40(N1507_6_r_2,n40_2,n53_2);
nor I_41(N1508_6_r_2,n33_2,n50_2);
DFFARX1 I_42(n4_7_r_2,blif_clk_net_7_r_2,n10_2,G42_7_r_2,);
nor I_43(n_572_7_r_2,n36_2,n37_2);
or I_44(n_573_7_r_2,n34_2,n35_2);
nor I_45(n_549_7_r_2,n40_2,n41_2);
nand I_46(n_569_7_r_2,n38_2,n39_2);
nor I_47(n_452_7_r_2,n59_2,n35_2);
nor I_48(n4_7_l_2,n_573_7_r_0,N1371_0_r_0);
not I_49(n10_2,blif_reset_net_7_r_2);
DFFARX1 I_50(n4_7_l_2,blif_clk_net_7_r_2,n10_2,n59_2,);
not I_51(n33_2,n59_2);
and I_52(N3_8_l_2,n49_2,N1508_0_r_0);
DFFARX1 I_53(N3_8_l_2,blif_clk_net_7_r_2,n10_2,n32_internal_2,);
not I_54(n32_2,n32_internal_2);
nor I_55(n4_7_r_2,n59_2,n36_2);
not I_56(n34_2,n39_2);
nor I_57(n35_2,n_576_5_r_0,n_572_7_r_0);
nor I_58(n36_2,n_429_or_0_5_r_0,n_573_7_r_0);
or I_59(n37_2,n_549_7_r_0,n_429_or_0_5_r_0);
not I_60(n38_2,n40_2);
nand I_61(n39_2,n45_2,n57_2);
nor I_62(n40_2,n47_2,G78_5_r_0);
nor I_63(n41_2,n32_2,n36_2);
not I_64(n42_2,n53_2);
nand I_65(n43_2,n44_2,n45_2);
nand I_66(n44_2,n38_2,n46_2);
not I_67(n45_2,n_429_or_0_5_r_0);
nand I_68(n46_2,n47_2,n48_2);
nand I_69(n47_2,n_547_5_r_0,G42_7_r_0);
or I_70(n48_2,N1371_0_r_0,N1508_0_r_0);
nand I_71(n49_2,n_576_5_r_0,G78_5_r_0);
nand I_72(n50_2,n51_2,n52_2);
not I_73(n51_2,n47_2);
nand I_74(n52_2,n38_2,n53_2);
nor I_75(n53_2,n_429_or_0_5_r_0,n_549_7_r_0);
nand I_76(n54_2,n42_2,n56_2);
nor I_77(n55_2,n34_2,n56_2);
nor I_78(n56_2,N1371_0_r_0,N1508_0_r_0);
nand I_79(n57_2,n58_2,n_569_7_r_0);
not I_80(n58_2,N1371_0_r_0);
endmodule


