module test_I1668(I1215,I1668);
input I1215;
output I1668;
wire I1637;
not I_0(I1637,I1215);
not I_1(I1668,I1637);
endmodule


