module test_I13508(I11361,I11542,I1477,I1470,I11395,I8848,I13508);
input I11361,I11542,I1477,I1470,I11395,I8848;
output I13508;
wire I11672,I11559,I11296,I11429,I13197,I11768,I11272,I11689,I13491,I11310,I11751;
DFFARX1 I_0(I1470,I11310,,,I11672,);
DFFARX1 I_1(I11542,I1470,I11310,,,I11559,);
nand I_2(I11296,I11559,I11689);
not I_3(I11429,I8848);
not I_4(I13197,I1477);
and I_5(I11768,I11429,I11751);
DFFARX1 I_6(I11768,I1470,I11310,,,I11272,);
nor I_7(I11689,I11672,I11395);
and I_8(I13508,I13491,I11272);
DFFARX1 I_9(I11296,I1470,I13197,,,I13491,);
not I_10(I11310,I1477);
nand I_11(I11751,I11672,I11361);
endmodule


