module test_I16792(I1477,I1470,I15126,I16792);
input I1477,I1470,I15126;
output I16792;
wire I14927,I16934,I17205,I14945,I16818,I16951,I14965,I15372,I15485,I15502;
DFFARX1 I_0(I15502,I1470,I14965,,,I14927,);
DFFARX1 I_1(I14945,I1470,I16818,,,I16934,);
nand I_2(I16792,I17205,I16951);
DFFARX1 I_3(I14927,I1470,I16818,,,I17205,);
nand I_4(I14945,I15372,I15126);
not I_5(I16818,I1477);
not I_6(I16951,I16934);
not I_7(I14965,I1477);
DFFARX1 I_8(I1470,I14965,,,I15372,);
DFFARX1 I_9(I1470,I14965,,,I15485,);
not I_10(I15502,I15485);
endmodule


