module test_final(IN_1_0_l_11,IN_2_0_l_11,IN_3_0_l_11,IN_4_0_l_11,IN_1_1_l_11,IN_2_1_l_11,IN_3_1_l_11,IN_1_3_l_11,IN_2_3_l_11,IN_3_3_l_11,IN_1_6_l_11,IN_2_6_l_11,IN_3_6_l_11,IN_4_6_l_11,IN_5_6_l_11,blif_clk_net_5_r_0,blif_reset_net_5_r_0,N1371_0_r_0,N1508_0_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_547_5_r_0,G42_7_r_0,n_572_7_r_0,n_573_7_r_0,n_549_7_r_0,n_569_7_r_0);
input IN_1_0_l_11,IN_2_0_l_11,IN_3_0_l_11,IN_4_0_l_11,IN_1_1_l_11,IN_2_1_l_11,IN_3_1_l_11,IN_1_3_l_11,IN_2_3_l_11,IN_3_3_l_11,IN_1_6_l_11,IN_2_6_l_11,IN_3_6_l_11,IN_4_6_l_11,IN_5_6_l_11,blif_clk_net_5_r_0,blif_reset_net_5_r_0;
output N1371_0_r_0,N1508_0_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_547_5_r_0,G42_7_r_0,n_572_7_r_0,n_573_7_r_0,n_549_7_r_0,n_569_7_r_0;
wire N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_102_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1372_10_r_11,N1508_10_r_11,n_431_5_r_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11,n43_11,n44_11,n45_11,n46_11,n47_11,n48_11,n49_11,n50_11,n51_11,n52_11,n53_11,n54_11,n55_11,n56_11,n57_11,n58_11,n59_11,n60_11,n61_11,n62_11,n63_11,n_102_5_r_0,n_452_7_r_0,n_431_5_r_0,n6_0,n4_7_r_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0,n37_0,n38_0,n39_0,n40_0,n41_0,n42_0,n43_0,n44_0,n45_0;
not I_0(N1372_1_r_11,n53_11);
nor I_1(N1508_1_r_11,n39_11,n53_11);
nor I_2(N6147_2_r_11,n48_11,n49_11);
nor I_3(N6147_3_r_11,n44_11,n45_11);
nand I_4(n_429_or_0_5_r_11,n42_11,n43_11);
DFFARX1 I_5(n_431_5_r_11,blif_clk_net_5_r_0,n6_0,G78_5_r_11,);
nand I_6(n_576_5_r_11,n_102_5_r_11,N1372_10_r_11);
not I_7(n_102_5_r_11,n39_11);
nand I_8(n_547_5_r_11,n36_11,n37_11);
nor I_9(N1507_6_r_11,n52_11,n57_11);
nor I_10(N1508_6_r_11,n46_11,n51_11);
nor I_11(N1372_10_r_11,n43_11,n47_11);
nor I_12(N1508_10_r_11,n55_11,n56_11);
nand I_13(n_431_5_r_11,n40_11,n41_11);
nor I_14(n36_11,n38_11,n39_11);
not I_15(n37_11,n40_11);
nor I_16(n38_11,IN_2_0_l_11,n60_11);
nor I_17(n39_11,IN_1_3_l_11,n54_11);
nand I_18(n40_11,IN_1_1_l_11,IN_2_1_l_11);
nand I_19(n41_11,n_102_5_r_11,n42_11);
and I_20(n42_11,IN_2_6_l_11,n58_11);
not I_21(n43_11,n44_11);
nor I_22(n44_11,IN_3_1_l_11,n40_11);
nand I_23(n45_11,n46_11,n47_11);
not I_24(n46_11,n38_11);
nand I_25(n47_11,n59_11,n62_11);
and I_26(n48_11,n37_11,n47_11);
or I_27(n49_11,n44_11,n50_11);
nor I_28(n50_11,n60_11,n61_11);
or I_29(n51_11,n_102_5_r_11,n52_11);
nor I_30(n52_11,n42_11,n57_11);
nand I_31(n53_11,n37_11,n50_11);
or I_32(n54_11,IN_2_3_l_11,IN_3_3_l_11);
nor I_33(n55_11,n38_11,n42_11);
not I_34(n56_11,N1372_10_r_11);
and I_35(n57_11,n38_11,n50_11);
and I_36(n58_11,IN_1_6_l_11,n59_11);
or I_37(n59_11,IN_5_6_l_11,n63_11);
not I_38(n60_11,IN_1_0_l_11);
nor I_39(n61_11,IN_3_0_l_11,IN_4_0_l_11);
nand I_40(n62_11,IN_3_6_l_11,IN_4_6_l_11);
and I_41(n63_11,IN_3_6_l_11,IN_4_6_l_11);
nor I_42(N1371_0_r_0,n_102_5_r_0,n29_0);
nor I_43(N1508_0_r_0,n_102_5_r_0,n_452_7_r_0);
or I_44(n_429_or_0_5_r_0,n38_0,n_547_5_r_11);
DFFARX1 I_45(n_431_5_r_0,blif_clk_net_5_r_0,n6_0,G78_5_r_0,);
nand I_46(n_576_5_r_0,n26_0,n_547_5_r_11);
not I_47(n_102_5_r_0,n27_0);
nand I_48(n_547_5_r_0,n30_0,n34_0);
DFFARX1 I_49(n4_7_r_0,blif_clk_net_5_r_0,n6_0,G42_7_r_0,);
nor I_50(n_572_7_r_0,n31_0,n_547_5_r_11);
or I_51(n_573_7_r_0,n29_0,n30_0);
nor I_52(n_549_7_r_0,n29_0,n33_0);
nand I_53(n_569_7_r_0,n28_0,n32_0);
nor I_54(n_452_7_r_0,n30_0,n31_0);
nand I_55(n_431_5_r_0,n_102_5_r_0,n35_0);
not I_56(n6_0,blif_reset_net_5_r_0);
nor I_57(n4_7_r_0,n31_0,n37_0);
nor I_58(n26_0,n27_0,n28_0);
nor I_59(n27_0,n28_0,n44_0);
nand I_60(n28_0,N1508_1_r_11,n_576_5_r_11);
not I_61(n29_0,n32_0);
nor I_62(n30_0,n39_0,G78_5_r_11);
not I_63(n31_0,n38_0);
nand I_64(n32_0,n41_0,n42_0);
nor I_65(n33_0,n_102_5_r_0,n_547_5_r_11);
nor I_66(n34_0,n27_0,n_547_5_r_11);
nand I_67(n35_0,n29_0,n36_0);
nor I_68(n36_0,n37_0,n38_0);
not I_69(n37_0,n28_0);
nand I_70(n38_0,n40_0,n_429_or_0_5_r_11);
nor I_71(n39_0,N1372_1_r_11,N6147_2_r_11);
or I_72(n40_0,N1372_1_r_11,N6147_2_r_11);
nor I_73(n41_0,N6147_3_r_11,N1508_1_r_11);
or I_74(n42_0,n43_0,N1372_1_r_11);
nor I_75(n43_0,N1508_6_r_11,N1508_10_r_11);
nor I_76(n44_0,n45_0,N6147_3_r_11);
and I_77(n45_0,N6147_2_r_11,N1507_6_r_11);
endmodule


