module test_final(IN_1_1_l_12,IN_2_1_l_12,IN_3_1_l_12,IN_1_2_l_12,IN_2_2_l_12,IN_3_2_l_12,IN_4_2_l_12,IN_5_2_l_12,IN_1_3_l_12,IN_2_3_l_12,IN_3_3_l_12,IN_1_10_l_12,IN_2_10_l_12,IN_3_10_l_12,IN_4_10_l_12,blif_clk_net_7_r_3,blif_reset_net_7_r_3,N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6134_9_r_3);
input IN_1_1_l_12,IN_2_1_l_12,IN_3_1_l_12,IN_1_2_l_12,IN_2_2_l_12,IN_3_2_l_12,IN_4_2_l_12,IN_5_2_l_12,IN_1_3_l_12,IN_2_3_l_12,IN_3_3_l_12,IN_1_10_l_12,IN_2_10_l_12,IN_3_10_l_12,IN_4_10_l_12,blif_clk_net_7_r_3,blif_reset_net_7_r_3;
output N1372_1_r_3,N1508_1_r_3,N1507_6_r_3,N1508_6_r_3,G42_7_r_3,n_573_7_r_3,n_549_7_r_3,n_569_7_r_3,n_452_7_r_3,N6134_9_r_3;
wire N1371_0_r_12,N1508_0_r_12,N1507_6_r_12,N1508_6_r_12,G42_7_r_12,n_572_7_r_12,n_573_7_r_12,n_549_7_r_12,n_569_7_r_12,n_452_7_r_12,N6147_9_r_12,N6134_9_r_12,I_BUFF_1_9_r_12,n1_12,n23_12,n24_12,n25_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12,n41_12,n42_12,n_572_7_r_3,N6147_9_r_3,I_BUFF_1_9_r_3,n4_7_r_3,n10_3,n30_3,n31_3,n32_3,n33_3,n34_3,n35_3,n36_3,n37_3,n38_3,n39_3,n40_3,n41_3,n42_3,n43_3,n44_3,n45_3,n46_3,n47_3,n48_3,n49_3,n50_3,n51_3;
nor I_0(N1371_0_r_12,I_BUFF_1_9_r_12,n36_12);
nand I_1(N1508_0_r_12,n30_12,n37_12);
nor I_2(N1507_6_r_12,n25_12,n39_12);
nor I_3(N1508_6_r_12,n25_12,n29_12);
DFFARX1 I_4(n1_12,blif_clk_net_7_r_3,n10_3,G42_7_r_12,);
nor I_5(n_572_7_r_12,n23_12,n24_12);
nand I_6(n_573_7_r_12,n_452_7_r_12,n25_12);
nand I_7(n_549_7_r_12,n27_12,n28_12);
nand I_8(n_569_7_r_12,n25_12,n26_12);
nand I_9(n_452_7_r_12,IN_1_1_l_12,IN_2_1_l_12);
nand I_10(N6147_9_r_12,n30_12,n31_12);
nor I_11(N6134_9_r_12,n35_12,n36_12);
not I_12(I_BUFF_1_9_r_12,n_452_7_r_12);
not I_13(n1_12,n_573_7_r_12);
not I_14(n23_12,n36_12);
nor I_15(n24_12,IN_3_1_l_12,n_452_7_r_12);
nand I_16(n25_12,n23_12,n40_12);
not I_17(n26_12,n35_12);
not I_18(n27_12,N6134_9_r_12);
nand I_19(n28_12,n26_12,n29_12);
not I_20(n29_12,n24_12);
nand I_21(n30_12,n33_12,n41_12);
nand I_22(n31_12,n32_12,n33_12);
nor I_23(n32_12,n26_12,n34_12);
nor I_24(n33_12,IN_1_2_l_12,IN_2_2_l_12);
nor I_25(n34_12,IN_5_2_l_12,n42_12);
nor I_26(n35_12,IN_1_3_l_12,n38_12);
nand I_27(n36_12,IN_1_10_l_12,IN_2_10_l_12);
nand I_28(n37_12,n23_12,n35_12);
or I_29(n38_12,IN_2_3_l_12,IN_3_3_l_12);
not I_30(n39_12,n30_12);
or I_31(n40_12,IN_3_10_l_12,IN_4_10_l_12);
nor I_32(n41_12,n34_12,n36_12);
nor I_33(n42_12,IN_3_2_l_12,IN_4_2_l_12);
not I_34(N1372_1_r_3,n40_3);
nor I_35(N1508_1_r_3,N6147_9_r_3,n40_3);
nor I_36(N1507_6_r_3,n31_3,n42_3);
nor I_37(N1508_6_r_3,n30_3,n38_3);
DFFARX1 I_38(n4_7_r_3,blif_clk_net_7_r_3,n10_3,G42_7_r_3,);
nor I_39(n_572_7_r_3,I_BUFF_1_9_r_3,n35_3);
nand I_40(n_573_7_r_3,n30_3,n31_3);
nor I_41(n_549_7_r_3,N6147_9_r_3,n33_3);
nand I_42(n_569_7_r_3,n30_3,n32_3);
nor I_43(n_452_7_r_3,n35_3,N6147_9_r_12);
not I_44(N6147_9_r_3,n32_3);
nor I_45(N6134_9_r_3,n36_3,n37_3);
not I_46(I_BUFF_1_9_r_3,n45_3);
nor I_47(n4_7_r_3,I_BUFF_1_9_r_3,N6147_9_r_12);
not I_48(n10_3,blif_reset_net_7_r_3);
not I_49(n30_3,n39_3);
not I_50(n31_3,n35_3);
nand I_51(n32_3,n41_3,G42_7_r_12);
nor I_52(n33_3,I_BUFF_1_9_r_3,n34_3);
nand I_53(n34_3,n46_3,n_569_7_r_12);
nor I_54(n35_3,n43_3,n44_3);
not I_55(n36_3,n34_3);
nor I_56(n37_3,N6147_9_r_3,N6147_9_r_12);
or I_57(n38_3,n_572_7_r_3,n34_3);
nor I_58(n39_3,n44_3,N1508_0_r_12);
nand I_59(n40_3,n39_3,N6147_9_r_12);
nand I_60(n41_3,N1507_6_r_12,N1508_6_r_12);
nor I_61(n42_3,n34_3,n45_3);
not I_62(n43_3,n_572_7_r_12);
nor I_63(n44_3,N1371_0_r_12,n_572_7_r_12);
nand I_64(n45_3,n49_3,n50_3);
and I_65(n46_3,n47_3,N1508_0_r_12);
nand I_66(n47_3,n41_3,n48_3);
not I_67(n48_3,G42_7_r_12);
nor I_68(n49_3,N1508_6_r_12,n_549_7_r_12);
or I_69(n50_3,n51_3,G42_7_r_12);
nor I_70(n51_3,N1371_0_r_12,n_549_7_r_12);
endmodule


