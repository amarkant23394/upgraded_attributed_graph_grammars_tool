module test_I14999(I1477,I10627,I1470,I10630,I12636,I14999);
input I1477,I10627,I1470,I10630,I12636;
output I14999;
wire I12619,I12670,I12783,I12590,I12584,I12752,I12735,I12653;
not I_0(I12619,I1477);
DFFARX1 I_1(I12653,I1470,I12619,,,I12670,);
DFFARX1 I_2(I12735,I1470,I12619,,,I12783,);
not I_3(I12590,I12752);
and I_4(I12584,I12670,I12783);
nor I_5(I14999,I12584,I12590);
DFFARX1 I_6(I12735,I1470,I12619,,,I12752,);
DFFARX1 I_7(I10630,I1470,I12619,,,I12735,);
and I_8(I12653,I12636,I10627);
endmodule


