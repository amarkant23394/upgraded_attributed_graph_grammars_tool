module test_final(IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_4_2_l_6,IN_5_2_l_6,IN_1_6_l_6,IN_2_6_l_6,IN_3_6_l_6,IN_4_6_l_6,IN_5_6_l_6,IN_1_9_l_6,IN_2_9_l_6,IN_3_9_l_6,IN_4_9_l_6,IN_5_9_l_6,blif_clk_net_7_r_4,blif_reset_net_7_r_4,N1371_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6134_9_r_4);
input IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_4_2_l_6,IN_5_2_l_6,IN_1_6_l_6,IN_2_6_l_6,IN_3_6_l_6,IN_4_6_l_6,IN_5_6_l_6,IN_1_9_l_6,IN_2_9_l_6,IN_3_9_l_6,IN_4_9_l_6,IN_5_9_l_6,blif_clk_net_7_r_4,blif_reset_net_7_r_4;
output N1371_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6134_9_r_4;
wire N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,I_BUFF_1_9_r_6,N1372_10_r_6,N1508_10_r_6,N3_8_r_6,n30_6,n31_6,n32_6,n33_6,n34_6,n35_6,n36_6,n37_6,n38_6,n39_6,n40_6,n41_6,n42_6,n43_6,n44_6,n45_6,n46_6,n47_6,n48_6,n49_6,n50_6,n51_6,n52_6,n53_6,n54_6,N1508_0_r_4,n_573_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4,n4_7_r_4,n6_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4,n38_4,n39_4,n40_4,n41_4;
nor I_0(N1371_0_r_6,n30_6,n33_6);
nor I_1(N1508_0_r_6,n33_6,n44_6);
not I_2(N1372_1_r_6,n41_6);
nor I_3(N1508_1_r_6,n40_6,n41_6);
nor I_4(N1507_6_r_6,n39_6,n45_6);
nor I_5(N1508_6_r_6,n37_6,n38_6);
nor I_6(n_42_8_r_6,n30_6,n31_6);
DFFARX1 I_7(N3_8_r_6,blif_clk_net_7_r_4,n6_4,G199_8_r_6,);
nor I_8(N6147_9_r_6,n32_6,n33_6);
nor I_9(N6134_9_r_6,I_BUFF_1_9_r_6,n35_6);
not I_10(I_BUFF_1_9_r_6,n37_6);
not I_11(N1372_10_r_6,n43_6);
nor I_12(N1508_10_r_6,n42_6,n43_6);
nor I_13(N3_8_r_6,IN_1_9_l_6,n36_6);
nor I_14(n30_6,IN_5_9_l_6,n53_6);
not I_15(n31_6,n36_6);
nor I_16(n32_6,I_BUFF_1_9_r_6,n34_6);
not I_17(n33_6,IN_1_9_l_6);
not I_18(n34_6,n35_6);
nand I_19(n35_6,IN_2_6_l_6,n49_6);
nand I_20(n36_6,IN_5_6_l_6,n51_6);
nand I_21(n37_6,IN_2_9_l_6,n54_6);
or I_22(n38_6,n35_6,n39_6);
nor I_23(n39_6,n40_6,n45_6);
and I_24(n40_6,n46_6,n47_6);
nand I_25(n41_6,n30_6,n31_6);
nor I_26(n42_6,n34_6,n40_6);
nand I_27(n43_6,IN_1_9_l_6,n30_6);
nor I_28(n44_6,n31_6,n40_6);
nor I_29(n45_6,n35_6,n36_6);
nor I_30(n46_6,IN_1_2_l_6,IN_2_2_l_6);
or I_31(n47_6,IN_5_2_l_6,n48_6);
nor I_32(n48_6,IN_3_2_l_6,IN_4_2_l_6);
and I_33(n49_6,IN_1_6_l_6,n50_6);
nand I_34(n50_6,n51_6,n52_6);
nand I_35(n51_6,IN_3_6_l_6,IN_4_6_l_6);
not I_36(n52_6,IN_5_6_l_6);
nor I_37(n53_6,IN_3_9_l_6,IN_4_9_l_6);
or I_38(n54_6,IN_3_9_l_6,IN_4_9_l_6);
nor I_39(N1371_0_r_4,n25_4,N1371_0_r_6);
not I_40(N1508_0_r_4,n25_4);
nor I_41(N1507_6_r_4,n32_4,n33_4);
nor I_42(N1508_6_r_4,n22_4,n29_4);
DFFARX1 I_43(n4_7_r_4,blif_clk_net_7_r_4,n6_4,G42_7_r_4,);
not I_44(n_572_7_r_4,n_573_7_r_4);
nand I_45(n_573_7_r_4,n21_4,n22_4);
nor I_46(n_549_7_r_4,n24_4,N1371_0_r_6);
nand I_47(n_569_7_r_4,n22_4,n23_4);
nor I_48(n_452_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4);
not I_49(N6147_9_r_4,n28_4);
nor I_50(N6134_9_r_4,N1508_0_r_4,n28_4);
not I_51(I_BUFF_1_9_r_4,n21_4);
nor I_52(n4_7_r_4,N6147_9_r_4,N1371_0_r_6);
not I_53(n6_4,blif_reset_net_7_r_4);
nand I_54(n21_4,n39_4,n40_4);
or I_55(n22_4,n31_4,N6134_9_r_6);
not I_56(n23_4,N1371_0_r_6);
nor I_57(n24_4,n25_4,n26_4);
nand I_58(n25_4,N1371_0_r_6,N1508_0_r_6);
nand I_59(n26_4,n21_4,n27_4);
nand I_60(n27_4,n36_4,n37_4);
nand I_61(n28_4,n38_4,N1507_6_r_6);
nand I_62(n29_4,N1508_0_r_4,n30_4);
nand I_63(n30_4,n34_4,n35_4);
nor I_64(n31_4,N1508_6_r_6,n_42_8_r_6);
not I_65(n32_4,n30_4);
nor I_66(n33_4,n21_4,n28_4);
nand I_67(n34_4,N6147_9_r_4,I_BUFF_1_9_r_4);
nand I_68(n35_4,N1508_0_r_4,n27_4);
not I_69(n36_4,N1372_1_r_6);
nand I_70(n37_4,N1372_10_r_6,N1508_10_r_6);
or I_71(n38_4,N1508_6_r_6,n_42_8_r_6);
nor I_72(n39_4,N1508_0_r_6,N1508_1_r_6);
or I_73(n40_4,n41_4,N1372_1_r_6);
nor I_74(n41_4,G199_8_r_6,N6147_9_r_6);
endmodule


