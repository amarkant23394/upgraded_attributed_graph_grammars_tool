module test_I5864(I1477,I2328,I2695,I2161,I2509,I2557,I1470,I5864);
input I1477,I2328,I2695,I2161,I2509,I2557,I1470;
output I5864;
wire I2167,I4629,I4595,I4544,I4869,I2149,I2633,I4536,I4561,I4578,I2173,I2181,I4515;
nand I_0(I2167,I2633,I2328);
nor I_1(I4629,I2167,I2173);
DFFARX1 I_2(I4578,I1470,I4544,,,I4595,);
not I_3(I4544,I1477);
DFFARX1 I_4(I2149,I1470,I4544,,,I4869,);
DFFARX1 I_5(I2695,I1470,I2181,,,I2149,);
DFFARX1 I_6(I1470,I2181,,,I2633,);
nor I_7(I4536,I4869,I4595);
nand I_8(I4561,I2173);
and I_9(I4578,I4561,I2161);
nor I_10(I5864,I4536,I4515);
nand I_11(I2173,I2557,I2509);
not I_12(I2181,I1477);
not I_13(I4515,I4629);
endmodule


