module test_I4401(I2878,I1477,I1470,I2793,I1335,I4401);
input I2878,I1477,I1470,I2793,I1335;
output I4401;
wire I2810,I3124,I2727,I3076,I4308,I3983;
nand I_0(I2810,I2793,I1335);
nor I_1(I3124,I3076,I2878);
nand I_2(I2727,I2810,I3124);
DFFARX1 I_3(I1470,,,I3076,);
not I_4(I4401,I4308);
DFFARX1 I_5(I2727,I1470,I3983,,,I4308,);
not I_6(I3983,I1477);
endmodule


