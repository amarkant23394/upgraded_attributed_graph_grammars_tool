module test_I14715(I1477,I1470,I13296,I13618,I14715);
input I1477,I1470,I13296,I13618;
output I14715;
wire I14667,I13189,I13197,I14650,I13165,I14370,I13635,I13248;
and I_0(I14667,I14650,I13189);
DFFARX1 I_1(I13635,I1470,I13197,,,I13189,);
not I_2(I13197,I1477);
DFFARX1 I_3(I13165,I1470,I14370,,,I14650,);
DFFARX1 I_4(I13248,I1470,I13197,,,I13165,);
not I_5(I14370,I1477);
and I_6(I13635,I13296,I13618);
DFFARX1 I_7(I1470,I13197,,,I13248,);
not I_8(I14715,I14667);
endmodule


