module test_final(IN_1_2_l_9,IN_2_2_l_9,IN_3_2_l_9,IN_6_2_l_9,IN_1_3_l_9,IN_2_3_l_9,IN_4_3_l_9,IN_1_4_l_9,IN_2_4_l_9,IN_3_4_l_9,IN_6_4_l_9,blif_clk_net_1_r_12,blif_reset_net_1_r_12,G42_1_r_12,n_572_1_r_12,n_573_1_r_12,n_549_1_r_12,n_42_2_r_12,G199_2_r_12,ACVQN1_5_r_12,P6_5_r_12);
input IN_1_2_l_9,IN_2_2_l_9,IN_3_2_l_9,IN_6_2_l_9,IN_1_3_l_9,IN_2_3_l_9,IN_4_3_l_9,IN_1_4_l_9,IN_2_4_l_9,IN_3_4_l_9,IN_6_4_l_9,blif_clk_net_1_r_12,blif_reset_net_1_r_12;
output G42_1_r_12,n_572_1_r_12,n_573_1_r_12,n_549_1_r_12,n_42_2_r_12,G199_2_r_12,ACVQN1_5_r_12,P6_5_r_12;
wire G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_452_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9,N3_2_l_9,n27_9,n16_9,n26_9,n15_9,n29_internal_9,n29_9,N1_4_l_9,n25_9,n28_internal_9,n28_9,n4_1_r_9,N3_2_r_9,N1_4_r_9,n_42_2_l_9,n17_9,n18_9,n19_9,n20_9,n21_9,n22_9,n23_9,n24_9,n_431_0_l_12,n8_12,n41_12,ACVQN1_5_l_12,n22_12,n42_12,n4_1_r_12,N3_2_r_12,n3_12,P6_5_r_internal_12,n26_12,n27_12,n28_12,n29_12,n30_12,n31_12,n32_12,n33_12,n34_12,n35_12,n36_12,n37_12,n38_12,n39_12,n40_12;
DFFARX1 I_0(n4_1_r_9,blif_clk_net_1_r_12,n8_12,G42_1_r_9,);
nor I_1(n_572_1_r_9,n27_9,n_42_2_l_9);
or I_2(n_573_1_r_9,n25_9,n_42_2_l_9);
nand I_3(n_549_1_r_9,n17_9,n18_9);
or I_4(n_569_1_r_9,n26_9,n_42_2_l_9);
nor I_5(n_452_1_r_9,n26_9,n25_9);
nor I_6(n_42_2_r_9,n25_9,n19_9);
DFFARX1 I_7(N3_2_r_9,blif_clk_net_1_r_12,n8_12,G199_2_r_9,);
DFFARX1 I_8(N1_4_r_9,blif_clk_net_1_r_12,n8_12,G199_4_r_9,);
DFFARX1 I_9(n_42_2_l_9,blif_clk_net_1_r_12,n8_12,G214_4_r_9,);
and I_10(N3_2_l_9,IN_6_2_l_9,n22_9);
DFFARX1 I_11(N3_2_l_9,blif_clk_net_1_r_12,n8_12,n27_9,);
not I_12(n16_9,n27_9);
DFFARX1 I_13(IN_1_3_l_9,blif_clk_net_1_r_12,n8_12,n26_9,);
not I_14(n15_9,n26_9);
DFFARX1 I_15(IN_2_3_l_9,blif_clk_net_1_r_12,n8_12,n29_internal_9,);
not I_16(n29_9,n29_internal_9);
and I_17(N1_4_l_9,IN_6_4_l_9,n24_9);
DFFARX1 I_18(N1_4_l_9,blif_clk_net_1_r_12,n8_12,n25_9,);
DFFARX1 I_19(IN_3_4_l_9,blif_clk_net_1_r_12,n8_12,n28_internal_9,);
not I_20(n28_9,n28_internal_9);
nor I_21(n4_1_r_9,n27_9,n26_9);
nor I_22(N3_2_r_9,n15_9,n21_9);
nor I_23(N1_4_r_9,n16_9,n21_9);
nor I_24(n_42_2_l_9,IN_1_2_l_9,IN_3_2_l_9);
not I_25(n17_9,n_452_1_r_9);
nand I_26(n18_9,n27_9,n15_9);
nor I_27(n19_9,n29_9,n20_9);
not I_28(n20_9,IN_4_3_l_9);
and I_29(n21_9,IN_4_3_l_9,n23_9);
nand I_30(n22_9,IN_2_2_l_9,IN_3_2_l_9);
nor I_31(n23_9,n29_9,n28_9);
nand I_32(n24_9,IN_1_4_l_9,IN_2_4_l_9);
DFFARX1 I_33(n4_1_r_12,blif_clk_net_1_r_12,n8_12,G42_1_r_12,);
nor I_34(n_572_1_r_12,n29_12,n30_12);
nand I_35(n_573_1_r_12,n26_12,n27_12);
nor I_36(n_549_1_r_12,n33_12,n34_12);
and I_37(n_42_2_r_12,n42_12,n39_12);
DFFARX1 I_38(N3_2_r_12,blif_clk_net_1_r_12,n8_12,G199_2_r_12,);
DFFARX1 I_39(n3_12,blif_clk_net_1_r_12,n8_12,ACVQN1_5_r_12,);
not I_40(P6_5_r_12,P6_5_r_internal_12);
or I_41(n_431_0_l_12,n36_12,n_573_1_r_9);
not I_42(n8_12,blif_reset_net_1_r_12);
DFFARX1 I_43(n_431_0_l_12,blif_clk_net_1_r_12,n8_12,n41_12,);
DFFARX1 I_44(G214_4_r_9,blif_clk_net_1_r_12,n8_12,ACVQN1_5_l_12,);
not I_45(n22_12,ACVQN1_5_l_12);
DFFARX1 I_46(G199_2_r_9,blif_clk_net_1_r_12,n8_12,n42_12,);
nor I_47(n4_1_r_12,n41_12,n31_12);
nor I_48(N3_2_r_12,n22_12,n40_12);
not I_49(n3_12,n39_12);
DFFARX1 I_50(ACVQN1_5_l_12,blif_clk_net_1_r_12,n8_12,P6_5_r_internal_12,);
and I_51(n26_12,n_569_1_r_9,G42_1_r_9);
nor I_52(n27_12,n28_12,n29_12);
not I_53(n28_12,n_572_1_r_9);
nand I_54(n29_12,n31_12,n32_12);
nand I_55(n30_12,n42_12,n_572_1_r_9);
not I_56(n31_12,n_572_1_r_9);
not I_57(n32_12,n_549_1_r_9);
nand I_58(n33_12,n31_12,n35_12);
nand I_59(n34_12,n_569_1_r_9,G42_1_r_9);
nand I_60(n35_12,n41_12,n42_12);
and I_61(n36_12,n37_12,G199_4_r_9);
nor I_62(n37_12,n38_12,n_42_2_r_9);
not I_63(n38_12,G42_1_r_9);
nor I_64(n39_12,n38_12,G42_1_r_9);
nor I_65(n40_12,n39_12,n_572_1_r_9);
endmodule


