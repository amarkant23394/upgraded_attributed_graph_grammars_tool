module test_I2022(I1475,I1207,I1294,I1279,I1301,I2022);
input I1475,I1207,I1294,I1279,I1301;
output I2022;
wire I2005,I1444,I1316,I1322,I1492,I1310,I1639,I1577,I1427,I1954,I1687,I1704,I1622,I1342,I1509;
nor I_0(I2005,I1954,I1310);
nand I_1(I2022,I2005,I1316);
nand I_2(I1444,I1427);
nand I_3(I1316,I1509,I1687);
nand I_4(I1322,I1427,I1704);
and I_5(I1492,I1475,I1279);
DFFARX1 I_6(I1577,I1294,I1342,,,I1310,);
and I_7(I1639,I1622,I1207);
and I_8(I1577,I1509,I1444);
DFFARX1 I_9(I1294,I1342,,,I1427,);
not I_10(I1954,I1322);
not I_11(I1687,I1639);
nor I_12(I1704,I1687);
DFFARX1 I_13(I1294,I1342,,,I1622,);
not I_14(I1342,I1301);
DFFARX1 I_15(I1492,I1294,I1342,,,I1509,);
endmodule


