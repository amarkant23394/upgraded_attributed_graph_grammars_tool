module test_I4742(I1477,I2574,I1470,I4742);
input I1477,I2574,I1470;
output I4742;
wire I2181,I4544,I2232,I4708,I4725,I2164,I2393,I2263,I2158,I2146;
not I_0(I2181,I1477);
not I_1(I4544,I1477);
DFFARX1 I_2(I1470,I2181,,,I2232,);
nand I_3(I4708,I2146,I2164);
and I_4(I4725,I4708,I2158);
DFFARX1 I_5(I4725,I1470,I4544,,,I4742,);
DFFARX1 I_6(I2574,I1470,I2181,,,I2164,);
DFFARX1 I_7(I1470,I2181,,,I2393,);
DFFARX1 I_8(I2232,I1470,I2181,,,I2263,);
not I_9(I2158,I2263);
and I_10(I2146,I2232,I2393);
endmodule


