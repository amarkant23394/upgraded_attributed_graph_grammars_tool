module test_I7833(I1477,I7765,I6363,I6843,I1470,I7833);
input I1477,I7765,I6363,I6843,I1470;
output I7833;
wire I7816,I6380,I6312,I6297,I7652,I6329,I6318,I7782,I7669,I6306,I7799,I7570,I7587,I6411,I6300;
DFFARX1 I_0(I7799,I1470,I7570,,,I7816,);
DFFARX1 I_1(I6363,I1470,I6329,,,I6380,);
DFFARX1 I_2(I1470,I6329,,,I6312,);
DFFARX1 I_3(I6843,I1470,I6329,,,I6297,);
nor I_4(I7652,I7587,I6297);
not I_5(I6329,I1477);
not I_6(I6318,I6380);
and I_7(I7782,I7765,I6312);
nor I_8(I7833,I7816,I7669);
nand I_9(I7669,I7652,I6318);
not I_10(I6306,I6411);
or I_11(I7799,I7782,I6306);
not I_12(I7570,I1477);
not I_13(I7587,I6300);
DFFARX1 I_14(I6380,I1470,I6329,,,I6411,);
DFFARX1 I_15(I1470,I6329,,,I6300,);
endmodule


