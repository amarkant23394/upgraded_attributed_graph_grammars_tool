module test_final(IN_1_2_l,IN_2_2_l,IN_3_2_l,IN_4_2_l,IN_5_2_l,IN_1_4_l,IN_2_4_l,IN_3_4_l,IN_4_4_l,IN_5_4_l,IN_1_9_l,IN_2_9_l,IN_3_9_l,IN_4_9_l,IN_5_9_l,blif_clk_net_7_r,blif_reset_net_7_r,N6147_2_r,N6147_3_r,N1507_6_r,N1508_6_r,G42_7_r,n_572_7_r,n_573_7_r,n_549_7_r,n_569_7_r,n_452_7_r,N6147_9_r,N6134_9_r,I_BUFF_1_9_r);
input IN_1_2_l,IN_2_2_l,IN_3_2_l,IN_4_2_l,IN_5_2_l,IN_1_4_l,IN_2_4_l,IN_3_4_l,IN_4_4_l,IN_5_4_l,IN_1_9_l,IN_2_9_l,IN_3_9_l,IN_4_9_l,IN_5_9_l,blif_clk_net_7_r,blif_reset_net_7_r;
output N6147_2_r,N6147_3_r,N1507_6_r,N1508_6_r,G42_7_r,n_572_7_r,n_573_7_r,n_549_7_r,n_569_7_r,n_452_7_r,N6147_9_r,N6134_9_r,I_BUFF_1_9_r;
wire N6147_2_l,n5_2_l,n6_2_l,N6138_2_l,n7_2_l,N1372_4_l,N1508_4_l,n6_4_l,n7_4_l,n8_4_l,N6150_9_l,N6147_9_l,N6134_9_l,n3_9_l,I_BUFF_1_9_l,n5_2_r,n6_2_r,N6138_2_r,n7_2_r,n3_3_r,N6138_3_r,n6_6_r,n7_6_r,n8_6_r,n9_6_r,n_87_7_r,n4_7_r,n2_7_r,n7_7_r,N6150_9_r,n3_9_r;
nor I_0(N6147_2_l,n5_2_l,n6_2_l);
nor I_1(n5_2_l,IN_5_2_l,n7_2_l);
not I_2(n6_2_l,N6138_2_l);
nor I_3(N6138_2_l,IN_1_2_l,IN_2_2_l);
nor I_4(n7_2_l,IN_3_2_l,IN_4_2_l);
not I_5(N1372_4_l,n7_4_l);
nor I_6(N1508_4_l,n6_4_l,n7_4_l);
nor I_7(n6_4_l,IN_5_4_l,n8_4_l);
nand I_8(n7_4_l,IN_1_4_l,IN_2_4_l);
and I_9(n8_4_l,IN_3_4_l,IN_4_4_l);
not I_10(N6150_9_l,IN_2_9_l);
nor I_11(N6147_9_l,N6150_9_l,n3_9_l);
nor I_12(N6134_9_l,IN_5_9_l,n3_9_l);
nor I_13(n3_9_l,IN_3_9_l,IN_4_9_l);
buf I_14(I_BUFF_1_9_l,IN_1_9_l);
nor I_15(N6147_2_r,n5_2_r,n6_2_r);
nor I_16(n5_2_r,n7_2_r,N6147_9_l);
not I_17(n6_2_r,N6138_2_r);
nor I_18(N6138_2_r,N6147_2_l,N6134_9_l);
nor I_19(n7_2_r,N1372_4_l,N1508_4_l);
nor I_20(N6147_3_r,n3_3_r,N6134_9_l);
not I_21(n3_3_r,N6138_3_r);
nor I_22(N6138_3_r,N6147_2_l,I_BUFF_1_9_l);
nor I_23(N1507_6_r,n8_6_r,n9_6_r);
and I_24(N1508_6_r,n6_6_r,N6147_9_l);
nor I_25(n6_6_r,n7_6_r,n8_6_r);
not I_26(n7_6_r,N6147_2_l);
nor I_27(n8_6_r,n9_6_r,N1508_4_l);
and I_28(n9_6_r,N6134_9_l,N1508_4_l);
DFFARX1 I_29(n4_7_r,blif_clk_net_7_r,n2_7_r,G42_7_r,);
not I_30(n_87_7_r,N6147_2_l);
nor I_31(n_572_7_r,I_BUFF_1_9_l,N6147_2_l);
or I_32(n_573_7_r,N1372_4_l,I_BUFF_1_9_l);
nor I_33(n_549_7_r,n7_7_r,N1508_4_l);
or I_34(n_569_7_r,N1508_4_l,N1372_4_l);
nor I_35(n_452_7_r,I_BUFF_1_9_l,N6147_2_l);
nor I_36(n4_7_r,I_BUFF_1_9_l,N1372_4_l);
not I_37(n2_7_r,blif_reset_net_7_r);
and I_38(n7_7_r,n_87_7_r,N1372_4_l);
not I_39(N6150_9_r,N6147_9_l);
nor I_40(N6147_9_r,N6150_9_r,n3_9_r);
nor I_41(N6134_9_r,n3_9_r,N6147_9_l);
nor I_42(n3_9_r,N6147_9_l,N6134_9_l);
buf I_43(I_BUFF_1_9_r,N1508_4_l);
endmodule


