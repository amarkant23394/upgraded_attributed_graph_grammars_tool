module test_final(IN_1_0_l_15,IN_2_0_l_15,IN_3_0_l_15,IN_4_0_l_15,IN_1_1_l_15,IN_2_1_l_15,IN_3_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_3_3_l_15,IN_1_6_l_15,IN_2_6_l_15,IN_3_6_l_15,IN_4_6_l_15,IN_5_6_l_15,blif_clk_net_8_r_8,blif_reset_net_8_r_8,N1371_0_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,N1508_10_r_8);
input IN_1_0_l_15,IN_2_0_l_15,IN_3_0_l_15,IN_4_0_l_15,IN_1_1_l_15,IN_2_1_l_15,IN_3_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_3_3_l_15,IN_1_6_l_15,IN_2_6_l_15,IN_3_6_l_15,IN_4_6_l_15,IN_5_6_l_15,blif_clk_net_8_r_8,blif_reset_net_8_r_8;
output N1371_0_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,N1508_10_r_8;
wire N1371_0_r_15,N1508_0_r_15,N1372_1_r_15,N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_102_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15,n_431_5_r_15,n31_15,n32_15,n33_15,n34_15,n35_15,n36_15,n37_15,n38_15,n39_15,n40_15,n41_15,n42_15,n43_15,n44_15,n45_15,n46_15,n47_15,n48_15,n49_15,n50_15,n51_15,n52_15,n53_15,n54_15,n55_15,N1508_0_r_8,N1372_1_r_8,I_BUFF_1_9_r_8,N1372_10_r_8,N3_8_l_8,n8_8,n53_8,n29_8,N3_8_r_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8,n38_8,n39_8,n40_8,n41_8,n42_8,n43_8,n44_8,n45_8,n46_8,n47_8,n48_8,n49_8,n50_8,n51_8,n52_8;
and I_0(N1371_0_r_15,N1508_0_r_15,n_102_5_r_15);
nor I_1(N1508_0_r_15,IN_2_0_l_15,n55_15);
nor I_2(N1372_1_r_15,n_102_5_r_15,n46_15);
nor I_3(N1508_1_r_15,N1508_0_r_15,n45_15);
not I_4(N1372_4_r_15,n39_15);
nor I_5(N1508_4_r_15,n39_15,n43_15);
nand I_6(n_429_or_0_5_r_15,n36_15,n38_15);
DFFARX1 I_7(n_431_5_r_15,blif_clk_net_8_r_8,n8_8,G78_5_r_15,);
nand I_8(n_576_5_r_15,n31_15,n32_15);
not I_9(n_102_5_r_15,n33_15);
nand I_10(n_547_5_r_15,N1371_0_r_15,n35_15);
nor I_11(N1507_6_r_15,n42_15,n46_15);
nand I_12(N1508_6_r_15,n39_15,n40_15);
nand I_13(n_431_5_r_15,n36_15,n37_15);
nor I_14(n31_15,n33_15,n34_15);
nor I_15(n32_15,IN_1_3_l_15,n44_15);
nor I_16(n33_15,n54_15,n55_15);
nand I_17(n34_15,IN_2_6_l_15,n49_15);
nand I_18(n35_15,IN_1_1_l_15,IN_2_1_l_15);
not I_19(n36_15,n32_15);
nand I_20(n37_15,n34_15,n38_15);
not I_21(n38_15,n46_15);
nand I_22(n39_15,n38_15,n41_15);
nand I_23(n40_15,n41_15,n42_15);
and I_24(n41_15,IN_5_6_l_15,n51_15);
and I_25(n42_15,IN_2_1_l_15,n47_15);
and I_26(n43_15,n34_15,n36_15);
or I_27(n44_15,IN_2_3_l_15,IN_3_3_l_15);
not I_28(n45_15,N1372_1_r_15);
nand I_29(n46_15,IN_2_1_l_15,n53_15);
nor I_30(n47_15,n34_15,n48_15);
not I_31(n48_15,IN_1_1_l_15);
and I_32(n49_15,IN_1_6_l_15,n50_15);
nand I_33(n50_15,n51_15,n52_15);
nand I_34(n51_15,IN_3_6_l_15,IN_4_6_l_15);
not I_35(n52_15,IN_5_6_l_15);
nor I_36(n53_15,IN_3_1_l_15,n48_15);
nor I_37(n54_15,IN_3_0_l_15,IN_4_0_l_15);
not I_38(n55_15,IN_1_0_l_15);
nor I_39(N1371_0_r_8,n46_8,n51_8);
not I_40(N1508_0_r_8,n46_8);
nor I_41(N1372_1_r_8,n37_8,n49_8);
and I_42(N1508_1_r_8,N1372_1_r_8,n29_8);
nor I_43(N1507_6_r_8,n47_8,n48_8);
nor I_44(N1508_6_r_8,n37_8,n38_8);
nor I_45(n_42_8_r_8,I_BUFF_1_9_r_8,n53_8);
DFFARX1 I_46(N3_8_r_8,blif_clk_net_8_r_8,n8_8,G199_8_r_8,);
nor I_47(N6147_9_r_8,n29_8,n30_8);
nor I_48(N6134_9_r_8,n30_8,n31_8);
not I_49(I_BUFF_1_9_r_8,n35_8);
nor I_50(N1372_10_r_8,n46_8,n49_8);
nor I_51(N1508_10_r_8,n40_8,n41_8);
and I_52(N3_8_l_8,n36_8,N1508_1_r_15);
not I_53(n8_8,blif_reset_net_8_r_8);
DFFARX1 I_54(N3_8_l_8,blif_clk_net_8_r_8,n8_8,n53_8,);
not I_55(n29_8,n53_8);
nor I_56(N3_8_r_8,n33_8,n34_8);
and I_57(n30_8,n32_8,n33_8);
nor I_58(n31_8,N1508_4_r_15,n_576_5_r_15);
nand I_59(n32_8,n42_8,n_576_5_r_15);
or I_60(n33_8,n46_8,N1508_1_r_15);
nor I_61(n34_8,n32_8,n35_8);
nand I_62(n35_8,n44_8,G78_5_r_15);
nand I_63(n36_8,N1507_6_r_15,n_576_5_r_15);
not I_64(n37_8,n31_8);
nand I_65(n38_8,N1508_0_r_8,n39_8);
nand I_66(n39_8,n33_8,n50_8);
and I_67(n40_8,n32_8,n35_8);
not I_68(n41_8,N1372_10_r_8);
and I_69(n42_8,n43_8,N1508_4_r_15);
nand I_70(n43_8,n44_8,n45_8);
nand I_71(n44_8,N1372_4_r_15,n_429_or_0_5_r_15);
not I_72(n45_8,G78_5_r_15);
nand I_73(n46_8,n_429_or_0_5_r_15,G78_5_r_15);
not I_74(n47_8,n39_8);
nor I_75(n48_8,n35_8,n49_8);
not I_76(n49_8,n51_8);
nand I_77(n50_8,I_BUFF_1_9_r_8,n51_8);
nor I_78(n51_8,n52_8,N1372_4_r_15);
or I_79(n52_8,n_547_5_r_15,N1508_6_r_15);
endmodule


