module test_I13023(I9638,I1477,I10664,I9771,I1470,I13023);
input I9638,I1477,I10664,I9771,I1470;
output I13023;
wire I12619,I10715,I9477,I9465,I9816,I10766,I10636,I9833,I10732;
not I_0(I12619,I1477);
nor I_1(I10715,I10664,I9477);
nor I_2(I9477,I9771,I9833);
DFFARX1 I_3(I10636,I1470,I12619,,,I13023,);
nand I_4(I9465,I9816,I9638);
DFFARX1 I_5(I1470,,,I9816,);
not I_6(I10766,I9477);
nor I_7(I10636,I10732,I10766);
and I_8(I9833,I9816);
nand I_9(I10732,I10715,I9465);
endmodule


