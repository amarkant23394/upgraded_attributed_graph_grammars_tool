module test_final(G1_0_l_11,G2_0_l_11,IN_2_0_l_11,IN_4_0_l_11,IN_5_0_l_11,IN_7_0_l_11,IN_8_0_l_11,IN_10_0_l_11,IN_11_0_l_11,IN_1_5_l_11,IN_2_5_l_11,blif_clk_net_1_r_8,blif_reset_net_1_r_8,G42_1_r_8,n_572_1_r_8,n_549_1_r_8,n_569_1_r_8,n_452_1_r_8,n_42_2_r_8,G199_2_r_8,G199_4_r_8,G214_4_r_8);
input G1_0_l_11,G2_0_l_11,IN_2_0_l_11,IN_4_0_l_11,IN_5_0_l_11,IN_7_0_l_11,IN_8_0_l_11,IN_10_0_l_11,IN_11_0_l_11,IN_1_5_l_11,IN_2_5_l_11,blif_clk_net_1_r_8,blif_reset_net_1_r_8;
output G42_1_r_8,n_572_1_r_8,n_549_1_r_8,n_569_1_r_8,n_452_1_r_8,n_42_2_r_8,G199_2_r_8,G199_4_r_8,G214_4_r_8;
wire G42_1_r_11,n_572_1_r_11,n_573_1_r_11,n_549_1_r_11,n_569_1_r_11,n_452_1_r_11,n_42_2_r_11,G199_2_r_11,ACVQN2_3_r_11,n_266_and_0_3_r_11,n_431_0_l_11,n43_11,n26_11,n44_11,n45_11,n27_11,n4_1_r_11,N3_2_r_11,n24_11,n25_11,n20_internal_11,n20_11,n28_11,n29_11,n30_11,n31_11,n32_11,n33_11,n34_11,n35_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11,n_431_0_l_8,n8_8,G78_0_l_8,n19_8,n39_8,n22_8,n38_8,n4_1_r_8,N3_2_r_8,N1_4_r_8,n23_8,n24_8,n25_8,n26_8,n27_8,n28_8,n29_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8;
DFFARX1 I_0(n4_1_r_11,blif_clk_net_1_r_8,n8_8,G42_1_r_11,);
nor I_1(n_572_1_r_11,n29_11,n30_11);
nand I_2(n_573_1_r_11,n26_11,n28_11);
nor I_3(n_549_1_r_11,n27_11,n32_11);
nand I_4(n_569_1_r_11,n45_11,n28_11);
nor I_5(n_452_1_r_11,n43_11,n44_11);
nor I_6(n_42_2_r_11,n35_11,n36_11);
DFFARX1 I_7(N3_2_r_11,blif_clk_net_1_r_8,n8_8,G199_2_r_11,);
DFFARX1 I_8(n24_11,blif_clk_net_1_r_8,n8_8,ACVQN2_3_r_11,);
nor I_9(n_266_and_0_3_r_11,n20_11,n37_11);
or I_10(n_431_0_l_11,IN_8_0_l_11,n33_11);
DFFARX1 I_11(n_431_0_l_11,blif_clk_net_1_r_8,n8_8,n43_11,);
not I_12(n26_11,n43_11);
DFFARX1 I_13(IN_2_5_l_11,blif_clk_net_1_r_8,n8_8,n44_11,);
DFFARX1 I_14(IN_1_5_l_11,blif_clk_net_1_r_8,n8_8,n45_11,);
not I_15(n27_11,n45_11);
nor I_16(n4_1_r_11,n44_11,n25_11);
nor I_17(N3_2_r_11,n45_11,n40_11);
nand I_18(n24_11,IN_11_0_l_11,n39_11);
nand I_19(n25_11,IN_7_0_l_11,n38_11);
DFFARX1 I_20(n25_11,blif_clk_net_1_r_8,n8_8,n20_internal_11,);
not I_21(n20_11,n20_internal_11);
not I_22(n28_11,n25_11);
not I_23(n29_11,G1_0_l_11);
nand I_24(n30_11,n26_11,n31_11);
not I_25(n31_11,IN_5_0_l_11);
and I_26(n32_11,n26_11,n44_11);
and I_27(n33_11,IN_2_0_l_11,n34_11);
nor I_28(n34_11,IN_4_0_l_11,n29_11);
not I_29(n35_11,G2_0_l_11);
nand I_30(n36_11,G1_0_l_11,n31_11);
nor I_31(n37_11,IN_5_0_l_11,n29_11);
nor I_32(n38_11,G2_0_l_11,n31_11);
nor I_33(n39_11,G2_0_l_11,IN_10_0_l_11);
nor I_34(n40_11,G2_0_l_11,n41_11);
nor I_35(n41_11,IN_10_0_l_11,n42_11);
not I_36(n42_11,IN_11_0_l_11);
DFFARX1 I_37(n4_1_r_8,blif_clk_net_1_r_8,n8_8,G42_1_r_8,);
nor I_38(n_572_1_r_8,n39_8,n23_8);
and I_39(n_549_1_r_8,n38_8,n23_8);
nand I_40(n_569_1_r_8,n38_8,n24_8);
nor I_41(n_452_1_r_8,n25_8,n26_8);
nor I_42(n_42_2_r_8,n23_8,n28_8);
DFFARX1 I_43(N3_2_r_8,blif_clk_net_1_r_8,n8_8,G199_2_r_8,);
DFFARX1 I_44(N1_4_r_8,blif_clk_net_1_r_8,n8_8,G199_4_r_8,);
DFFARX1 I_45(G78_0_l_8,blif_clk_net_1_r_8,n8_8,G214_4_r_8,);
or I_46(n_431_0_l_8,n29_8,G42_1_r_11);
not I_47(n8_8,blif_reset_net_1_r_8);
DFFARX1 I_48(n_431_0_l_8,blif_clk_net_1_r_8,n8_8,G78_0_l_8,);
not I_49(n19_8,G78_0_l_8);
DFFARX1 I_50(n_573_1_r_11,blif_clk_net_1_r_8,n8_8,n39_8,);
not I_51(n22_8,n39_8);
DFFARX1 I_52(n_572_1_r_11,blif_clk_net_1_r_8,n8_8,n38_8,);
nor I_53(n4_1_r_8,G78_0_l_8,n33_8);
nor I_54(N3_2_r_8,n22_8,n35_8);
nor I_55(N1_4_r_8,n27_8,n37_8);
nand I_56(n23_8,n32_8,n_569_1_r_11);
not I_57(n24_8,n23_8);
nand I_58(n25_8,n36_8,n_266_and_0_3_r_11);
nand I_59(n26_8,n27_8,n28_8);
nor I_60(n27_8,n31_8,G199_2_r_11);
not I_61(n28_8,n_452_1_r_11);
and I_62(n29_8,n30_8,n_42_2_r_11);
nor I_63(n30_8,n31_8,ACVQN2_3_r_11);
not I_64(n31_8,n_549_1_r_11);
and I_65(n32_8,n28_8,G199_2_r_11);
nand I_66(n33_8,n28_8,n34_8);
not I_67(n34_8,n25_8);
nor I_68(n35_8,n34_8,n_452_1_r_11);
not I_69(n36_8,G42_1_r_11);
nor I_70(n37_8,n19_8,n38_8);
endmodule


