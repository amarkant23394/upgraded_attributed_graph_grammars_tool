module test_I5716(I4629,I1477,I1470,I4530,I5716);
input I4629,I1477,I1470,I4530;
output I5716;
wire I5963,I5751,I4515,I4524,I4527,I4595,I5785,I5915,I5802,I5768,I4742;
and I_0(I5716,I5802,I5963);
DFFARX1 I_1(I5915,I1470,I5751,,,I5963,);
not I_2(I5751,I1477);
not I_3(I4515,I4629);
nor I_4(I4524,I4742,I4595);
or I_5(I4527,I4629,I4595);
DFFARX1 I_6(I1470,,,I4595,);
and I_7(I5785,I5768,I4524);
DFFARX1 I_8(I4527,I1470,I5751,,,I5915,);
DFFARX1 I_9(I5785,I1470,I5751,,,I5802,);
nand I_10(I5768,I4530,I4515);
DFFARX1 I_11(I1470,,,I4742,);
endmodule


