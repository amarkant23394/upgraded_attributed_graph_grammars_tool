module test_final(IN_1_1_l_7,IN_2_1_l_7,IN_3_1_l_7,G18_7_l_7,G15_7_l_7,IN_1_7_l_7,IN_4_7_l_7,IN_5_7_l_7,IN_7_7_l_7,IN_9_7_l_7,IN_10_7_l_7,IN_1_8_l_7,IN_2_8_l_7,IN_3_8_l_7,IN_6_8_l_7,blif_clk_net_7_r_4,blif_reset_net_7_r_4,N1371_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6134_9_r_4);
input IN_1_1_l_7,IN_2_1_l_7,IN_3_1_l_7,G18_7_l_7,G15_7_l_7,IN_1_7_l_7,IN_4_7_l_7,IN_5_7_l_7,IN_7_7_l_7,IN_9_7_l_7,IN_10_7_l_7,IN_1_8_l_7,IN_2_8_l_7,IN_3_8_l_7,IN_6_8_l_7,blif_clk_net_7_r_4,blif_reset_net_7_r_4;
output N1371_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6134_9_r_4;
wire N1371_0_r_7,N1508_0_r_7,n_429_or_0_5_r_7,G78_5_r_7,n_576_5_r_7,n_102_5_r_7,n_547_5_r_7,G42_7_r_7,n_572_7_r_7,n_573_7_r_7,n_549_7_r_7,n_569_7_r_7,n_452_7_r_7,n4_7_l_7,n53_7,n30_7,N3_8_l_7,n54_7,n_431_5_r_7,n4_7_r_7,n31_7,n32_7,n33_7,n34_7,n35_7,n36_7,n37_7,n38_7,n39_7,n40_7,n41_7,n42_7,n43_7,n44_7,n45_7,n46_7,n47_7,n48_7,n49_7,n50_7,n51_7,n52_7,N1508_0_r_4,n_573_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4,n4_7_r_4,n6_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4,n38_4,n39_4,n40_4,n41_4;
nor I_0(N1371_0_r_7,n53_7,n52_7);
nor I_1(N1508_0_r_7,n51_7,n52_7);
nand I_2(n_429_or_0_5_r_7,n43_7,n48_7);
DFFARX1 I_3(n_431_5_r_7,blif_clk_net_7_r_4,n6_4,G78_5_r_7,);
nand I_4(n_576_5_r_7,n31_7,n32_7);
nor I_5(n_102_5_r_7,IN_5_7_l_7,IN_9_7_l_7);
nand I_6(n_547_5_r_7,n31_7,n38_7);
DFFARX1 I_7(n4_7_r_7,blif_clk_net_7_r_4,n6_4,G42_7_r_7,);
nor I_8(n_572_7_r_7,n54_7,n33_7);
nand I_9(n_573_7_r_7,n_102_5_r_7,n_452_7_r_7);
nor I_10(n_549_7_r_7,n53_7,n36_7);
nand I_11(n_569_7_r_7,n_102_5_r_7,n30_7);
nand I_12(n_452_7_r_7,IN_1_1_l_7,IN_2_1_l_7);
nor I_13(n4_7_l_7,G18_7_l_7,IN_1_7_l_7);
DFFARX1 I_14(n4_7_l_7,blif_clk_net_7_r_4,n6_4,n53_7,);
not I_15(n30_7,n53_7);
and I_16(N3_8_l_7,IN_6_8_l_7,n50_7);
DFFARX1 I_17(N3_8_l_7,blif_clk_net_7_r_4,n6_4,n54_7,);
nand I_18(n_431_5_r_7,n40_7,n41_7);
nor I_19(n4_7_r_7,n54_7,n49_7);
and I_20(n31_7,n_102_5_r_7,n39_7);
not I_21(n32_7,G18_7_l_7);
nor I_22(n33_7,IN_10_7_l_7,n34_7);
and I_23(n34_7,IN_4_7_l_7,n35_7);
not I_24(n35_7,G15_7_l_7);
nor I_25(n36_7,G18_7_l_7,n37_7);
or I_26(n37_7,IN_5_7_l_7,n54_7);
or I_27(n38_7,IN_1_8_l_7,IN_3_8_l_7);
nor I_28(n39_7,IN_3_1_l_7,n_452_7_r_7);
nand I_29(n40_7,n46_7,n47_7);
nand I_30(n41_7,n42_7,n43_7);
nor I_31(n42_7,n44_7,n45_7);
nor I_32(n43_7,IN_1_8_l_7,IN_3_8_l_7);
nor I_33(n44_7,G15_7_l_7,IN_7_7_l_7);
nor I_34(n45_7,IN_9_7_l_7,IN_10_7_l_7);
nand I_35(n46_7,IN_4_7_l_7,n35_7);
not I_36(n47_7,IN_10_7_l_7);
or I_37(n48_7,IN_3_1_l_7,n_452_7_r_7);
not I_38(n49_7,n_452_7_r_7);
nand I_39(n50_7,IN_2_8_l_7,IN_3_8_l_7);
and I_40(n51_7,n_452_7_r_7,n45_7);
not I_41(n52_7,n44_7);
nor I_42(N1371_0_r_4,n25_4,N1371_0_r_7);
not I_43(N1508_0_r_4,n25_4);
nor I_44(N1507_6_r_4,n32_4,n33_4);
nor I_45(N1508_6_r_4,n22_4,n29_4);
DFFARX1 I_46(n4_7_r_4,blif_clk_net_7_r_4,n6_4,G42_7_r_4,);
not I_47(n_572_7_r_4,n_573_7_r_4);
nand I_48(n_573_7_r_4,n21_4,n22_4);
nor I_49(n_549_7_r_4,n24_4,N1371_0_r_7);
nand I_50(n_569_7_r_4,n22_4,n23_4);
nor I_51(n_452_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4);
not I_52(N6147_9_r_4,n28_4);
nor I_53(N6134_9_r_4,N1508_0_r_4,n28_4);
not I_54(I_BUFF_1_9_r_4,n21_4);
nor I_55(n4_7_r_4,N6147_9_r_4,N1371_0_r_7);
not I_56(n6_4,blif_reset_net_7_r_4);
nand I_57(n21_4,n39_4,n40_4);
or I_58(n22_4,n31_4,n_549_7_r_7);
not I_59(n23_4,N1371_0_r_7);
nor I_60(n24_4,n25_4,n26_4);
nand I_61(n25_4,n_547_5_r_7,G42_7_r_7);
nand I_62(n26_4,n21_4,n27_4);
nand I_63(n27_4,n36_4,n37_4);
nand I_64(n28_4,n38_4,n_576_5_r_7);
nand I_65(n29_4,N1508_0_r_4,n30_4);
nand I_66(n30_4,n34_4,n35_4);
nor I_67(n31_4,N1508_0_r_7,G78_5_r_7);
not I_68(n32_4,n30_4);
nor I_69(n33_4,n21_4,n28_4);
nand I_70(n34_4,N6147_9_r_4,I_BUFF_1_9_r_4);
nand I_71(n35_4,N1508_0_r_4,n27_4);
not I_72(n36_4,n_572_7_r_7);
nand I_73(n37_4,n_569_7_r_7,G78_5_r_7);
or I_74(n38_4,N1508_0_r_7,G78_5_r_7);
nor I_75(n39_4,n_573_7_r_7,n_429_or_0_5_r_7);
or I_76(n40_4,n41_4,N1508_0_r_7);
nor I_77(n41_4,N1371_0_r_7,n_429_or_0_5_r_7);
endmodule


