module test_final(G18_1_l_13,G15_1_l_13,IN_1_1_l_13,IN_4_1_l_13,IN_5_1_l_13,IN_7_1_l_13,IN_9_1_l_13,IN_10_1_l_13,IN_1_3_l_13,IN_2_3_l_13,IN_4_3_l_13,blif_clk_net_1_r_0,blif_reset_net_1_r_0,G42_1_r_0,n_572_1_r_0,n_573_1_r_0,n_549_1_r_0,n_42_2_r_0,G199_2_r_0,G199_4_r_0,G214_4_r_0);
input G18_1_l_13,G15_1_l_13,IN_1_1_l_13,IN_4_1_l_13,IN_5_1_l_13,IN_7_1_l_13,IN_9_1_l_13,IN_10_1_l_13,IN_1_3_l_13,IN_2_3_l_13,IN_4_3_l_13,blif_clk_net_1_r_0,blif_reset_net_1_r_0;
output G42_1_r_0,n_572_1_r_0,n_573_1_r_0,n_549_1_r_0,n_42_2_r_0,G199_2_r_0,G199_4_r_0,G214_4_r_0;
wire G42_1_r_13,n_572_1_r_13,n_573_1_r_13,n_549_1_r_13,n_569_1_r_13,n_452_1_r_13,ACVQN2_3_r_13,n_266_and_0_3_r_13,ACVQN1_5_r_13,P6_5_r_13,n4_1_l_13,n17_internal_13,n17_13,n28_13,ACVQN1_3_l_13,n4_1_r_13,n_266_and_0_3_l_13,n_573_1_l_13,n14_internal_13,n14_13,n_549_1_l_13,n_569_1_l_13,P6_5_r_internal_13,n18_13,n19_13,n20_13,n21_13,n22_13,n23_13,n24_13,n25_13,n26_13,n27_13,n_569_1_r_0,n4_1_l_0,n6_0,n37_0,n38_0,n20_0,ACVQN1_3_l_0,n4_1_r_0,N3_2_r_0,N1_4_r_0,n2_0,n21_0,n22_0,n23_0,n24_0,n25_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0;
DFFARX1 I_0(n4_1_r_13,blif_clk_net_1_r_0,n6_0,G42_1_r_13,);
nor I_1(n_572_1_r_13,n28_13,n_569_1_l_13);
nand I_2(n_573_1_r_13,n18_13,n19_13);
nand I_3(n_549_1_r_13,n_569_1_r_13,n22_13);
nand I_4(n_569_1_r_13,n17_13,n18_13);
nor I_5(n_452_1_r_13,n_573_1_l_13,n25_13);
DFFARX1 I_6(n_266_and_0_3_l_13,blif_clk_net_1_r_0,n6_0,ACVQN2_3_r_13,);
nor I_7(n_266_and_0_3_r_13,n17_13,n14_13);
DFFARX1 I_8(n_549_1_l_13,blif_clk_net_1_r_0,n6_0,ACVQN1_5_r_13,);
not I_9(P6_5_r_13,P6_5_r_internal_13);
nor I_10(n4_1_l_13,G18_1_l_13,IN_1_1_l_13);
DFFARX1 I_11(n4_1_l_13,blif_clk_net_1_r_0,n6_0,n17_internal_13,);
not I_12(n17_13,n17_internal_13);
DFFARX1 I_13(IN_1_3_l_13,blif_clk_net_1_r_0,n6_0,n28_13,);
DFFARX1 I_14(IN_2_3_l_13,blif_clk_net_1_r_0,n6_0,ACVQN1_3_l_13,);
nor I_15(n4_1_r_13,n_573_1_l_13,n_549_1_l_13);
and I_16(n_266_and_0_3_l_13,IN_4_3_l_13,ACVQN1_3_l_13);
nand I_17(n_573_1_l_13,n20_13,n24_13);
DFFARX1 I_18(n_573_1_l_13,blif_clk_net_1_r_0,n6_0,n14_internal_13,);
not I_19(n14_13,n14_internal_13);
and I_20(n_549_1_l_13,n21_13,n26_13);
nand I_21(n_569_1_l_13,n20_13,n21_13);
DFFARX1 I_22(n_569_1_l_13,blif_clk_net_1_r_0,n6_0,P6_5_r_internal_13,);
nand I_23(n18_13,n23_13,n24_13);
or I_24(n19_13,G15_1_l_13,IN_7_1_l_13);
not I_25(n20_13,IN_9_1_l_13);
not I_26(n21_13,IN_10_1_l_13);
nand I_27(n22_13,n17_13,n28_13);
not I_28(n23_13,G18_1_l_13);
not I_29(n24_13,IN_5_1_l_13);
nor I_30(n25_13,G15_1_l_13,IN_7_1_l_13);
nand I_31(n26_13,IN_4_1_l_13,n27_13);
not I_32(n27_13,G15_1_l_13);
DFFARX1 I_33(n4_1_r_0,blif_clk_net_1_r_0,n6_0,G42_1_r_0,);
nor I_34(n_572_1_r_0,n23_0,n_549_1_r_13);
nand I_35(n_573_1_r_0,n21_0,n22_0);
nand I_36(n_549_1_r_0,n_569_1_r_0,n24_0);
nand I_37(n_569_1_r_0,n21_0,n26_0);
nor I_38(n_42_2_r_0,n27_0,n28_0);
DFFARX1 I_39(N3_2_r_0,blif_clk_net_1_r_0,n6_0,G199_2_r_0,);
DFFARX1 I_40(N1_4_r_0,blif_clk_net_1_r_0,n6_0,G199_4_r_0,);
DFFARX1 I_41(n2_0,blif_clk_net_1_r_0,n6_0,G214_4_r_0,);
nor I_42(n4_1_l_0,n_452_1_r_13,ACVQN2_3_r_13);
not I_43(n6_0,blif_reset_net_1_r_0);
DFFARX1 I_44(n4_1_l_0,blif_clk_net_1_r_0,n6_0,n37_0,);
DFFARX1 I_45(n_266_and_0_3_r_13,blif_clk_net_1_r_0,n6_0,n38_0,);
not I_46(n20_0,n38_0);
DFFARX1 I_47(n_572_1_r_13,blif_clk_net_1_r_0,n6_0,ACVQN1_3_l_0,);
nor I_48(n4_1_r_0,n23_0,n_572_1_r_13);
nor I_49(N3_2_r_0,n31_0,n32_0);
nor I_50(N1_4_r_0,n29_0,n32_0);
not I_51(n2_0,n31_0);
nor I_52(n21_0,n37_0,n_573_1_r_13);
not I_53(n22_0,n_549_1_r_13);
nand I_54(n23_0,n20_0,n30_0);
nand I_55(n24_0,n38_0,n25_0);
nor I_56(n25_0,n_573_1_r_13,n_572_1_r_13);
not I_57(n26_0,n_572_1_r_13);
not I_58(n27_0,n29_0);
nor I_59(n28_0,G42_1_r_13,P6_5_r_13);
nand I_60(n29_0,n26_0,n33_0);
not I_61(n30_0,n_573_1_r_13);
nand I_62(n31_0,ACVQN1_3_l_0,ACVQN1_5_r_13);
and I_63(n32_0,n35_0,n36_0);
nand I_64(n33_0,n34_0,G42_1_r_13);
not I_65(n34_0,P6_5_r_13);
nor I_66(n35_0,ACVQN2_3_r_13,P6_5_r_13);
nor I_67(n36_0,G42_1_r_13,n_549_1_r_13);
endmodule


