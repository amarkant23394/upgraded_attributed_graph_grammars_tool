module test_final(IN_1_0_l_15,IN_2_0_l_15,IN_3_0_l_15,IN_4_0_l_15,IN_1_1_l_15,IN_2_1_l_15,IN_3_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_3_3_l_15,IN_1_6_l_15,IN_2_6_l_15,IN_3_6_l_15,IN_4_6_l_15,IN_5_6_l_15,blif_clk_net_5_r_13,blif_reset_net_5_r_13,N1371_0_r_13,N1508_0_r_13,n_429_or_0_5_r_13,G78_5_r_13,n_576_5_r_13,n_547_5_r_13,G42_7_r_13,n_572_7_r_13,n_573_7_r_13,n_549_7_r_13,n_569_7_r_13,n_452_7_r_13);
input IN_1_0_l_15,IN_2_0_l_15,IN_3_0_l_15,IN_4_0_l_15,IN_1_1_l_15,IN_2_1_l_15,IN_3_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_3_3_l_15,IN_1_6_l_15,IN_2_6_l_15,IN_3_6_l_15,IN_4_6_l_15,IN_5_6_l_15,blif_clk_net_5_r_13,blif_reset_net_5_r_13;
output N1371_0_r_13,N1508_0_r_13,n_429_or_0_5_r_13,G78_5_r_13,n_576_5_r_13,n_547_5_r_13,G42_7_r_13,n_572_7_r_13,n_573_7_r_13,n_549_7_r_13,n_569_7_r_13,n_452_7_r_13;
wire N1371_0_r_15,N1508_0_r_15,N1372_1_r_15,N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_102_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15,n_431_5_r_15,n31_15,n32_15,n33_15,n34_15,n35_15,n36_15,n37_15,n38_15,n39_15,n40_15,n41_15,n42_15,n43_15,n44_15,n45_15,n46_15,n47_15,n48_15,n49_15,n50_15,n51_15,n52_15,n53_15,n54_15,n55_15,n_102_5_r_13,n4_7_l_13,n9_13,n62_13,n33_13,n_431_5_r_13,n1_13,n34_13,n35_13,n36_13,n37_13,n38_13,n39_13,n40_13,n41_13,n42_13,n43_13,n44_13,n45_13,n46_13,n47_13,n48_13,n49_13,n50_13,n51_13,n52_13,n53_13,n54_13,n55_13,n56_13,n57_13,n58_13,n59_13,n60_13,n61_13;
and I_0(N1371_0_r_15,N1508_0_r_15,n_102_5_r_15);
nor I_1(N1508_0_r_15,IN_2_0_l_15,n55_15);
nor I_2(N1372_1_r_15,n_102_5_r_15,n46_15);
nor I_3(N1508_1_r_15,N1508_0_r_15,n45_15);
not I_4(N1372_4_r_15,n39_15);
nor I_5(N1508_4_r_15,n39_15,n43_15);
nand I_6(n_429_or_0_5_r_15,n36_15,n38_15);
DFFARX1 I_7(n_431_5_r_15,blif_clk_net_5_r_13,n9_13,G78_5_r_15,);
nand I_8(n_576_5_r_15,n31_15,n32_15);
not I_9(n_102_5_r_15,n33_15);
nand I_10(n_547_5_r_15,N1371_0_r_15,n35_15);
nor I_11(N1507_6_r_15,n42_15,n46_15);
nand I_12(N1508_6_r_15,n39_15,n40_15);
nand I_13(n_431_5_r_15,n36_15,n37_15);
nor I_14(n31_15,n33_15,n34_15);
nor I_15(n32_15,IN_1_3_l_15,n44_15);
nor I_16(n33_15,n54_15,n55_15);
nand I_17(n34_15,IN_2_6_l_15,n49_15);
nand I_18(n35_15,IN_1_1_l_15,IN_2_1_l_15);
not I_19(n36_15,n32_15);
nand I_20(n37_15,n34_15,n38_15);
not I_21(n38_15,n46_15);
nand I_22(n39_15,n38_15,n41_15);
nand I_23(n40_15,n41_15,n42_15);
and I_24(n41_15,IN_5_6_l_15,n51_15);
and I_25(n42_15,IN_2_1_l_15,n47_15);
and I_26(n43_15,n34_15,n36_15);
or I_27(n44_15,IN_2_3_l_15,IN_3_3_l_15);
not I_28(n45_15,N1372_1_r_15);
nand I_29(n46_15,IN_2_1_l_15,n53_15);
nor I_30(n47_15,n34_15,n48_15);
not I_31(n48_15,IN_1_1_l_15);
and I_32(n49_15,IN_1_6_l_15,n50_15);
nand I_33(n50_15,n51_15,n52_15);
nand I_34(n51_15,IN_3_6_l_15,IN_4_6_l_15);
not I_35(n52_15,IN_5_6_l_15);
nor I_36(n53_15,IN_3_1_l_15,n48_15);
nor I_37(n54_15,IN_3_0_l_15,IN_4_0_l_15);
not I_38(n55_15,IN_1_0_l_15);
nor I_39(N1371_0_r_13,n59_13,n61_13);
nor I_40(N1508_0_r_13,n59_13,n60_13);
not I_41(n_429_or_0_5_r_13,n46_13);
DFFARX1 I_42(n_431_5_r_13,blif_clk_net_5_r_13,n9_13,G78_5_r_13,);
nand I_43(n_576_5_r_13,n_102_5_r_13,n34_13);
nor I_44(n_102_5_r_13,n_429_or_0_5_r_15,N1507_6_r_15);
nand I_45(n_547_5_r_13,n48_13,n49_13);
DFFARX1 I_46(n1_13,blif_clk_net_5_r_13,n9_13,G42_7_r_13,);
nor I_47(n_572_7_r_13,n40_13,n41_13);
nand I_48(n_573_7_r_13,n37_13,n38_13);
nor I_49(n_549_7_r_13,n46_13,n47_13);
nand I_50(n_569_7_r_13,n37_13,n43_13);
nand I_51(n_452_7_r_13,n52_13,n53_13);
nor I_52(n4_7_l_13,N1372_4_r_15,n_429_or_0_5_r_15);
not I_53(n9_13,blif_reset_net_5_r_13);
DFFARX1 I_54(n4_7_l_13,blif_clk_net_5_r_13,n9_13,n62_13,);
not I_55(n33_13,n62_13);
nand I_56(n_431_5_r_13,n54_13,n55_13);
not I_57(n1_13,n52_13);
nor I_58(n34_13,n35_13,n36_13);
nor I_59(n35_13,n42_13,n_576_5_r_15);
nand I_60(n36_13,n50_13,n58_13);
nand I_61(n37_13,n44_13,n45_13);
or I_62(n38_13,n39_13,N1508_4_r_15);
nand I_63(n39_13,G78_5_r_15,N1372_4_r_15);
not I_64(n40_13,n36_13);
nor I_65(n41_13,n35_13,N1507_6_r_15);
not I_66(n42_13,G78_5_r_15);
or I_67(n43_13,n_429_or_0_5_r_15,n_576_5_r_15);
not I_68(n44_13,n_576_5_r_15);
not I_69(n45_13,N1508_1_r_15);
nor I_70(n46_13,n39_13,n40_13);
nor I_71(n47_13,n_429_or_0_5_r_15,n_576_5_r_15);
nor I_72(n48_13,n50_13,n51_13);
nor I_73(n49_13,N1508_1_r_15,n_576_5_r_15);
not I_74(n50_13,n59_13);
not I_75(n51_13,n_102_5_r_13);
nand I_76(n52_13,n33_13,n39_13);
nand I_77(n53_13,n33_13,N1508_4_r_15);
nor I_78(n54_13,n_429_or_0_5_r_15,n_576_5_r_15);
nand I_79(n55_13,n62_13,n56_13);
nor I_80(n56_13,n39_13,n57_13);
not I_81(n57_13,n_429_or_0_5_r_15);
or I_82(n58_13,N1508_1_r_15,N1508_4_r_15);
nand I_83(n59_13,n_547_5_r_15,N1508_6_r_15);
nor I_84(n60_13,n51_13,n_576_5_r_15);
nor I_85(n61_13,n39_13,N1508_4_r_15);
endmodule


