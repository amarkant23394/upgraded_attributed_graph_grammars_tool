module test_I2170(I1343,I1231,I1477,I1470,I1271,I2170);
input I1343,I1231,I1477,I1470,I1271;
output I2170;
wire I2181,I2232,I2198,I2215;
not I_0(I2181,I1477);
not I_1(I2170,I2232);
DFFARX1 I_2(I2215,I1470,I2181,,,I2232,);
nand I_3(I2198,I1343,I1231);
and I_4(I2215,I2198,I1271);
endmodule


