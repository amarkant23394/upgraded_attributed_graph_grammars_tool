module test_final(IN_1_2_l_0,IN_2_2_l_0,IN_3_2_l_0,IN_4_2_l_0,IN_5_2_l_0,IN_1_4_l_0,IN_2_4_l_0,IN_3_4_l_0,IN_4_4_l_0,IN_5_4_l_0,IN_1_9_l_0,IN_2_9_l_0,IN_3_9_l_0,IN_4_9_l_0,IN_5_9_l_0,blif_clk_net_5_r_9,blif_reset_net_5_r_9,N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,G78_5_r_9,n_576_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9);
input IN_1_2_l_0,IN_2_2_l_0,IN_3_2_l_0,IN_4_2_l_0,IN_5_2_l_0,IN_1_4_l_0,IN_2_4_l_0,IN_3_4_l_0,IN_4_4_l_0,IN_5_4_l_0,IN_1_9_l_0,IN_2_9_l_0,IN_3_9_l_0,IN_4_9_l_0,IN_5_9_l_0,blif_clk_net_5_r_9,blif_reset_net_5_r_9;
output N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,G78_5_r_9,n_576_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9;
wire N1371_0_r_0,N1508_0_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_102_5_r_0,n_547_5_r_0,G42_7_r_0,n_572_7_r_0,n_573_7_r_0,n_549_7_r_0,n_569_7_r_0,n_452_7_r_0,n_431_5_r_0,n4_7_r_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0,n37_0,n38_0,n39_0,n40_0,n41_0,n42_0,n43_0,n44_0,n45_0,n_429_or_0_5_r_9,n_102_5_r_9,I_BUFF_1_9_r_9,n4_7_l_9,n10_9,n62_9,N3_8_l_9,n63_9,n38_9,n_431_5_r_9,N3_8_r_9,n39_9,n40_9,n41_9,n42_9,n43_9,n44_9,n45_9,n46_9,n47_9,n48_9,n49_9,n50_9,n51_9,n52_9,n53_9,n54_9,n55_9,n56_9,n57_9,n58_9,n59_9,n60_9,n61_9;
nor I_0(N1371_0_r_0,n_102_5_r_0,n29_0);
nor I_1(N1508_0_r_0,n_102_5_r_0,n_452_7_r_0);
or I_2(n_429_or_0_5_r_0,IN_1_9_l_0,n38_0);
DFFARX1 I_3(n_431_5_r_0,blif_clk_net_5_r_9,n10_9,G78_5_r_0,);
nand I_4(n_576_5_r_0,IN_1_9_l_0,n26_0);
not I_5(n_102_5_r_0,n27_0);
nand I_6(n_547_5_r_0,n30_0,n34_0);
DFFARX1 I_7(n4_7_r_0,blif_clk_net_5_r_9,n10_9,G42_7_r_0,);
nor I_8(n_572_7_r_0,IN_1_9_l_0,n31_0);
or I_9(n_573_7_r_0,n29_0,n30_0);
nor I_10(n_549_7_r_0,n29_0,n33_0);
nand I_11(n_569_7_r_0,n28_0,n32_0);
nor I_12(n_452_7_r_0,n30_0,n31_0);
nand I_13(n_431_5_r_0,n_102_5_r_0,n35_0);
nor I_14(n4_7_r_0,n31_0,n37_0);
nor I_15(n26_0,n27_0,n28_0);
nor I_16(n27_0,n28_0,n44_0);
nand I_17(n28_0,IN_1_4_l_0,IN_2_4_l_0);
not I_18(n29_0,n32_0);
nor I_19(n30_0,IN_5_9_l_0,n39_0);
not I_20(n31_0,n38_0);
nand I_21(n32_0,n41_0,n42_0);
nor I_22(n33_0,IN_1_9_l_0,n_102_5_r_0);
nor I_23(n34_0,IN_1_9_l_0,n27_0);
nand I_24(n35_0,n29_0,n36_0);
nor I_25(n36_0,n37_0,n38_0);
not I_26(n37_0,n28_0);
nand I_27(n38_0,IN_2_9_l_0,n40_0);
nor I_28(n39_0,IN_3_9_l_0,IN_4_9_l_0);
or I_29(n40_0,IN_3_9_l_0,IN_4_9_l_0);
nor I_30(n41_0,IN_1_2_l_0,IN_2_2_l_0);
or I_31(n42_0,IN_5_2_l_0,n43_0);
nor I_32(n43_0,IN_3_2_l_0,IN_4_2_l_0);
nor I_33(n44_0,IN_5_4_l_0,n45_0);
and I_34(n45_0,IN_3_4_l_0,IN_4_4_l_0);
nor I_35(N6147_2_r_9,n62_9,n46_9);
not I_36(N1372_4_r_9,n59_9);
nor I_37(N1508_4_r_9,n58_9,n59_9);
nand I_38(n_429_or_0_5_r_9,n_431_5_r_9,n42_9);
DFFARX1 I_39(n_431_5_r_9,blif_clk_net_5_r_9,n10_9,G78_5_r_9,);
nand I_40(n_576_5_r_9,n39_9,n40_9);
not I_41(n_102_5_r_9,I_BUFF_1_9_r_9);
nand I_42(n_547_5_r_9,n43_9,n_429_or_0_5_r_0);
and I_43(n_42_8_r_9,n44_9,n_429_or_0_5_r_0);
DFFARX1 I_44(N3_8_r_9,blif_clk_net_5_r_9,n10_9,G199_8_r_9,);
nor I_45(N6147_9_r_9,n41_9,n45_9);
nor I_46(N6134_9_r_9,n45_9,n51_9);
nor I_47(I_BUFF_1_9_r_9,n41_9,n_429_or_0_5_r_0);
nor I_48(n4_7_l_9,G78_5_r_0,n_429_or_0_5_r_0);
not I_49(n10_9,blif_reset_net_5_r_9);
DFFARX1 I_50(n4_7_l_9,blif_clk_net_5_r_9,n10_9,n62_9,);
and I_51(N3_8_l_9,n57_9,n_547_5_r_0);
DFFARX1 I_52(N3_8_l_9,blif_clk_net_5_r_9,n10_9,n63_9,);
not I_53(n38_9,n63_9);
nor I_54(n_431_5_r_9,n_549_7_r_0,G78_5_r_0);
nor I_55(N3_8_r_9,n_102_5_r_9,n53_9);
nor I_56(n39_9,I_BUFF_1_9_r_9,n42_9);
not I_57(n40_9,n41_9);
nand I_58(n41_9,n_576_5_r_0,n_569_7_r_0);
nor I_59(n42_9,G42_7_r_0,n_573_7_r_0);
nor I_60(n43_9,n63_9,n41_9);
nor I_61(n44_9,G42_7_r_0,N1371_0_r_0);
and I_62(n45_9,n52_9,N1508_0_r_0);
nor I_63(n46_9,n47_9,n48_9);
nor I_64(n47_9,n49_9,n50_9);
not I_65(n48_9,n_429_or_0_5_r_9);
not I_66(n49_9,n42_9);
or I_67(n50_9,n63_9,n51_9);
nor I_68(n51_9,N1371_0_r_0,N1508_0_r_0);
nor I_69(n52_9,n49_9,n_549_7_r_0);
nor I_70(n53_9,n54_9,n55_9);
nor I_71(n54_9,n56_9,n_549_7_r_0);
or I_72(n55_9,n44_9,n_573_7_r_0);
not I_73(n56_9,N1508_0_r_0);
nand I_74(n57_9,N1371_0_r_0,n_572_7_r_0);
nor I_75(n58_9,n62_9,n60_9);
nand I_76(n59_9,n51_9,n61_9);
nor I_77(n60_9,n38_9,n44_9);
nor I_78(n61_9,N1371_0_r_0,n_429_or_0_5_r_0);
endmodule


