module test_final(IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_6_2_l_6,IN_1_3_l_6,IN_2_3_l_6,IN_4_3_l_6,IN_1_4_l_6,IN_2_4_l_6,IN_3_4_l_6,IN_6_4_l_6,blif_clk_net_1_r_17,blif_reset_net_1_r_17,G42_1_r_17,n_572_1_r_17,n_573_1_r_17,n_549_1_r_17,n_569_1_r_17,n_452_1_r_17,ACVQN2_3_r_17,n_266_and_0_3_r_17,G199_4_r_17,G214_4_r_17);
input IN_1_2_l_6,IN_2_2_l_6,IN_3_2_l_6,IN_6_2_l_6,IN_1_3_l_6,IN_2_3_l_6,IN_4_3_l_6,IN_1_4_l_6,IN_2_4_l_6,IN_3_4_l_6,IN_6_4_l_6,blif_clk_net_1_r_17,blif_reset_net_1_r_17;
output G42_1_r_17,n_572_1_r_17,n_573_1_r_17,n_549_1_r_17,n_569_1_r_17,n_452_1_r_17,ACVQN2_3_r_17,n_266_and_0_3_r_17,G199_4_r_17,G214_4_r_17;
wire G42_1_r_6,n_572_1_r_6,n_573_1_r_6,n_549_1_r_6,n_569_1_r_6,n_452_1_r_6,G199_4_r_6,G214_4_r_6,ACVQN1_5_r_6,P6_5_r_6,N3_2_l_6,n27_6,n17_6,n28_6,n26_6,N1_4_l_6,n29_6,n18_6,G214_4_l_6,n12_6,n4_1_r_6,N1_4_r_6,n_42_2_l_6,P6_5_r_internal_6,n19_6,n20_6,n21_6,n22_6,n23_6,n24_6,n25_6,n_431_0_l_17,n6_17,n20_internal_17,n20_17,ACVQN1_5_l_17,n19_internal_17,n19_17,n4_1_r_17,n2_17,n17_internal_17,n17_17,N1_4_r_17,n5_17,n21_17,n22_17,n23_17,n24_17,n25_17,n26_17,n27_17,n28_17,n29_17,n30_17,n31_17,n32_17;
DFFARX1 I_0(n4_1_r_6,blif_clk_net_1_r_17,n6_17,G42_1_r_6,);
nor I_1(n_572_1_r_6,n27_6,n28_6);
nand I_2(n_573_1_r_6,n18_6,n19_6);
nor I_3(n_549_1_r_6,n_42_2_l_6,n21_6);
nand I_4(n_569_1_r_6,n19_6,n20_6);
nor I_5(n_452_1_r_6,n28_6,n29_6);
DFFARX1 I_6(N1_4_r_6,blif_clk_net_1_r_17,n6_17,G199_4_r_6,);
DFFARX1 I_7(n_42_2_l_6,blif_clk_net_1_r_17,n6_17,G214_4_r_6,);
DFFARX1 I_8(n_42_2_l_6,blif_clk_net_1_r_17,n6_17,ACVQN1_5_r_6,);
not I_9(P6_5_r_6,P6_5_r_internal_6);
and I_10(N3_2_l_6,IN_6_2_l_6,n23_6);
DFFARX1 I_11(N3_2_l_6,blif_clk_net_1_r_17,n6_17,n27_6,);
not I_12(n17_6,n27_6);
DFFARX1 I_13(IN_1_3_l_6,blif_clk_net_1_r_17,n6_17,n28_6,);
DFFARX1 I_14(IN_2_3_l_6,blif_clk_net_1_r_17,n6_17,n26_6,);
and I_15(N1_4_l_6,IN_6_4_l_6,n25_6);
DFFARX1 I_16(N1_4_l_6,blif_clk_net_1_r_17,n6_17,n29_6,);
not I_17(n18_6,n29_6);
DFFARX1 I_18(IN_3_4_l_6,blif_clk_net_1_r_17,n6_17,G214_4_l_6,);
not I_19(n12_6,G214_4_l_6);
nor I_20(n4_1_r_6,n28_6,n22_6);
nor I_21(N1_4_r_6,n12_6,n24_6);
nor I_22(n_42_2_l_6,IN_1_2_l_6,IN_3_2_l_6);
DFFARX1 I_23(G214_4_l_6,blif_clk_net_1_r_17,n6_17,P6_5_r_internal_6,);
nand I_24(n19_6,IN_4_3_l_6,n26_6);
not I_25(n20_6,n_42_2_l_6);
nor I_26(n21_6,n17_6,n28_6);
and I_27(n22_6,IN_4_3_l_6,n26_6);
nand I_28(n23_6,IN_2_2_l_6,IN_3_2_l_6);
nor I_29(n24_6,n17_6,n18_6);
nand I_30(n25_6,IN_1_4_l_6,IN_2_4_l_6);
DFFARX1 I_31(n4_1_r_17,blif_clk_net_1_r_17,n6_17,G42_1_r_17,);
nor I_32(n_572_1_r_17,ACVQN1_5_l_17,n19_17);
nand I_33(n_573_1_r_17,n20_17,n21_17);
nand I_34(n_549_1_r_17,n23_17,n24_17);
nand I_35(n_569_1_r_17,n21_17,n22_17);
not I_36(n_452_1_r_17,n23_17);
DFFARX1 I_37(n19_17,blif_clk_net_1_r_17,n6_17,ACVQN2_3_r_17,);
nor I_38(n_266_and_0_3_r_17,n17_17,n29_17);
DFFARX1 I_39(N1_4_r_17,blif_clk_net_1_r_17,n6_17,G199_4_r_17,);
DFFARX1 I_40(n5_17,blif_clk_net_1_r_17,n6_17,G214_4_r_17,);
or I_41(n_431_0_l_17,n26_17,G199_4_r_6);
not I_42(n6_17,blif_reset_net_1_r_17);
DFFARX1 I_43(n_431_0_l_17,blif_clk_net_1_r_17,n6_17,n20_internal_17,);
not I_44(n20_17,n20_internal_17);
DFFARX1 I_45(G42_1_r_6,blif_clk_net_1_r_17,n6_17,ACVQN1_5_l_17,);
DFFARX1 I_46(n_573_1_r_6,blif_clk_net_1_r_17,n6_17,n19_internal_17,);
not I_47(n19_17,n19_internal_17);
nor I_48(n4_1_r_17,n5_17,n25_17);
not I_49(n2_17,n29_17);
DFFARX1 I_50(n2_17,blif_clk_net_1_r_17,n6_17,n17_internal_17,);
not I_51(n17_17,n17_internal_17);
nor I_52(N1_4_r_17,n29_17,n31_17);
not I_53(n5_17,n_452_1_r_6);
and I_54(n21_17,n32_17,P6_5_r_6);
not I_55(n22_17,n25_17);
nand I_56(n23_17,n20_17,n22_17);
nand I_57(n24_17,n19_17,n22_17);
nand I_58(n25_17,n30_17,ACVQN1_5_r_6);
and I_59(n26_17,n27_17,G214_4_r_6);
nor I_60(n27_17,n28_17,n_549_1_r_6);
not I_61(n28_17,n_569_1_r_6);
nor I_62(n29_17,n28_17,n_572_1_r_6);
and I_63(n30_17,n5_17,n_572_1_r_6);
nor I_64(n31_17,n21_17,n_452_1_r_6);
nor I_65(n32_17,G42_1_r_6,n_452_1_r_6);
endmodule


