module test_I7365(I5385,I1477,I5416,I5156,I5094,I3380,I5642,I1470,I7365);
input I5385,I1477,I5416,I5156,I5094,I3380,I5642,I1470;
output I7365;
wire I6941,I5067,I6907,I5249,I5481,I5091,I7269,I6958,I5070,I7026,I5105,I7348;
nor I_0(I6941,I5070,I5094);
and I_1(I7365,I7026,I7348);
DFFARX1 I_2(I5642,I1470,I5105,,,I5067,);
not I_3(I6907,I1477);
not I_4(I5249,I3380);
DFFARX1 I_5(I5416,I1470,I5105,,,I5481,);
nand I_6(I5091,I5156,I5385);
DFFARX1 I_7(I5067,I1470,I6907,,,I7269,);
nand I_8(I6958,I6941,I5091);
and I_9(I5070,I5249,I5481);
not I_10(I7026,I5070);
not I_11(I5105,I1477);
nand I_12(I7348,I7269,I6958);
endmodule


