module test_I13171(I13392,I11720,I1477,I11281,I11830,I1470,I13171);
input I13392,I11720,I1477,I11281,I11830,I1470;
output I13171;
wire I13214,I13231,I11290,I13197,I13426,I11275,I11302,I13460,I13248,I13409;
nand I_0(I13214,I11275,I11302);
and I_1(I13231,I13214,I11290);
nand I_2(I11290,I11830,I11720);
not I_3(I13197,I1477);
DFFARX1 I_4(I13409,I1470,I13197,,,I13426,);
DFFARX1 I_5(I1470,,,I11275,);
DFFARX1 I_6(I1470,,,I11302,);
not I_7(I13460,I13426);
nand I_8(I13171,I13248,I13460);
DFFARX1 I_9(I13231,I1470,I13197,,,I13248,);
and I_10(I13409,I13392,I11281);
endmodule


