module test_final(IN_1_0_l_15,IN_2_0_l_15,IN_3_0_l_15,IN_4_0_l_15,IN_1_1_l_15,IN_2_1_l_15,IN_3_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_3_3_l_15,IN_1_6_l_15,IN_2_6_l_15,IN_3_6_l_15,IN_4_6_l_15,IN_5_6_l_15,blif_clk_net_8_r_6,blif_reset_net_8_r_6,N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,N1372_10_r_6,N1508_10_r_6);
input IN_1_0_l_15,IN_2_0_l_15,IN_3_0_l_15,IN_4_0_l_15,IN_1_1_l_15,IN_2_1_l_15,IN_3_1_l_15,IN_1_3_l_15,IN_2_3_l_15,IN_3_3_l_15,IN_1_6_l_15,IN_2_6_l_15,IN_3_6_l_15,IN_4_6_l_15,IN_5_6_l_15,blif_clk_net_8_r_6,blif_reset_net_8_r_6;
output N1371_0_r_6,N1508_0_r_6,N1372_1_r_6,N1508_1_r_6,N1507_6_r_6,N1508_6_r_6,n_42_8_r_6,G199_8_r_6,N6147_9_r_6,N6134_9_r_6,N1372_10_r_6,N1508_10_r_6;
wire N1371_0_r_15,N1508_0_r_15,N1372_1_r_15,N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_102_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15,n_431_5_r_15,n31_15,n32_15,n33_15,n34_15,n35_15,n36_15,n37_15,n38_15,n39_15,n40_15,n41_15,n42_15,n43_15,n44_15,n45_15,n46_15,n47_15,n48_15,n49_15,n50_15,n51_15,n52_15,n53_15,n54_15,n55_15,I_BUFF_1_9_r_6,N3_8_r_6,n9_6,n30_6,n31_6,n32_6,n33_6,n34_6,n35_6,n36_6,n37_6,n38_6,n39_6,n40_6,n41_6,n42_6,n43_6,n44_6,n45_6,n46_6,n47_6,n48_6,n49_6,n50_6,n51_6,n52_6,n53_6,n54_6;
and I_0(N1371_0_r_15,N1508_0_r_15,n_102_5_r_15);
nor I_1(N1508_0_r_15,IN_2_0_l_15,n55_15);
nor I_2(N1372_1_r_15,n_102_5_r_15,n46_15);
nor I_3(N1508_1_r_15,N1508_0_r_15,n45_15);
not I_4(N1372_4_r_15,n39_15);
nor I_5(N1508_4_r_15,n39_15,n43_15);
nand I_6(n_429_or_0_5_r_15,n36_15,n38_15);
DFFARX1 I_7(n_431_5_r_15,blif_clk_net_8_r_6,n9_6,G78_5_r_15,);
nand I_8(n_576_5_r_15,n31_15,n32_15);
not I_9(n_102_5_r_15,n33_15);
nand I_10(n_547_5_r_15,N1371_0_r_15,n35_15);
nor I_11(N1507_6_r_15,n42_15,n46_15);
nand I_12(N1508_6_r_15,n39_15,n40_15);
nand I_13(n_431_5_r_15,n36_15,n37_15);
nor I_14(n31_15,n33_15,n34_15);
nor I_15(n32_15,IN_1_3_l_15,n44_15);
nor I_16(n33_15,n54_15,n55_15);
nand I_17(n34_15,IN_2_6_l_15,n49_15);
nand I_18(n35_15,IN_1_1_l_15,IN_2_1_l_15);
not I_19(n36_15,n32_15);
nand I_20(n37_15,n34_15,n38_15);
not I_21(n38_15,n46_15);
nand I_22(n39_15,n38_15,n41_15);
nand I_23(n40_15,n41_15,n42_15);
and I_24(n41_15,IN_5_6_l_15,n51_15);
and I_25(n42_15,IN_2_1_l_15,n47_15);
and I_26(n43_15,n34_15,n36_15);
or I_27(n44_15,IN_2_3_l_15,IN_3_3_l_15);
not I_28(n45_15,N1372_1_r_15);
nand I_29(n46_15,IN_2_1_l_15,n53_15);
nor I_30(n47_15,n34_15,n48_15);
not I_31(n48_15,IN_1_1_l_15);
and I_32(n49_15,IN_1_6_l_15,n50_15);
nand I_33(n50_15,n51_15,n52_15);
nand I_34(n51_15,IN_3_6_l_15,IN_4_6_l_15);
not I_35(n52_15,IN_5_6_l_15);
nor I_36(n53_15,IN_3_1_l_15,n48_15);
nor I_37(n54_15,IN_3_0_l_15,IN_4_0_l_15);
not I_38(n55_15,IN_1_0_l_15);
nor I_39(N1371_0_r_6,n30_6,n33_6);
nor I_40(N1508_0_r_6,n33_6,n44_6);
not I_41(N1372_1_r_6,n41_6);
nor I_42(N1508_1_r_6,n40_6,n41_6);
nor I_43(N1507_6_r_6,n39_6,n45_6);
nor I_44(N1508_6_r_6,n37_6,n38_6);
nor I_45(n_42_8_r_6,n30_6,n31_6);
DFFARX1 I_46(N3_8_r_6,blif_clk_net_8_r_6,n9_6,G199_8_r_6,);
nor I_47(N6147_9_r_6,n32_6,n33_6);
nor I_48(N6134_9_r_6,I_BUFF_1_9_r_6,n35_6);
not I_49(I_BUFF_1_9_r_6,n37_6);
not I_50(N1372_10_r_6,n43_6);
nor I_51(N1508_10_r_6,n42_6,n43_6);
nor I_52(N3_8_r_6,n36_6,N1508_6_r_15);
not I_53(n9_6,blif_reset_net_8_r_6);
nor I_54(n30_6,n53_6,N1508_4_r_15);
not I_55(n31_6,n36_6);
nor I_56(n32_6,I_BUFF_1_9_r_6,n34_6);
not I_57(n33_6,N1508_6_r_15);
not I_58(n34_6,n35_6);
nand I_59(n35_6,n49_6,N1508_4_r_15);
nand I_60(n36_6,n51_6,N1508_1_r_15);
nand I_61(n37_6,n54_6,N1507_6_r_15);
or I_62(n38_6,n35_6,n39_6);
nor I_63(n39_6,n40_6,n45_6);
and I_64(n40_6,n46_6,n47_6);
nand I_65(n41_6,n30_6,n31_6);
nor I_66(n42_6,n34_6,n40_6);
nand I_67(n43_6,n30_6,N1508_6_r_15);
nor I_68(n44_6,n31_6,n40_6);
nor I_69(n45_6,n35_6,n36_6);
nor I_70(n46_6,N1372_4_r_15,n_429_or_0_5_r_15);
or I_71(n47_6,n48_6,N1372_4_r_15);
nor I_72(n48_6,n_576_5_r_15,G78_5_r_15);
and I_73(n49_6,n50_6,n_547_5_r_15);
nand I_74(n50_6,n51_6,n52_6);
nand I_75(n51_6,G78_5_r_15,n_429_or_0_5_r_15);
not I_76(n52_6,N1508_1_r_15);
nor I_77(n53_6,N1508_1_r_15,n_576_5_r_15);
or I_78(n54_6,N1508_1_r_15,n_576_5_r_15);
endmodule


