module test_I1828(I1231,I1215,I1294,I1301,I1287,I1239,I1828);
input I1231,I1215,I1294,I1301,I1287,I1239;
output I1828;
wire I1376,I1342,I1359,I1393,I1780;
and I_0(I1376,I1359,I1231);
not I_1(I1342,I1301);
nand I_2(I1359,I1287,I1239);
nor I_3(I1828,I1780,I1393);
DFFARX1 I_4(I1376,I1294,I1342,,,I1393,);
DFFARX1 I_5(I1215,I1294,I1342,,,I1780,);
endmodule


