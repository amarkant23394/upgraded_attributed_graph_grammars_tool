module test_I7541(I1477,I6843,I1470,I6363,I7541);
input I1477,I6843,I1470,I6363;
output I7541;
wire I6297,I6300,I7652,I7570,I7587,I6380,I6329,I6318,I7669;
DFFARX1 I_0(I6843,I1470,I6329,,,I6297,);
DFFARX1 I_1(I1470,I6329,,,I6300,);
nor I_2(I7652,I7587,I6297);
not I_3(I7570,I1477);
not I_4(I7587,I6300);
DFFARX1 I_5(I6363,I1470,I6329,,,I6380,);
not I_6(I6329,I1477);
not I_7(I6318,I6380);
DFFARX1 I_8(I7669,I1470,I7570,,,I7541,);
nand I_9(I7669,I7652,I6318);
endmodule


