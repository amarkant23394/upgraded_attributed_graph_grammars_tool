module test_final(IN_1_1_l_16,IN_2_1_l_16,IN_3_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_3_3_l_16,IN_1_6_l_16,IN_2_6_l_16,IN_3_6_l_16,IN_4_6_l_16,IN_5_6_l_16,IN_1_8_l_16,IN_2_8_l_16,IN_3_8_l_16,IN_6_8_l_16,blif_clk_net_5_r_9,blif_reset_net_5_r_9,N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,G78_5_r_9,n_576_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9);
input IN_1_1_l_16,IN_2_1_l_16,IN_3_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_3_3_l_16,IN_1_6_l_16,IN_2_6_l_16,IN_3_6_l_16,IN_4_6_l_16,IN_5_6_l_16,IN_1_8_l_16,IN_2_8_l_16,IN_3_8_l_16,IN_6_8_l_16,blif_clk_net_5_r_9,blif_reset_net_5_r_9;
output N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,G78_5_r_9,n_576_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9;
wire N1371_0_r_16,N1508_0_r_16,N1372_1_r_16,N1508_1_r_16,N6147_2_r_16,N1507_6_r_16,N1508_6_r_16,G42_7_r_16,n_572_7_r_16,n_573_7_r_16,n_549_7_r_16,n_569_7_r_16,n_452_7_r_16,N3_8_l_16,n53_16,n29_16,n4_7_r_16,n30_16,n31_16,n32_16,n33_16,n34_16,n35_16,n36_16,n37_16,n38_16,n39_16,n40_16,n41_16,n42_16,n43_16,n44_16,n45_16,n46_16,n47_16,n48_16,n49_16,n50_16,n51_16,n52_16,n_429_or_0_5_r_9,n_102_5_r_9,I_BUFF_1_9_r_9,n4_7_l_9,n10_9,n62_9,N3_8_l_9,n63_9,n38_9,n_431_5_r_9,N3_8_r_9,n39_9,n40_9,n41_9,n42_9,n43_9,n44_9,n45_9,n46_9,n47_9,n48_9,n49_9,n50_9,n51_9,n52_9,n53_9,n54_9,n55_9,n56_9,n57_9,n58_9,n59_9,n60_9,n61_9;
nor I_0(N1371_0_r_16,n35_16,n39_16);
nor I_1(N1508_0_r_16,n39_16,n46_16);
not I_2(N1372_1_r_16,n45_16);
nor I_3(N1508_1_r_16,n53_16,n45_16);
nor I_4(N6147_2_r_16,n37_16,n38_16);
nor I_5(N1507_6_r_16,n44_16,n49_16);
nor I_6(N1508_6_r_16,n29_16,n42_16);
DFFARX1 I_7(n4_7_r_16,blif_clk_net_5_r_9,n10_9,G42_7_r_16,);
nor I_8(n_572_7_r_16,n32_16,n33_16);
nand I_9(n_573_7_r_16,n30_16,n31_16);
nand I_10(n_549_7_r_16,IN_5_6_l_16,n47_16);
nand I_11(n_569_7_r_16,n_549_7_r_16,n30_16);
nor I_12(n_452_7_r_16,n34_16,n35_16);
and I_13(N3_8_l_16,IN_6_8_l_16,n41_16);
DFFARX1 I_14(N3_8_l_16,blif_clk_net_5_r_9,n10_9,n53_16,);
not I_15(n29_16,n53_16);
nor I_16(n4_7_r_16,n35_16,n36_16);
nand I_17(n30_16,IN_1_1_l_16,IN_2_1_l_16);
not I_18(n31_16,n34_16);
nor I_19(n32_16,IN_3_1_l_16,n30_16);
not I_20(n33_16,n_549_7_r_16);
nor I_21(n34_16,IN_1_3_l_16,n48_16);
and I_22(n35_16,IN_2_6_l_16,n50_16);
not I_23(n36_16,n30_16);
nor I_24(n37_16,n31_16,n40_16);
nand I_25(n38_16,n29_16,n39_16);
not I_26(n39_16,n32_16);
nor I_27(n40_16,IN_1_8_l_16,IN_3_8_l_16);
nand I_28(n41_16,IN_2_8_l_16,IN_3_8_l_16);
nand I_29(n42_16,n35_16,n43_16);
not I_30(n43_16,n44_16);
nor I_31(n44_16,n32_16,n49_16);
nand I_32(n45_16,n36_16,n40_16);
nor I_33(n46_16,n33_16,n34_16);
nand I_34(n47_16,IN_3_6_l_16,IN_4_6_l_16);
or I_35(n48_16,IN_2_3_l_16,IN_3_3_l_16);
and I_36(n49_16,n35_16,n36_16);
and I_37(n50_16,IN_1_6_l_16,n51_16);
nand I_38(n51_16,n47_16,n52_16);
not I_39(n52_16,IN_5_6_l_16);
nor I_40(N6147_2_r_9,n62_9,n46_9);
not I_41(N1372_4_r_9,n59_9);
nor I_42(N1508_4_r_9,n58_9,n59_9);
nand I_43(n_429_or_0_5_r_9,n_431_5_r_9,n42_9);
DFFARX1 I_44(n_431_5_r_9,blif_clk_net_5_r_9,n10_9,G78_5_r_9,);
nand I_45(n_576_5_r_9,n39_9,n40_9);
not I_46(n_102_5_r_9,I_BUFF_1_9_r_9);
nand I_47(n_547_5_r_9,n43_9,N1371_0_r_16);
and I_48(n_42_8_r_9,n44_9,G42_7_r_16);
DFFARX1 I_49(N3_8_r_9,blif_clk_net_5_r_9,n10_9,G199_8_r_9,);
nor I_50(N6147_9_r_9,n41_9,n45_9);
nor I_51(N6134_9_r_9,n45_9,n51_9);
nor I_52(I_BUFF_1_9_r_9,n41_9,N1371_0_r_16);
nor I_53(n4_7_l_9,N1507_6_r_16,G42_7_r_16);
not I_54(n10_9,blif_reset_net_5_r_9);
DFFARX1 I_55(n4_7_l_9,blif_clk_net_5_r_9,n10_9,n62_9,);
and I_56(N3_8_l_9,n57_9,n_572_7_r_16);
DFFARX1 I_57(N3_8_l_9,blif_clk_net_5_r_9,n10_9,n63_9,);
not I_58(n38_9,n63_9);
nor I_59(n_431_5_r_9,N1508_0_r_16,n_452_7_r_16);
nor I_60(N3_8_r_9,n_102_5_r_9,n53_9);
nor I_61(n39_9,I_BUFF_1_9_r_9,n42_9);
not I_62(n40_9,n41_9);
nand I_63(n41_9,N1508_6_r_16,n_569_7_r_16);
nor I_64(n42_9,N1508_1_r_16,n_573_7_r_16);
nor I_65(n43_9,n63_9,n41_9);
nor I_66(n44_9,n_573_7_r_16,N1372_1_r_16);
and I_67(n45_9,n52_9,N1372_1_r_16);
nor I_68(n46_9,n47_9,n48_9);
nor I_69(n47_9,n49_9,n50_9);
not I_70(n48_9,n_429_or_0_5_r_9);
not I_71(n49_9,n42_9);
or I_72(n50_9,n63_9,n51_9);
nor I_73(n51_9,N1371_0_r_16,N6147_2_r_16);
nor I_74(n52_9,n49_9,N1508_0_r_16);
nor I_75(n53_9,n54_9,n55_9);
nor I_76(n54_9,n56_9,N1508_0_r_16);
or I_77(n55_9,n44_9,N1508_1_r_16);
not I_78(n56_9,N1372_1_r_16);
nand I_79(n57_9,N1371_0_r_16,N1508_0_r_16);
nor I_80(n58_9,n62_9,n60_9);
nand I_81(n59_9,n51_9,n61_9);
nor I_82(n60_9,n38_9,n44_9);
nor I_83(n61_9,G42_7_r_16,N1372_1_r_16);
endmodule


