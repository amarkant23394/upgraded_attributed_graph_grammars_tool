module test_final(IN_1_2_l_0,IN_2_2_l_0,IN_3_2_l_0,IN_4_2_l_0,IN_5_2_l_0,IN_1_4_l_0,IN_2_4_l_0,IN_3_4_l_0,IN_4_4_l_0,IN_5_4_l_0,IN_1_9_l_0,IN_2_9_l_0,IN_3_9_l_0,IN_4_9_l_0,IN_5_9_l_0,blif_clk_net_5_r_15,blif_reset_net_5_r_15,N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15);
input IN_1_2_l_0,IN_2_2_l_0,IN_3_2_l_0,IN_4_2_l_0,IN_5_2_l_0,IN_1_4_l_0,IN_2_4_l_0,IN_3_4_l_0,IN_4_4_l_0,IN_5_4_l_0,IN_1_9_l_0,IN_2_9_l_0,IN_3_9_l_0,IN_4_9_l_0,IN_5_9_l_0,blif_clk_net_5_r_15,blif_reset_net_5_r_15;
output N1508_1_r_15,N1372_4_r_15,N1508_4_r_15,n_429_or_0_5_r_15,G78_5_r_15,n_576_5_r_15,n_547_5_r_15,N1507_6_r_15,N1508_6_r_15;
wire N1371_0_r_0,N1508_0_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_102_5_r_0,n_547_5_r_0,G42_7_r_0,n_572_7_r_0,n_573_7_r_0,n_549_7_r_0,n_569_7_r_0,n_452_7_r_0,n_431_5_r_0,n4_7_r_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0,n37_0,n38_0,n39_0,n40_0,n41_0,n42_0,n43_0,n44_0,n45_0,N1371_0_r_15,N1508_0_r_15,N1372_1_r_15,n_102_5_r_15,n_431_5_r_15,n9_15,n31_15,n32_15,n33_15,n34_15,n35_15,n36_15,n37_15,n38_15,n39_15,n40_15,n41_15,n42_15,n43_15,n44_15,n45_15,n46_15,n47_15,n48_15,n49_15,n50_15,n51_15,n52_15,n53_15,n54_15,n55_15;
nor I_0(N1371_0_r_0,n_102_5_r_0,n29_0);
nor I_1(N1508_0_r_0,n_102_5_r_0,n_452_7_r_0);
or I_2(n_429_or_0_5_r_0,IN_1_9_l_0,n38_0);
DFFARX1 I_3(n_431_5_r_0,blif_clk_net_5_r_15,n9_15,G78_5_r_0,);
nand I_4(n_576_5_r_0,IN_1_9_l_0,n26_0);
not I_5(n_102_5_r_0,n27_0);
nand I_6(n_547_5_r_0,n30_0,n34_0);
DFFARX1 I_7(n4_7_r_0,blif_clk_net_5_r_15,n9_15,G42_7_r_0,);
nor I_8(n_572_7_r_0,IN_1_9_l_0,n31_0);
or I_9(n_573_7_r_0,n29_0,n30_0);
nor I_10(n_549_7_r_0,n29_0,n33_0);
nand I_11(n_569_7_r_0,n28_0,n32_0);
nor I_12(n_452_7_r_0,n30_0,n31_0);
nand I_13(n_431_5_r_0,n_102_5_r_0,n35_0);
nor I_14(n4_7_r_0,n31_0,n37_0);
nor I_15(n26_0,n27_0,n28_0);
nor I_16(n27_0,n28_0,n44_0);
nand I_17(n28_0,IN_1_4_l_0,IN_2_4_l_0);
not I_18(n29_0,n32_0);
nor I_19(n30_0,IN_5_9_l_0,n39_0);
not I_20(n31_0,n38_0);
nand I_21(n32_0,n41_0,n42_0);
nor I_22(n33_0,IN_1_9_l_0,n_102_5_r_0);
nor I_23(n34_0,IN_1_9_l_0,n27_0);
nand I_24(n35_0,n29_0,n36_0);
nor I_25(n36_0,n37_0,n38_0);
not I_26(n37_0,n28_0);
nand I_27(n38_0,IN_2_9_l_0,n40_0);
nor I_28(n39_0,IN_3_9_l_0,IN_4_9_l_0);
or I_29(n40_0,IN_3_9_l_0,IN_4_9_l_0);
nor I_30(n41_0,IN_1_2_l_0,IN_2_2_l_0);
or I_31(n42_0,IN_5_2_l_0,n43_0);
nor I_32(n43_0,IN_3_2_l_0,IN_4_2_l_0);
nor I_33(n44_0,IN_5_4_l_0,n45_0);
and I_34(n45_0,IN_3_4_l_0,IN_4_4_l_0);
and I_35(N1371_0_r_15,N1508_0_r_15,n_102_5_r_15);
nor I_36(N1508_0_r_15,n55_15,N1508_0_r_0);
nor I_37(N1372_1_r_15,n_102_5_r_15,n46_15);
nor I_38(N1508_1_r_15,N1508_0_r_15,n45_15);
not I_39(N1372_4_r_15,n39_15);
nor I_40(N1508_4_r_15,n39_15,n43_15);
nand I_41(n_429_or_0_5_r_15,n36_15,n38_15);
DFFARX1 I_42(n_431_5_r_15,blif_clk_net_5_r_15,n9_15,G78_5_r_15,);
nand I_43(n_576_5_r_15,n31_15,n32_15);
not I_44(n_102_5_r_15,n33_15);
nand I_45(n_547_5_r_15,N1371_0_r_15,n35_15);
nor I_46(N1507_6_r_15,n42_15,n46_15);
nand I_47(N1508_6_r_15,n39_15,n40_15);
nand I_48(n_431_5_r_15,n36_15,n37_15);
not I_49(n9_15,blif_reset_net_5_r_15);
nor I_50(n31_15,n33_15,n34_15);
nor I_51(n32_15,n44_15,n_572_7_r_0);
nor I_52(n33_15,n54_15,n55_15);
nand I_53(n34_15,n49_15,G42_7_r_0);
nand I_54(n35_15,G78_5_r_0,n_569_7_r_0);
not I_55(n36_15,n32_15);
nand I_56(n37_15,n34_15,n38_15);
not I_57(n38_15,n46_15);
nand I_58(n39_15,n38_15,n41_15);
nand I_59(n40_15,n41_15,n42_15);
and I_60(n41_15,n51_15,n_576_5_r_0);
and I_61(n42_15,n47_15,G78_5_r_0);
and I_62(n43_15,n34_15,n36_15);
or I_63(n44_15,N1508_0_r_0,n_573_7_r_0);
not I_64(n45_15,N1372_1_r_15);
nand I_65(n46_15,n53_15,G78_5_r_0);
nor I_66(n47_15,n34_15,n48_15);
not I_67(n48_15,n_569_7_r_0);
and I_68(n49_15,n50_15,n_547_5_r_0);
nand I_69(n50_15,n51_15,n52_15);
nand I_70(n51_15,N1371_0_r_0,n_429_or_0_5_r_0);
not I_71(n52_15,n_576_5_r_0);
nor I_72(n53_15,n48_15,n_549_7_r_0);
nor I_73(n54_15,N1371_0_r_0,n_429_or_0_5_r_0);
not I_74(n55_15,G78_5_r_0);
endmodule


