module test_I17967(I1477,I15662,I15832,I15897,I1470,I17967);
input I1477,I15662,I15832,I15897,I1470;
output I17967;
wire I17413,I16007,I15600,I15815,I15579,I15611,I17498,I15928,I15597,I17727,I17430,I17916,I15576,I17950,I15603,I17933,I15976,I17481;
not I_0(I17413,I1477);
or I_1(I16007,I15928,I15897);
or I_2(I15600,I15832,I15815);
DFFARX1 I_3(I1470,I15611,,,I15815,);
nand I_4(I15579,I15662,I15976);
not I_5(I15611,I1477);
nand I_6(I17498,I17481,I15600);
DFFARX1 I_7(I1470,I15611,,,I15928,);
and I_8(I17967,I17727,I17950);
nor I_9(I15597,I15832);
nand I_10(I17727,I17430,I15576);
not I_11(I17430,I15579);
DFFARX1 I_12(I15603,I1470,I17413,,,I17916,);
DFFARX1 I_13(I16007,I1470,I15611,,,I15576,);
nand I_14(I17950,I17933,I17498);
nor I_15(I15603,I15928);
not I_16(I17933,I17916);
nor I_17(I15976,I15928);
nor I_18(I17481,I17430,I15597);
endmodule


