module test_I11429(I9320,I6884,I6992,I7057,I6887,I11429);
input I9320,I6884,I6992,I7057,I6887;
output I11429;
wire I9396,I8930,I6881,I8879,I8848,I9083,I9413,I8947;
not I_0(I9396,I9320);
not I_1(I11429,I8848);
nor I_2(I8930,I8879);
nand I_3(I6881,I6992,I7057);
not I_4(I8879,I6887);
nor I_5(I8848,I9083,I9413);
nand I_6(I9083,I8879,I6881);
and I_7(I9413,I8947,I9396);
nand I_8(I8947,I8930,I6884);
endmodule


