module test_final(IN_1_2_l_0,IN_2_2_l_0,IN_3_2_l_0,IN_4_2_l_0,IN_5_2_l_0,IN_1_4_l_0,IN_2_4_l_0,IN_3_4_l_0,IN_4_4_l_0,IN_5_4_l_0,IN_1_9_l_0,IN_2_9_l_0,IN_3_9_l_0,IN_4_9_l_0,IN_5_9_l_0,blif_clk_net_7_r_5,blif_reset_net_7_r_5,N1371_0_r_5,N1508_0_r_5,N1372_1_r_5,N1508_1_r_5,N6147_2_r_5,N1507_6_r_5,N1508_6_r_5,G42_7_r_5,n_572_7_r_5,n_573_7_r_5,n_569_7_r_5,n_452_7_r_5);
input IN_1_2_l_0,IN_2_2_l_0,IN_3_2_l_0,IN_4_2_l_0,IN_5_2_l_0,IN_1_4_l_0,IN_2_4_l_0,IN_3_4_l_0,IN_4_4_l_0,IN_5_4_l_0,IN_1_9_l_0,IN_2_9_l_0,IN_3_9_l_0,IN_4_9_l_0,IN_5_9_l_0,blif_clk_net_7_r_5,blif_reset_net_7_r_5;
output N1371_0_r_5,N1508_0_r_5,N1372_1_r_5,N1508_1_r_5,N6147_2_r_5,N1507_6_r_5,N1508_6_r_5,G42_7_r_5,n_572_7_r_5,n_573_7_r_5,n_569_7_r_5,n_452_7_r_5;
wire N1371_0_r_0,N1508_0_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_102_5_r_0,n_547_5_r_0,G42_7_r_0,n_572_7_r_0,n_573_7_r_0,n_549_7_r_0,n_569_7_r_0,n_452_7_r_0,n_431_5_r_0,n4_7_r_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0,n37_0,n38_0,n39_0,n40_0,n41_0,n42_0,n43_0,n44_0,n45_0,n_549_7_r_5,n4_7_r_5,n7_5,n26_5,n27_5,n28_5,n29_5,n30_5,n31_5,n32_5,n33_5,n34_5,n35_5,n36_5,n37_5,n38_5,n39_5,n40_5,n41_5,n42_5,n43_5,n44_5,n45_5,n46_5,n47_5;
nor I_0(N1371_0_r_0,n_102_5_r_0,n29_0);
nor I_1(N1508_0_r_0,n_102_5_r_0,n_452_7_r_0);
or I_2(n_429_or_0_5_r_0,IN_1_9_l_0,n38_0);
DFFARX1 I_3(n_431_5_r_0,blif_clk_net_7_r_5,n7_5,G78_5_r_0,);
nand I_4(n_576_5_r_0,IN_1_9_l_0,n26_0);
not I_5(n_102_5_r_0,n27_0);
nand I_6(n_547_5_r_0,n30_0,n34_0);
DFFARX1 I_7(n4_7_r_0,blif_clk_net_7_r_5,n7_5,G42_7_r_0,);
nor I_8(n_572_7_r_0,IN_1_9_l_0,n31_0);
or I_9(n_573_7_r_0,n29_0,n30_0);
nor I_10(n_549_7_r_0,n29_0,n33_0);
nand I_11(n_569_7_r_0,n28_0,n32_0);
nor I_12(n_452_7_r_0,n30_0,n31_0);
nand I_13(n_431_5_r_0,n_102_5_r_0,n35_0);
nor I_14(n4_7_r_0,n31_0,n37_0);
nor I_15(n26_0,n27_0,n28_0);
nor I_16(n27_0,n28_0,n44_0);
nand I_17(n28_0,IN_1_4_l_0,IN_2_4_l_0);
not I_18(n29_0,n32_0);
nor I_19(n30_0,IN_5_9_l_0,n39_0);
not I_20(n31_0,n38_0);
nand I_21(n32_0,n41_0,n42_0);
nor I_22(n33_0,IN_1_9_l_0,n_102_5_r_0);
nor I_23(n34_0,IN_1_9_l_0,n27_0);
nand I_24(n35_0,n29_0,n36_0);
nor I_25(n36_0,n37_0,n38_0);
not I_26(n37_0,n28_0);
nand I_27(n38_0,IN_2_9_l_0,n40_0);
nor I_28(n39_0,IN_3_9_l_0,IN_4_9_l_0);
or I_29(n40_0,IN_3_9_l_0,IN_4_9_l_0);
nor I_30(n41_0,IN_1_2_l_0,IN_2_2_l_0);
or I_31(n42_0,IN_5_2_l_0,n43_0);
nor I_32(n43_0,IN_3_2_l_0,IN_4_2_l_0);
nor I_33(n44_0,IN_5_4_l_0,n45_0);
and I_34(n45_0,IN_3_4_l_0,IN_4_4_l_0);
nor I_35(N1371_0_r_5,n28_5,n46_5);
nand I_36(N1508_0_r_5,n26_5,n43_5);
not I_37(N1372_1_r_5,n43_5);
nor I_38(N1508_1_r_5,n30_5,n43_5);
nor I_39(N6147_2_r_5,n29_5,n32_5);
nor I_40(N1507_6_r_5,n26_5,n44_5);
nor I_41(N1508_6_r_5,n27_5,n37_5);
DFFARX1 I_42(n4_7_r_5,blif_clk_net_7_r_5,n7_5,G42_7_r_5,);
and I_43(n_572_7_r_5,n27_5,n28_5);
nand I_44(n_573_7_r_5,n26_5,n27_5);
nand I_45(n_549_7_r_5,G42_7_r_0,n_569_7_r_0);
nand I_46(n_569_7_r_5,n_549_7_r_5,n26_5);
not I_47(n_452_7_r_5,n29_5);
nor I_48(n4_7_r_5,n30_5,n31_5);
not I_49(n7_5,blif_reset_net_7_r_5);
not I_50(n26_5,n35_5);
nand I_51(n27_5,n40_5,n41_5);
nand I_52(n28_5,G78_5_r_0,n_429_or_0_5_r_0);
nand I_53(n29_5,n27_5,n33_5);
nor I_54(n30_5,n45_5,N1371_0_r_0);
not I_55(n31_5,n_549_7_r_5);
nor I_56(n32_5,n34_5,n35_5);
not I_57(n33_5,n30_5);
nor I_58(n34_5,n31_5,n36_5);
nor I_59(n35_5,n28_5,n_549_7_r_0);
not I_60(n36_5,n28_5);
nand I_61(n37_5,n36_5,n38_5);
nand I_62(n38_5,n26_5,n39_5);
nand I_63(n39_5,n30_5,n31_5);
nor I_64(n40_5,N1371_0_r_0,G78_5_r_0);
or I_65(n41_5,n42_5,n_429_or_0_5_r_0);
nor I_66(n42_5,n_573_7_r_0,N1508_0_r_0);
nand I_67(n43_5,n36_5,n46_5);
nor I_68(n44_5,n_549_7_r_5,n33_5);
or I_69(n45_5,N1508_0_r_0,n_547_5_r_0);
and I_70(n46_5,n31_5,n47_5);
or I_71(n47_5,n_576_5_r_0,n_572_7_r_0);
endmodule


