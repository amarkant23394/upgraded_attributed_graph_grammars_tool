module test_final(IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_4_2_l_10,IN_5_2_l_10,IN_1_6_l_10,IN_2_6_l_10,IN_3_6_l_10,IN_4_6_l_10,IN_5_6_l_10,IN_1_9_l_10,IN_2_9_l_10,IN_3_9_l_10,IN_4_9_l_10,IN_5_9_l_10,blif_clk_net_7_r_4,blif_reset_net_7_r_4,N1371_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6134_9_r_4);
input IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_4_2_l_10,IN_5_2_l_10,IN_1_6_l_10,IN_2_6_l_10,IN_3_6_l_10,IN_4_6_l_10,IN_5_6_l_10,IN_1_9_l_10,IN_2_9_l_10,IN_3_9_l_10,IN_4_9_l_10,IN_5_9_l_10,blif_clk_net_7_r_4,blif_reset_net_7_r_4;
output N1371_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6134_9_r_4;
wire N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1372_4_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10,I_BUFF_1_9_r_10,N3_8_r_10,n35_10,n36_10,n37_10,n38_10,n39_10,n40_10,n41_10,n42_10,n43_10,n44_10,n45_10,n46_10,n47_10,n48_10,n49_10,n50_10,n51_10,n52_10,n53_10,n54_10,n55_10,n56_10,n57_10,n58_10,n59_10,n60_10,n61_10,n62_10,n63_10,n64_10,N1508_0_r_4,n_573_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4,n4_7_r_4,n6_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4,n38_4,n39_4,n40_4,n41_4;
nor I_0(N1371_0_r_10,n37_10,n38_10);
nor I_1(N1508_0_r_10,n37_10,n58_10);
nand I_2(N6147_2_r_10,n39_10,n40_10);
not I_3(N6147_3_r_10,n39_10);
nor I_4(N1372_4_r_10,n46_10,n49_10);
nor I_5(N1508_4_r_10,n51_10,n52_10);
nor I_6(N1507_6_r_10,n49_10,n60_10);
nor I_7(N1508_6_r_10,n49_10,n50_10);
nor I_8(n_42_8_r_10,I_BUFF_1_9_r_10,n35_10);
DFFARX1 I_9(N3_8_r_10,blif_clk_net_7_r_4,n6_4,G199_8_r_10,);
nor I_10(N6147_9_r_10,n36_10,n37_10);
nor I_11(N6134_9_r_10,I_BUFF_1_9_r_10,n46_10);
not I_12(I_BUFF_1_9_r_10,n48_10);
nor I_13(N3_8_r_10,n44_10,n47_10);
not I_14(n35_10,n49_10);
nor I_15(n36_10,I_BUFF_1_9_r_10,n38_10);
not I_16(n37_10,IN_1_9_l_10);
not I_17(n38_10,n46_10);
nand I_18(n39_10,n43_10,n44_10);
nand I_19(n40_10,I_BUFF_1_9_r_10,n41_10);
nor I_20(n41_10,IN_1_9_l_10,n42_10);
not I_21(n42_10,n44_10);
nor I_22(n43_10,IN_1_9_l_10,n45_10);
nand I_23(n44_10,IN_2_6_l_10,n54_10);
nor I_24(n45_10,IN_5_9_l_10,n59_10);
nand I_25(n46_10,IN_2_9_l_10,n61_10);
nor I_26(n47_10,n46_10,n48_10);
nand I_27(n48_10,n62_10,n63_10);
nand I_28(n49_10,IN_5_6_l_10,n56_10);
not I_29(n50_10,n45_10);
nor I_30(n51_10,n42_10,n53_10);
not I_31(n52_10,N1372_4_r_10);
nor I_32(n53_10,n48_10,n50_10);
and I_33(n54_10,IN_1_6_l_10,n55_10);
nand I_34(n55_10,n56_10,n57_10);
nand I_35(n56_10,IN_3_6_l_10,IN_4_6_l_10);
not I_36(n57_10,IN_5_6_l_10);
nor I_37(n58_10,n35_10,n45_10);
nor I_38(n59_10,IN_3_9_l_10,IN_4_9_l_10);
nor I_39(n60_10,n37_10,n46_10);
or I_40(n61_10,IN_3_9_l_10,IN_4_9_l_10);
nor I_41(n62_10,IN_1_2_l_10,IN_2_2_l_10);
or I_42(n63_10,IN_5_2_l_10,n64_10);
nor I_43(n64_10,IN_3_2_l_10,IN_4_2_l_10);
nor I_44(N1371_0_r_4,n25_4,N1507_6_r_10);
not I_45(N1508_0_r_4,n25_4);
nor I_46(N1507_6_r_4,n32_4,n33_4);
nor I_47(N1508_6_r_4,n22_4,n29_4);
DFFARX1 I_48(n4_7_r_4,blif_clk_net_7_r_4,n6_4,G42_7_r_4,);
not I_49(n_572_7_r_4,n_573_7_r_4);
nand I_50(n_573_7_r_4,n21_4,n22_4);
nor I_51(n_549_7_r_4,n24_4,N1507_6_r_10);
nand I_52(n_569_7_r_4,n22_4,n23_4);
nor I_53(n_452_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4);
not I_54(N6147_9_r_4,n28_4);
nor I_55(N6134_9_r_4,N1508_0_r_4,n28_4);
not I_56(I_BUFF_1_9_r_4,n21_4);
nor I_57(n4_7_r_4,N6147_9_r_4,N1507_6_r_10);
not I_58(n6_4,blif_reset_net_7_r_4);
nand I_59(n21_4,n39_4,n40_4);
or I_60(n22_4,n31_4,N1371_0_r_10);
not I_61(n23_4,N1507_6_r_10);
nor I_62(n24_4,n25_4,n26_4);
nand I_63(n25_4,N6147_3_r_10,N1508_0_r_10);
nand I_64(n26_4,n21_4,n27_4);
nand I_65(n27_4,n36_4,n37_4);
nand I_66(n28_4,n38_4,N1371_0_r_10);
nand I_67(n29_4,N1508_0_r_4,n30_4);
nand I_68(n30_4,n34_4,n35_4);
nor I_69(n31_4,N6147_2_r_10,N6147_3_r_10);
not I_70(n32_4,n30_4);
nor I_71(n33_4,n21_4,n28_4);
nand I_72(n34_4,N6147_9_r_4,I_BUFF_1_9_r_4);
nand I_73(n35_4,N1508_0_r_4,n27_4);
not I_74(n36_4,N1508_6_r_10);
nand I_75(n37_4,N6147_9_r_10,N1508_4_r_10);
or I_76(n38_4,N6147_2_r_10,N6147_3_r_10);
nor I_77(n39_4,N1508_4_r_10,N6134_9_r_10);
or I_78(n40_4,n41_4,G199_8_r_10);
nor I_79(n41_4,N1508_0_r_10,n_42_8_r_10);
endmodule


