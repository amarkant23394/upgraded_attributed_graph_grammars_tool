module test_I15177(I13040,I12831,I12718,I10627,I12636,I1470_clk,I1477_rst,I15177);
input I13040,I12831,I12718,I10627,I12636,I1470_clk,I1477_rst;
output I15177;
wire I12599,I12653,I15143,I13057,I12619_rst,I15160,I12611,I12670,I12882,I12964,I12848,I12593;
nand I_0(I12599,I12718,I12964);
and I_1(I15177,I15160,I12593);
and I_2(I12653,I12636,I10627);
not I_3(I15143,I12599);
and I_4(I13057,I12718,I13040);
not I_5(I12619_rst,I1477_rst);
nor I_6(I15160,I15143,I12611);
DFFARX1 I_7 (I13057,I1470_clk,I12619_rst,I12611);
DFFARX1 I_8 (I12653,I1470_clk,I12619_rst,I12670);
not I_9(I12882,I12848);
nor I_10(I12964,I12882);
DFFARX1 I_11 (I12831,I1470_clk,I12619_rst,I12848);
nand I_12(I12593,I12670,I12882);
endmodule



//DFF Module (with asynch reset)
module DFFARX1(d, clock, reset, q);
	input d, clock, reset;
	output q;
	wire clock_inv, l1_x, l1_y, l1, l1_inv;
	wire l2_x, l2_y, q_inv, q_sync;
	not  dff0 (clock_inv, clock);
	nand dff1 (l1_x, d, clock_inv);
	nand dff2 (l1_y, l1_x, clock_inv);
	nand dff3 (l1, l1_x, l1_inv);
	nand dff4 (l1_inv, l1_y, l1);
	nand dff5 (l2_x, l1, clock);
	nand dff6 (l2_y, l2_x, clock);
	nand dff7 (q_sync, l2_x, q_inv);
	nand dff8 (q_inv, l2_y, q_sync);
	and  dff9 (q, q_sync, reset);
	and dff10 (q, q_sync, reset);
endmodule