module test_I10041(I8107,I1477,I7881,I6321,I1470,I10041);
input I8107,I1477,I7881,I6321,I1470;
output I10041;
wire I10120,I6297,I7538,I7731,I10052,I7977,I10349,I7898,I7714,I7946,I7535,I10332,I7550,I7570,I7915,I7532;
nor I_0(I10120,I7538,I7535);
DFFARX1 I_1(I1470,,,I6297,);
DFFARX1 I_2(I7915,I1470,I7570,,,I7538,);
nor I_3(I10041,I10349,I10120);
not I_4(I7731,I7714);
not I_5(I10052,I1477);
DFFARX1 I_6(I6321,I1470,I7570,,,I7977,);
and I_7(I10349,I10332,I7550);
nand I_8(I7898,I7881);
not I_9(I7714,I6297);
DFFARX1 I_10(I7881,I1470,I7570,,,I7946,);
and I_11(I7535,I7714,I7946);
DFFARX1 I_12(I7532,I1470,I10052,,,I10332,);
nand I_13(I7550,I7977,I7731);
not I_14(I7570,I1477);
and I_15(I7915,I7881,I7898);
DFFARX1 I_16(I8107,I1470,I7570,,,I7532,);
endmodule


