module test_I15897(I1477,I13749,I15781,I13843,I11944,I15628,I1470,I15897);
input I1477,I13749,I15781,I13843,I11944,I15628,I1470;
output I15897;
wire I13860,I13891,I15832,I15815,I15880,I13775,I15611,I13761,I15713,I13826,I13767,I15863,I15798;
nor I_0(I13860,I13843,I13826);
DFFARX1 I_1(I11944,I1470,I13775,,,I13891,);
nand I_2(I15832,I15628,I13749);
DFFARX1 I_3(I15798,I1470,I15611,,,I15815,);
nor I_4(I15880,I15815,I15863);
not I_5(I13775,I1477);
not I_6(I15611,I1477);
and I_7(I15897,I15713,I15880);
nand I_8(I13761,I13891,I13860);
not I_9(I15713,I13761);
DFFARX1 I_10(I1470,I13775,,,I13826,);
DFFARX1 I_11(I1470,I13775,,,I13767,);
not I_12(I15863,I15832);
or I_13(I15798,I15781,I13767);
endmodule


