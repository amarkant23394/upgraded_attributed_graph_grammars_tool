module test_I11412(I8830,I9049,I1470,I6881,I8879,I8862,I9413,I11412);
input I8830,I9049,I1470,I6881,I8879,I8862,I9413;
output I11412;
wire I11378,I9066,I11395,I8848,I11327,I9083,I8851;
nor I_0(I11378,I11327,I8848);
not I_1(I11412,I11395);
DFFARX1 I_2(I9049,I1470,I8862,,,I9066,);
nand I_3(I11395,I11378,I8851);
nor I_4(I8848,I9083,I9413);
not I_5(I11327,I8830);
nand I_6(I9083,I8879,I6881);
or I_7(I8851,I9083,I9066);
endmodule


