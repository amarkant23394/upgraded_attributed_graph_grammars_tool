module test_final(IN_1_0_l_11,IN_2_0_l_11,IN_3_0_l_11,IN_4_0_l_11,IN_1_1_l_11,IN_2_1_l_11,IN_3_1_l_11,IN_1_3_l_11,IN_2_3_l_11,IN_3_3_l_11,IN_1_6_l_11,IN_2_6_l_11,IN_3_6_l_11,IN_4_6_l_11,IN_5_6_l_11,blif_clk_net_5_r_9,blif_reset_net_5_r_9,N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,G78_5_r_9,n_576_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9);
input IN_1_0_l_11,IN_2_0_l_11,IN_3_0_l_11,IN_4_0_l_11,IN_1_1_l_11,IN_2_1_l_11,IN_3_1_l_11,IN_1_3_l_11,IN_2_3_l_11,IN_3_3_l_11,IN_1_6_l_11,IN_2_6_l_11,IN_3_6_l_11,IN_4_6_l_11,IN_5_6_l_11,blif_clk_net_5_r_9,blif_reset_net_5_r_9;
output N6147_2_r_9,N1372_4_r_9,N1508_4_r_9,G78_5_r_9,n_576_5_r_9,n_547_5_r_9,n_42_8_r_9,G199_8_r_9,N6147_9_r_9,N6134_9_r_9;
wire N1372_1_r_11,N1508_1_r_11,N6147_2_r_11,N6147_3_r_11,n_429_or_0_5_r_11,G78_5_r_11,n_576_5_r_11,n_102_5_r_11,n_547_5_r_11,N1507_6_r_11,N1508_6_r_11,N1372_10_r_11,N1508_10_r_11,n_431_5_r_11,n36_11,n37_11,n38_11,n39_11,n40_11,n41_11,n42_11,n43_11,n44_11,n45_11,n46_11,n47_11,n48_11,n49_11,n50_11,n51_11,n52_11,n53_11,n54_11,n55_11,n56_11,n57_11,n58_11,n59_11,n60_11,n61_11,n62_11,n63_11,n_429_or_0_5_r_9,n_102_5_r_9,I_BUFF_1_9_r_9,n4_7_l_9,n10_9,n62_9,N3_8_l_9,n63_9,n38_9,n_431_5_r_9,N3_8_r_9,n39_9,n40_9,n41_9,n42_9,n43_9,n44_9,n45_9,n46_9,n47_9,n48_9,n49_9,n50_9,n51_9,n52_9,n53_9,n54_9,n55_9,n56_9,n57_9,n58_9,n59_9,n60_9,n61_9;
not I_0(N1372_1_r_11,n53_11);
nor I_1(N1508_1_r_11,n39_11,n53_11);
nor I_2(N6147_2_r_11,n48_11,n49_11);
nor I_3(N6147_3_r_11,n44_11,n45_11);
nand I_4(n_429_or_0_5_r_11,n42_11,n43_11);
DFFARX1 I_5(n_431_5_r_11,blif_clk_net_5_r_9,n10_9,G78_5_r_11,);
nand I_6(n_576_5_r_11,n_102_5_r_11,N1372_10_r_11);
not I_7(n_102_5_r_11,n39_11);
nand I_8(n_547_5_r_11,n36_11,n37_11);
nor I_9(N1507_6_r_11,n52_11,n57_11);
nor I_10(N1508_6_r_11,n46_11,n51_11);
nor I_11(N1372_10_r_11,n43_11,n47_11);
nor I_12(N1508_10_r_11,n55_11,n56_11);
nand I_13(n_431_5_r_11,n40_11,n41_11);
nor I_14(n36_11,n38_11,n39_11);
not I_15(n37_11,n40_11);
nor I_16(n38_11,IN_2_0_l_11,n60_11);
nor I_17(n39_11,IN_1_3_l_11,n54_11);
nand I_18(n40_11,IN_1_1_l_11,IN_2_1_l_11);
nand I_19(n41_11,n_102_5_r_11,n42_11);
and I_20(n42_11,IN_2_6_l_11,n58_11);
not I_21(n43_11,n44_11);
nor I_22(n44_11,IN_3_1_l_11,n40_11);
nand I_23(n45_11,n46_11,n47_11);
not I_24(n46_11,n38_11);
nand I_25(n47_11,n59_11,n62_11);
and I_26(n48_11,n37_11,n47_11);
or I_27(n49_11,n44_11,n50_11);
nor I_28(n50_11,n60_11,n61_11);
or I_29(n51_11,n_102_5_r_11,n52_11);
nor I_30(n52_11,n42_11,n57_11);
nand I_31(n53_11,n37_11,n50_11);
or I_32(n54_11,IN_2_3_l_11,IN_3_3_l_11);
nor I_33(n55_11,n38_11,n42_11);
not I_34(n56_11,N1372_10_r_11);
and I_35(n57_11,n38_11,n50_11);
and I_36(n58_11,IN_1_6_l_11,n59_11);
or I_37(n59_11,IN_5_6_l_11,n63_11);
not I_38(n60_11,IN_1_0_l_11);
nor I_39(n61_11,IN_3_0_l_11,IN_4_0_l_11);
nand I_40(n62_11,IN_3_6_l_11,IN_4_6_l_11);
and I_41(n63_11,IN_3_6_l_11,IN_4_6_l_11);
nor I_42(N6147_2_r_9,n62_9,n46_9);
not I_43(N1372_4_r_9,n59_9);
nor I_44(N1508_4_r_9,n58_9,n59_9);
nand I_45(n_429_or_0_5_r_9,n_431_5_r_9,n42_9);
DFFARX1 I_46(n_431_5_r_9,blif_clk_net_5_r_9,n10_9,G78_5_r_9,);
nand I_47(n_576_5_r_9,n39_9,n40_9);
not I_48(n_102_5_r_9,I_BUFF_1_9_r_9);
nand I_49(n_547_5_r_9,n43_9,N1507_6_r_11);
and I_50(n_42_8_r_9,n44_9,N6147_2_r_11);
DFFARX1 I_51(N3_8_r_9,blif_clk_net_5_r_9,n10_9,G199_8_r_9,);
nor I_52(N6147_9_r_9,n41_9,n45_9);
nor I_53(N6134_9_r_9,n45_9,n51_9);
nor I_54(I_BUFF_1_9_r_9,n41_9,N1507_6_r_11);
nor I_55(n4_7_l_9,N6147_2_r_11,N1508_1_r_11);
not I_56(n10_9,blif_reset_net_5_r_9);
DFFARX1 I_57(n4_7_l_9,blif_clk_net_5_r_9,n10_9,n62_9,);
and I_58(N3_8_l_9,n57_9,N1372_1_r_11);
DFFARX1 I_59(N3_8_l_9,blif_clk_net_5_r_9,n10_9,n63_9,);
not I_60(n38_9,n63_9);
nor I_61(n_431_5_r_9,N6147_3_r_11,n_547_5_r_11);
nor I_62(N3_8_r_9,n_102_5_r_9,n53_9);
nor I_63(n39_9,I_BUFF_1_9_r_9,n42_9);
not I_64(n40_9,n41_9);
nand I_65(n41_9,n_429_or_0_5_r_11,n_576_5_r_11);
nor I_66(n42_9,N1372_1_r_11,N1508_6_r_11);
nor I_67(n43_9,n63_9,n41_9);
nor I_68(n44_9,N1508_6_r_11,N1508_10_r_11);
and I_69(n45_9,n52_9,G78_5_r_11);
nor I_70(n46_9,n47_9,n48_9);
nor I_71(n47_9,n49_9,n50_9);
not I_72(n48_9,n_429_or_0_5_r_9);
not I_73(n49_9,n42_9);
or I_74(n50_9,n63_9,n51_9);
nor I_75(n51_9,N1508_1_r_11,N6147_3_r_11);
nor I_76(n52_9,n49_9,n_547_5_r_11);
nor I_77(n53_9,n54_9,n55_9);
nor I_78(n54_9,n56_9,n_547_5_r_11);
or I_79(n55_9,n44_9,N1372_1_r_11);
not I_80(n56_9,G78_5_r_11);
nand I_81(n57_9,N1508_1_r_11,N6147_2_r_11);
nor I_82(n58_9,n62_9,n60_9);
nand I_83(n59_9,n51_9,n61_9);
nor I_84(n60_9,n38_9,n44_9);
nor I_85(n61_9,N6147_2_r_11,N1508_10_r_11);
endmodule


