module test_final(IN_1_0_l_1,IN_2_0_l_1,IN_3_0_l_1,IN_4_0_l_1,IN_1_1_l_1,IN_2_1_l_1,IN_3_1_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_3_3_l_1,IN_1_6_l_1,IN_2_6_l_1,IN_3_6_l_1,IN_4_6_l_1,IN_5_6_l_1,blif_clk_net_5_r_0,blif_reset_net_5_r_0,N1371_0_r_0,N1508_0_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_547_5_r_0,G42_7_r_0,n_572_7_r_0,n_573_7_r_0,n_549_7_r_0,n_569_7_r_0);
input IN_1_0_l_1,IN_2_0_l_1,IN_3_0_l_1,IN_4_0_l_1,IN_1_1_l_1,IN_2_1_l_1,IN_3_1_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_3_3_l_1,IN_1_6_l_1,IN_2_6_l_1,IN_3_6_l_1,IN_4_6_l_1,IN_5_6_l_1,blif_clk_net_5_r_0,blif_reset_net_5_r_0;
output N1371_0_r_0,N1508_0_r_0,n_429_or_0_5_r_0,G78_5_r_0,n_576_5_r_0,n_547_5_r_0,G42_7_r_0,n_572_7_r_0,n_573_7_r_0,n_549_7_r_0,n_569_7_r_0;
wire N1371_0_r_1,N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,n_452_7_r_1,N6147_9_r_1,N6134_9_r_1,I_BUFF_1_9_r_1,n4_7_r_1,n29_1,n30_1,n31_1,n32_1,n33_1,n34_1,n35_1,n36_1,n37_1,n38_1,n39_1,n40_1,n41_1,n42_1,n43_1,n44_1,n45_1,n46_1,n47_1,n48_1,n49_1,n50_1,n51_1,n52_1,n53_1,n54_1,n55_1,n_102_5_r_0,n_452_7_r_0,n_431_5_r_0,n6_0,n4_7_r_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0,n37_0,n38_0,n39_0,n40_0,n41_0,n42_0,n43_0,n44_0,n45_0;
and I_0(N1371_0_r_1,I_BUFF_1_9_r_1,n55_1);
nor I_1(N1508_0_r_1,n40_1,n44_1);
nor I_2(N1507_6_r_1,n43_1,n49_1);
nor I_3(N1508_6_r_1,n41_1,n42_1);
DFFARX1 I_4(n4_7_r_1,blif_clk_net_5_r_0,n6_0,G42_7_r_1,);
nor I_5(n_572_7_r_1,n29_1,n30_1);
not I_6(n_573_7_r_1,n_452_7_r_1);
nor I_7(n_549_7_r_1,N1371_0_r_1,n31_1);
or I_8(n_569_7_r_1,n30_1,n31_1);
nor I_9(n_452_7_r_1,n30_1,n32_1);
nor I_10(N6147_9_r_1,n35_1,n36_1);
nand I_11(N6134_9_r_1,n38_1,n39_1);
not I_12(I_BUFF_1_9_r_1,n40_1);
nor I_13(n4_7_r_1,I_BUFF_1_9_r_1,n30_1);
nor I_14(n29_1,IN_2_0_l_1,n34_1);
nor I_15(n30_1,n33_1,n34_1);
nor I_16(n31_1,IN_1_3_l_1,n54_1);
not I_17(n32_1,n48_1);
nor I_18(n33_1,IN_3_0_l_1,IN_4_0_l_1);
not I_19(n34_1,IN_1_0_l_1);
nor I_20(n35_1,I_BUFF_1_9_r_1,n37_1);
not I_21(n36_1,n29_1);
not I_22(n37_1,n41_1);
nand I_23(n38_1,IN_3_1_l_1,I_BUFF_1_9_r_1);
nand I_24(n39_1,n37_1,n40_1);
nand I_25(n40_1,IN_1_1_l_1,IN_2_1_l_1);
nand I_26(n41_1,IN_5_6_l_1,n52_1);
or I_27(n42_1,n36_1,n43_1);
nor I_28(n43_1,n32_1,n49_1);
nand I_29(n44_1,n45_1,n46_1);
nand I_30(n45_1,n47_1,n48_1);
not I_31(n46_1,IN_3_1_l_1);
not I_32(n47_1,n31_1);
nand I_33(n48_1,IN_2_6_l_1,n50_1);
nor I_34(n49_1,n41_1,n47_1);
and I_35(n50_1,IN_1_6_l_1,n51_1);
nand I_36(n51_1,n52_1,n53_1);
nand I_37(n52_1,IN_3_6_l_1,IN_4_6_l_1);
not I_38(n53_1,IN_5_6_l_1);
or I_39(n54_1,IN_2_3_l_1,IN_3_3_l_1);
nor I_40(n55_1,IN_3_1_l_1,n29_1);
nor I_41(N1371_0_r_0,n_102_5_r_0,n29_0);
nor I_42(N1508_0_r_0,n_102_5_r_0,n_452_7_r_0);
or I_43(n_429_or_0_5_r_0,n38_0,N1508_6_r_1);
DFFARX1 I_44(n_431_5_r_0,blif_clk_net_5_r_0,n6_0,G78_5_r_0,);
nand I_45(n_576_5_r_0,n26_0,N1508_6_r_1);
not I_46(n_102_5_r_0,n27_0);
nand I_47(n_547_5_r_0,n30_0,n34_0);
DFFARX1 I_48(n4_7_r_0,blif_clk_net_5_r_0,n6_0,G42_7_r_0,);
nor I_49(n_572_7_r_0,n31_0,N1508_6_r_1);
or I_50(n_573_7_r_0,n29_0,n30_0);
nor I_51(n_549_7_r_0,n29_0,n33_0);
nand I_52(n_569_7_r_0,n28_0,n32_0);
nor I_53(n_452_7_r_0,n30_0,n31_0);
nand I_54(n_431_5_r_0,n_102_5_r_0,n35_0);
not I_55(n6_0,blif_reset_net_5_r_0);
nor I_56(n4_7_r_0,n31_0,n37_0);
nor I_57(n26_0,n27_0,n28_0);
nor I_58(n27_0,n28_0,n44_0);
nand I_59(n28_0,G42_7_r_1,n_573_7_r_1);
not I_60(n29_0,n32_0);
nor I_61(n30_0,n39_0,G42_7_r_1);
not I_62(n31_0,n38_0);
nand I_63(n32_0,n41_0,n42_0);
nor I_64(n33_0,n_102_5_r_0,N1508_6_r_1);
nor I_65(n34_0,n27_0,N1508_6_r_1);
nand I_66(n35_0,n29_0,n36_0);
nor I_67(n36_0,n37_0,n38_0);
not I_68(n37_0,n28_0);
nand I_69(n38_0,n40_0,N1507_6_r_1);
nor I_70(n39_0,N1508_0_r_1,n_549_7_r_1);
or I_71(n40_0,N1508_0_r_1,n_549_7_r_1);
nor I_72(n41_0,N6134_9_r_1,N1508_0_r_1);
or I_73(n42_0,n43_0,N6147_9_r_1);
nor I_74(n43_0,n_572_7_r_1,N1508_6_r_1);
nor I_75(n44_0,n45_0,n_572_7_r_1);
and I_76(n45_0,n_569_7_r_1,N1507_6_r_1);
endmodule


