module test_I3028(I1415,I1391,I1263,I1477,I1470,I2912,I1407,I3028);
input I1415,I1391,I1263,I1477,I1470,I2912,I1407;
output I3028;
wire I3011,I2759,I2946,I2929,I2963,I2980,I2776;
not I_0(I3011,I2980);
not I_1(I2759,I1477);
or I_2(I2946,I2929,I1263);
and I_3(I2929,I2912,I1391);
nor I_4(I3028,I2963,I3011);
DFFARX1 I_5(I2946,I1470,I2759,,,I2963,);
nand I_6(I2980,I2776,I1415);
not I_7(I2776,I1407);
endmodule


