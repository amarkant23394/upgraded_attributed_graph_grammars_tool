module test_final(IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_4_l_4,IN_2_4_l_4,IN_3_4_l_4,IN_4_4_l_4,IN_5_4_l_4,IN_1_9_l_4,IN_2_9_l_4,IN_3_9_l_4,IN_4_9_l_4,IN_5_9_l_4,blif_clk_net_7_r_14,blif_reset_net_7_r_14,N1371_0_r_14,N1508_0_r_14,N1507_6_r_14,N1508_6_r_14,G42_7_r_14,n_572_7_r_14,n_573_7_r_14,n_549_7_r_14,n_569_7_r_14,n_452_7_r_14,N6147_9_r_14,N6134_9_r_14);
input IN_1_2_l_4,IN_2_2_l_4,IN_3_2_l_4,IN_4_2_l_4,IN_5_2_l_4,IN_1_4_l_4,IN_2_4_l_4,IN_3_4_l_4,IN_4_4_l_4,IN_5_4_l_4,IN_1_9_l_4,IN_2_9_l_4,IN_3_9_l_4,IN_4_9_l_4,IN_5_9_l_4,blif_clk_net_7_r_14,blif_reset_net_7_r_14;
output N1371_0_r_14,N1508_0_r_14,N1507_6_r_14,N1508_6_r_14,G42_7_r_14,n_572_7_r_14,n_573_7_r_14,n_549_7_r_14,n_569_7_r_14,n_452_7_r_14,N6147_9_r_14,N6134_9_r_14;
wire N1371_0_r_4,N1508_0_r_4,N1507_6_r_4,N1508_6_r_4,G42_7_r_4,n_572_7_r_4,n_573_7_r_4,n_549_7_r_4,n_569_7_r_4,n_452_7_r_4,N6147_9_r_4,N6134_9_r_4,I_BUFF_1_9_r_4,n4_7_r_4,n21_4,n22_4,n23_4,n24_4,n25_4,n26_4,n27_4,n28_4,n29_4,n30_4,n31_4,n32_4,n33_4,n34_4,n35_4,n36_4,n37_4,n38_4,n39_4,n40_4,n41_4,I_BUFF_1_9_r_14,N3_8_l_14,n8_14,n47_14,n4_7_r_14,n26_14,n27_14,n28_14,n29_14,n30_14,n31_14,n32_14,n33_14,n34_14,n35_14,n36_14,n37_14,n38_14,n39_14,n40_14,n41_14,n42_14,n43_14,n44_14,n45_14,n46_14;
nor I_0(N1371_0_r_4,IN_1_9_l_4,n25_4);
not I_1(N1508_0_r_4,n25_4);
nor I_2(N1507_6_r_4,n32_4,n33_4);
nor I_3(N1508_6_r_4,n22_4,n29_4);
DFFARX1 I_4(n4_7_r_4,blif_clk_net_7_r_14,n8_14,G42_7_r_4,);
not I_5(n_572_7_r_4,n_573_7_r_4);
nand I_6(n_573_7_r_4,n21_4,n22_4);
nor I_7(n_549_7_r_4,IN_1_9_l_4,n24_4);
nand I_8(n_569_7_r_4,n22_4,n23_4);
nor I_9(n_452_7_r_4,N6147_9_r_4,I_BUFF_1_9_r_4);
not I_10(N6147_9_r_4,n28_4);
nor I_11(N6134_9_r_4,N1508_0_r_4,n28_4);
not I_12(I_BUFF_1_9_r_4,n21_4);
nor I_13(n4_7_r_4,IN_1_9_l_4,N6147_9_r_4);
nand I_14(n21_4,n39_4,n40_4);
or I_15(n22_4,IN_5_9_l_4,n31_4);
not I_16(n23_4,IN_1_9_l_4);
nor I_17(n24_4,n25_4,n26_4);
nand I_18(n25_4,IN_1_4_l_4,IN_2_4_l_4);
nand I_19(n26_4,n21_4,n27_4);
nand I_20(n27_4,n36_4,n37_4);
nand I_21(n28_4,IN_2_9_l_4,n38_4);
nand I_22(n29_4,N1508_0_r_4,n30_4);
nand I_23(n30_4,n34_4,n35_4);
nor I_24(n31_4,IN_3_9_l_4,IN_4_9_l_4);
not I_25(n32_4,n30_4);
nor I_26(n33_4,n21_4,n28_4);
nand I_27(n34_4,N6147_9_r_4,I_BUFF_1_9_r_4);
nand I_28(n35_4,N1508_0_r_4,n27_4);
not I_29(n36_4,IN_5_4_l_4);
nand I_30(n37_4,IN_3_4_l_4,IN_4_4_l_4);
or I_31(n38_4,IN_3_9_l_4,IN_4_9_l_4);
nor I_32(n39_4,IN_1_2_l_4,IN_2_2_l_4);
or I_33(n40_4,IN_5_2_l_4,n41_4);
nor I_34(n41_4,IN_3_2_l_4,IN_4_2_l_4);
nor I_35(N1371_0_r_14,n47_14,n30_14);
nor I_36(N1508_0_r_14,n30_14,n41_14);
nor I_37(N1507_6_r_14,n37_14,n44_14);
nor I_38(N1508_6_r_14,n30_14,n39_14);
DFFARX1 I_39(n4_7_r_14,blif_clk_net_7_r_14,n8_14,G42_7_r_14,);
nor I_40(n_572_7_r_14,n28_14,n29_14);
nand I_41(n_573_7_r_14,n26_14,n27_14);
nor I_42(n_549_7_r_14,n31_14,n32_14);
nand I_43(n_569_7_r_14,n26_14,n30_14);
nor I_44(n_452_7_r_14,n47_14,n28_14);
nor I_45(N6147_9_r_14,n36_14,n37_14);
nor I_46(N6134_9_r_14,n28_14,n36_14);
not I_47(I_BUFF_1_9_r_14,n26_14);
and I_48(N3_8_l_14,n38_14,G42_7_r_4);
not I_49(n8_14,blif_reset_net_7_r_14);
DFFARX1 I_50(N3_8_l_14,blif_clk_net_7_r_14,n8_14,n47_14,);
nor I_51(n4_7_r_14,n47_14,n35_14);
nand I_52(n26_14,N1507_6_r_4,G42_7_r_4);
not I_53(n27_14,n28_14);
nor I_54(n28_14,n43_14,n_452_7_r_4);
not I_55(n29_14,n33_14);
not I_56(n30_14,n31_14);
nor I_57(n31_14,n46_14,n_572_7_r_4);
and I_58(n32_14,n33_14,n34_14);
nand I_59(n33_14,I_BUFF_1_9_r_14,n45_14);
nor I_60(n34_14,n42_14,n43_14);
nor I_61(n35_14,n_572_7_r_4,n_569_7_r_4);
nor I_62(n36_14,n47_14,n34_14);
not I_63(n37_14,n35_14);
nand I_64(n38_14,n_572_7_r_4,N1371_0_r_4);
nand I_65(n39_14,n29_14,n40_14);
nand I_66(n40_14,n27_14,n37_14);
nor I_67(n41_14,I_BUFF_1_9_r_14,n34_14);
nor I_68(n42_14,N1371_0_r_4,N1507_6_r_4);
not I_69(n43_14,N1508_6_r_4);
nor I_70(n44_14,n27_14,n33_14);
or I_71(n45_14,N1508_6_r_4,n_549_7_r_4);
or I_72(n46_14,n_549_7_r_4,N6134_9_r_4);
endmodule


