module test_I15502(I12930,I1477,I1470,I10636,I15502);
input I12930,I1477,I1470,I10636;
output I15502;
wire I12619,I13023,I12605,I12947,I14965,I12848,I15485;
not I_0(I12619,I1477);
DFFARX1 I_1(I10636,I1470,I12619,,,I13023,);
nand I_2(I12605,I13023,I12947);
nor I_3(I12947,I12930,I12848);
not I_4(I14965,I1477);
DFFARX1 I_5(I1470,I12619,,,I12848,);
DFFARX1 I_6(I12605,I1470,I14965,,,I15485,);
not I_7(I15502,I15485);
endmodule


