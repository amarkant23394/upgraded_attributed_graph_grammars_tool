module test_I2198(I1343,I1231,I2198);
input I1343,I1231;
output I2198;
wire ;
nand I_0(I2198,I1343,I1231);
endmodule


