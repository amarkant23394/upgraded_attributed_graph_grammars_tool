module test_final(IN_1_0_l_7,IN_2_0_l_7,IN_4_0_l_7,G18_4_l_7,G15_4_l_7,IN_1_4_l_7,IN_4_4_l_7,IN_5_4_l_7,IN_7_4_l_7,IN_9_4_l_7,IN_10_4_l_7,blif_clk_net_3_r_0,blif_reset_net_3_r_0,n_429_or_0_3_r_0,G78_3_r_0,n_576_3_r_0,n_102_3_r_0,n_547_3_r_0,G42_4_r_0,n_572_4_r_0,n_573_4_r_0,n_549_4_r_0,n_569_4_r_0,n_452_4_r_0);
input IN_1_0_l_7,IN_2_0_l_7,IN_4_0_l_7,G18_4_l_7,G15_4_l_7,IN_1_4_l_7,IN_4_4_l_7,IN_5_4_l_7,IN_7_4_l_7,IN_9_4_l_7,IN_10_4_l_7,blif_clk_net_3_r_0,blif_reset_net_3_r_0;
output n_429_or_0_3_r_0,G78_3_r_0,n_576_3_r_0,n_102_3_r_0,n_547_3_r_0,G42_4_r_0,n_572_4_r_0,n_573_4_r_0,n_549_4_r_0,n_569_4_r_0,n_452_4_r_0;
wire ACVQN2_0_r_7,n_266_and_0_0_r_7,G199_1_r_7,G214_1_r_7,n_429_or_0_3_r_7,G78_3_r_7,n_576_3_r_7,n_102_3_r_7,n_547_3_r_7,n_42_5_r_7,G199_5_r_7,ACVQN2_0_l_7,n_266_and_0_0_l_7,ACVQN1_0_l_7,n4_4_l_7,G42_4_l_7,n_87_4_l_7,n_572_4_l_7,n_573_4_l_7,n_549_4_l_7,n7_4_l_7,n_569_4_l_7,n_452_4_l_7,ACVQN1_0_r_7,N1_1_r_7,n3_1_r_7,n12_3_r_7,n_431_3_r_7,n11_3_r_7,n13_3_r_7,n14_3_r_7,n15_3_r_7,n16_3_r_7,N3_5_r_7,n3_5_r_7,n2_3_r_0,ACVQN2_0_l_0,n_266_and_0_0_l_0,ACVQN1_0_l_0,N1_1_l_0,G199_1_l_0,G214_1_l_0,n3_1_l_0,n_42_5_l_0,N3_5_l_0,G199_5_l_0,n3_5_l_0,n12_3_r_0,n_431_3_r_0,n11_3_r_0,n13_3_r_0,n14_3_r_0,n15_3_r_0,n16_3_r_0,n4_4_r_0,n_87_4_r_0,n7_4_r_0;
DFFARX1 I_0(n_572_4_l_7,blif_clk_net_3_r_0,n2_3_r_0,ACVQN2_0_r_7,);
and I_1(n_266_and_0_0_r_7,n_452_4_l_7,ACVQN1_0_r_7);
DFFARX1 I_2(N1_1_r_7,blif_clk_net_3_r_0,n2_3_r_0,G199_1_r_7,);
DFFARX1 I_3(G42_4_l_7,blif_clk_net_3_r_0,n2_3_r_0,G214_1_r_7,);
nand I_4(n_429_or_0_3_r_7,n_266_and_0_0_l_7,n12_3_r_7);
DFFARX1 I_5(n_431_3_r_7,blif_clk_net_3_r_0,n2_3_r_0,G78_3_r_7,);
nand I_6(n_576_3_r_7,ACVQN2_0_l_7,n11_3_r_7);
not I_7(n_102_3_r_7,n_266_and_0_0_l_7);
nand I_8(n_547_3_r_7,n_573_4_l_7,n13_3_r_7);
nor I_9(n_42_5_r_7,n_266_and_0_0_l_7,n_549_4_l_7);
DFFARX1 I_10(N3_5_r_7,blif_clk_net_3_r_0,n2_3_r_0,G199_5_r_7,);
DFFARX1 I_11(IN_1_0_l_7,blif_clk_net_3_r_0,n2_3_r_0,ACVQN2_0_l_7,);
and I_12(n_266_and_0_0_l_7,IN_4_0_l_7,ACVQN1_0_l_7);
DFFARX1 I_13(IN_2_0_l_7,blif_clk_net_3_r_0,n2_3_r_0,ACVQN1_0_l_7,);
nor I_14(n4_4_l_7,G18_4_l_7,IN_1_4_l_7);
DFFARX1 I_15(n4_4_l_7,blif_clk_net_3_r_0,n2_3_r_0,G42_4_l_7,);
not I_16(n_87_4_l_7,G15_4_l_7);
nor I_17(n_572_4_l_7,G15_4_l_7,IN_7_4_l_7);
or I_18(n_573_4_l_7,IN_5_4_l_7,IN_9_4_l_7);
nor I_19(n_549_4_l_7,IN_10_4_l_7,n7_4_l_7);
and I_20(n7_4_l_7,IN_4_4_l_7,n_87_4_l_7);
or I_21(n_569_4_l_7,IN_9_4_l_7,IN_10_4_l_7);
nor I_22(n_452_4_l_7,G18_4_l_7,IN_5_4_l_7);
DFFARX1 I_23(n_572_4_l_7,blif_clk_net_3_r_0,n2_3_r_0,ACVQN1_0_r_7,);
and I_24(N1_1_r_7,n_572_4_l_7,n3_1_r_7);
nand I_25(n3_1_r_7,ACVQN2_0_l_7,n_549_4_l_7);
not I_26(n12_3_r_7,G42_4_l_7);
or I_27(n_431_3_r_7,n_569_4_l_7,n14_3_r_7);
nor I_28(n11_3_r_7,n_266_and_0_0_l_7,n12_3_r_7);
nor I_29(n13_3_r_7,n_266_and_0_0_l_7,n_452_4_l_7);
and I_30(n14_3_r_7,ACVQN2_0_l_7,n15_3_r_7);
nor I_31(n15_3_r_7,n_569_4_l_7,n16_3_r_7);
not I_32(n16_3_r_7,n_266_and_0_0_l_7);
and I_33(N3_5_r_7,G42_4_l_7,n3_5_r_7);
nand I_34(n3_5_r_7,n_266_and_0_0_l_7,n_573_4_l_7);
nand I_35(n_429_or_0_3_r_0,ACVQN2_0_l_0,n12_3_r_0);
DFFARX1 I_36(n_431_3_r_0,blif_clk_net_3_r_0,n2_3_r_0,G78_3_r_0,);
nand I_37(n_576_3_r_0,n_266_and_0_0_l_0,n11_3_r_0);
not I_38(n_102_3_r_0,n_42_5_l_0);
nand I_39(n_547_3_r_0,ACVQN2_0_l_0,n13_3_r_0);
DFFARX1 I_40(n4_4_r_0,blif_clk_net_3_r_0,n2_3_r_0,G42_4_r_0,);
nor I_41(n_572_4_r_0,G199_1_l_0,G199_5_l_0);
or I_42(n_573_4_r_0,n_42_5_l_0,G199_5_l_0);
nor I_43(n_549_4_r_0,n_266_and_0_0_l_0,n7_4_r_0);
or I_44(n_569_4_r_0,n_266_and_0_0_l_0,n_42_5_l_0);
nor I_45(n_452_4_r_0,ACVQN2_0_l_0,G199_5_l_0);
not I_46(n2_3_r_0,blif_reset_net_3_r_0);
DFFARX1 I_47(n_429_or_0_3_r_7,blif_clk_net_3_r_0,n2_3_r_0,ACVQN2_0_l_0,);
and I_48(n_266_and_0_0_l_0,ACVQN1_0_l_0,ACVQN2_0_r_7);
DFFARX1 I_49(G199_5_r_7,blif_clk_net_3_r_0,n2_3_r_0,ACVQN1_0_l_0,);
and I_50(N1_1_l_0,n3_1_l_0,G199_1_r_7);
DFFARX1 I_51(N1_1_l_0,blif_clk_net_3_r_0,n2_3_r_0,G199_1_l_0,);
DFFARX1 I_52(n_266_and_0_0_r_7,blif_clk_net_3_r_0,n2_3_r_0,G214_1_l_0,);
nand I_53(n3_1_l_0,G214_1_r_7,n_576_3_r_7);
nor I_54(n_42_5_l_0,G78_3_r_7,n_547_3_r_7);
and I_55(N3_5_l_0,n3_5_l_0,n_42_5_r_7);
DFFARX1 I_56(N3_5_l_0,blif_clk_net_3_r_0,n2_3_r_0,G199_5_l_0,);
nand I_57(n3_5_l_0,G78_3_r_7,n_102_3_r_7);
not I_58(n12_3_r_0,G199_1_l_0);
or I_59(n_431_3_r_0,n_266_and_0_0_l_0,n14_3_r_0);
nor I_60(n11_3_r_0,G214_1_l_0,n12_3_r_0);
nor I_61(n13_3_r_0,G214_1_l_0,n_42_5_l_0);
and I_62(n14_3_r_0,n_42_5_l_0,n15_3_r_0);
nor I_63(n15_3_r_0,G199_1_l_0,n16_3_r_0);
not I_64(n16_3_r_0,ACVQN2_0_l_0);
nor I_65(n4_4_r_0,ACVQN2_0_l_0,G214_1_l_0);
not I_66(n_87_4_r_0,G199_5_l_0);
and I_67(n7_4_r_0,ACVQN2_0_l_0,n_87_4_r_0);
endmodule


