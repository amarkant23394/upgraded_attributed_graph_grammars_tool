module test_I17109(I14982,I1477,I1470,I12599,I17109);
input I14982,I1477,I1470,I12599;
output I17109;
wire I14933,I12587,I15047,I15064,I15276,I15293,I14954,I17092,I16818,I15310,I15211,I14965;
DFFARX1 I_0(I15310,I1470,I14965,,,I14933,);
DFFARX1 I_1(I1470,,,I12587,);
nor I_2(I15047,I14982);
nand I_3(I15064,I15047,I12587);
nand I_4(I15276,I14982,I12599);
nand I_5(I15293,I15276,I15211);
not I_6(I14954,I15064);
DFFARX1 I_7(I14954,I1470,I16818,,,I17092,);
not I_8(I16818,I1477);
and I_9(I15310,I15276,I15293);
DFFARX1 I_10(I1470,I14965,,,I15211,);
not I_11(I14965,I1477);
and I_12(I17109,I17092,I14933);
endmodule


