module test_I7348(I1477,I5249,I5204,I5139,I1470,I7348);
input I1477,I5249,I5204,I5139,I1470;
output I7348;
wire I5266,I6941,I5385,I5067,I6907,I5481,I5156,I5091,I7269,I5094,I6958,I3371,I5625,I5070,I5105,I5642,I5351;
not I_0(I5266,I5249);
nor I_1(I6941,I5070,I5094);
nor I_2(I5385,I5351,I5266);
DFFARX1 I_3(I5642,I1470,I5105,,,I5067,);
not I_4(I6907,I1477);
DFFARX1 I_5(I1470,I5105,,,I5481,);
nand I_6(I5156,I5139,I3371);
nand I_7(I5091,I5156,I5385);
DFFARX1 I_8(I5067,I1470,I6907,,,I7269,);
not I_9(I5094,I5204);
nand I_10(I6958,I6941,I5091);
DFFARX1 I_11(I1470,,,I3371,);
DFFARX1 I_12(I1470,I5105,,,I5625,);
and I_13(I5070,I5249,I5481);
not I_14(I5105,I1477);
not I_15(I5642,I5625);
DFFARX1 I_16(I1470,I5105,,,I5351,);
nand I_17(I7348,I7269,I6958);
endmodule


