module test_final(IN_1_2_l,IN_2_2_l,G1_3_l,G2_3_l,IN_2_3_l,IN_4_3_l,IN_5_3_l,IN_7_3_l,IN_8_3_l,IN_10_3_l,IN_11_3_l,blif_reset_net_0_r,blif_clk_net_0_r,ACVQN2_0_r,n_266_and_0_0_r,G199_1_r,G214_1_r,ACVQN1_2_r,P6_2_r,n_429_or_0_3_r,G78_3_r,n_576_3_r,n_102_3_r,n_547_3_r);
input IN_1_2_l,IN_2_2_l,G1_3_l,G2_3_l,IN_2_3_l,IN_4_3_l,IN_5_3_l,IN_7_3_l,IN_8_3_l,IN_10_3_l,IN_11_3_l,blif_reset_net_0_r,blif_clk_net_0_r;
output ACVQN2_0_r,n_266_and_0_0_r,G199_1_r,G214_1_r,ACVQN1_2_r,P6_2_r,n_429_or_0_3_r,G78_3_r,n_576_3_r,n_102_3_r,n_547_3_r;
wire ACVQN1_2_l,P6_2_l,P6_internal_2_l,n_429_or_0_3_l,G78_3_l,n_576_3_l,n_102_3_l,n_547_3_l,n_431_3_l,n11_3_l,n12_3_l,n13_3_l,n14_3_l,n15_3_l,n16_3_l,n1_0_r,ACVQN1_0_r,N1_1_r,n3_1_r,P6_internal_2_r,n_431_3_r,n11_3_r,n12_3_r,n13_3_r,n14_3_r,n15_3_r,n16_3_r;
DFFARX1 I_0(IN_2_2_l,blif_clk_net_0_r,n1_0_r,ACVQN1_2_l,);
not I_1(P6_2_l,P6_internal_2_l);
DFFARX1 I_2(IN_1_2_l,blif_clk_net_0_r,n1_0_r,P6_internal_2_l,);
nand I_3(n_429_or_0_3_l,G1_3_l,n12_3_l);
DFFARX1 I_4(n_431_3_l,blif_clk_net_0_r,n1_0_r,G78_3_l,);
nand I_5(n_576_3_l,IN_7_3_l,n11_3_l);
not I_6(n_102_3_l,G2_3_l);
nand I_7(n_547_3_l,IN_11_3_l,n13_3_l);
or I_8(n_431_3_l,IN_8_3_l,n14_3_l);
nor I_9(n11_3_l,G2_3_l,n12_3_l);
not I_10(n12_3_l,IN_5_3_l);
nor I_11(n13_3_l,G2_3_l,IN_10_3_l);
and I_12(n14_3_l,IN_2_3_l,n15_3_l);
nor I_13(n15_3_l,IN_4_3_l,n16_3_l);
not I_14(n16_3_l,G1_3_l);
DFFARX1 I_15(P6_2_l,blif_clk_net_0_r,n1_0_r,ACVQN2_0_r,);
and I_16(n_266_and_0_0_r,ACVQN1_0_r,n_102_3_l);
not I_17(n1_0_r,blif_reset_net_0_r);
DFFARX1 I_18(n_429_or_0_3_l,blif_clk_net_0_r,n1_0_r,ACVQN1_0_r,);
DFFARX1 I_19(N1_1_r,blif_clk_net_0_r,n1_0_r,G199_1_r,);
DFFARX1 I_20(n_576_3_l,blif_clk_net_0_r,n1_0_r,G214_1_r,);
and I_21(N1_1_r,n3_1_r,n_429_or_0_3_l);
nand I_22(n3_1_r,G78_3_l,n_429_or_0_3_l);
DFFARX1 I_23(n_547_3_l,blif_clk_net_0_r,n1_0_r,ACVQN1_2_r,);
not I_24(P6_2_r,P6_internal_2_r);
DFFARX1 I_25(ACVQN1_2_l,blif_clk_net_0_r,n1_0_r,P6_internal_2_r,);
nand I_26(n_429_or_0_3_r,n12_3_r,ACVQN1_2_l);
DFFARX1 I_27(n_431_3_r,blif_clk_net_0_r,n1_0_r,G78_3_r,);
nand I_28(n_576_3_r,n11_3_r,n_547_3_l);
not I_29(n_102_3_r,n_576_3_l);
nand I_30(n_547_3_r,n13_3_r,P6_2_l);
or I_31(n_431_3_r,n14_3_r,P6_2_l);
nor I_32(n11_3_r,n12_3_r,G78_3_l);
not I_33(n12_3_r,n_102_3_l);
nor I_34(n13_3_r,G78_3_l,n_576_3_l);
and I_35(n14_3_r,n15_3_r,ACVQN1_2_l);
nor I_36(n15_3_r,n16_3_r,n_576_3_l);
not I_37(n16_3_r,ACVQN1_2_l);
endmodule


