module test_final(IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_4_2_l_10,IN_5_2_l_10,IN_1_6_l_10,IN_2_6_l_10,IN_3_6_l_10,IN_4_6_l_10,IN_5_6_l_10,IN_1_9_l_10,IN_2_9_l_10,IN_3_9_l_10,IN_4_9_l_10,IN_5_9_l_10,blif_clk_net_8_r_8,blif_reset_net_8_r_8,N1371_0_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,N1508_10_r_8);
input IN_1_2_l_10,IN_2_2_l_10,IN_3_2_l_10,IN_4_2_l_10,IN_5_2_l_10,IN_1_6_l_10,IN_2_6_l_10,IN_3_6_l_10,IN_4_6_l_10,IN_5_6_l_10,IN_1_9_l_10,IN_2_9_l_10,IN_3_9_l_10,IN_4_9_l_10,IN_5_9_l_10,blif_clk_net_8_r_8,blif_reset_net_8_r_8;
output N1371_0_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,N1508_10_r_8;
wire N1371_0_r_10,N1508_0_r_10,N6147_2_r_10,N6147_3_r_10,N1372_4_r_10,N1508_4_r_10,N1507_6_r_10,N1508_6_r_10,n_42_8_r_10,G199_8_r_10,N6147_9_r_10,N6134_9_r_10,I_BUFF_1_9_r_10,N3_8_r_10,n35_10,n36_10,n37_10,n38_10,n39_10,n40_10,n41_10,n42_10,n43_10,n44_10,n45_10,n46_10,n47_10,n48_10,n49_10,n50_10,n51_10,n52_10,n53_10,n54_10,n55_10,n56_10,n57_10,n58_10,n59_10,n60_10,n61_10,n62_10,n63_10,n64_10,N1508_0_r_8,N1372_1_r_8,I_BUFF_1_9_r_8,N1372_10_r_8,N3_8_l_8,n8_8,n53_8,n29_8,N3_8_r_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8,n38_8,n39_8,n40_8,n41_8,n42_8,n43_8,n44_8,n45_8,n46_8,n47_8,n48_8,n49_8,n50_8,n51_8,n52_8;
nor I_0(N1371_0_r_10,n37_10,n38_10);
nor I_1(N1508_0_r_10,n37_10,n58_10);
nand I_2(N6147_2_r_10,n39_10,n40_10);
not I_3(N6147_3_r_10,n39_10);
nor I_4(N1372_4_r_10,n46_10,n49_10);
nor I_5(N1508_4_r_10,n51_10,n52_10);
nor I_6(N1507_6_r_10,n49_10,n60_10);
nor I_7(N1508_6_r_10,n49_10,n50_10);
nor I_8(n_42_8_r_10,I_BUFF_1_9_r_10,n35_10);
DFFARX1 I_9(N3_8_r_10,blif_clk_net_8_r_8,n8_8,G199_8_r_10,);
nor I_10(N6147_9_r_10,n36_10,n37_10);
nor I_11(N6134_9_r_10,I_BUFF_1_9_r_10,n46_10);
not I_12(I_BUFF_1_9_r_10,n48_10);
nor I_13(N3_8_r_10,n44_10,n47_10);
not I_14(n35_10,n49_10);
nor I_15(n36_10,I_BUFF_1_9_r_10,n38_10);
not I_16(n37_10,IN_1_9_l_10);
not I_17(n38_10,n46_10);
nand I_18(n39_10,n43_10,n44_10);
nand I_19(n40_10,I_BUFF_1_9_r_10,n41_10);
nor I_20(n41_10,IN_1_9_l_10,n42_10);
not I_21(n42_10,n44_10);
nor I_22(n43_10,IN_1_9_l_10,n45_10);
nand I_23(n44_10,IN_2_6_l_10,n54_10);
nor I_24(n45_10,IN_5_9_l_10,n59_10);
nand I_25(n46_10,IN_2_9_l_10,n61_10);
nor I_26(n47_10,n46_10,n48_10);
nand I_27(n48_10,n62_10,n63_10);
nand I_28(n49_10,IN_5_6_l_10,n56_10);
not I_29(n50_10,n45_10);
nor I_30(n51_10,n42_10,n53_10);
not I_31(n52_10,N1372_4_r_10);
nor I_32(n53_10,n48_10,n50_10);
and I_33(n54_10,IN_1_6_l_10,n55_10);
nand I_34(n55_10,n56_10,n57_10);
nand I_35(n56_10,IN_3_6_l_10,IN_4_6_l_10);
not I_36(n57_10,IN_5_6_l_10);
nor I_37(n58_10,n35_10,n45_10);
nor I_38(n59_10,IN_3_9_l_10,IN_4_9_l_10);
nor I_39(n60_10,n37_10,n46_10);
or I_40(n61_10,IN_3_9_l_10,IN_4_9_l_10);
nor I_41(n62_10,IN_1_2_l_10,IN_2_2_l_10);
or I_42(n63_10,IN_5_2_l_10,n64_10);
nor I_43(n64_10,IN_3_2_l_10,IN_4_2_l_10);
nor I_44(N1371_0_r_8,n46_8,n51_8);
not I_45(N1508_0_r_8,n46_8);
nor I_46(N1372_1_r_8,n37_8,n49_8);
and I_47(N1508_1_r_8,N1372_1_r_8,n29_8);
nor I_48(N1507_6_r_8,n47_8,n48_8);
nor I_49(N1508_6_r_8,n37_8,n38_8);
nor I_50(n_42_8_r_8,I_BUFF_1_9_r_8,n53_8);
DFFARX1 I_51(N3_8_r_8,blif_clk_net_8_r_8,n8_8,G199_8_r_8,);
nor I_52(N6147_9_r_8,n29_8,n30_8);
nor I_53(N6134_9_r_8,n30_8,n31_8);
not I_54(I_BUFF_1_9_r_8,n35_8);
nor I_55(N1372_10_r_8,n46_8,n49_8);
nor I_56(N1508_10_r_8,n40_8,n41_8);
and I_57(N3_8_l_8,n36_8,G199_8_r_10);
not I_58(n8_8,blif_reset_net_8_r_8);
DFFARX1 I_59(N3_8_l_8,blif_clk_net_8_r_8,n8_8,n53_8,);
not I_60(n29_8,n53_8);
nor I_61(N3_8_r_8,n33_8,n34_8);
and I_62(n30_8,n32_8,n33_8);
nor I_63(n31_8,N1508_6_r_10,N6147_2_r_10);
nand I_64(n32_8,n42_8,N1371_0_r_10);
or I_65(n33_8,n46_8,N6147_3_r_10);
nor I_66(n34_8,n32_8,n35_8);
nand I_67(n35_8,n44_8,N6147_9_r_10);
nand I_68(n36_8,N1508_0_r_10,N1508_6_r_10);
not I_69(n37_8,n31_8);
nand I_70(n38_8,N1508_0_r_8,n39_8);
nand I_71(n39_8,n33_8,n50_8);
and I_72(n40_8,n32_8,n35_8);
not I_73(n41_8,N1372_10_r_8);
and I_74(n42_8,n43_8,n_42_8_r_10);
nand I_75(n43_8,n44_8,n45_8);
nand I_76(n44_8,N1507_6_r_10,N1508_0_r_10);
not I_77(n45_8,N6147_9_r_10);
nand I_78(n46_8,N1371_0_r_10,N1508_4_r_10);
not I_79(n47_8,n39_8);
nor I_80(n48_8,n35_8,n49_8);
not I_81(n49_8,n51_8);
nand I_82(n50_8,I_BUFF_1_9_r_8,n51_8);
nor I_83(n51_8,n52_8,N6134_9_r_10);
or I_84(n52_8,N6147_2_r_10,N6147_3_r_10);
endmodule


