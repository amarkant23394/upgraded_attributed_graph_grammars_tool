module test_I11167(I8202,I8181,I1477,I1470,I9525,I11167);
input I8202,I8181,I1477,I1470,I9525;
output I11167;
wire I10647,I9576,I9542,I9474,I11150,I9491;
not I_0(I10647,I1477);
nor I_1(I9576,I8181,I8202);
DFFARX1 I_2(I9525,I1470,I9491,,,I9542,);
not I_3(I11167,I11150);
or I_4(I9474,I9576,I9542);
DFFARX1 I_5(I9474,I1470,I10647,,,I11150,);
not I_6(I9491,I1477);
endmodule


