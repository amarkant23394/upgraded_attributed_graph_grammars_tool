module test_final(IN_1_2_l_1,IN_2_2_l_1,IN_3_2_l_1,IN_6_2_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_4_3_l_1,IN_1_4_l_1,IN_2_4_l_1,IN_3_4_l_1,IN_6_4_l_1,blif_clk_net_1_r_2,blif_reset_net_1_r_2,G42_1_r_2,n_572_1_r_2,n_549_1_r_2,n_569_1_r_2,n_452_1_r_2,n_42_2_r_2,G199_2_r_2,ACVQN1_5_r_2,P6_5_r_2);
input IN_1_2_l_1,IN_2_2_l_1,IN_3_2_l_1,IN_6_2_l_1,IN_1_3_l_1,IN_2_3_l_1,IN_4_3_l_1,IN_1_4_l_1,IN_2_4_l_1,IN_3_4_l_1,IN_6_4_l_1,blif_clk_net_1_r_2,blif_reset_net_1_r_2;
output G42_1_r_2,n_572_1_r_2,n_549_1_r_2,n_569_1_r_2,n_452_1_r_2,n_42_2_r_2,G199_2_r_2,ACVQN1_5_r_2,P6_5_r_2;
wire G42_1_r_1,n_572_1_r_1,n_573_1_r_1,n_549_1_r_1,n_452_1_r_1,ACVQN2_3_r_1,n_266_and_0_3_r_1,G199_4_r_1,G214_4_r_1,N3_2_l_1,n26_1,n17_1,n16_internal_1,n16_1,ACVQN1_3_l_1,N1_4_l_1,G199_4_l_1,G214_4_l_1,n4_1_r_1,n14_internal_1,n14_1,N1_4_r_1,n18_1,n19_1,n20_1,n21_1,n22_1,n23_1,n24_1,n25_1,n_573_1_r_2,N3_2_l_2,n5_2,G199_2_l_2,n13_2,ACVQN2_3_l_2,n16_2,N1_4_l_2,n26_2,n17_internal_2,n17_2,n4_1_r_2,N3_2_r_2,P6_5_r_internal_2,n18_2,n19_2,n20_2,n21_2,n22_2,n23_2,n24_2,n25_2;
DFFARX1 I_0(n4_1_r_1,blif_clk_net_1_r_2,n5_2,G42_1_r_1,);
nor I_1(n_572_1_r_1,n26_1,n19_1);
nand I_2(n_573_1_r_1,n16_1,n18_1);
nor I_3(n_549_1_r_1,n20_1,n21_1);
nor I_4(n_452_1_r_1,G214_4_l_1,n20_1);
DFFARX1 I_5(G199_4_l_1,blif_clk_net_1_r_2,n5_2,ACVQN2_3_r_1,);
nor I_6(n_266_and_0_3_r_1,n16_1,n14_1);
DFFARX1 I_7(N1_4_r_1,blif_clk_net_1_r_2,n5_2,G199_4_r_1,);
DFFARX1 I_8(G199_4_l_1,blif_clk_net_1_r_2,n5_2,G214_4_r_1,);
and I_9(N3_2_l_1,IN_6_2_l_1,n23_1);
DFFARX1 I_10(N3_2_l_1,blif_clk_net_1_r_2,n5_2,n26_1,);
not I_11(n17_1,n26_1);
DFFARX1 I_12(IN_1_3_l_1,blif_clk_net_1_r_2,n5_2,n16_internal_1,);
not I_13(n16_1,n16_internal_1);
DFFARX1 I_14(IN_2_3_l_1,blif_clk_net_1_r_2,n5_2,ACVQN1_3_l_1,);
and I_15(N1_4_l_1,IN_6_4_l_1,n25_1);
DFFARX1 I_16(N1_4_l_1,blif_clk_net_1_r_2,n5_2,G199_4_l_1,);
DFFARX1 I_17(IN_3_4_l_1,blif_clk_net_1_r_2,n5_2,G214_4_l_1,);
nor I_18(n4_1_r_1,n26_1,G214_4_l_1);
DFFARX1 I_19(G214_4_l_1,blif_clk_net_1_r_2,n5_2,n14_internal_1,);
not I_20(n14_1,n14_internal_1);
nor I_21(N1_4_r_1,n17_1,n24_1);
nand I_22(n18_1,IN_4_3_l_1,ACVQN1_3_l_1);
nor I_23(n19_1,IN_1_2_l_1,IN_3_2_l_1);
not I_24(n20_1,n18_1);
nor I_25(n21_1,n26_1,n22_1);
not I_26(n22_1,n19_1);
nand I_27(n23_1,IN_2_2_l_1,IN_3_2_l_1);
nor I_28(n24_1,n18_1,n22_1);
nand I_29(n25_1,IN_1_4_l_1,IN_2_4_l_1);
DFFARX1 I_30(n4_1_r_2,blif_clk_net_1_r_2,n5_2,G42_1_r_2,);
nor I_31(n_572_1_r_2,n26_2,n18_2);
nand I_32(n_573_1_r_2,n17_2,n19_2);
nor I_33(n_549_1_r_2,G199_2_l_2,n20_2);
nand I_34(n_569_1_r_2,n13_2,n19_2);
not I_35(n_452_1_r_2,n_573_1_r_2);
nor I_36(n_42_2_r_2,ACVQN2_3_l_2,n18_2);
DFFARX1 I_37(N3_2_r_2,blif_clk_net_1_r_2,n5_2,G199_2_r_2,);
DFFARX1 I_38(ACVQN2_3_l_2,blif_clk_net_1_r_2,n5_2,ACVQN1_5_r_2,);
not I_39(P6_5_r_2,P6_5_r_internal_2);
and I_40(N3_2_l_2,n24_2,n_572_1_r_1);
not I_41(n5_2,blif_reset_net_1_r_2);
DFFARX1 I_42(N3_2_l_2,blif_clk_net_1_r_2,n5_2,G199_2_l_2,);
not I_43(n13_2,G199_2_l_2);
DFFARX1 I_44(G42_1_r_1,blif_clk_net_1_r_2,n5_2,ACVQN2_3_l_2,);
DFFARX1 I_45(n_573_1_r_1,blif_clk_net_1_r_2,n5_2,n16_2,);
and I_46(N1_4_l_2,n25_2,n_452_1_r_1);
DFFARX1 I_47(N1_4_l_2,blif_clk_net_1_r_2,n5_2,n26_2,);
DFFARX1 I_48(n_572_1_r_1,blif_clk_net_1_r_2,n5_2,n17_internal_2,);
not I_49(n17_2,n17_internal_2);
nor I_50(n4_1_r_2,n26_2,n22_2);
nor I_51(N3_2_r_2,n17_2,n23_2);
DFFARX1 I_52(G199_2_l_2,blif_clk_net_1_r_2,n5_2,P6_5_r_internal_2,);
nor I_53(n18_2,n_549_1_r_1,ACVQN2_3_r_1);
nand I_54(n19_2,n16_2,n_266_and_0_3_r_1);
nor I_55(n20_2,n26_2,n21_2);
not I_56(n21_2,n18_2);
and I_57(n22_2,n16_2,n_266_and_0_3_r_1);
nor I_58(n23_2,n13_2,n21_2);
nand I_59(n24_2,ACVQN2_3_r_1,G214_4_r_1);
nand I_60(n25_2,G199_4_r_1,G42_1_r_1);
endmodule


