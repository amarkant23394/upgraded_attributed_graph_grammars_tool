module test_I8178(I1477,I1470,I5881,I8178);
input I1477,I1470,I5881;
output I8178;
wire I8216,I8753,I5915,I5731,I8736;
not I_0(I8216,I1477);
not I_1(I8753,I8736);
DFFARX1 I_2(I8753,I1470,I8216,,,I8178,);
DFFARX1 I_3(I1470,,,I5915,);
nand I_4(I5731,I5915,I5881);
DFFARX1 I_5(I5731,I1470,I8216,,,I8736,);
endmodule


