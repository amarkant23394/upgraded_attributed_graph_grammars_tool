module test_final(IN_1_2_l_9,IN_2_2_l_9,IN_3_2_l_9,IN_6_2_l_9,IN_1_3_l_9,IN_2_3_l_9,IN_4_3_l_9,IN_1_4_l_9,IN_2_4_l_9,IN_3_4_l_9,IN_6_4_l_9,blif_clk_net_1_r_0,blif_reset_net_1_r_0,G42_1_r_0,n_572_1_r_0,n_573_1_r_0,n_549_1_r_0,n_42_2_r_0,G199_2_r_0,G199_4_r_0,G214_4_r_0);
input IN_1_2_l_9,IN_2_2_l_9,IN_3_2_l_9,IN_6_2_l_9,IN_1_3_l_9,IN_2_3_l_9,IN_4_3_l_9,IN_1_4_l_9,IN_2_4_l_9,IN_3_4_l_9,IN_6_4_l_9,blif_clk_net_1_r_0,blif_reset_net_1_r_0;
output G42_1_r_0,n_572_1_r_0,n_573_1_r_0,n_549_1_r_0,n_42_2_r_0,G199_2_r_0,G199_4_r_0,G214_4_r_0;
wire G42_1_r_9,n_572_1_r_9,n_573_1_r_9,n_549_1_r_9,n_569_1_r_9,n_452_1_r_9,n_42_2_r_9,G199_2_r_9,G199_4_r_9,G214_4_r_9,N3_2_l_9,n27_9,n16_9,n26_9,n15_9,n29_internal_9,n29_9,N1_4_l_9,n25_9,n28_internal_9,n28_9,n4_1_r_9,N3_2_r_9,N1_4_r_9,n_42_2_l_9,n17_9,n18_9,n19_9,n20_9,n21_9,n22_9,n23_9,n24_9,n_569_1_r_0,n4_1_l_0,n6_0,n37_0,n38_0,n20_0,ACVQN1_3_l_0,n4_1_r_0,N3_2_r_0,N1_4_r_0,n2_0,n21_0,n22_0,n23_0,n24_0,n25_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0;
DFFARX1 I_0(n4_1_r_9,blif_clk_net_1_r_0,n6_0,G42_1_r_9,);
nor I_1(n_572_1_r_9,n27_9,n_42_2_l_9);
or I_2(n_573_1_r_9,n25_9,n_42_2_l_9);
nand I_3(n_549_1_r_9,n17_9,n18_9);
or I_4(n_569_1_r_9,n26_9,n_42_2_l_9);
nor I_5(n_452_1_r_9,n26_9,n25_9);
nor I_6(n_42_2_r_9,n25_9,n19_9);
DFFARX1 I_7(N3_2_r_9,blif_clk_net_1_r_0,n6_0,G199_2_r_9,);
DFFARX1 I_8(N1_4_r_9,blif_clk_net_1_r_0,n6_0,G199_4_r_9,);
DFFARX1 I_9(n_42_2_l_9,blif_clk_net_1_r_0,n6_0,G214_4_r_9,);
and I_10(N3_2_l_9,IN_6_2_l_9,n22_9);
DFFARX1 I_11(N3_2_l_9,blif_clk_net_1_r_0,n6_0,n27_9,);
not I_12(n16_9,n27_9);
DFFARX1 I_13(IN_1_3_l_9,blif_clk_net_1_r_0,n6_0,n26_9,);
not I_14(n15_9,n26_9);
DFFARX1 I_15(IN_2_3_l_9,blif_clk_net_1_r_0,n6_0,n29_internal_9,);
not I_16(n29_9,n29_internal_9);
and I_17(N1_4_l_9,IN_6_4_l_9,n24_9);
DFFARX1 I_18(N1_4_l_9,blif_clk_net_1_r_0,n6_0,n25_9,);
DFFARX1 I_19(IN_3_4_l_9,blif_clk_net_1_r_0,n6_0,n28_internal_9,);
not I_20(n28_9,n28_internal_9);
nor I_21(n4_1_r_9,n27_9,n26_9);
nor I_22(N3_2_r_9,n15_9,n21_9);
nor I_23(N1_4_r_9,n16_9,n21_9);
nor I_24(n_42_2_l_9,IN_1_2_l_9,IN_3_2_l_9);
not I_25(n17_9,n_452_1_r_9);
nand I_26(n18_9,n27_9,n15_9);
nor I_27(n19_9,n29_9,n20_9);
not I_28(n20_9,IN_4_3_l_9);
and I_29(n21_9,IN_4_3_l_9,n23_9);
nand I_30(n22_9,IN_2_2_l_9,IN_3_2_l_9);
nor I_31(n23_9,n29_9,n28_9);
nand I_32(n24_9,IN_1_4_l_9,IN_2_4_l_9);
DFFARX1 I_33(n4_1_r_0,blif_clk_net_1_r_0,n6_0,G42_1_r_0,);
nor I_34(n_572_1_r_0,n23_0,n_573_1_r_9);
nand I_35(n_573_1_r_0,n21_0,n22_0);
nand I_36(n_549_1_r_0,n_569_1_r_0,n24_0);
nand I_37(n_569_1_r_0,n21_0,n26_0);
nor I_38(n_42_2_r_0,n27_0,n28_0);
DFFARX1 I_39(N3_2_r_0,blif_clk_net_1_r_0,n6_0,G199_2_r_0,);
DFFARX1 I_40(N1_4_r_0,blif_clk_net_1_r_0,n6_0,G199_4_r_0,);
DFFARX1 I_41(n2_0,blif_clk_net_1_r_0,n6_0,G214_4_r_0,);
nor I_42(n4_1_l_0,G42_1_r_9,n_549_1_r_9);
not I_43(n6_0,blif_reset_net_1_r_0);
DFFARX1 I_44(n4_1_l_0,blif_clk_net_1_r_0,n6_0,n37_0,);
DFFARX1 I_45(n_569_1_r_9,blif_clk_net_1_r_0,n6_0,n38_0,);
not I_46(n20_0,n38_0);
DFFARX1 I_47(G214_4_r_9,blif_clk_net_1_r_0,n6_0,ACVQN1_3_l_0,);
nor I_48(n4_1_r_0,n23_0,G199_2_r_9);
nor I_49(N3_2_r_0,n31_0,n32_0);
nor I_50(N1_4_r_0,n29_0,n32_0);
not I_51(n2_0,n31_0);
nor I_52(n21_0,n37_0,n_42_2_r_9);
not I_53(n22_0,n_573_1_r_9);
nand I_54(n23_0,n20_0,n30_0);
nand I_55(n24_0,n38_0,n25_0);
nor I_56(n25_0,n_42_2_r_9,G199_2_r_9);
not I_57(n26_0,G199_2_r_9);
not I_58(n27_0,n29_0);
nor I_59(n28_0,G199_4_r_9,G42_1_r_9);
nand I_60(n29_0,n26_0,n33_0);
not I_61(n30_0,n_42_2_r_9);
nand I_62(n31_0,ACVQN1_3_l_0,n_572_1_r_9);
and I_63(n32_0,n35_0,n36_0);
nand I_64(n33_0,n34_0,n_572_1_r_9);
not I_65(n34_0,G199_4_r_9);
nor I_66(n35_0,n_549_1_r_9,G199_4_r_9);
nor I_67(n36_0,n_573_1_r_9,G42_1_r_9);
endmodule


