module test_final(G18_1_l_16,G15_1_l_16,IN_1_1_l_16,IN_4_1_l_16,IN_5_1_l_16,IN_7_1_l_16,IN_9_1_l_16,IN_10_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_4_3_l_16,blif_clk_net_1_r_0,blif_reset_net_1_r_0,G42_1_r_0,n_572_1_r_0,n_573_1_r_0,n_549_1_r_0,n_42_2_r_0,G199_2_r_0,G199_4_r_0,G214_4_r_0);
input G18_1_l_16,G15_1_l_16,IN_1_1_l_16,IN_4_1_l_16,IN_5_1_l_16,IN_7_1_l_16,IN_9_1_l_16,IN_10_1_l_16,IN_1_3_l_16,IN_2_3_l_16,IN_4_3_l_16,blif_clk_net_1_r_0,blif_reset_net_1_r_0;
output G42_1_r_0,n_572_1_r_0,n_573_1_r_0,n_549_1_r_0,n_42_2_r_0,G199_2_r_0,G199_4_r_0,G214_4_r_0;
wire G42_1_r_16,n_572_1_r_16,n_573_1_r_16,n_549_1_r_16,n_569_1_r_16,n_452_1_r_16,G199_4_r_16,G214_4_r_16,ACVQN1_5_r_16,P6_5_r_16,n4_1_l_16,n29_16,n16_internal_16,n16_16,ACVQN1_3_l_16,n4_1_r_16,N1_4_r_16,n6_16,n_573_1_l_16,n_452_1_l_16,P6_5_r_internal_16,n18_16,n19_16,n20_16,n21_16,n22_16,n23_16,n24_16,n25_16,n26_16,n27_16,n28_16,n_569_1_r_0,n4_1_l_0,n6_0,n37_0,n38_0,n20_0,ACVQN1_3_l_0,n4_1_r_0,N3_2_r_0,N1_4_r_0,n2_0,n21_0,n22_0,n23_0,n24_0,n25_0,n26_0,n27_0,n28_0,n29_0,n30_0,n31_0,n32_0,n33_0,n34_0,n35_0,n36_0;
DFFARX1 I_0(n4_1_r_16,blif_clk_net_1_r_0,n6_0,G42_1_r_16,);
nor I_1(n_572_1_r_16,n20_16,n21_16);
nand I_2(n_573_1_r_16,n18_16,n19_16);
nor I_3(n_549_1_r_16,n23_16,n24_16);
nand I_4(n_569_1_r_16,n18_16,n22_16);
nor I_5(n_452_1_r_16,n29_16,n6_16);
DFFARX1 I_6(N1_4_r_16,blif_clk_net_1_r_0,n6_0,G199_4_r_16,);
DFFARX1 I_7(n6_16,blif_clk_net_1_r_0,n6_0,G214_4_r_16,);
DFFARX1 I_8(n_573_1_l_16,blif_clk_net_1_r_0,n6_0,ACVQN1_5_r_16,);
not I_9(P6_5_r_16,P6_5_r_internal_16);
nor I_10(n4_1_l_16,G18_1_l_16,IN_1_1_l_16);
DFFARX1 I_11(n4_1_l_16,blif_clk_net_1_r_0,n6_0,n29_16,);
DFFARX1 I_12(IN_1_3_l_16,blif_clk_net_1_r_0,n6_0,n16_internal_16,);
not I_13(n16_16,n16_internal_16);
DFFARX1 I_14(IN_2_3_l_16,blif_clk_net_1_r_0,n6_0,ACVQN1_3_l_16,);
nor I_15(n4_1_r_16,n29_16,n21_16);
nor I_16(N1_4_r_16,n27_16,n28_16);
not I_17(n6_16,n19_16);
or I_18(n_573_1_l_16,IN_5_1_l_16,IN_9_1_l_16);
nor I_19(n_452_1_l_16,G18_1_l_16,IN_5_1_l_16);
DFFARX1 I_20(n_452_1_l_16,blif_clk_net_1_r_0,n6_0,P6_5_r_internal_16,);
not I_21(n18_16,n20_16);
nor I_22(n19_16,IN_9_1_l_16,IN_10_1_l_16);
nor I_23(n20_16,G15_1_l_16,IN_7_1_l_16);
nor I_24(n21_16,IN_10_1_l_16,n25_16);
nand I_25(n22_16,IN_4_3_l_16,ACVQN1_3_l_16);
not I_26(n23_16,n22_16);
nor I_27(n24_16,n16_16,n20_16);
nor I_28(n25_16,G15_1_l_16,n26_16);
not I_29(n26_16,IN_4_1_l_16);
and I_30(n27_16,IN_9_1_l_16,n29_16);
not I_31(n28_16,n_452_1_l_16);
DFFARX1 I_32(n4_1_r_0,blif_clk_net_1_r_0,n6_0,G42_1_r_0,);
nor I_33(n_572_1_r_0,n23_0,G42_1_r_16);
nand I_34(n_573_1_r_0,n21_0,n22_0);
nand I_35(n_549_1_r_0,n_569_1_r_0,n24_0);
nand I_36(n_569_1_r_0,n21_0,n26_0);
nor I_37(n_42_2_r_0,n27_0,n28_0);
DFFARX1 I_38(N3_2_r_0,blif_clk_net_1_r_0,n6_0,G199_2_r_0,);
DFFARX1 I_39(N1_4_r_0,blif_clk_net_1_r_0,n6_0,G199_4_r_0,);
DFFARX1 I_40(n2_0,blif_clk_net_1_r_0,n6_0,G214_4_r_0,);
nor I_41(n4_1_l_0,n_569_1_r_16,G199_4_r_16);
not I_42(n6_0,blif_reset_net_1_r_0);
DFFARX1 I_43(n4_1_l_0,blif_clk_net_1_r_0,n6_0,n37_0,);
DFFARX1 I_44(G42_1_r_16,blif_clk_net_1_r_0,n6_0,n38_0,);
not I_45(n20_0,n38_0);
DFFARX1 I_46(n_549_1_r_16,blif_clk_net_1_r_0,n6_0,ACVQN1_3_l_0,);
nor I_47(n4_1_r_0,n23_0,P6_5_r_16);
nor I_48(N3_2_r_0,n31_0,n32_0);
nor I_49(N1_4_r_0,n29_0,n32_0);
not I_50(n2_0,n31_0);
nor I_51(n21_0,n37_0,n_573_1_r_16);
not I_52(n22_0,G42_1_r_16);
nand I_53(n23_0,n20_0,n30_0);
nand I_54(n24_0,n38_0,n25_0);
nor I_55(n25_0,n_573_1_r_16,P6_5_r_16);
not I_56(n26_0,P6_5_r_16);
not I_57(n27_0,n29_0);
nor I_58(n28_0,G214_4_r_16,ACVQN1_5_r_16);
nand I_59(n29_0,n26_0,n33_0);
not I_60(n30_0,n_573_1_r_16);
nand I_61(n31_0,ACVQN1_3_l_0,n_572_1_r_16);
and I_62(n32_0,n35_0,n36_0);
nand I_63(n33_0,n34_0,n_452_1_r_16);
not I_64(n34_0,ACVQN1_5_r_16);
nor I_65(n35_0,n_569_1_r_16,ACVQN1_5_r_16);
nor I_66(n36_0,G214_4_r_16,G42_1_r_16);
endmodule


