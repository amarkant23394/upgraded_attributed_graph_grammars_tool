module test_final(IN_1_1_l_8,IN_2_1_l_8,IN_3_1_l_8,IN_1_3_l_8,IN_2_3_l_8,IN_3_3_l_8,IN_1_6_l_8,IN_2_6_l_8,IN_3_6_l_8,IN_4_6_l_8,IN_5_6_l_8,IN_1_8_l_8,IN_2_8_l_8,IN_3_8_l_8,IN_6_8_l_8,blif_clk_net_7_r_1,blif_reset_net_7_r_1,N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,N6147_9_r_1,N6134_9_r_1);
input IN_1_1_l_8,IN_2_1_l_8,IN_3_1_l_8,IN_1_3_l_8,IN_2_3_l_8,IN_3_3_l_8,IN_1_6_l_8,IN_2_6_l_8,IN_3_6_l_8,IN_4_6_l_8,IN_5_6_l_8,IN_1_8_l_8,IN_2_8_l_8,IN_3_8_l_8,IN_6_8_l_8,blif_clk_net_7_r_1,blif_reset_net_7_r_1;
output N1508_0_r_1,N1507_6_r_1,N1508_6_r_1,G42_7_r_1,n_572_7_r_1,n_573_7_r_1,n_549_7_r_1,n_569_7_r_1,N6147_9_r_1,N6134_9_r_1;
wire N1371_0_r_8,N1508_0_r_8,N1372_1_r_8,N1508_1_r_8,N1507_6_r_8,N1508_6_r_8,n_42_8_r_8,G199_8_r_8,N6147_9_r_8,N6134_9_r_8,I_BUFF_1_9_r_8,N1372_10_r_8,N1508_10_r_8,N3_8_l_8,n53_8,n29_8,N3_8_r_8,n30_8,n31_8,n32_8,n33_8,n34_8,n35_8,n36_8,n37_8,n38_8,n39_8,n40_8,n41_8,n42_8,n43_8,n44_8,n45_8,n46_8,n47_8,n48_8,n49_8,n50_8,n51_8,n52_8,N1371_0_r_1,n_452_7_r_1,I_BUFF_1_9_r_1,n4_7_r_1,n9_1,n29_1,n30_1,n31_1,n32_1,n33_1,n34_1,n35_1,n36_1,n37_1,n38_1,n39_1,n40_1,n41_1,n42_1,n43_1,n44_1,n45_1,n46_1,n47_1,n48_1,n49_1,n50_1,n51_1,n52_1,n53_1,n54_1,n55_1;
nor I_0(N1371_0_r_8,n46_8,n51_8);
not I_1(N1508_0_r_8,n46_8);
nor I_2(N1372_1_r_8,n37_8,n49_8);
and I_3(N1508_1_r_8,N1372_1_r_8,n29_8);
nor I_4(N1507_6_r_8,n47_8,n48_8);
nor I_5(N1508_6_r_8,n37_8,n38_8);
nor I_6(n_42_8_r_8,I_BUFF_1_9_r_8,n53_8);
DFFARX1 I_7(N3_8_r_8,blif_clk_net_7_r_1,n9_1,G199_8_r_8,);
nor I_8(N6147_9_r_8,n29_8,n30_8);
nor I_9(N6134_9_r_8,n30_8,n31_8);
not I_10(I_BUFF_1_9_r_8,n35_8);
nor I_11(N1372_10_r_8,n46_8,n49_8);
nor I_12(N1508_10_r_8,n40_8,n41_8);
and I_13(N3_8_l_8,IN_6_8_l_8,n36_8);
DFFARX1 I_14(N3_8_l_8,blif_clk_net_7_r_1,n9_1,n53_8,);
not I_15(n29_8,n53_8);
nor I_16(N3_8_r_8,n33_8,n34_8);
and I_17(n30_8,n32_8,n33_8);
nor I_18(n31_8,IN_1_8_l_8,IN_3_8_l_8);
nand I_19(n32_8,IN_2_6_l_8,n42_8);
or I_20(n33_8,IN_3_1_l_8,n46_8);
nor I_21(n34_8,n32_8,n35_8);
nand I_22(n35_8,IN_5_6_l_8,n44_8);
nand I_23(n36_8,IN_2_8_l_8,IN_3_8_l_8);
not I_24(n37_8,n31_8);
nand I_25(n38_8,N1508_0_r_8,n39_8);
nand I_26(n39_8,n33_8,n50_8);
and I_27(n40_8,n32_8,n35_8);
not I_28(n41_8,N1372_10_r_8);
and I_29(n42_8,IN_1_6_l_8,n43_8);
nand I_30(n43_8,n44_8,n45_8);
nand I_31(n44_8,IN_3_6_l_8,IN_4_6_l_8);
not I_32(n45_8,IN_5_6_l_8);
nand I_33(n46_8,IN_1_1_l_8,IN_2_1_l_8);
not I_34(n47_8,n39_8);
nor I_35(n48_8,n35_8,n49_8);
not I_36(n49_8,n51_8);
nand I_37(n50_8,I_BUFF_1_9_r_8,n51_8);
nor I_38(n51_8,IN_1_3_l_8,n52_8);
or I_39(n52_8,IN_2_3_l_8,IN_3_3_l_8);
and I_40(N1371_0_r_1,I_BUFF_1_9_r_1,n55_1);
nor I_41(N1508_0_r_1,n40_1,n44_1);
nor I_42(N1507_6_r_1,n43_1,n49_1);
nor I_43(N1508_6_r_1,n41_1,n42_1);
DFFARX1 I_44(n4_7_r_1,blif_clk_net_7_r_1,n9_1,G42_7_r_1,);
nor I_45(n_572_7_r_1,n29_1,n30_1);
not I_46(n_573_7_r_1,n_452_7_r_1);
nor I_47(n_549_7_r_1,N1371_0_r_1,n31_1);
or I_48(n_569_7_r_1,n30_1,n31_1);
nor I_49(n_452_7_r_1,n30_1,n32_1);
nor I_50(N6147_9_r_1,n35_1,n36_1);
nand I_51(N6134_9_r_1,n38_1,n39_1);
not I_52(I_BUFF_1_9_r_1,n40_1);
nor I_53(n4_7_r_1,I_BUFF_1_9_r_1,n30_1);
not I_54(n9_1,blif_reset_net_7_r_1);
nor I_55(n29_1,n34_1,n_42_8_r_8);
nor I_56(n30_1,n33_1,n34_1);
nor I_57(n31_1,n54_1,N1508_1_r_8);
not I_58(n32_1,n48_1);
nor I_59(n33_1,N1508_6_r_8,N6134_9_r_8);
not I_60(n34_1,G199_8_r_8);
nor I_61(n35_1,I_BUFF_1_9_r_1,n37_1);
not I_62(n36_1,n29_1);
not I_63(n37_1,n41_1);
nand I_64(n38_1,I_BUFF_1_9_r_1,N1508_1_r_8);
nand I_65(n39_1,n37_1,n40_1);
nand I_66(n40_1,N1508_10_r_8,N1507_6_r_8);
nand I_67(n41_1,n52_1,N1508_6_r_8);
or I_68(n42_1,n36_1,n43_1);
nor I_69(n43_1,n32_1,n49_1);
nand I_70(n44_1,n45_1,n46_1);
nand I_71(n45_1,n47_1,n48_1);
not I_72(n46_1,N1508_1_r_8);
not I_73(n47_1,n31_1);
nand I_74(n48_1,n50_1,N6147_9_r_8);
nor I_75(n49_1,n41_1,n47_1);
and I_76(n50_1,n51_1,N1371_0_r_8);
nand I_77(n51_1,n52_1,n53_1);
nand I_78(n52_1,N1371_0_r_8,G199_8_r_8);
not I_79(n53_1,N1508_6_r_8);
or I_80(n54_1,N1507_6_r_8,n_42_8_r_8);
nor I_81(n55_1,n29_1,N1508_1_r_8);
endmodule


