module test_I14965(I1477,I14965);
input I1477;
output I14965;
wire ;
not I_0(I14965,I1477);
endmodule


