module test_I2861(I1351,I2861);
input I1351;
output I2861;
wire ;
not I_0(I2861,I1351);
endmodule


