module test_I9320(I1477,I1470,I6924,I9320);
input I1477,I1470,I6924;
output I9320;
wire I6875,I5088,I9303,I8862,I6907,I7221;
not I_0(I9320,I9303);
DFFARX1 I_1(I7221,I1470,I6907,,,I6875,);
DFFARX1 I_2(I1470,,,I5088,);
DFFARX1 I_3(I6875,I1470,I8862,,,I9303,);
not I_4(I8862,I1477);
not I_5(I6907,I1477);
nand I_6(I7221,I6924,I5088);
endmodule


