module test_I2776(I1407,I2776);
input I1407;
output I2776;
wire ;
not I_0(I2776,I1407);
endmodule


